// Benchmark "top" written by ABC on Mon Nov 27 17:21:25 2023

module top ( 
    A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15,
    A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28, A29,
    A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42, A43,
    A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56, A57,
    A58, A59, A60, A61, A62, A63, A64, A65, A66, A67, A68, A69, A70, A71,
    A72, A73, A74, A75, A76, A77, A78, A79, A80, A81, A82, A83, A84, A85,
    A86, A87, A88, A89, A90, A91, A92, A93, A94, A95, A96, A97, A98, A99,
    A100, A101, A102, A103, A104, A105, A106, A107, A108, A109, A110, A111,
    A112, A113, A114, A115, A116, A117, A118, A119, A120, A121, A122, A123,
    A124, A125, A126, A127,
    P0, P1, P2, P3, P4, P5, P6, F  );
  input  A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14,
    A15, A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28,
    A29, A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42,
    A43, A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56,
    A57, A58, A59, A60, A61, A62, A63, A64, A65, A66, A67, A68, A69, A70,
    A71, A72, A73, A74, A75, A76, A77, A78, A79, A80, A81, A82, A83, A84,
    A85, A86, A87, A88, A89, A90, A91, A92, A93, A94, A95, A96, A97, A98,
    A99, A100, A101, A102, A103, A104, A105, A106, A107, A108, A109, A110,
    A111, A112, A113, A114, A115, A116, A117, A118, A119, A120, A121, A122,
    A123, A124, A125, A126, A127;
  output P0, P1, P2, P3, P4, P5, P6, F;
  wire new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536;
  assign new_n137 = A116 & ~A117;
  assign new_n138 = ~A118 & ~new_n137;
  assign new_n139 = ~A119 & ~new_n138;
  assign new_n140 = ~A120 & ~new_n139;
  assign new_n141 = ~A121 & ~new_n140;
  assign new_n142 = ~A122 & ~new_n141;
  assign new_n143 = ~A123 & ~new_n142;
  assign new_n144 = ~A124 & ~new_n143;
  assign new_n145 = ~A125 & ~new_n144;
  assign new_n146 = ~A126 & ~new_n145;
  assign new_n147 = ~A127 & ~new_n146;
  assign new_n148 = ~A90 & ~A91;
  assign new_n149 = ~A88 & ~A89;
  assign new_n150 = new_n148 & new_n149;
  assign new_n151 = ~A94 & ~A95;
  assign new_n152 = ~A92 & ~A93;
  assign new_n153 = new_n151 & new_n152;
  assign new_n154 = new_n150 & new_n153;
  assign new_n155 = ~A80 & ~A81;
  assign new_n156 = ~A82 & ~A83;
  assign new_n157 = new_n155 & new_n156;
  assign new_n158 = ~A84 & ~A85;
  assign new_n159 = ~A86 & ~A87;
  assign new_n160 = new_n158 & new_n159;
  assign new_n161 = new_n157 & new_n160;
  assign new_n162 = new_n154 & new_n161;
  assign new_n163 = A74 & ~A75;
  assign new_n164 = ~A76 & ~new_n163;
  assign new_n165 = ~A77 & ~new_n164;
  assign new_n166 = ~A78 & ~new_n165;
  assign new_n167 = ~A79 & ~new_n166;
  assign new_n168 = new_n162 & ~new_n167;
  assign new_n169 = A81 & ~A82;
  assign new_n170 = ~A83 & ~new_n169;
  assign new_n171 = ~A84 & ~new_n170;
  assign new_n172 = ~A85 & ~new_n171;
  assign new_n173 = ~A86 & ~new_n172;
  assign new_n174 = ~A87 & ~new_n173;
  assign new_n175 = ~A88 & ~new_n174;
  assign new_n176 = ~A89 & ~new_n175;
  assign new_n177 = ~A90 & ~new_n176;
  assign new_n178 = ~A99 & ~A101;
  assign new_n179 = ~A91 & ~A93;
  assign new_n180 = ~A95 & ~A97;
  assign new_n181 = new_n179 & new_n180;
  assign new_n182 = new_n178 & new_n181;
  assign new_n183 = ~new_n177 & new_n182;
  assign new_n184 = ~new_n168 & new_n183;
  assign new_n185 = A92 & ~A93;
  assign new_n186 = ~A94 & ~new_n185;
  assign new_n187 = ~A95 & ~new_n186;
  assign new_n188 = ~A96 & ~new_n187;
  assign new_n189 = ~A97 & ~new_n188;
  assign new_n190 = ~A98 & ~new_n189;
  assign new_n191 = new_n178 & ~new_n190;
  assign new_n192 = A100 & ~A101;
  assign new_n193 = ~A112 & ~A114;
  assign new_n194 = A56 & ~A57;
  assign new_n195 = ~A58 & ~new_n194;
  assign new_n196 = ~A59 & ~new_n195;
  assign new_n197 = ~A60 & ~new_n196;
  assign new_n198 = ~A61 & ~new_n197;
  assign new_n199 = ~A62 & ~new_n198;
  assign new_n200 = ~A63 & ~new_n199;
  assign new_n201 = ~A64 & ~new_n200;
  assign new_n202 = ~A65 & ~new_n201;
  assign new_n203 = ~A66 & ~new_n202;
  assign new_n204 = ~A67 & ~new_n203;
  assign new_n205 = ~A68 & ~A70;
  assign new_n206 = ~A52 & ~A53;
  assign new_n207 = ~A54 & ~A55;
  assign new_n208 = new_n206 & new_n207;
  assign new_n209 = ~A50 & ~A51;
  assign new_n210 = ~A48 & ~A49;
  assign new_n211 = new_n209 & new_n210;
  assign new_n212 = new_n208 & new_n211;
  assign new_n213 = ~A24 & ~A26;
  assign new_n214 = A1 & ~A2;
  assign new_n215 = ~A3 & ~new_n214;
  assign new_n216 = ~A4 & ~new_n215;
  assign new_n217 = ~A5 & ~new_n216;
  assign new_n218 = ~A6 & ~new_n217;
  assign new_n219 = ~A7 & ~new_n218;
  assign new_n220 = ~A8 & ~new_n219;
  assign new_n221 = ~A9 & ~new_n220;
  assign new_n222 = ~A10 & ~new_n221;
  assign new_n223 = ~A11 & ~new_n222;
  assign new_n224 = ~A12 & ~new_n223;
  assign new_n225 = ~A13 & ~new_n224;
  assign new_n226 = ~A14 & ~new_n225;
  assign new_n227 = ~A15 & ~new_n226;
  assign new_n228 = ~A16 & ~new_n227;
  assign new_n229 = ~A17 & ~new_n228;
  assign new_n230 = ~A18 & ~new_n229;
  assign new_n231 = ~A19 & ~new_n230;
  assign new_n232 = ~A20 & ~new_n231;
  assign new_n233 = ~A21 & ~new_n232;
  assign new_n234 = ~A22 & ~new_n233;
  assign new_n235 = ~A23 & ~new_n234;
  assign new_n236 = new_n213 & ~new_n235;
  assign new_n237 = A25 & ~A26;
  assign new_n238 = ~A27 & ~new_n237;
  assign new_n239 = ~new_n236 & new_n238;
  assign new_n240 = ~A28 & ~new_n239;
  assign new_n241 = ~A29 & ~new_n240;
  assign new_n242 = ~A30 & ~new_n241;
  assign new_n243 = ~A31 & ~new_n242;
  assign new_n244 = ~A32 & ~new_n243;
  assign new_n245 = ~A33 & ~new_n244;
  assign new_n246 = ~A34 & ~new_n245;
  assign new_n247 = ~A35 & ~new_n246;
  assign new_n248 = ~A36 & ~new_n247;
  assign new_n249 = ~A37 & ~new_n248;
  assign new_n250 = ~A38 & ~new_n249;
  assign new_n251 = ~A39 & ~new_n250;
  assign new_n252 = ~A40 & ~new_n251;
  assign new_n253 = ~A41 & ~new_n252;
  assign new_n254 = ~A42 & ~new_n253;
  assign new_n255 = ~A43 & ~new_n254;
  assign new_n256 = ~A44 & ~new_n255;
  assign new_n257 = ~A45 & ~new_n256;
  assign new_n258 = ~A46 & ~new_n257;
  assign new_n259 = ~A47 & ~new_n258;
  assign new_n260 = new_n212 & ~new_n259;
  assign new_n261 = A49 & ~A50;
  assign new_n262 = ~A51 & ~new_n261;
  assign new_n263 = ~A52 & ~new_n262;
  assign new_n264 = ~A53 & ~new_n263;
  assign new_n265 = ~A54 & ~new_n264;
  assign new_n266 = ~A55 & ~A57;
  assign new_n267 = ~A59 & ~A61;
  assign new_n268 = ~A63 & ~A65;
  assign new_n269 = ~A67 & new_n268;
  assign new_n270 = new_n266 & new_n267;
  assign new_n271 = new_n269 & new_n270;
  assign new_n272 = ~new_n265 & new_n271;
  assign new_n273 = ~new_n260 & new_n272;
  assign new_n274 = ~A72 & new_n205;
  assign new_n275 = ~new_n204 & new_n274;
  assign new_n276 = ~new_n273 & new_n275;
  assign new_n277 = A69 & ~A70;
  assign new_n278 = ~A71 & ~new_n277;
  assign new_n279 = ~A72 & ~new_n278;
  assign new_n280 = ~A73 & ~A75;
  assign new_n281 = ~A77 & ~A79;
  assign new_n282 = new_n280 & new_n281;
  assign new_n283 = ~new_n279 & new_n282;
  assign new_n284 = new_n183 & new_n283;
  assign new_n285 = ~new_n276 & new_n284;
  assign new_n286 = ~A102 & ~A104;
  assign new_n287 = ~A106 & ~A108;
  assign new_n288 = ~A110 & new_n287;
  assign new_n289 = ~new_n192 & new_n286;
  assign new_n290 = new_n193 & new_n289;
  assign new_n291 = new_n288 & new_n290;
  assign new_n292 = ~new_n191 & new_n291;
  assign new_n293 = ~new_n184 & new_n292;
  assign new_n294 = ~new_n285 & new_n293;
  assign new_n295 = ~A124 & ~A125;
  assign new_n296 = ~A126 & ~A127;
  assign new_n297 = new_n295 & new_n296;
  assign new_n298 = ~A122 & ~A123;
  assign new_n299 = ~A120 & ~A121;
  assign new_n300 = new_n298 & new_n299;
  assign new_n301 = new_n297 & new_n300;
  assign new_n302 = A103 & ~A104;
  assign new_n303 = ~A105 & ~new_n302;
  assign new_n304 = ~A106 & ~new_n303;
  assign new_n305 = ~A107 & ~new_n304;
  assign new_n306 = ~A108 & ~new_n305;
  assign new_n307 = ~A109 & ~new_n306;
  assign new_n308 = ~A110 & ~new_n307;
  assign new_n309 = ~A111 & ~new_n308;
  assign new_n310 = new_n193 & ~new_n309;
  assign new_n311 = A113 & ~A114;
  assign new_n312 = ~A115 & ~A117;
  assign new_n313 = ~A119 & new_n312;
  assign new_n314 = ~new_n311 & new_n313;
  assign new_n315 = new_n301 & new_n314;
  assign new_n316 = ~new_n310 & new_n315;
  assign new_n317 = ~new_n294 & new_n316;
  assign P0 = ~new_n147 & ~new_n317;
  assign new_n319 = new_n295 & ~new_n298;
  assign new_n320 = ~A112 & ~A113;
  assign new_n321 = ~A110 & ~A111;
  assign new_n322 = ~A78 & ~A79;
  assign new_n323 = ~A74 & ~A75;
  assign new_n324 = ~A72 & ~A73;
  assign new_n325 = ~A64 & ~A65;
  assign new_n326 = ~A60 & ~A61;
  assign new_n327 = ~A58 & ~A59;
  assign new_n328 = ~A56 & ~A57;
  assign new_n329 = ~new_n206 & new_n207;
  assign new_n330 = ~A44 & ~A45;
  assign new_n331 = ~A40 & ~A41;
  assign new_n332 = ~A36 & ~A37;
  assign new_n333 = ~A30 & ~A31;
  assign new_n334 = ~A28 & ~A29;
  assign new_n335 = ~A20 & ~A21;
  assign new_n336 = ~A16 & ~A17;
  assign new_n337 = ~A12 & ~A13;
  assign new_n338 = ~A8 & ~A9;
  assign new_n339 = ~A2 & ~A3;
  assign new_n340 = ~A4 & ~A5;
  assign new_n341 = ~new_n339 & new_n340;
  assign new_n342 = ~A6 & ~A7;
  assign new_n343 = ~new_n341 & new_n342;
  assign new_n344 = new_n338 & ~new_n343;
  assign new_n345 = ~A10 & ~A11;
  assign new_n346 = ~new_n344 & new_n345;
  assign new_n347 = new_n337 & ~new_n346;
  assign new_n348 = ~A14 & ~A15;
  assign new_n349 = ~new_n347 & new_n348;
  assign new_n350 = new_n336 & ~new_n349;
  assign new_n351 = ~A18 & ~A19;
  assign new_n352 = ~new_n350 & new_n351;
  assign new_n353 = new_n335 & ~new_n352;
  assign new_n354 = ~A22 & ~A23;
  assign new_n355 = ~new_n353 & new_n354;
  assign new_n356 = ~A24 & ~A25;
  assign new_n357 = ~new_n355 & new_n356;
  assign new_n358 = ~A26 & ~A27;
  assign new_n359 = ~new_n357 & new_n358;
  assign new_n360 = new_n334 & ~new_n359;
  assign new_n361 = new_n333 & ~new_n360;
  assign new_n362 = ~A32 & ~A33;
  assign new_n363 = ~new_n361 & new_n362;
  assign new_n364 = ~A34 & ~A35;
  assign new_n365 = ~new_n363 & new_n364;
  assign new_n366 = new_n332 & ~new_n365;
  assign new_n367 = ~A38 & ~A39;
  assign new_n368 = ~new_n366 & new_n367;
  assign new_n369 = new_n331 & ~new_n368;
  assign new_n370 = ~A42 & ~A43;
  assign new_n371 = ~new_n369 & new_n370;
  assign new_n372 = new_n330 & ~new_n371;
  assign new_n373 = ~A46 & ~A47;
  assign new_n374 = ~new_n372 & new_n373;
  assign new_n375 = new_n210 & ~new_n374;
  assign new_n376 = new_n207 & new_n209;
  assign new_n377 = ~new_n375 & new_n376;
  assign new_n378 = new_n328 & ~new_n329;
  assign new_n379 = ~new_n377 & new_n378;
  assign new_n380 = new_n327 & ~new_n379;
  assign new_n381 = new_n326 & ~new_n380;
  assign new_n382 = ~A62 & ~A63;
  assign new_n383 = ~new_n381 & new_n382;
  assign new_n384 = new_n325 & ~new_n383;
  assign new_n385 = ~A66 & ~A67;
  assign new_n386 = ~new_n384 & new_n385;
  assign new_n387 = ~A68 & ~A69;
  assign new_n388 = ~new_n386 & new_n387;
  assign new_n389 = ~A70 & ~A71;
  assign new_n390 = ~new_n388 & new_n389;
  assign new_n391 = new_n324 & ~new_n390;
  assign new_n392 = new_n322 & new_n323;
  assign new_n393 = ~new_n391 & new_n392;
  assign new_n394 = ~A76 & ~A77;
  assign new_n395 = new_n322 & ~new_n394;
  assign new_n396 = new_n155 & new_n158;
  assign new_n397 = ~new_n395 & new_n396;
  assign new_n398 = ~new_n393 & new_n397;
  assign new_n399 = ~new_n156 & new_n158;
  assign new_n400 = new_n148 & new_n159;
  assign new_n401 = ~new_n399 & new_n400;
  assign new_n402 = ~new_n398 & new_n401;
  assign new_n403 = new_n148 & ~new_n149;
  assign new_n404 = ~A100 & ~A101;
  assign new_n405 = ~A96 & ~A97;
  assign new_n406 = new_n404 & new_n405;
  assign new_n407 = new_n152 & ~new_n403;
  assign new_n408 = new_n406 & new_n407;
  assign new_n409 = ~new_n402 & new_n408;
  assign new_n410 = ~A98 & ~A99;
  assign new_n411 = new_n404 & ~new_n410;
  assign new_n412 = ~A106 & ~A107;
  assign new_n413 = ~new_n151 & new_n406;
  assign new_n414 = ~A102 & ~A103;
  assign new_n415 = new_n412 & new_n414;
  assign new_n416 = ~new_n411 & new_n415;
  assign new_n417 = ~new_n413 & new_n416;
  assign new_n418 = ~new_n409 & new_n417;
  assign new_n419 = ~A104 & ~A105;
  assign new_n420 = new_n412 & ~new_n419;
  assign new_n421 = ~A108 & ~A109;
  assign new_n422 = ~new_n420 & new_n421;
  assign new_n423 = ~new_n418 & new_n422;
  assign new_n424 = new_n321 & ~new_n423;
  assign new_n425 = new_n320 & ~new_n424;
  assign new_n426 = ~A114 & ~A115;
  assign new_n427 = ~new_n425 & new_n426;
  assign new_n428 = ~A116 & ~A117;
  assign new_n429 = ~new_n427 & new_n428;
  assign new_n430 = ~A118 & ~A119;
  assign new_n431 = ~new_n429 & new_n430;
  assign new_n432 = new_n301 & ~new_n431;
  assign new_n433 = new_n296 & ~new_n319;
  assign P1 = new_n432 | ~new_n433;
  assign new_n435 = new_n321 & new_n421;
  assign new_n436 = new_n412 & new_n419;
  assign new_n437 = new_n404 & new_n414;
  assign new_n438 = new_n405 & new_n410;
  assign new_n439 = new_n325 & new_n385;
  assign new_n440 = new_n326 & new_n382;
  assign new_n441 = new_n330 & new_n373;
  assign new_n442 = new_n331 & new_n370;
  assign new_n443 = new_n332 & new_n367;
  assign new_n444 = new_n333 & new_n334;
  assign new_n445 = new_n335 & new_n354;
  assign new_n446 = new_n336 & new_n351;
  assign new_n447 = new_n337 & new_n348;
  assign new_n448 = new_n340 & new_n342;
  assign new_n449 = new_n338 & new_n345;
  assign new_n450 = ~new_n448 & new_n449;
  assign new_n451 = new_n447 & ~new_n450;
  assign new_n452 = new_n446 & ~new_n451;
  assign new_n453 = new_n445 & ~new_n452;
  assign new_n454 = new_n213 & new_n238;
  assign new_n455 = ~new_n453 & new_n454;
  assign new_n456 = new_n444 & ~new_n455;
  assign new_n457 = new_n362 & new_n364;
  assign new_n458 = ~new_n456 & new_n457;
  assign new_n459 = new_n443 & ~new_n458;
  assign new_n460 = new_n442 & ~new_n459;
  assign new_n461 = new_n441 & ~new_n460;
  assign new_n462 = new_n211 & ~new_n461;
  assign new_n463 = new_n208 & ~new_n462;
  assign new_n464 = new_n327 & new_n328;
  assign new_n465 = ~new_n463 & new_n464;
  assign new_n466 = new_n440 & ~new_n465;
  assign new_n467 = new_n439 & ~new_n466;
  assign new_n468 = new_n205 & new_n278;
  assign new_n469 = ~new_n467 & new_n468;
  assign new_n470 = new_n323 & new_n324;
  assign new_n471 = ~new_n469 & new_n470;
  assign new_n472 = new_n322 & new_n394;
  assign new_n473 = ~new_n471 & new_n472;
  assign new_n474 = new_n157 & ~new_n473;
  assign new_n475 = new_n160 & ~new_n474;
  assign new_n476 = new_n150 & ~new_n475;
  assign new_n477 = new_n153 & ~new_n476;
  assign new_n478 = new_n438 & ~new_n477;
  assign new_n479 = new_n437 & ~new_n478;
  assign new_n480 = new_n436 & ~new_n479;
  assign new_n481 = new_n435 & ~new_n480;
  assign new_n482 = new_n320 & new_n426;
  assign new_n483 = ~new_n481 & new_n482;
  assign new_n484 = new_n428 & new_n430;
  assign new_n485 = ~new_n483 & new_n484;
  assign new_n486 = new_n300 & ~new_n485;
  assign P2 = ~new_n297 | new_n486;
  assign new_n488 = new_n482 & new_n484;
  assign new_n489 = new_n435 & new_n436;
  assign new_n490 = new_n488 & ~new_n489;
  assign new_n491 = new_n301 & new_n488;
  assign new_n492 = new_n437 & new_n438;
  assign new_n493 = new_n489 & new_n492;
  assign new_n494 = new_n491 & new_n493;
  assign new_n495 = new_n470 & new_n472;
  assign new_n496 = new_n439 & new_n468;
  assign new_n497 = new_n440 & new_n464;
  assign new_n498 = new_n441 & new_n442;
  assign new_n499 = new_n443 & new_n457;
  assign new_n500 = new_n444 & new_n454;
  assign new_n501 = new_n447 & new_n449;
  assign new_n502 = new_n445 & new_n446;
  assign new_n503 = ~new_n501 & new_n502;
  assign new_n504 = new_n500 & ~new_n503;
  assign new_n505 = new_n499 & ~new_n504;
  assign new_n506 = new_n498 & ~new_n505;
  assign new_n507 = new_n212 & ~new_n506;
  assign new_n508 = new_n497 & ~new_n507;
  assign new_n509 = new_n496 & ~new_n508;
  assign new_n510 = new_n495 & ~new_n509;
  assign new_n511 = new_n161 & ~new_n510;
  assign new_n512 = new_n154 & ~new_n511;
  assign new_n513 = new_n494 & ~new_n512;
  assign new_n514 = new_n301 & ~new_n490;
  assign P3 = new_n513 | ~new_n514;
  assign new_n516 = new_n495 & new_n496;
  assign new_n517 = new_n212 & new_n497;
  assign new_n518 = new_n500 & new_n502;
  assign new_n519 = new_n498 & new_n499;
  assign new_n520 = ~new_n518 & new_n519;
  assign new_n521 = new_n517 & ~new_n520;
  assign new_n522 = new_n516 & ~new_n521;
  assign new_n523 = new_n162 & ~new_n522;
  assign new_n524 = new_n493 & ~new_n523;
  assign P4 = ~new_n491 | new_n524;
  assign new_n526 = new_n517 & new_n519;
  assign new_n527 = new_n162 & new_n516;
  assign new_n528 = ~new_n526 & new_n527;
  assign P5 = ~new_n494 | new_n528;
  assign P6 = ~new_n494 | ~new_n527;
  assign new_n531 = ~A0 & ~A1;
  assign new_n532 = new_n339 & new_n531;
  assign new_n533 = new_n448 & new_n532;
  assign new_n534 = new_n501 & new_n533;
  assign new_n535 = new_n518 & new_n534;
  assign new_n536 = new_n526 & new_n535;
  assign F = P6 | ~new_n536;
endmodule


