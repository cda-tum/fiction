// Benchmark "top" written by ABC on Mon Nov 27 16:50:38 2023

module top ( 
    \1 , \4 , \11 , \14 , \17 , \20 , \23 , \24 , \25 , \26 , \27 , \31 ,
    \34 , \37 , \40 , \43 , \46 , \49 , \52 , \53 , \54 , \61 , \64 , \67 ,
    \70 , \73 , \76 , \79 , \80 , \81 , \82 , \83 , \86 , \87 , \88 , \91 ,
    \94 , \97 , \100 , \103 , \106 , \109 , \112 , \113 , \114 , \115 ,
    \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 , \126 , \127 ,
    \128 , \129 , \130 , \131 , \132 , \135 , \136 , \137 , \140 , \141 ,
    \145 , \146 , \149 , \152 , \155 , \158 , \161 , \164 , \167 , \170 ,
    \173 , \176 , \179 , \182 , \185 , \188 , \191 , \194 , \197 , \200 ,
    \203 , \206 , \209 , \210 , \217 , \218 , \225 , \226 , \233 , \234 ,
    \241 , \242 , \245 , \248 , \251 , \254 , \257 , \264 , \265 , \272 ,
    \273 , \280 , \281 , \288 , \289 , \292 , \293 , \299 , \302 , \307 ,
    \308 , \315 , \316 , \323 , \324 , \331 , \332 , \335 , \338 , \341 ,
    \348 , \351 , \358 , \361 , \366 , \369 , \372 , \373 , \374 , \386 ,
    \389 , \400 , \411 , \422 , \435 , \446 , \457 , \468 , \479 , \490 ,
    \503 , \514 , \523 , \534 , \545 , \549 , \552 , \556 , \559 , \562 ,
    \566 , \571 , \574 , \577 , \580 , \583 , \588 , \591 , \592 , \595 ,
    \596 , \597 , \598 , \599 , \603 , \607 , \610 , \613 , \616 , \619 ,
    \625 , \631 ,
    \709 , \816 , \1066 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
    \1143 , \1144 , \1145 , \1147 , \1152 , \1153 , \1154 , \1155 , \1972 ,
    \2054 , \2060 , \2061 , \2139 , \2142 , \2309 , \2387 , \2527 , \2584 ,
    \2590 , \2623 , \3357 , \3358 , \3359 , \3360 , \3604 , \3613 , \4272 ,
    \4275 , \4278 , \4279 , \4737 , \4738 , \4739 , \4740 , \5240 , \5388 ,
    \6641 , \6643 , \6646 , \6648 , \6716 , \6877 , \6924 , \6925 , \6926 ,
    \6927 , \7015 , \7363 , \7365 , \7432 , \7449 , \7465 , \7466 , \7467 ,
    \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7476 , \7503 , \7504 ,
    \7506 , \7511 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
    \7522 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
    \7626 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 ,
    \7706 , \7707 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 ,
    \7742 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
    \8075 , \8076 , \8123 , \8124 , \8127 , \8128   );
  input  \1 , \4 , \11 , \14 , \17 , \20 , \23 , \24 , \25 , \26 , \27 ,
    \31 , \34 , \37 , \40 , \43 , \46 , \49 , \52 , \53 , \54 , \61 , \64 ,
    \67 , \70 , \73 , \76 , \79 , \80 , \81 , \82 , \83 , \86 , \87 , \88 ,
    \91 , \94 , \97 , \100 , \103 , \106 , \109 , \112 , \113 , \114 ,
    \115 , \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 , \126 ,
    \127 , \128 , \129 , \130 , \131 , \132 , \135 , \136 , \137 , \140 ,
    \141 , \145 , \146 , \149 , \152 , \155 , \158 , \161 , \164 , \167 ,
    \170 , \173 , \176 , \179 , \182 , \185 , \188 , \191 , \194 , \197 ,
    \200 , \203 , \206 , \209 , \210 , \217 , \218 , \225 , \226 , \233 ,
    \234 , \241 , \242 , \245 , \248 , \251 , \254 , \257 , \264 , \265 ,
    \272 , \273 , \280 , \281 , \288 , \289 , \292 , \293 , \299 , \302 ,
    \307 , \308 , \315 , \316 , \323 , \324 , \331 , \332 , \335 , \338 ,
    \341 , \348 , \351 , \358 , \361 , \366 , \369 , \372 , \373 , \374 ,
    \386 , \389 , \400 , \411 , \422 , \435 , \446 , \457 , \468 , \479 ,
    \490 , \503 , \514 , \523 , \534 , \545 , \549 , \552 , \556 , \559 ,
    \562 , \566 , \571 , \574 , \577 , \580 , \583 , \588 , \591 , \592 ,
    \595 , \596 , \597 , \598 , \599 , \603 , \607 , \610 , \613 , \616 ,
    \619 , \625 , \631 ;
  output \709 , \816 , \1066 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
    \1143 , \1144 , \1145 , \1147 , \1152 , \1153 , \1154 , \1155 , \1972 ,
    \2054 , \2060 , \2061 , \2139 , \2142 , \2309 , \2387 , \2527 , \2584 ,
    \2590 , \2623 , \3357 , \3358 , \3359 , \3360 , \3604 , \3613 , \4272 ,
    \4275 , \4278 , \4279 , \4737 , \4738 , \4739 , \4740 , \5240 , \5388 ,
    \6641 , \6643 , \6646 , \6648 , \6716 , \6877 , \6924 , \6925 , \6926 ,
    \6927 , \7015 , \7363 , \7365 , \7432 , \7449 , \7465 , \7466 , \7467 ,
    \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7476 , \7503 , \7504 ,
    \7506 , \7511 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
    \7522 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
    \7626 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 ,
    \7706 , \7707 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 ,
    \7742 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
    \8075 , \8076 , \8123 , \8124 , \8127 , \8128 ;
  wire new_n310, new_n311, new_n312, new_n313, new_n315, new_n316, new_n319,
    new_n320, new_n321, new_n323, new_n324, new_n325, new_n327, new_n328,
    new_n329, new_n331, new_n332, new_n333, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1116, new_n1117, new_n1118, new_n1119, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495, new_n1496, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1501, new_n1502, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556;
  assign \1140  = \552  & \562 ;
  assign \1147  = \141  & \145 ;
  assign \1972  = \1  & \373 ;
  assign \2054  = \136  & ~\592 ;
  assign \2060  = ~\27  | \591 ;
  assign \2061  = ~\386  | ~\556 ;
  assign \2623  = ~\27  | ~\31 ;
  assign \2590  = ~\140  | \2623 ;
  assign new_n310 = \588  & ~\2623 ;
  assign new_n311 = \87  & new_n310;
  assign new_n312 = ~\588  & ~\2623 ;
  assign new_n313 = \86  & new_n312;
  assign \4272  = ~new_n311 & ~new_n313;
  assign new_n315 = \88  & new_n312;
  assign new_n316 = \34  & new_n310;
  assign \4275  = ~new_n315 & ~new_n316;
  assign \4279  = ~\83  | \2623 ;
  assign new_n319 = ~\25  & new_n310;
  assign new_n320 = ~\24  & new_n312;
  assign new_n321 = \141  & ~new_n319;
  assign \4737  = ~new_n320 & new_n321;
  assign new_n323 = ~\81  & new_n310;
  assign new_n324 = ~\26  & new_n312;
  assign new_n325 = \141  & ~new_n323;
  assign \4738  = ~new_n324 & new_n325;
  assign new_n327 = ~\79  & new_n312;
  assign new_n328 = ~\23  & new_n310;
  assign new_n329 = \141  & ~new_n327;
  assign \4739  = ~new_n328 & new_n329;
  assign new_n331 = ~\82  & new_n312;
  assign new_n332 = ~\80  & new_n310;
  assign new_n333 = \141  & ~new_n331;
  assign \4740  = ~new_n332 & new_n333;
  assign new_n335 = \503  & ~\598 ;
  assign new_n336 = ~\503  & \595 ;
  assign new_n337 = \324  & ~new_n335;
  assign new_n338 = ~new_n336 & new_n337;
  assign new_n339 = \503  & ~\597 ;
  assign new_n340 = ~\503  & \596 ;
  assign new_n341 = ~\324  & ~new_n339;
  assign new_n342 = ~new_n340 & new_n341;
  assign new_n343 = ~new_n338 & ~new_n342;
  assign new_n344 = \523  & ~\598 ;
  assign new_n345 = ~\523  & \595 ;
  assign new_n346 = \341  & ~new_n344;
  assign new_n347 = ~new_n345 & new_n346;
  assign new_n348 = \523  & ~\597 ;
  assign new_n349 = ~\523  & \596 ;
  assign new_n350 = ~\341  & ~new_n348;
  assign new_n351 = ~new_n349 & new_n350;
  assign new_n352 = ~new_n347 & ~new_n351;
  assign new_n353 = \534  & ~\598 ;
  assign new_n354 = ~\534  & \595 ;
  assign new_n355 = \351  & ~new_n353;
  assign new_n356 = ~new_n354 & new_n355;
  assign new_n357 = \534  & ~\597 ;
  assign new_n358 = ~\534  & \596 ;
  assign new_n359 = ~\351  & ~new_n357;
  assign new_n360 = ~new_n358 & new_n359;
  assign new_n361 = ~new_n356 & ~new_n360;
  assign new_n362 = ~\248  & \490 ;
  assign new_n363 = \242  & ~\490 ;
  assign new_n364 = \316  & ~new_n362;
  assign new_n365 = ~new_n363 & new_n364;
  assign new_n366 = ~\251  & \490 ;
  assign new_n367 = \254  & ~\490 ;
  assign new_n368 = ~\316  & ~new_n366;
  assign new_n369 = ~new_n367 & new_n368;
  assign new_n370 = ~new_n365 & ~new_n369;
  assign new_n371 = ~\248  & \479 ;
  assign new_n372 = \242  & ~\479 ;
  assign new_n373 = \308  & ~new_n371;
  assign new_n374 = ~new_n372 & new_n373;
  assign new_n375 = ~\251  & \479 ;
  assign new_n376 = \254  & ~\479 ;
  assign new_n377 = ~\308  & ~new_n375;
  assign new_n378 = ~new_n376 & new_n377;
  assign new_n379 = ~new_n374 & ~new_n378;
  assign new_n380 = ~new_n370 & ~new_n379;
  assign new_n381 = ~\251  & ~\302 ;
  assign new_n382 = ~\248  & \302 ;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = ~\254  & ~\293 ;
  assign new_n385 = ~\242  & \293 ;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = ~\251  & ~\361 ;
  assign new_n388 = ~\248  & \361 ;
  assign new_n389 = ~new_n387 & ~new_n388;
  assign new_n390 = ~new_n386 & new_n389;
  assign new_n391 = \514  & ~\598 ;
  assign new_n392 = ~\514  & \595 ;
  assign new_n393 = ~new_n391 & ~new_n392;
  assign new_n394 = new_n383 & ~new_n393;
  assign new_n395 = new_n390 & new_n394;
  assign new_n396 = new_n343 & new_n395;
  assign new_n397 = new_n352 & new_n361;
  assign new_n398 = new_n396 & new_n397;
  assign \5240  = new_n380 & new_n398;
  assign new_n400 = \374  & ~\598 ;
  assign new_n401 = ~\374  & \595 ;
  assign new_n402 = \281  & ~new_n400;
  assign new_n403 = ~new_n401 & new_n402;
  assign new_n404 = \374  & ~\597 ;
  assign new_n405 = ~\374  & \596 ;
  assign new_n406 = ~\281  & ~new_n404;
  assign new_n407 = ~new_n405 & new_n406;
  assign new_n408 = ~new_n403 & ~new_n407;
  assign new_n409 = \400  & ~\598 ;
  assign new_n410 = ~\400  & \595 ;
  assign new_n411 = \265  & ~new_n409;
  assign new_n412 = ~new_n410 & new_n411;
  assign new_n413 = \400  & ~\597 ;
  assign new_n414 = ~\400  & \596 ;
  assign new_n415 = ~\265  & ~new_n413;
  assign new_n416 = ~new_n414 & new_n415;
  assign new_n417 = ~new_n412 & ~new_n416;
  assign new_n418 = \422  & ~\598 ;
  assign new_n419 = ~\422  & \595 ;
  assign new_n420 = \226  & ~new_n418;
  assign new_n421 = ~new_n419 & new_n420;
  assign new_n422 = \422  & ~\597 ;
  assign new_n423 = ~\422  & \596 ;
  assign new_n424 = ~\226  & ~new_n422;
  assign new_n425 = ~new_n423 & new_n424;
  assign new_n426 = ~new_n421 & ~new_n425;
  assign new_n427 = \457  & ~\598 ;
  assign new_n428 = ~\457  & \595 ;
  assign new_n429 = \210  & ~new_n427;
  assign new_n430 = ~new_n428 & new_n429;
  assign new_n431 = \457  & ~\597 ;
  assign new_n432 = ~\457  & \596 ;
  assign new_n433 = ~\210  & ~new_n431;
  assign new_n434 = ~new_n432 & new_n433;
  assign new_n435 = ~new_n430 & ~new_n434;
  assign new_n436 = \468  & ~\598 ;
  assign new_n437 = ~\468  & \595 ;
  assign new_n438 = \218  & ~new_n436;
  assign new_n439 = ~new_n437 & new_n438;
  assign new_n440 = \468  & ~\597 ;
  assign new_n441 = ~\468  & \596 ;
  assign new_n442 = ~\218  & ~new_n440;
  assign new_n443 = ~new_n441 & new_n442;
  assign new_n444 = ~new_n439 & ~new_n443;
  assign new_n445 = \435  & ~\598 ;
  assign new_n446 = ~\435  & \595 ;
  assign new_n447 = \234  & ~new_n445;
  assign new_n448 = ~new_n446 & new_n447;
  assign new_n449 = \435  & ~\597 ;
  assign new_n450 = ~\435  & \596 ;
  assign new_n451 = ~\234  & ~new_n449;
  assign new_n452 = ~new_n450 & new_n451;
  assign new_n453 = ~new_n448 & ~new_n452;
  assign new_n454 = ~\248  & \446 ;
  assign new_n455 = \242  & ~\446 ;
  assign new_n456 = \206  & ~new_n454;
  assign new_n457 = ~new_n455 & new_n456;
  assign new_n458 = ~\251  & \446 ;
  assign new_n459 = \254  & ~\446 ;
  assign new_n460 = ~\206  & ~new_n458;
  assign new_n461 = ~new_n459 & new_n460;
  assign new_n462 = ~new_n457 & ~new_n461;
  assign new_n463 = \411  & ~\598 ;
  assign new_n464 = ~\411  & \595 ;
  assign new_n465 = \273  & ~new_n463;
  assign new_n466 = ~new_n464 & new_n465;
  assign new_n467 = \411  & ~\597 ;
  assign new_n468 = ~\411  & \596 ;
  assign new_n469 = ~\273  & ~new_n467;
  assign new_n470 = ~new_n468 & new_n469;
  assign new_n471 = ~new_n466 & ~new_n470;
  assign new_n472 = \389  & ~\598 ;
  assign new_n473 = ~\389  & \595 ;
  assign new_n474 = \257  & ~new_n472;
  assign new_n475 = ~new_n473 & new_n474;
  assign new_n476 = \389  & ~\597 ;
  assign new_n477 = ~\389  & \596 ;
  assign new_n478 = ~\257  & ~new_n476;
  assign new_n479 = ~new_n477 & new_n478;
  assign new_n480 = ~new_n475 & ~new_n479;
  assign new_n481 = new_n408 & new_n417;
  assign new_n482 = new_n426 & new_n435;
  assign new_n483 = new_n444 & new_n453;
  assign new_n484 = ~new_n462 & new_n471;
  assign new_n485 = new_n480 & new_n484;
  assign new_n486 = new_n482 & new_n483;
  assign new_n487 = new_n481 & new_n486;
  assign \5388  = new_n485 & new_n487;
  assign new_n489 = ~\217  & \335 ;
  assign new_n490 = ~\210  & ~\335 ;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = ~\457  & ~new_n491;
  assign new_n493 = ~\225  & \335 ;
  assign new_n494 = ~\218  & ~\335 ;
  assign new_n495 = ~new_n493 & ~new_n494;
  assign new_n496 = ~\468  & ~new_n495;
  assign new_n497 = \468  & new_n495;
  assign new_n498 = ~\233  & \335 ;
  assign new_n499 = ~\226  & ~\335 ;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = ~\422  & ~new_n500;
  assign new_n502 = ~new_n497 & new_n501;
  assign new_n503 = ~new_n496 & ~new_n502;
  assign new_n504 = ~new_n492 & new_n503;
  assign new_n505 = ~\264  & \335 ;
  assign new_n506 = ~\257  & ~\335 ;
  assign new_n507 = ~new_n505 & ~new_n506;
  assign new_n508 = ~\389  & ~new_n507;
  assign new_n509 = ~\272  & \335 ;
  assign new_n510 = ~\265  & ~\335 ;
  assign new_n511 = ~new_n509 & ~new_n510;
  assign new_n512 = ~\400  & ~new_n511;
  assign new_n513 = ~new_n508 & ~new_n512;
  assign new_n514 = ~\280  & \335 ;
  assign new_n515 = ~\273  & ~\335 ;
  assign new_n516 = ~new_n514 & ~new_n515;
  assign new_n517 = ~\411  & ~new_n516;
  assign new_n518 = new_n513 & ~new_n517;
  assign new_n519 = ~\241  & \335 ;
  assign new_n520 = ~\234  & ~\335 ;
  assign new_n521 = ~new_n519 & ~new_n520;
  assign new_n522 = ~\435  & ~new_n521;
  assign new_n523 = \435  & new_n521;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = ~\288  & \335 ;
  assign new_n526 = ~\281  & ~\335 ;
  assign new_n527 = ~new_n525 & ~new_n526;
  assign new_n528 = \374  & new_n527;
  assign new_n529 = ~\374  & ~new_n527;
  assign new_n530 = ~new_n528 & ~new_n529;
  assign new_n531 = new_n524 & new_n530;
  assign new_n532 = \389  & new_n507;
  assign new_n533 = \400  & new_n511;
  assign new_n534 = \411  & new_n516;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536 = new_n513 & ~new_n535;
  assign new_n537 = ~new_n532 & ~new_n536;
  assign new_n538 = new_n518 & new_n531;
  assign new_n539 = new_n537 & new_n538;
  assign new_n540 = \422  & new_n500;
  assign new_n541 = ~new_n497 & ~new_n540;
  assign new_n542 = new_n504 & ~new_n541;
  assign new_n543 = \457  & new_n491;
  assign new_n544 = ~new_n503 & ~new_n543;
  assign new_n545 = ~new_n504 & ~new_n544;
  assign new_n546 = new_n540 & new_n545;
  assign new_n547 = ~new_n497 & ~new_n543;
  assign new_n548 = ~new_n542 & ~new_n547;
  assign new_n549 = ~new_n546 & ~new_n548;
  assign new_n550 = ~new_n542 & new_n549;
  assign new_n551 = ~\209  & \335 ;
  assign new_n552 = ~\206  & ~\335 ;
  assign new_n553 = ~new_n551 & ~new_n552;
  assign new_n554 = ~\446  & ~new_n553;
  assign new_n555 = \446  & new_n553;
  assign new_n556 = ~new_n554 & ~new_n555;
  assign new_n557 = new_n504 & new_n556;
  assign new_n558 = new_n539 & new_n557;
  assign \6641  = new_n550 & new_n558;
  assign new_n560 = \332  & ~\366 ;
  assign new_n561 = ~\332  & ~\361 ;
  assign new_n562 = ~new_n560 & ~new_n561;
  assign new_n563 = ~\315  & \332 ;
  assign new_n564 = ~\308  & ~\332 ;
  assign new_n565 = ~new_n563 & ~new_n564;
  assign new_n566 = \479  & new_n565;
  assign new_n567 = ~\307  & \332 ;
  assign new_n568 = ~\302  & ~\332 ;
  assign new_n569 = ~new_n567 & ~new_n568;
  assign new_n570 = new_n566 & new_n569;
  assign new_n571 = ~\479  & ~new_n565;
  assign new_n572 = ~new_n566 & ~new_n571;
  assign new_n573 = ~\323  & \332 ;
  assign new_n574 = ~\316  & ~\332 ;
  assign new_n575 = ~new_n573 & ~new_n574;
  assign new_n576 = ~\490  & ~new_n575;
  assign new_n577 = new_n569 & ~new_n576;
  assign new_n578 = new_n572 & ~new_n577;
  assign new_n579 = ~new_n570 & ~new_n578;
  assign new_n580 = ~\299  & \332 ;
  assign new_n581 = ~\293  & ~\332 ;
  assign new_n582 = ~new_n580 & ~new_n581;
  assign new_n583 = new_n579 & ~new_n582;
  assign new_n584 = ~new_n579 & new_n582;
  assign new_n585 = ~new_n583 & ~new_n584;
  assign new_n586 = ~\331  & \332 ;
  assign new_n587 = ~\324  & ~\332 ;
  assign new_n588 = ~new_n586 & ~new_n587;
  assign new_n589 = ~\503  & ~new_n588;
  assign new_n590 = \503  & new_n588;
  assign new_n591 = ~new_n589 & ~new_n590;
  assign new_n592 = \332  & ~\338 ;
  assign new_n593 = \514  & ~new_n592;
  assign new_n594 = ~\514  & new_n592;
  assign new_n595 = ~new_n593 & ~new_n594;
  assign new_n596 = new_n591 & new_n595;
  assign new_n597 = \332  & \348 ;
  assign new_n598 = ~\332  & \341 ;
  assign new_n599 = ~new_n597 & ~new_n598;
  assign new_n600 = ~\523  & new_n599;
  assign new_n601 = \523  & ~new_n599;
  assign new_n602 = ~new_n600 & ~new_n601;
  assign new_n603 = \332  & ~\358 ;
  assign new_n604 = ~\332  & ~\351 ;
  assign new_n605 = ~new_n603 & ~new_n604;
  assign new_n606 = \534  & new_n605;
  assign new_n607 = ~\534  & ~new_n605;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = new_n602 & new_n608;
  assign new_n610 = new_n596 & new_n609;
  assign new_n611 = \490  & new_n575;
  assign new_n612 = ~new_n576 & ~new_n611;
  assign new_n613 = new_n572 & ~new_n582;
  assign new_n614 = new_n612 & new_n613;
  assign new_n615 = new_n610 & new_n614;
  assign new_n616 = new_n585 & new_n615;
  assign \6643  = ~new_n562 & new_n616;
  assign new_n618 = \308  & ~\324 ;
  assign new_n619 = ~\308  & \324 ;
  assign new_n620 = ~new_n618 & ~new_n619;
  assign new_n621 = ~\302  & ~\316 ;
  assign new_n622 = \302  & \316 ;
  assign new_n623 = ~new_n621 & ~new_n622;
  assign new_n624 = ~\293  & ~\361 ;
  assign new_n625 = \293  & \361 ;
  assign new_n626 = ~new_n624 & ~new_n625;
  assign new_n627 = \341  & new_n626;
  assign new_n628 = ~\341  & ~new_n626;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = \351  & ~\369 ;
  assign new_n631 = ~\351  & \369 ;
  assign new_n632 = ~new_n630 & ~new_n631;
  assign new_n633 = new_n629 & new_n632;
  assign new_n634 = ~new_n629 & ~new_n632;
  assign new_n635 = ~new_n633 & ~new_n634;
  assign new_n636 = new_n623 & ~new_n635;
  assign new_n637 = ~new_n623 & new_n635;
  assign new_n638 = ~new_n636 & ~new_n637;
  assign new_n639 = new_n620 & new_n638;
  assign new_n640 = ~new_n620 & ~new_n638;
  assign \6716  = ~new_n639 & ~new_n640;
  assign new_n642 = ~\281  & ~\289 ;
  assign new_n643 = \281  & \289 ;
  assign new_n644 = ~new_n642 & ~new_n643;
  assign new_n645 = ~\206  & ~\210 ;
  assign new_n646 = \206  & \210 ;
  assign new_n647 = ~new_n645 & ~new_n646;
  assign new_n648 = new_n644 & ~new_n647;
  assign new_n649 = ~new_n644 & new_n647;
  assign new_n650 = ~new_n648 & ~new_n649;
  assign new_n651 = ~\218  & ~\226 ;
  assign new_n652 = \218  & \226 ;
  assign new_n653 = ~new_n651 & ~new_n652;
  assign new_n654 = \265  & ~\273 ;
  assign new_n655 = ~\265  & \273 ;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = new_n653 & new_n656;
  assign new_n658 = ~new_n653 & ~new_n656;
  assign new_n659 = ~new_n657 & ~new_n658;
  assign new_n660 = \234  & ~\257 ;
  assign new_n661 = ~\234  & \257 ;
  assign new_n662 = ~new_n660 & ~new_n661;
  assign new_n663 = new_n659 & ~new_n662;
  assign new_n664 = ~new_n659 & new_n662;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = new_n650 & new_n665;
  assign new_n667 = ~new_n650 & ~new_n665;
  assign \6877  = ~new_n666 & ~new_n667;
  assign new_n669 = ~new_n492 & ~new_n550;
  assign new_n670 = new_n518 & new_n528;
  assign new_n671 = new_n537 & ~new_n670;
  assign new_n672 = new_n524 & ~new_n671;
  assign new_n673 = ~new_n523 & ~new_n672;
  assign new_n674 = new_n504 & ~new_n673;
  assign new_n675 = ~new_n555 & ~new_n674;
  assign new_n676 = ~new_n669 & new_n675;
  assign \6924  = ~new_n554 & ~new_n676;
  assign new_n678 = ~new_n569 & ~new_n582;
  assign new_n679 = ~new_n566 & new_n678;
  assign new_n680 = ~new_n601 & ~new_n606;
  assign new_n681 = new_n562 & ~new_n607;
  assign new_n682 = new_n680 & ~new_n681;
  assign new_n683 = ~new_n600 & ~new_n682;
  assign new_n684 = ~new_n593 & ~new_n683;
  assign new_n685 = ~new_n589 & ~new_n594;
  assign new_n686 = ~new_n684 & new_n685;
  assign new_n687 = ~new_n590 & ~new_n686;
  assign new_n688 = ~new_n611 & new_n687;
  assign new_n689 = new_n572 & ~new_n576;
  assign new_n690 = ~new_n688 & new_n689;
  assign \6925  = ~new_n679 | new_n690;
  assign new_n692 = ~\619  & ~\625 ;
  assign new_n693 = ~new_n389 & new_n692;
  assign new_n694 = \619  & ~\625 ;
  assign new_n695 = ~\54  & ~new_n562;
  assign new_n696 = \54  & new_n562;
  assign new_n697 = ~new_n695 & ~new_n696;
  assign new_n698 = new_n694 & ~new_n697;
  assign new_n699 = ~\619  & \625 ;
  assign new_n700 = \131  & new_n699;
  assign new_n701 = ~new_n693 & ~new_n700;
  assign \7015  = ~new_n698 & new_n701;
  assign new_n703 = ~new_n361 & new_n692;
  assign new_n704 = \129  & new_n699;
  assign new_n705 = new_n608 & ~new_n695;
  assign new_n706 = ~new_n608 & new_n695;
  assign new_n707 = new_n694 & ~new_n705;
  assign new_n708 = ~new_n706 & new_n707;
  assign new_n709 = ~new_n703 & ~new_n704;
  assign \7363  = ~new_n708 & new_n709;
  assign new_n711 = ~new_n408 & new_n692;
  assign new_n712 = \4  & ~new_n530;
  assign new_n713 = ~\4  & new_n530;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = new_n694 & ~new_n714;
  assign new_n716 = \117  & new_n699;
  assign new_n717 = ~new_n711 & ~new_n716;
  assign \7365  = ~new_n715 & new_n717;
  assign new_n719 = ~new_n606 & ~new_n705;
  assign new_n720 = new_n602 & ~new_n719;
  assign new_n721 = ~new_n683 & ~new_n720;
  assign new_n722 = new_n595 & ~new_n721;
  assign new_n723 = ~new_n593 & ~new_n722;
  assign new_n724 = new_n591 & ~new_n723;
  assign new_n725 = new_n687 & ~new_n724;
  assign new_n726 = new_n612 & ~new_n725;
  assign new_n727 = ~new_n611 & ~new_n726;
  assign new_n728 = new_n572 & ~new_n727;
  assign new_n729 = ~new_n566 & ~new_n728;
  assign new_n730 = ~new_n569 & new_n729;
  assign new_n731 = new_n582 & ~new_n730;
  assign new_n732 = new_n679 & ~new_n728;
  assign \7432  = ~new_n731 & ~new_n732;
  assign new_n734 = ~\607  & ~\610 ;
  assign new_n735 = \7015  & new_n734;
  assign new_n736 = \607  & ~\610 ;
  assign new_n737 = ~\11  & new_n736;
  assign new_n738 = \607  & \610 ;
  assign new_n739 = ~\61  & new_n738;
  assign new_n740 = ~\607  & \610 ;
  assign new_n741 = \7365  & new_n740;
  assign new_n742 = ~new_n737 & ~new_n739;
  assign new_n743 = ~new_n735 & new_n742;
  assign \7449  = ~new_n741 & new_n743;
  assign new_n745 = ~new_n343 & new_n692;
  assign new_n746 = \52  & new_n699;
  assign new_n747 = ~new_n591 & new_n723;
  assign new_n748 = new_n694 & ~new_n724;
  assign new_n749 = ~new_n747 & new_n748;
  assign new_n750 = ~new_n745 & ~new_n746;
  assign \7465  = ~new_n749 & new_n750;
  assign new_n752 = new_n393 & new_n692;
  assign new_n753 = \130  & new_n699;
  assign new_n754 = ~new_n595 & new_n721;
  assign new_n755 = new_n694 & ~new_n722;
  assign new_n756 = ~new_n754 & new_n755;
  assign new_n757 = ~new_n752 & ~new_n753;
  assign \7466  = ~new_n756 & new_n757;
  assign new_n759 = ~new_n352 & new_n692;
  assign new_n760 = \119  & new_n699;
  assign new_n761 = ~new_n602 & new_n719;
  assign new_n762 = new_n694 & ~new_n720;
  assign new_n763 = ~new_n761 & new_n762;
  assign new_n764 = ~new_n759 & ~new_n760;
  assign \7467  = ~new_n763 & new_n764;
  assign new_n766 = ~\613  & ~\616 ;
  assign new_n767 = ~\7015  & new_n766;
  assign new_n768 = ~\613  & \616 ;
  assign new_n769 = \11  & new_n768;
  assign new_n770 = \613  & \616 ;
  assign new_n771 = \61  & new_n770;
  assign new_n772 = \613  & ~\616 ;
  assign new_n773 = ~\7365  & new_n772;
  assign new_n774 = ~new_n769 & ~new_n771;
  assign new_n775 = ~new_n767 & new_n774;
  assign \7469  = new_n773 | ~new_n775;
  assign new_n777 = ~new_n453 & new_n692;
  assign new_n778 = ~new_n529 & ~new_n713;
  assign new_n779 = ~new_n517 & ~new_n534;
  assign new_n780 = ~new_n778 & new_n779;
  assign new_n781 = ~new_n517 & ~new_n780;
  assign new_n782 = ~new_n512 & ~new_n533;
  assign new_n783 = new_n781 & new_n782;
  assign new_n784 = ~new_n533 & ~new_n783;
  assign new_n785 = ~new_n508 & ~new_n532;
  assign new_n786 = new_n784 & new_n785;
  assign new_n787 = ~new_n508 & ~new_n786;
  assign new_n788 = ~new_n524 & new_n787;
  assign new_n789 = new_n524 & ~new_n787;
  assign new_n790 = ~new_n788 & ~new_n789;
  assign new_n791 = new_n694 & ~new_n790;
  assign new_n792 = \122  & new_n699;
  assign new_n793 = ~new_n777 & ~new_n792;
  assign \7470  = ~new_n791 & new_n793;
  assign new_n795 = ~new_n480 & new_n692;
  assign new_n796 = ~new_n784 & ~new_n785;
  assign new_n797 = ~new_n786 & ~new_n796;
  assign new_n798 = new_n694 & ~new_n797;
  assign new_n799 = \128  & new_n699;
  assign new_n800 = ~new_n795 & ~new_n799;
  assign \7471  = ~new_n798 & new_n800;
  assign new_n802 = ~new_n417 & new_n692;
  assign new_n803 = ~new_n781 & ~new_n782;
  assign new_n804 = ~new_n783 & ~new_n803;
  assign new_n805 = new_n694 & new_n804;
  assign new_n806 = \127  & new_n699;
  assign new_n807 = ~new_n802 & ~new_n806;
  assign \7472  = ~new_n805 & new_n807;
  assign new_n809 = ~new_n471 & new_n692;
  assign new_n810 = new_n778 & ~new_n779;
  assign new_n811 = ~new_n780 & ~new_n810;
  assign new_n812 = new_n694 & ~new_n811;
  assign new_n813 = \126  & new_n699;
  assign new_n814 = ~new_n809 & ~new_n813;
  assign \7473  = ~new_n812 & new_n814;
  assign new_n816 = new_n588 & ~new_n605;
  assign new_n817 = ~new_n588 & new_n605;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = new_n565 & new_n818;
  assign new_n820 = ~new_n565 & ~new_n818;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = \348  & new_n821;
  assign new_n823 = ~\348  & ~new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = \338  & ~new_n824;
  assign new_n826 = ~\338  & new_n824;
  assign new_n827 = ~new_n825 & ~new_n826;
  assign new_n828 = \332  & ~new_n827;
  assign new_n829 = \341  & new_n821;
  assign new_n830 = ~\341  & ~new_n821;
  assign new_n831 = ~new_n829 & ~new_n830;
  assign new_n832 = ~\332  & ~new_n831;
  assign new_n833 = ~new_n828 & ~new_n832;
  assign new_n834 = new_n569 & new_n582;
  assign new_n835 = ~new_n678 & ~new_n834;
  assign new_n836 = \332  & ~\372 ;
  assign new_n837 = ~\332  & ~\369 ;
  assign new_n838 = ~new_n836 & ~new_n837;
  assign new_n839 = new_n562 & ~new_n575;
  assign new_n840 = ~new_n562 & new_n575;
  assign new_n841 = ~new_n839 & ~new_n840;
  assign new_n842 = new_n838 & new_n841;
  assign new_n843 = ~new_n838 & ~new_n841;
  assign new_n844 = ~new_n842 & ~new_n843;
  assign new_n845 = new_n835 & ~new_n844;
  assign new_n846 = ~new_n835 & new_n844;
  assign new_n847 = ~new_n845 & ~new_n846;
  assign new_n848 = new_n833 & new_n847;
  assign new_n849 = ~new_n833 & ~new_n847;
  assign \7474  = ~new_n848 & ~new_n849;
  assign new_n851 = new_n491 & ~new_n495;
  assign new_n852 = ~new_n491 & new_n495;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = new_n507 & new_n853;
  assign new_n855 = ~new_n507 & ~new_n853;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = ~\292  & \335 ;
  assign new_n858 = ~\289  & ~\335 ;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = new_n500 & ~new_n553;
  assign new_n861 = ~new_n500 & new_n553;
  assign new_n862 = ~new_n860 & ~new_n861;
  assign new_n863 = new_n859 & new_n862;
  assign new_n864 = ~new_n859 & ~new_n862;
  assign new_n865 = ~new_n863 & ~new_n864;
  assign new_n866 = new_n521 & ~new_n865;
  assign new_n867 = ~new_n521 & new_n865;
  assign new_n868 = ~new_n866 & ~new_n867;
  assign new_n869 = ~new_n516 & new_n527;
  assign new_n870 = new_n516 & ~new_n527;
  assign new_n871 = ~new_n869 & ~new_n870;
  assign new_n872 = new_n868 & new_n871;
  assign new_n873 = ~new_n868 & ~new_n871;
  assign new_n874 = ~new_n872 & ~new_n873;
  assign new_n875 = new_n511 & ~new_n874;
  assign new_n876 = ~new_n511 & new_n874;
  assign new_n877 = ~new_n875 & ~new_n876;
  assign new_n878 = new_n856 & new_n877;
  assign new_n879 = ~new_n856 & ~new_n877;
  assign \7476  = new_n878 | new_n879;
  assign new_n881 = ~new_n492 & ~new_n543;
  assign new_n882 = ~new_n496 & ~new_n497;
  assign new_n883 = ~new_n523 & ~new_n787;
  assign new_n884 = ~new_n522 & ~new_n883;
  assign new_n885 = ~new_n501 & ~new_n540;
  assign new_n886 = ~new_n884 & new_n885;
  assign new_n887 = ~new_n501 & ~new_n886;
  assign new_n888 = new_n882 & ~new_n887;
  assign new_n889 = ~new_n496 & ~new_n888;
  assign new_n890 = new_n881 & ~new_n889;
  assign new_n891 = ~new_n881 & new_n889;
  assign new_n892 = ~new_n890 & ~new_n891;
  assign new_n893 = new_n504 & new_n884;
  assign new_n894 = ~new_n669 & ~new_n893;
  assign new_n895 = new_n556 & ~new_n894;
  assign new_n896 = ~new_n556 & new_n894;
  assign new_n897 = ~new_n895 & ~new_n896;
  assign new_n898 = ~new_n882 & new_n887;
  assign new_n899 = ~new_n888 & ~new_n898;
  assign new_n900 = new_n883 & new_n885;
  assign new_n901 = ~new_n522 & ~new_n885;
  assign new_n902 = new_n714 & ~new_n901;
  assign new_n903 = new_n811 & new_n902;
  assign new_n904 = ~new_n804 & new_n903;
  assign new_n905 = new_n797 & new_n904;
  assign new_n906 = ~new_n788 & new_n905;
  assign new_n907 = ~new_n900 & new_n906;
  assign new_n908 = ~new_n897 & new_n907;
  assign new_n909 = new_n899 & new_n908;
  assign \7503  = new_n892 & new_n909;
  assign \7504  = new_n616 & new_n697;
  assign new_n912 = ~\571  & ~\574 ;
  assign new_n913 = ~\7015  & new_n912;
  assign new_n914 = ~\571  & \574 ;
  assign new_n915 = \182  & new_n914;
  assign new_n916 = \571  & \574 ;
  assign new_n917 = \185  & new_n916;
  assign new_n918 = \571  & ~\574 ;
  assign new_n919 = ~\7365  & new_n918;
  assign new_n920 = ~new_n915 & ~new_n917;
  assign new_n921 = ~new_n913 & new_n920;
  assign new_n922 = ~new_n919 & new_n921;
  assign \7506  = \137  & ~new_n922;
  assign new_n924 = ~\577  & ~\580 ;
  assign new_n925 = ~\7015  & new_n924;
  assign new_n926 = ~\577  & \580 ;
  assign new_n927 = \182  & new_n926;
  assign new_n928 = \577  & \580 ;
  assign new_n929 = \185  & new_n928;
  assign new_n930 = \577  & ~\580 ;
  assign new_n931 = ~\7365  & new_n930;
  assign new_n932 = ~new_n927 & ~new_n929;
  assign new_n933 = ~new_n925 & new_n932;
  assign new_n934 = ~new_n931 & new_n933;
  assign \7511  = \137  & ~new_n934;
  assign new_n936 = new_n734 & ~\7465 ;
  assign new_n937 = \37  & new_n738;
  assign new_n938 = \43  & new_n736;
  assign new_n939 = new_n740 & ~\7470 ;
  assign new_n940 = ~new_n937 & ~new_n938;
  assign new_n941 = ~new_n936 & new_n940;
  assign \7515  = new_n939 | ~new_n941;
  assign new_n943 = new_n734 & ~\7466 ;
  assign new_n944 = \20  & new_n738;
  assign new_n945 = \76  & new_n736;
  assign new_n946 = new_n740 & ~\7471 ;
  assign new_n947 = ~new_n944 & ~new_n945;
  assign new_n948 = ~new_n943 & new_n947;
  assign \7516  = new_n946 | ~new_n948;
  assign new_n950 = new_n734 & ~\7467 ;
  assign new_n951 = \17  & new_n738;
  assign new_n952 = \73  & new_n736;
  assign new_n953 = new_n740 & ~\7472 ;
  assign new_n954 = ~new_n951 & ~new_n952;
  assign new_n955 = ~new_n950 & new_n954;
  assign \7517  = new_n953 | ~new_n955;
  assign new_n957 = ~\7363  & new_n734;
  assign new_n958 = \67  & new_n736;
  assign new_n959 = \70  & new_n738;
  assign new_n960 = new_n740 & ~\7473 ;
  assign new_n961 = ~new_n958 & ~new_n959;
  assign new_n962 = ~new_n957 & new_n961;
  assign \7518  = new_n960 | ~new_n962;
  assign new_n964 = ~\7465  & new_n766;
  assign new_n965 = \37  & new_n770;
  assign new_n966 = \43  & new_n768;
  assign new_n967 = new_n772 & ~\7470 ;
  assign new_n968 = ~new_n965 & ~new_n966;
  assign new_n969 = ~new_n964 & new_n968;
  assign \7519  = new_n967 | ~new_n969;
  assign new_n971 = ~\7466  & new_n766;
  assign new_n972 = \20  & new_n770;
  assign new_n973 = \76  & new_n768;
  assign new_n974 = new_n772 & ~\7471 ;
  assign new_n975 = ~new_n972 & ~new_n973;
  assign new_n976 = ~new_n971 & new_n975;
  assign \7520  = new_n974 | ~new_n976;
  assign new_n978 = ~\7467  & new_n766;
  assign new_n979 = \17  & new_n770;
  assign new_n980 = \73  & new_n768;
  assign new_n981 = new_n772 & ~\7472 ;
  assign new_n982 = ~new_n979 & ~new_n980;
  assign new_n983 = ~new_n978 & new_n982;
  assign \7521  = new_n981 | ~new_n983;
  assign new_n985 = ~\7363  & new_n766;
  assign new_n986 = \67  & new_n768;
  assign new_n987 = \70  & new_n770;
  assign new_n988 = new_n772 & ~\7473 ;
  assign new_n989 = ~new_n986 & ~new_n987;
  assign new_n990 = ~new_n985 & new_n989;
  assign \7522  = new_n988 | ~new_n990;
  assign new_n992 = ~\7465  & new_n912;
  assign new_n993 = \170  & new_n916;
  assign new_n994 = \200  & new_n914;
  assign new_n995 = ~\7470  & new_n918;
  assign new_n996 = ~new_n993 & ~new_n994;
  assign new_n997 = ~new_n992 & new_n996;
  assign new_n998 = ~new_n995 & new_n997;
  assign \7600  = \137  & ~new_n998;
  assign new_n1000 = ~\7363  & new_n912;
  assign new_n1001 = \158  & new_n916;
  assign new_n1002 = \188  & new_n914;
  assign new_n1003 = ~\7473  & new_n918;
  assign new_n1004 = ~new_n1001 & ~new_n1002;
  assign new_n1005 = ~new_n1000 & new_n1004;
  assign new_n1006 = ~new_n1003 & new_n1005;
  assign \7601  = \137  & ~new_n1006;
  assign new_n1008 = ~\7467  & new_n912;
  assign new_n1009 = \152  & new_n916;
  assign new_n1010 = \155  & new_n914;
  assign new_n1011 = ~\7472  & new_n918;
  assign new_n1012 = ~new_n1009 & ~new_n1010;
  assign new_n1013 = ~new_n1008 & new_n1012;
  assign new_n1014 = ~new_n1011 & new_n1013;
  assign \7602  = \137  & ~new_n1014;
  assign new_n1016 = ~\7466  & new_n912;
  assign new_n1017 = \146  & new_n916;
  assign new_n1018 = \149  & new_n914;
  assign new_n1019 = ~\7471  & new_n918;
  assign new_n1020 = ~new_n1017 & ~new_n1018;
  assign new_n1021 = ~new_n1016 & new_n1020;
  assign new_n1022 = ~new_n1019 & new_n1021;
  assign \7603  = \137  & ~new_n1022;
  assign new_n1024 = ~\7465  & new_n924;
  assign new_n1025 = \170  & new_n928;
  assign new_n1026 = \200  & new_n926;
  assign new_n1027 = ~\7470  & new_n930;
  assign new_n1028 = ~new_n1025 & ~new_n1026;
  assign new_n1029 = ~new_n1024 & new_n1028;
  assign new_n1030 = ~new_n1027 & new_n1029;
  assign \7604  = \137  & ~new_n1030;
  assign new_n1032 = ~\7363  & new_n924;
  assign new_n1033 = \158  & new_n928;
  assign new_n1034 = \188  & new_n926;
  assign new_n1035 = ~\7473  & new_n930;
  assign new_n1036 = ~new_n1033 & ~new_n1034;
  assign new_n1037 = ~new_n1032 & new_n1036;
  assign new_n1038 = ~new_n1035 & new_n1037;
  assign \7605  = \137  & ~new_n1038;
  assign new_n1040 = ~\7467  & new_n924;
  assign new_n1041 = \152  & new_n928;
  assign new_n1042 = \155  & new_n926;
  assign new_n1043 = ~\7472  & new_n930;
  assign new_n1044 = ~new_n1041 & ~new_n1042;
  assign new_n1045 = ~new_n1040 & new_n1044;
  assign new_n1046 = ~new_n1043 & new_n1045;
  assign \7606  = \137  & ~new_n1046;
  assign new_n1048 = ~\7466  & new_n924;
  assign new_n1049 = \146  & new_n928;
  assign new_n1050 = \149  & new_n926;
  assign new_n1051 = ~\7471  & new_n930;
  assign new_n1052 = ~new_n1049 & ~new_n1050;
  assign new_n1053 = ~new_n1048 & new_n1052;
  assign new_n1054 = ~new_n1051 & new_n1053;
  assign \7607  = \137  & ~new_n1054;
  assign new_n1056 = \135  & \631 ;
  assign new_n1057 = ~\603  & new_n386;
  assign new_n1058 = ~\132  & ~new_n582;
  assign new_n1059 = \132  & new_n582;
  assign new_n1060 = ~new_n1058 & ~new_n1059;
  assign new_n1061 = \603  & ~new_n1060;
  assign new_n1062 = ~\599  & ~new_n1057;
  assign new_n1063 = ~new_n1061 & new_n1062;
  assign new_n1064 = \123  & ~\603 ;
  assign new_n1065 = \603  & ~\7432 ;
  assign new_n1066 = \599  & ~new_n1064;
  assign new_n1067 = ~new_n1065 & new_n1066;
  assign new_n1068 = ~new_n1056 & ~new_n1063;
  assign \7626  = ~new_n1067 & new_n1068;
  assign new_n1070 = ~\132  & ~new_n730;
  assign new_n1071 = \132  & new_n730;
  assign \7698  = new_n1070 | new_n1071;
  assign new_n1073 = new_n386 & new_n692;
  assign new_n1074 = \123  & new_n699;
  assign new_n1075 = new_n694 & ~\7432 ;
  assign new_n1076 = ~new_n1073 & ~new_n1074;
  assign \7699  = ~new_n1075 & new_n1076;
  assign new_n1078 = ~new_n383 & new_n692;
  assign new_n1079 = new_n569 & ~new_n729;
  assign new_n1080 = ~new_n730 & ~new_n1079;
  assign new_n1081 = new_n694 & ~new_n1080;
  assign new_n1082 = \121  & new_n699;
  assign new_n1083 = ~new_n1078 & ~new_n1082;
  assign \7700  = ~new_n1081 & new_n1083;
  assign new_n1085 = new_n379 & new_n692;
  assign new_n1086 = \116  & new_n699;
  assign new_n1087 = ~new_n572 & new_n727;
  assign new_n1088 = new_n694 & ~new_n728;
  assign new_n1089 = ~new_n1087 & new_n1088;
  assign new_n1090 = ~new_n1085 & ~new_n1086;
  assign \7701  = ~new_n1089 & new_n1090;
  assign new_n1092 = new_n370 & new_n692;
  assign new_n1093 = \112  & new_n699;
  assign new_n1094 = ~new_n612 & new_n725;
  assign new_n1095 = new_n694 & ~new_n726;
  assign new_n1096 = ~new_n1094 & new_n1095;
  assign new_n1097 = ~new_n1092 & ~new_n1093;
  assign \7702  = ~new_n1096 & new_n1097;
  assign new_n1099 = \245  & \559 ;
  assign new_n1100 = \1140  & new_n1099;
  assign new_n1101 = ~\2061  & new_n1100;
  assign new_n1102 = ~\6877  & new_n1101;
  assign new_n1103 = ~\6716  & new_n1102;
  assign new_n1104 = ~\7474  & new_n1103;
  assign \7703  = ~\7476  & new_n1104;
  assign new_n1106 = new_n462 & new_n692;
  assign new_n1107 = new_n694 & new_n897;
  assign new_n1108 = \115  & new_n699;
  assign new_n1109 = ~new_n1106 & ~new_n1108;
  assign \7704  = ~new_n1107 & new_n1109;
  assign new_n1111 = ~new_n435 & new_n692;
  assign new_n1112 = new_n694 & ~new_n892;
  assign new_n1113 = \114  & new_n699;
  assign new_n1114 = ~new_n1111 & ~new_n1113;
  assign \7705  = ~new_n1112 & new_n1114;
  assign new_n1116 = ~new_n444 & new_n692;
  assign new_n1117 = new_n694 & ~new_n899;
  assign new_n1118 = \53  & new_n699;
  assign new_n1119 = ~new_n1116 & ~new_n1118;
  assign \7706  = ~new_n1117 & new_n1119;
  assign new_n1121 = ~new_n426 & new_n692;
  assign new_n1122 = new_n884 & ~new_n885;
  assign new_n1123 = ~new_n886 & ~new_n1122;
  assign new_n1124 = new_n694 & ~new_n1123;
  assign new_n1125 = \113  & new_n699;
  assign new_n1126 = ~new_n1121 & ~new_n1125;
  assign \7707  = ~new_n1124 & new_n1126;
  assign new_n1128 = new_n766 & ~\7699 ;
  assign new_n1129 = \106  & new_n770;
  assign new_n1130 = \109  & new_n768;
  assign new_n1131 = new_n772 & ~\7704 ;
  assign new_n1132 = ~new_n1129 & ~new_n1130;
  assign new_n1133 = ~new_n1131 & new_n1132;
  assign \7735  = new_n1128 | ~new_n1133;
  assign new_n1135 = new_n734 & ~\7699 ;
  assign new_n1136 = \106  & new_n738;
  assign new_n1137 = \109  & new_n736;
  assign new_n1138 = new_n740 & ~\7704 ;
  assign new_n1139 = ~new_n1136 & ~new_n1137;
  assign new_n1140 = ~new_n1138 & new_n1139;
  assign \7736  = new_n1135 | ~new_n1140;
  assign new_n1142 = new_n734 & ~\7700 ;
  assign new_n1143 = \46  & new_n736;
  assign new_n1144 = \49  & new_n738;
  assign new_n1145 = new_n740 & ~\7705 ;
  assign new_n1146 = ~new_n1143 & ~new_n1144;
  assign new_n1147 = ~new_n1142 & new_n1146;
  assign \7737  = new_n1145 | ~new_n1147;
  assign new_n1149 = new_n734 & \7701 ;
  assign new_n1150 = ~\100  & new_n736;
  assign new_n1151 = ~\103  & new_n738;
  assign new_n1152 = new_n740 & \7706 ;
  assign new_n1153 = ~new_n1150 & ~new_n1151;
  assign new_n1154 = ~new_n1149 & new_n1153;
  assign \7738  = ~new_n1152 & new_n1154;
  assign new_n1156 = new_n734 & ~\7702 ;
  assign new_n1157 = \40  & new_n738;
  assign new_n1158 = \91  & new_n736;
  assign new_n1159 = new_n740 & ~\7707 ;
  assign new_n1160 = ~new_n1157 & ~new_n1158;
  assign new_n1161 = ~new_n1156 & new_n1160;
  assign \7739  = new_n1159 | ~new_n1161;
  assign new_n1163 = new_n766 & \7700 ;
  assign new_n1164 = ~\46  & new_n768;
  assign new_n1165 = ~\49  & new_n770;
  assign new_n1166 = new_n772 & \7705 ;
  assign new_n1167 = ~new_n1164 & ~new_n1165;
  assign new_n1168 = ~new_n1163 & new_n1167;
  assign \7740  = ~new_n1166 & new_n1168;
  assign new_n1170 = new_n766 & ~\7701 ;
  assign new_n1171 = \100  & new_n768;
  assign new_n1172 = \103  & new_n770;
  assign new_n1173 = new_n772 & ~\7706 ;
  assign new_n1174 = ~new_n1171 & ~new_n1172;
  assign new_n1175 = ~new_n1170 & new_n1174;
  assign \7741  = new_n1173 | ~new_n1175;
  assign new_n1177 = new_n766 & ~\7702 ;
  assign new_n1178 = \40  & new_n770;
  assign new_n1179 = \91  & new_n768;
  assign new_n1180 = new_n772 & ~\7707 ;
  assign new_n1181 = ~new_n1178 & ~new_n1179;
  assign new_n1182 = ~new_n1177 & new_n1181;
  assign \7742  = new_n1180 | ~new_n1182;
  assign new_n1184 = new_n912 & ~\7702 ;
  assign new_n1185 = \173  & new_n916;
  assign new_n1186 = \203  & new_n914;
  assign new_n1187 = new_n918 & ~\7707 ;
  assign new_n1188 = ~new_n1185 & ~new_n1186;
  assign new_n1189 = ~new_n1184 & new_n1188;
  assign new_n1190 = ~new_n1187 & new_n1189;
  assign \7754  = \137  & ~new_n1190;
  assign new_n1192 = new_n912 & ~\7701 ;
  assign new_n1193 = \167  & new_n916;
  assign new_n1194 = \197  & new_n914;
  assign new_n1195 = new_n918 & ~\7706 ;
  assign new_n1196 = ~new_n1193 & ~new_n1194;
  assign new_n1197 = ~new_n1192 & new_n1196;
  assign new_n1198 = ~new_n1195 & new_n1197;
  assign \7755  = \137  & ~new_n1198;
  assign new_n1200 = new_n912 & ~\7700 ;
  assign new_n1201 = \164  & new_n916;
  assign new_n1202 = \194  & new_n914;
  assign new_n1203 = new_n918 & ~\7705 ;
  assign new_n1204 = ~new_n1201 & ~new_n1202;
  assign new_n1205 = ~new_n1200 & new_n1204;
  assign new_n1206 = ~new_n1203 & new_n1205;
  assign \7756  = \137  & ~new_n1206;
  assign new_n1208 = new_n918 & ~\7704 ;
  assign new_n1209 = \161  & new_n916;
  assign new_n1210 = \191  & new_n914;
  assign new_n1211 = new_n912 & ~\7699 ;
  assign new_n1212 = ~new_n1209 & ~new_n1210;
  assign new_n1213 = ~new_n1208 & new_n1212;
  assign new_n1214 = ~new_n1211 & new_n1213;
  assign \7757  = \137  & ~new_n1214;
  assign new_n1216 = new_n924 & ~\7702 ;
  assign new_n1217 = \173  & new_n928;
  assign new_n1218 = \203  & new_n926;
  assign new_n1219 = new_n930 & ~\7707 ;
  assign new_n1220 = ~new_n1217 & ~new_n1218;
  assign new_n1221 = ~new_n1216 & new_n1220;
  assign new_n1222 = ~new_n1219 & new_n1221;
  assign \7758  = \137  & ~new_n1222;
  assign new_n1224 = new_n924 & ~\7701 ;
  assign new_n1225 = \167  & new_n928;
  assign new_n1226 = \197  & new_n926;
  assign new_n1227 = new_n930 & ~\7706 ;
  assign new_n1228 = ~new_n1225 & ~new_n1226;
  assign new_n1229 = ~new_n1224 & new_n1228;
  assign new_n1230 = ~new_n1227 & new_n1229;
  assign \7759  = \137  & ~new_n1230;
  assign new_n1232 = new_n924 & ~\7700 ;
  assign new_n1233 = \164  & new_n928;
  assign new_n1234 = \194  & new_n926;
  assign new_n1235 = new_n930 & ~\7705 ;
  assign new_n1236 = ~new_n1233 & ~new_n1234;
  assign new_n1237 = ~new_n1232 & new_n1236;
  assign new_n1238 = ~new_n1235 & new_n1237;
  assign \7760  = \137  & ~new_n1238;
  assign new_n1240 = new_n924 & ~\7699 ;
  assign new_n1241 = \161  & new_n928;
  assign new_n1242 = \191  & new_n926;
  assign new_n1243 = new_n930 & ~\7704 ;
  assign new_n1244 = ~new_n1241 & ~new_n1242;
  assign new_n1245 = ~new_n1243 & new_n1244;
  assign new_n1246 = ~new_n1240 & new_n1245;
  assign \7761  = \137  & ~new_n1246;
  assign new_n1248 = new_n576 & ~new_n585;
  assign new_n1249 = new_n585 & new_n611;
  assign new_n1250 = ~new_n614 & ~new_n1248;
  assign new_n1251 = ~new_n1249 & new_n1250;
  assign new_n1252 = new_n572 & new_n1251;
  assign new_n1253 = new_n585 & new_n612;
  assign new_n1254 = ~new_n1252 & new_n1253;
  assign new_n1255 = \583  & new_n610;
  assign new_n1256 = new_n687 & ~new_n1255;
  assign new_n1257 = ~new_n1251 & new_n1256;
  assign new_n1258 = ~new_n585 & new_n612;
  assign new_n1259 = ~new_n1256 & ~new_n1258;
  assign new_n1260 = new_n1251 & new_n1259;
  assign new_n1261 = ~new_n1257 & ~new_n1260;
  assign new_n1262 = ~new_n1254 & new_n1261;
  assign new_n1263 = ~new_n591 & ~new_n595;
  assign new_n1264 = ~new_n596 & ~new_n1263;
  assign new_n1265 = ~new_n609 & new_n684;
  assign new_n1266 = ~new_n594 & ~new_n1265;
  assign new_n1267 = new_n601 & new_n606;
  assign new_n1268 = ~new_n680 & ~new_n1267;
  assign new_n1269 = ~new_n600 & new_n607;
  assign new_n1270 = ~new_n1268 & ~new_n1269;
  assign new_n1271 = new_n562 & ~new_n1270;
  assign new_n1272 = ~new_n562 & new_n1270;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = new_n1266 & ~new_n1273;
  assign new_n1275 = ~new_n1266 & new_n1273;
  assign new_n1276 = ~new_n1274 & ~new_n1275;
  assign new_n1277 = \583  & ~new_n1276;
  assign new_n1278 = ~new_n594 & new_n683;
  assign new_n1279 = ~new_n684 & ~new_n1278;
  assign new_n1280 = ~new_n562 & ~new_n607;
  assign new_n1281 = ~new_n606 & ~new_n1280;
  assign new_n1282 = new_n602 & ~new_n1281;
  assign new_n1283 = ~new_n602 & new_n1281;
  assign new_n1284 = ~new_n1282 & ~new_n1283;
  assign new_n1285 = new_n1279 & ~new_n1284;
  assign new_n1286 = ~new_n1279 & new_n1284;
  assign new_n1287 = ~new_n1285 & ~new_n1286;
  assign new_n1288 = ~\583  & ~new_n1287;
  assign new_n1289 = ~new_n1277 & ~new_n1288;
  assign new_n1290 = new_n1264 & ~new_n1289;
  assign new_n1291 = ~new_n1264 & new_n1289;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = ~new_n1262 & ~new_n1292;
  assign new_n1294 = new_n1262 & new_n1292;
  assign new_n1295 = new_n694 & ~new_n1293;
  assign new_n1296 = ~new_n1294 & new_n1295;
  assign new_n1297 = new_n370 & new_n379;
  assign new_n1298 = ~new_n380 & ~new_n1297;
  assign new_n1299 = ~\248  & \514 ;
  assign new_n1300 = \242  & ~\514 ;
  assign new_n1301 = ~new_n1299 & ~new_n1300;
  assign new_n1302 = ~\254  & ~\534 ;
  assign new_n1303 = \251  & \534 ;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = new_n1301 & ~new_n1304;
  assign new_n1306 = ~new_n1301 & new_n1304;
  assign new_n1307 = ~\351  & ~new_n1305;
  assign new_n1308 = ~new_n1306 & new_n1307;
  assign new_n1309 = ~\242  & ~\248 ;
  assign new_n1310 = \242  & \248 ;
  assign new_n1311 = ~new_n1309 & ~new_n1310;
  assign new_n1312 = ~\514  & ~\534 ;
  assign new_n1313 = \514  & \534 ;
  assign new_n1314 = \351  & ~new_n1312;
  assign new_n1315 = ~new_n1313 & new_n1314;
  assign new_n1316 = ~new_n1311 & new_n1315;
  assign new_n1317 = ~new_n1308 & ~new_n1316;
  assign new_n1318 = new_n1298 & ~new_n1317;
  assign new_n1319 = ~new_n1298 & new_n1317;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = ~\248  & \523 ;
  assign new_n1322 = \242  & ~\523 ;
  assign new_n1323 = \341  & ~new_n1321;
  assign new_n1324 = ~new_n1322 & new_n1323;
  assign new_n1325 = ~\251  & \523 ;
  assign new_n1326 = \254  & ~\523 ;
  assign new_n1327 = ~\341  & ~new_n1325;
  assign new_n1328 = ~new_n1326 & new_n1327;
  assign new_n1329 = ~new_n1324 & ~new_n1328;
  assign new_n1330 = new_n383 & ~new_n1329;
  assign new_n1331 = ~new_n383 & new_n1329;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = new_n386 & ~new_n389;
  assign new_n1334 = ~new_n390 & ~new_n1333;
  assign new_n1335 = ~\248  & \503 ;
  assign new_n1336 = \242  & ~\503 ;
  assign new_n1337 = \324  & ~new_n1335;
  assign new_n1338 = ~new_n1336 & new_n1337;
  assign new_n1339 = ~\251  & \503 ;
  assign new_n1340 = \254  & ~\503 ;
  assign new_n1341 = ~\324  & ~new_n1339;
  assign new_n1342 = ~new_n1340 & new_n1341;
  assign new_n1343 = ~new_n1338 & ~new_n1342;
  assign new_n1344 = new_n1334 & ~new_n1343;
  assign new_n1345 = ~new_n1334 & new_n1343;
  assign new_n1346 = ~new_n1344 & ~new_n1345;
  assign new_n1347 = new_n1332 & new_n1346;
  assign new_n1348 = ~new_n1332 & ~new_n1346;
  assign new_n1349 = ~new_n1347 & ~new_n1348;
  assign new_n1350 = ~new_n1320 & ~new_n1349;
  assign new_n1351 = new_n1320 & new_n1349;
  assign new_n1352 = new_n692 & ~new_n1350;
  assign new_n1353 = ~new_n1351 & new_n1352;
  assign new_n1354 = ~new_n1296 & ~new_n1353;
  assign new_n1355 = ~\120  & new_n699;
  assign \8075  = new_n1354 & ~new_n1355;
  assign new_n1357 = ~\248  & \389 ;
  assign new_n1358 = \242  & ~\389 ;
  assign new_n1359 = \257  & ~new_n1357;
  assign new_n1360 = ~new_n1358 & new_n1359;
  assign new_n1361 = ~\251  & \389 ;
  assign new_n1362 = \254  & ~\389 ;
  assign new_n1363 = ~\257  & ~new_n1361;
  assign new_n1364 = ~new_n1362 & new_n1363;
  assign new_n1365 = ~new_n1360 & ~new_n1364;
  assign new_n1366 = ~\248  & \435 ;
  assign new_n1367 = \242  & ~\435 ;
  assign new_n1368 = \234  & ~new_n1366;
  assign new_n1369 = ~new_n1367 & new_n1368;
  assign new_n1370 = ~\251  & \435 ;
  assign new_n1371 = \254  & ~\435 ;
  assign new_n1372 = ~\234  & ~new_n1370;
  assign new_n1373 = ~new_n1371 & new_n1372;
  assign new_n1374 = ~new_n1369 & ~new_n1373;
  assign new_n1375 = new_n1365 & ~new_n1374;
  assign new_n1376 = ~new_n1365 & new_n1374;
  assign new_n1377 = ~new_n1375 & ~new_n1376;
  assign new_n1378 = ~\248  & \411 ;
  assign new_n1379 = \242  & ~\411 ;
  assign new_n1380 = \273  & ~new_n1378;
  assign new_n1381 = ~new_n1379 & new_n1380;
  assign new_n1382 = ~\251  & \411 ;
  assign new_n1383 = \254  & ~\411 ;
  assign new_n1384 = ~\273  & ~new_n1382;
  assign new_n1385 = ~new_n1383 & new_n1384;
  assign new_n1386 = ~new_n1381 & ~new_n1385;
  assign new_n1387 = ~\248  & \374 ;
  assign new_n1388 = \242  & ~\374 ;
  assign new_n1389 = \281  & ~new_n1387;
  assign new_n1390 = ~new_n1388 & new_n1389;
  assign new_n1391 = ~\251  & \374 ;
  assign new_n1392 = \254  & ~\374 ;
  assign new_n1393 = ~\281  & ~new_n1391;
  assign new_n1394 = ~new_n1392 & new_n1393;
  assign new_n1395 = ~new_n1390 & ~new_n1394;
  assign new_n1396 = new_n1386 & ~new_n1395;
  assign new_n1397 = ~new_n1386 & new_n1395;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = new_n1377 & new_n1398;
  assign new_n1400 = ~new_n1377 & ~new_n1398;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = ~\248  & \457 ;
  assign new_n1403 = \242  & ~\457 ;
  assign new_n1404 = \210  & ~new_n1402;
  assign new_n1405 = ~new_n1403 & new_n1404;
  assign new_n1406 = ~\251  & \457 ;
  assign new_n1407 = \254  & ~\457 ;
  assign new_n1408 = ~\210  & ~new_n1406;
  assign new_n1409 = ~new_n1407 & new_n1408;
  assign new_n1410 = ~new_n1405 & ~new_n1409;
  assign new_n1411 = new_n462 & ~new_n1410;
  assign new_n1412 = ~new_n462 & new_n1410;
  assign new_n1413 = ~new_n1411 & ~new_n1412;
  assign new_n1414 = ~\248  & \400 ;
  assign new_n1415 = \242  & ~\400 ;
  assign new_n1416 = \265  & ~new_n1414;
  assign new_n1417 = ~new_n1415 & new_n1416;
  assign new_n1418 = ~\251  & \400 ;
  assign new_n1419 = \254  & ~\400 ;
  assign new_n1420 = ~\265  & ~new_n1418;
  assign new_n1421 = ~new_n1419 & new_n1420;
  assign new_n1422 = ~new_n1417 & ~new_n1421;
  assign new_n1423 = ~\248  & \468 ;
  assign new_n1424 = \242  & ~\468 ;
  assign new_n1425 = \218  & ~new_n1423;
  assign new_n1426 = ~new_n1424 & new_n1425;
  assign new_n1427 = ~\251  & \468 ;
  assign new_n1428 = \254  & ~\468 ;
  assign new_n1429 = ~\218  & ~new_n1427;
  assign new_n1430 = ~new_n1428 & new_n1429;
  assign new_n1431 = ~new_n1426 & ~new_n1430;
  assign new_n1432 = ~new_n1422 & new_n1431;
  assign new_n1433 = new_n1422 & ~new_n1431;
  assign new_n1434 = ~new_n1432 & ~new_n1433;
  assign new_n1435 = ~\248  & \422 ;
  assign new_n1436 = \242  & ~\422 ;
  assign new_n1437 = \226  & ~new_n1435;
  assign new_n1438 = ~new_n1436 & new_n1437;
  assign new_n1439 = ~\251  & \422 ;
  assign new_n1440 = \254  & ~\422 ;
  assign new_n1441 = ~\226  & ~new_n1439;
  assign new_n1442 = ~new_n1440 & new_n1441;
  assign new_n1443 = ~new_n1438 & ~new_n1442;
  assign new_n1444 = new_n1434 & ~new_n1443;
  assign new_n1445 = ~new_n1434 & new_n1443;
  assign new_n1446 = ~new_n1444 & ~new_n1445;
  assign new_n1447 = new_n1413 & new_n1446;
  assign new_n1448 = ~new_n1413 & ~new_n1446;
  assign new_n1449 = ~new_n1447 & ~new_n1448;
  assign new_n1450 = new_n1401 & new_n1449;
  assign new_n1451 = ~new_n1401 & ~new_n1449;
  assign new_n1452 = new_n692 & ~new_n1450;
  assign new_n1453 = ~new_n1451 & new_n1452;
  assign new_n1454 = ~\457  & ~\468 ;
  assign new_n1455 = \457  & \468 ;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = ~\389  & ~new_n556;
  assign new_n1458 = \389  & new_n556;
  assign new_n1459 = ~new_n1457 & ~new_n1458;
  assign new_n1460 = new_n1456 & ~new_n1459;
  assign new_n1461 = ~new_n1456 & new_n1459;
  assign new_n1462 = ~new_n1460 & ~new_n1461;
  assign new_n1463 = new_n856 & new_n1462;
  assign new_n1464 = ~new_n856 & ~new_n1462;
  assign new_n1465 = ~new_n1463 & ~new_n1464;
  assign new_n1466 = \566  & new_n539;
  assign new_n1467 = new_n673 & ~new_n1466;
  assign new_n1468 = ~new_n501 & new_n549;
  assign new_n1469 = new_n501 & new_n548;
  assign new_n1470 = new_n1467 & ~new_n1469;
  assign new_n1471 = ~new_n1468 & new_n1470;
  assign new_n1472 = ~new_n540 & ~new_n545;
  assign new_n1473 = ~new_n546 & ~new_n1472;
  assign new_n1474 = ~new_n1467 & new_n1473;
  assign new_n1475 = ~new_n1471 & ~new_n1474;
  assign new_n1476 = new_n518 & ~new_n529;
  assign new_n1477 = new_n537 & ~new_n1476;
  assign new_n1478 = ~new_n524 & ~new_n530;
  assign new_n1479 = ~new_n531 & ~new_n1478;
  assign new_n1480 = new_n779 & ~new_n1479;
  assign new_n1481 = ~new_n779 & new_n1479;
  assign new_n1482 = ~new_n1480 & ~new_n1481;
  assign new_n1483 = new_n1477 & new_n1482;
  assign new_n1484 = ~new_n1477 & ~new_n1482;
  assign new_n1485 = ~new_n1483 & ~new_n1484;
  assign new_n1486 = ~new_n512 & new_n517;
  assign new_n1487 = ~new_n533 & new_n534;
  assign new_n1488 = new_n512 & ~new_n517;
  assign new_n1489 = ~new_n1486 & ~new_n1487;
  assign new_n1490 = ~new_n1488 & new_n1489;
  assign new_n1491 = new_n529 & new_n1490;
  assign new_n1492 = ~new_n529 & ~new_n1490;
  assign new_n1493 = ~new_n1491 & ~new_n1492;
  assign new_n1494 = ~new_n779 & ~new_n1493;
  assign new_n1495 = ~new_n517 & new_n535;
  assign new_n1496 = ~new_n1491 & new_n1495;
  assign new_n1497 = ~new_n1494 & ~new_n1496;
  assign new_n1498 = ~new_n1485 & new_n1497;
  assign new_n1499 = new_n1485 & ~new_n1497;
  assign new_n1500 = ~new_n1498 & ~new_n1499;
  assign new_n1501 = \566  & ~new_n1500;
  assign new_n1502 = ~new_n524 & new_n671;
  assign new_n1503 = ~new_n672 & ~new_n1502;
  assign new_n1504 = new_n528 & new_n779;
  assign new_n1505 = ~new_n1493 & ~new_n1504;
  assign new_n1506 = new_n533 & new_n1504;
  assign new_n1507 = ~new_n1505 & ~new_n1506;
  assign new_n1508 = new_n1503 & new_n1507;
  assign new_n1509 = ~new_n1503 & ~new_n1507;
  assign new_n1510 = ~new_n1508 & ~new_n1509;
  assign new_n1511 = ~\566  & ~new_n1510;
  assign new_n1512 = ~new_n1501 & ~new_n1511;
  assign new_n1513 = new_n1475 & ~new_n1512;
  assign new_n1514 = ~new_n1475 & new_n1512;
  assign new_n1515 = ~new_n1513 & ~new_n1514;
  assign new_n1516 = ~new_n1465 & ~new_n1515;
  assign new_n1517 = new_n1465 & new_n1515;
  assign new_n1518 = new_n694 & ~new_n1516;
  assign new_n1519 = ~new_n1517 & new_n1518;
  assign new_n1520 = ~new_n1453 & ~new_n1519;
  assign new_n1521 = ~\118  & new_n699;
  assign \8076  = new_n1520 & ~new_n1521;
  assign new_n1523 = \94  & \625 ;
  assign new_n1524 = new_n1354 & ~new_n1523;
  assign new_n1525 = new_n734 & ~new_n1524;
  assign new_n1526 = \14  & new_n736;
  assign new_n1527 = \64  & new_n738;
  assign new_n1528 = \97  & \625 ;
  assign new_n1529 = new_n1520 & ~new_n1528;
  assign new_n1530 = new_n740 & ~new_n1529;
  assign new_n1531 = ~new_n1526 & ~new_n1527;
  assign new_n1532 = ~new_n1525 & new_n1531;
  assign \8123  = new_n1530 | ~new_n1532;
  assign new_n1534 = new_n766 & ~new_n1524;
  assign new_n1535 = \14  & new_n768;
  assign new_n1536 = \64  & new_n770;
  assign new_n1537 = new_n772 & ~new_n1529;
  assign new_n1538 = ~new_n1535 & ~new_n1536;
  assign new_n1539 = ~new_n1534 & new_n1538;
  assign \8124  = new_n1537 | ~new_n1539;
  assign new_n1541 = new_n912 & ~new_n1524;
  assign new_n1542 = new_n918 & ~new_n1529;
  assign new_n1543 = ~\176  & ~\571 ;
  assign new_n1544 = ~\179  & \571 ;
  assign new_n1545 = \574  & ~new_n1543;
  assign new_n1546 = ~new_n1544 & new_n1545;
  assign new_n1547 = ~new_n1541 & ~new_n1546;
  assign new_n1548 = ~new_n1542 & new_n1547;
  assign \8127  = ~\137  | new_n1548;
  assign new_n1550 = new_n924 & ~new_n1524;
  assign new_n1551 = \176  & new_n926;
  assign new_n1552 = \179  & new_n928;
  assign new_n1553 = new_n930 & ~new_n1529;
  assign new_n1554 = ~new_n1551 & ~new_n1552;
  assign new_n1555 = ~new_n1550 & new_n1554;
  assign new_n1556 = ~new_n1553 & new_n1555;
  assign \8128  = ~\137  | new_n1556;
  assign \1137  = ~\545 ;
  assign \1138  = ~\348 ;
  assign \1139  = ~\366 ;
  assign \1141  = ~\549 ;
  assign \1144  = ~\338 ;
  assign \1145  = ~\358 ;
  assign \1152  = ~\245 ;
  assign \1153  = ~\552 ;
  assign \1154  = ~\562 ;
  assign \1155  = ~\559 ;
  assign \3613  = ~\299 ;
  assign \709  = \141 ;
  assign \816  = \293 ;
  assign \1066  = \592 ;
  assign \1142  = \1137 ;
  assign \1143  = \1137 ;
  assign \2139  = \137 ;
  assign \2142  = \141 ;
  assign \2309  = \1 ;
  assign \2387  = \549 ;
  assign \2527  = \299 ;
  assign \2584  = \1141 ;
  assign \3357  = \1 ;
  assign \3358  = \1 ;
  assign \3359  = \1 ;
  assign \3360  = \1 ;
  assign \3604  = \299 ;
  assign \4278  = \4275 ;
  assign \6646  = \6643 ;
  assign \6648  = \6641 ;
  assign \6926  = \6924 ;
  assign \6927  = \6925 ;
endmodule


