// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    p_50_15_, p_133_66_, p_169_92_, p_182_105_, p_12_3_, p_94_49_,
    p_205_128_, p_212_135_, p_1197_165_, p_2211_176_, p_4432_203_,
    p_4526_205_, p_26_7_, p_53_16_, p_54_17_, p_192_115_, p_1496_173_,
    p_2208_175_, p_113_58_, p_153_76_, p_222_145_, p_4393_195_, p_103_52_,
    p_195_118_, p_3749_194_, p_4405_198_, p_4528_206_, p_114_59_,
    p_166_89_, p_176_99_, p_179_102_, p_197_120_, p_232_155_, p_3737_192_,
    p_4394_196_, p_23_6_, p_55_18_, p_56_19_, p_60_23_, p_61_24_,
    p_115_60_, p_159_82_, p_185_108_, p_163_86_, p_189_112_, p_1492_172_,
    p_2204_174_, p_3698_185_, p_186_109_, p_193_116_, p_207_130_, p_18_5_,
    p_69_30_, p_150_73_, p_152_75_, p_156_79_, p_177_100_, p_199_122_,
    p_201_124_, p_216_139_, p_223_146_, p_230_153_, p_2236_180_, p_62_25_,
    p_63_26_, p_66_29_, p_73_32_, p_74_33_, p_130_65_, p_147_72_,
    p_183_106_, p_196_119_, p_217_140_, p_187_110_, p_204_127_, p_213_136_,
    p_226_149_, p_240_163_, p_3717_189_, p_3729_191_, p_35_10_, p_70_31_,
    p_227_150_, p_3711_188_, p_15_4_, p_110_55_, p_162_85_, p_172_95_,
    p_210_133_, p_236_159_, p_1469_169_, p_2224_178_, p_2239_181_, p_1_0_,
    p_38_11_, p_64_27_, p_65_28_, p_237_160_, p_127_64_, p_175_98_,
    p_220_143_, p_233_156_, p_1455_166_, p_3701_186_, p_9_2_, p_135_68_,
    p_144_71_, p_167_90_, p_218_141_, p_1480_170_, p_3723_190_, p_188_111_,
    p_234_157_, p_82_41_, p_83_42_, p_86_45_, p_87_46_, p_157_80_,
    p_208_131_, p_3705_187_, p_41_12_, p_47_14_, p_58_21_, p_124_63_,
    p_161_84_, p_165_88_, p_178_101_, p_200_123_, p_231_154_, p_97_50_,
    p_118_61_, p_180_103_, p_238_161_, p_1459_167_, p_59_22_, p_160_83_,
    p_174_97_, p_203_126_, p_214_137_, p_221_144_, p_1462_168_,
    p_2230_179_, p_75_34_, p_76_35_, p_81_40_, p_88_47_, p_89_48_,
    p_100_51_, p_190_113_, p_228_151_, p_4420_201_, p_44_13_, p_111_56_,
    p_121_62_, p_155_78_, p_171_94_, p_206_129_, p_211_134_, p_224_147_,
    p_2247_182_, p_109_54_, p_134_67_, p_168_91_, p_229_152_, p_154_77_,
    p_2218_177_, p_77_36_, p_78_37_, p_141_70_, p_239_162_, p_173_96_,
    p_235_158_, p_2256_184_, p_4437_204_, p_184_107_, p_191_114_,
    p_209_132_, p_5_1_, p_32_9_, p_57_20_, p_112_57_, p_164_87_, p_170_93_,
    p_225_148_, p_3743_193_, p_4410_199_, p_29_8_, p_79_38_, p_84_43_,
    p_85_44_, p_106_53_, p_138_69_, p_158_81_, p_181_104_, p_194_117_,
    p_219_142_, p_4400_197_, p_4427_202_, p_80_39_, p_151_74_, p_198_121_,
    p_202_125_, p_215_138_, p_339_164_, p_1486_171_, p_2253_183_,
    p_4415_200_,
    p_279_304_, p_382_3148_, p_432_428_, p_450_288_, p_440_277_,
    p_444_282_, p_488_260_, p_494_267_, p_524_210_, p_246_3110_,
    p_373_2994_, p_376_3206_, p_530_216_, p_560_248_, p_316_3397_,
    p_534_220_, p_278_536_, p_370_3718_, p_544_230_, p_252_3450_,
    p_273_3402_, p_327_3408_, p_338_3716_, p_406_388_, p_422_3451_,
    p_484_256_, p_550_236_, p_321_3715_, p_368_3431_, p_448_284_,
    p_453_596_, p_540_227_, p_554_240_, p_3_312_, p_264_3121_, p_307_3389_,
    p_353_3425_, p_391_3094_, p_480_250_, p_301_3388_, p_388_3093_,
    p_438_274_, p_490_263_, p_528_214_, p_333_3416_, p_410_387_,
    p_469_3452_, p_486_258_, p_359_3426_, p_385_3151_, p_397_3097_,
    p_471_3445_, p_538_224_, p_281_547_, p_292_392_, p_310_3393_,
    p_324_3363_, p_412_3369_, p_548_234_, p_289_383_, p_379_3207_,
    p_418_3449_, p_404_390_, p_558_244_, p_2_313_, p_542_246_, p_313_3396_,
    p_319_3398_, p_546_232_, p_552_238_, p_270_3109_, p_556_242_,
    p_276_3401_, p_446_393_, p_496_271_, p_522_226_, p_304_3390_,
    p_336_3412_, p_341_420_, p_365_3430_, p_492_265_, p_526_212_,
    p_330_3411_, p_344_3382_, p_347_3420_, p_399_3717_, p_436_286_,
    p_532_218_, p_286_419_, p_408_385_, p_536_222_, p_362_3429_,
    p_394_3095_, p_416_3368_, p_414_3338_, p_478_269_, p_284_384_,
    p_402_395_, p_419_3444_, p_350_3421_, p_249_3418_, p_258_3122_,
    p_298_3387_, p_442_280_, p_482_253_, p_295_3352_, p_356_3424_  );
  input  p_50_15_, p_133_66_, p_169_92_, p_182_105_, p_12_3_, p_94_49_,
    p_205_128_, p_212_135_, p_1197_165_, p_2211_176_, p_4432_203_,
    p_4526_205_, p_26_7_, p_53_16_, p_54_17_, p_192_115_, p_1496_173_,
    p_2208_175_, p_113_58_, p_153_76_, p_222_145_, p_4393_195_, p_103_52_,
    p_195_118_, p_3749_194_, p_4405_198_, p_4528_206_, p_114_59_,
    p_166_89_, p_176_99_, p_179_102_, p_197_120_, p_232_155_, p_3737_192_,
    p_4394_196_, p_23_6_, p_55_18_, p_56_19_, p_60_23_, p_61_24_,
    p_115_60_, p_159_82_, p_185_108_, p_163_86_, p_189_112_, p_1492_172_,
    p_2204_174_, p_3698_185_, p_186_109_, p_193_116_, p_207_130_, p_18_5_,
    p_69_30_, p_150_73_, p_152_75_, p_156_79_, p_177_100_, p_199_122_,
    p_201_124_, p_216_139_, p_223_146_, p_230_153_, p_2236_180_, p_62_25_,
    p_63_26_, p_66_29_, p_73_32_, p_74_33_, p_130_65_, p_147_72_,
    p_183_106_, p_196_119_, p_217_140_, p_187_110_, p_204_127_, p_213_136_,
    p_226_149_, p_240_163_, p_3717_189_, p_3729_191_, p_35_10_, p_70_31_,
    p_227_150_, p_3711_188_, p_15_4_, p_110_55_, p_162_85_, p_172_95_,
    p_210_133_, p_236_159_, p_1469_169_, p_2224_178_, p_2239_181_, p_1_0_,
    p_38_11_, p_64_27_, p_65_28_, p_237_160_, p_127_64_, p_175_98_,
    p_220_143_, p_233_156_, p_1455_166_, p_3701_186_, p_9_2_, p_135_68_,
    p_144_71_, p_167_90_, p_218_141_, p_1480_170_, p_3723_190_, p_188_111_,
    p_234_157_, p_82_41_, p_83_42_, p_86_45_, p_87_46_, p_157_80_,
    p_208_131_, p_3705_187_, p_41_12_, p_47_14_, p_58_21_, p_124_63_,
    p_161_84_, p_165_88_, p_178_101_, p_200_123_, p_231_154_, p_97_50_,
    p_118_61_, p_180_103_, p_238_161_, p_1459_167_, p_59_22_, p_160_83_,
    p_174_97_, p_203_126_, p_214_137_, p_221_144_, p_1462_168_,
    p_2230_179_, p_75_34_, p_76_35_, p_81_40_, p_88_47_, p_89_48_,
    p_100_51_, p_190_113_, p_228_151_, p_4420_201_, p_44_13_, p_111_56_,
    p_121_62_, p_155_78_, p_171_94_, p_206_129_, p_211_134_, p_224_147_,
    p_2247_182_, p_109_54_, p_134_67_, p_168_91_, p_229_152_, p_154_77_,
    p_2218_177_, p_77_36_, p_78_37_, p_141_70_, p_239_162_, p_173_96_,
    p_235_158_, p_2256_184_, p_4437_204_, p_184_107_, p_191_114_,
    p_209_132_, p_5_1_, p_32_9_, p_57_20_, p_112_57_, p_164_87_, p_170_93_,
    p_225_148_, p_3743_193_, p_4410_199_, p_29_8_, p_79_38_, p_84_43_,
    p_85_44_, p_106_53_, p_138_69_, p_158_81_, p_181_104_, p_194_117_,
    p_219_142_, p_4400_197_, p_4427_202_, p_80_39_, p_151_74_, p_198_121_,
    p_202_125_, p_215_138_, p_339_164_, p_1486_171_, p_2253_183_,
    p_4415_200_;
  output p_279_304_, p_382_3148_, p_432_428_, p_450_288_, p_440_277_,
    p_444_282_, p_488_260_, p_494_267_, p_524_210_, p_246_3110_,
    p_373_2994_, p_376_3206_, p_530_216_, p_560_248_, p_316_3397_,
    p_534_220_, p_278_536_, p_370_3718_, p_544_230_, p_252_3450_,
    p_273_3402_, p_327_3408_, p_338_3716_, p_406_388_, p_422_3451_,
    p_484_256_, p_550_236_, p_321_3715_, p_368_3431_, p_448_284_,
    p_453_596_, p_540_227_, p_554_240_, p_3_312_, p_264_3121_, p_307_3389_,
    p_353_3425_, p_391_3094_, p_480_250_, p_301_3388_, p_388_3093_,
    p_438_274_, p_490_263_, p_528_214_, p_333_3416_, p_410_387_,
    p_469_3452_, p_486_258_, p_359_3426_, p_385_3151_, p_397_3097_,
    p_471_3445_, p_538_224_, p_281_547_, p_292_392_, p_310_3393_,
    p_324_3363_, p_412_3369_, p_548_234_, p_289_383_, p_379_3207_,
    p_418_3449_, p_404_390_, p_558_244_, p_2_313_, p_542_246_, p_313_3396_,
    p_319_3398_, p_546_232_, p_552_238_, p_270_3109_, p_556_242_,
    p_276_3401_, p_446_393_, p_496_271_, p_522_226_, p_304_3390_,
    p_336_3412_, p_341_420_, p_365_3430_, p_492_265_, p_526_212_,
    p_330_3411_, p_344_3382_, p_347_3420_, p_399_3717_, p_436_286_,
    p_532_218_, p_286_419_, p_408_385_, p_536_222_, p_362_3429_,
    p_394_3095_, p_416_3368_, p_414_3338_, p_478_269_, p_284_384_,
    p_402_395_, p_419_3444_, p_350_3421_, p_249_3418_, p_258_3122_,
    p_298_3387_, p_442_280_, p_482_253_, p_295_3352_, p_356_3424_;
  wire new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378, new_n379, new_n380, new_n381, new_n382, new_n383, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1357, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1378,
    new_n1379, new_n1380, new_n1381, new_n1382, new_n1383, new_n1384,
    new_n1385, new_n1386, new_n1387, new_n1388, new_n1389, new_n1390,
    new_n1391, new_n1392, new_n1393, new_n1394, new_n1395, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1409, new_n1410, new_n1411, new_n1412, new_n1413, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1418, new_n1419, new_n1420,
    new_n1421, new_n1422, new_n1423, new_n1424, new_n1425, new_n1426,
    new_n1427, new_n1428, new_n1429, new_n1430, new_n1431, new_n1432,
    new_n1433, new_n1434, new_n1435, new_n1436, new_n1437, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1452, new_n1453, new_n1454, new_n1455, new_n1456,
    new_n1457, new_n1458, new_n1459, new_n1460, new_n1461, new_n1462,
    new_n1463, new_n1464, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1469, new_n1470, new_n1471, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1761, new_n1762, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1775, new_n1776, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1783, new_n1784, new_n1786, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1799, new_n1800, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1957, new_n1958, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2251, new_n2252, new_n2254, new_n2255,
    new_n2256, new_n2257, new_n2258, new_n2259, new_n2260, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278, new_n2279, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2295, new_n2296,
    new_n2297, new_n2298, new_n2300, new_n2301, new_n2302, new_n2303,
    new_n2304, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2314, new_n2315, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2454, new_n2455, new_n2456, new_n2457, new_n2458,
    new_n2459, new_n2460, new_n2462, new_n2463, new_n2464, new_n2465,
    new_n2466, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2507, new_n2508, new_n2510, new_n2511;
  assign new_n315 = ~p_18_5_ & p_127_64_;
  assign new_n316 = p_18_5_ & p_233_156_;
  assign new_n317 = ~new_n315 & ~new_n316;
  assign new_n318 = ~p_3737_192_ & new_n317;
  assign new_n319 = p_3737_192_ & ~new_n317;
  assign new_n320 = ~new_n318 & ~new_n319;
  assign new_n321 = ~p_18_5_ & p_130_65_;
  assign new_n322 = p_18_5_ & p_234_157_;
  assign new_n323 = ~new_n321 & ~new_n322;
  assign new_n324 = p_3729_191_ & new_n323;
  assign new_n325 = new_n320 & new_n324;
  assign new_n326 = ~new_n320 & ~new_n324;
  assign new_n327 = ~new_n325 & ~new_n326;
  assign new_n328 = p_103_52_ & ~p_18_5_;
  assign new_n329 = p_18_5_ & p_235_158_;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = ~p_3723_190_ & new_n330;
  assign new_n332 = p_3723_190_ & ~new_n330;
  assign new_n333 = ~new_n331 & ~new_n332;
  assign new_n334 = ~p_18_5_ & p_29_8_;
  assign new_n335 = p_18_5_ & p_238_161_;
  assign new_n336 = ~new_n334 & ~new_n335;
  assign new_n337 = ~p_3705_187_ & new_n336;
  assign new_n338 = p_3705_187_ & ~new_n336;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = ~p_18_5_ & p_41_12_;
  assign new_n341 = p_18_5_ & p_229_152_;
  assign new_n342 = ~new_n340 & ~new_n341;
  assign new_n343 = ~p_18_5_ & ~new_n342;
  assign new_n344 = ~p_18_5_ & ~p_3701_186_;
  assign new_n345 = ~p_18_5_ & ~new_n344;
  assign new_n346 = ~new_n343 & ~new_n345;
  assign new_n347 = new_n343 & new_n345;
  assign new_n348 = ~new_n346 & ~new_n347;
  assign new_n349 = p_26_7_ & ~p_18_5_;
  assign new_n350 = p_18_5_ & p_237_160_;
  assign new_n351 = ~new_n349 & ~new_n350;
  assign new_n352 = ~p_3711_188_ & new_n351;
  assign new_n353 = p_3711_188_ & ~new_n351;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = p_23_6_ & ~p_18_5_;
  assign new_n356 = p_18_5_ & p_236_159_;
  assign new_n357 = ~new_n355 & ~new_n356;
  assign new_n358 = ~p_3717_189_ & new_n357;
  assign new_n359 = p_3717_189_ & ~new_n357;
  assign new_n360 = ~new_n358 & ~new_n359;
  assign new_n361 = ~new_n333 & ~new_n339;
  assign new_n362 = ~new_n348 & new_n361;
  assign new_n363 = ~new_n354 & new_n362;
  assign new_n364 = ~new_n360 & new_n363;
  assign new_n365 = p_4526_205_ & new_n364;
  assign new_n366 = ~p_3705_187_ & ~new_n336;
  assign new_n367 = ~new_n333 & ~new_n360;
  assign new_n368 = new_n366 & new_n367;
  assign new_n369 = ~new_n354 & new_n368;
  assign new_n370 = new_n343 & ~new_n345;
  assign new_n371 = ~new_n360 & new_n370;
  assign new_n372 = ~new_n354 & new_n371;
  assign new_n373 = ~new_n333 & new_n372;
  assign new_n374 = ~new_n339 & new_n373;
  assign new_n375 = ~p_3717_189_ & ~new_n357;
  assign new_n376 = ~new_n333 & new_n375;
  assign new_n377 = ~p_3711_188_ & ~new_n351;
  assign new_n378 = ~new_n333 & new_n377;
  assign new_n379 = ~new_n360 & new_n378;
  assign new_n380 = ~p_3723_190_ & ~new_n330;
  assign new_n381 = ~new_n369 & ~new_n374;
  assign new_n382 = ~new_n376 & new_n381;
  assign new_n383 = ~new_n379 & new_n382;
  assign new_n384 = ~new_n380 & new_n383;
  assign new_n385 = ~new_n365 & new_n384;
  assign new_n386 = new_n327 & ~new_n385;
  assign new_n387 = ~p_3729_191_ & ~new_n323;
  assign new_n388 = new_n320 & new_n387;
  assign new_n389 = ~new_n320 & ~new_n387;
  assign new_n390 = ~new_n388 & ~new_n389;
  assign new_n391 = new_n385 & ~new_n390;
  assign p_382_3148_ = new_n386 | new_n391;
  assign new_n393 = p_12_3_ & p_9_2_;
  assign new_n394 = p_18_5_ & p_213_136_;
  assign new_n395 = p_18_5_ & ~new_n394;
  assign new_n396 = ~new_n393 & ~new_n395;
  assign new_n397 = ~p_1486_171_ & ~new_n396;
  assign new_n398 = p_1486_171_ & new_n396;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = p_18_5_ & p_216_139_;
  assign new_n401 = p_18_5_ & ~new_n400;
  assign new_n402 = ~new_n393 & ~new_n401;
  assign new_n403 = ~p_1469_169_ & ~new_n402;
  assign new_n404 = p_1469_169_ & new_n402;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = p_18_5_ & p_209_132_;
  assign new_n407 = p_18_5_ & ~new_n406;
  assign new_n408 = ~new_n393 & ~new_n407;
  assign new_n409 = ~p_1462_168_ & ~new_n408;
  assign new_n410 = p_1462_168_ & new_n408;
  assign new_n411 = ~new_n409 & ~new_n410;
  assign new_n412 = p_18_5_ & p_215_138_;
  assign new_n413 = p_18_5_ & ~new_n412;
  assign new_n414 = ~new_n393 & ~new_n413;
  assign new_n415 = ~p_106_53_ & ~new_n414;
  assign new_n416 = p_106_53_ & new_n414;
  assign new_n417 = ~new_n415 & ~new_n416;
  assign new_n418 = p_18_5_ & p_214_137_;
  assign new_n419 = p_18_5_ & ~new_n418;
  assign new_n420 = ~new_n393 & ~new_n419;
  assign new_n421 = ~p_1480_170_ & ~new_n420;
  assign new_n422 = p_1480_170_ & new_n420;
  assign new_n423 = ~new_n421 & ~new_n422;
  assign new_n424 = ~new_n399 & ~new_n405;
  assign new_n425 = ~new_n411 & new_n424;
  assign new_n426 = ~new_n417 & new_n425;
  assign new_n427 = ~new_n423 & new_n426;
  assign new_n428 = p_1496_173_ & p_4528_206_;
  assign new_n429 = ~p_38_11_ & ~new_n428;
  assign new_n430 = p_38_11_ & new_n428;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = p_4528_206_ & p_1492_172_;
  assign new_n433 = ~p_38_11_ & ~new_n432;
  assign new_n434 = p_38_11_ & new_n432;
  assign new_n435 = ~new_n433 & ~new_n434;
  assign new_n436 = ~new_n431 & ~new_n435;
  assign new_n437 = new_n427 & new_n436;
  assign new_n438 = ~p_18_5_ & p_47_14_;
  assign new_n439 = p_18_5_ & p_223_146_;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = ~p_4415_200_ & new_n440;
  assign new_n442 = p_4415_200_ & ~new_n440;
  assign new_n443 = ~new_n441 & ~new_n442;
  assign new_n444 = ~p_18_5_ & p_97_50_;
  assign new_n445 = p_18_5_ & p_226_149_;
  assign new_n446 = ~new_n444 & ~new_n445;
  assign new_n447 = ~p_4400_197_ & new_n446;
  assign new_n448 = p_4400_197_ & ~new_n446;
  assign new_n449 = ~new_n447 & ~new_n448;
  assign new_n450 = ~p_18_5_ & p_118_61_;
  assign new_n451 = p_18_5_ & p_217_140_;
  assign new_n452 = ~new_n450 & ~new_n451;
  assign new_n453 = ~p_4394_196_ & new_n452;
  assign new_n454 = p_4394_196_ & ~new_n452;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = p_94_49_ & ~p_18_5_;
  assign new_n457 = p_18_5_ & p_225_148_;
  assign new_n458 = ~new_n456 & ~new_n457;
  assign new_n459 = ~p_4405_198_ & new_n458;
  assign new_n460 = p_4405_198_ & ~new_n458;
  assign new_n461 = ~new_n459 & ~new_n460;
  assign new_n462 = ~p_18_5_ & p_121_62_;
  assign new_n463 = p_18_5_ & p_224_147_;
  assign new_n464 = ~new_n462 & ~new_n463;
  assign new_n465 = ~p_4410_199_ & new_n464;
  assign new_n466 = p_4410_199_ & ~new_n464;
  assign new_n467 = ~new_n465 & ~new_n466;
  assign new_n468 = ~new_n443 & ~new_n449;
  assign new_n469 = ~new_n455 & new_n468;
  assign new_n470 = ~new_n461 & new_n469;
  assign new_n471 = ~new_n467 & new_n470;
  assign new_n472 = ~p_18_5_ & p_66_29_;
  assign new_n473 = p_18_5_ & p_219_142_;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign new_n475 = ~p_4437_204_ & new_n474;
  assign new_n476 = p_4437_204_ & ~new_n474;
  assign new_n477 = ~new_n475 & ~new_n476;
  assign new_n478 = ~p_18_5_ & p_35_10_;
  assign new_n479 = p_222_145_ & p_18_5_;
  assign new_n480 = ~new_n478 & ~new_n479;
  assign new_n481 = ~p_4420_201_ & new_n480;
  assign new_n482 = p_4420_201_ & ~new_n480;
  assign new_n483 = ~new_n481 & ~new_n482;
  assign new_n484 = ~p_18_5_ & p_32_9_;
  assign new_n485 = p_18_5_ & p_221_144_;
  assign new_n486 = ~new_n484 & ~new_n485;
  assign new_n487 = ~p_4427_202_ & new_n486;
  assign new_n488 = p_4427_202_ & ~new_n486;
  assign new_n489 = ~new_n487 & ~new_n488;
  assign new_n490 = p_50_15_ & ~p_18_5_;
  assign new_n491 = p_18_5_ & p_220_143_;
  assign new_n492 = ~new_n490 & ~new_n491;
  assign new_n493 = ~p_4432_203_ & new_n492;
  assign new_n494 = p_4432_203_ & ~new_n492;
  assign new_n495 = ~new_n493 & ~new_n494;
  assign new_n496 = ~new_n477 & ~new_n483;
  assign new_n497 = ~new_n489 & new_n496;
  assign new_n498 = ~new_n495 & new_n497;
  assign new_n499 = new_n471 & new_n498;
  assign new_n500 = p_18_5_ & p_157_80_;
  assign new_n501 = p_18_5_ & ~new_n500;
  assign new_n502 = ~new_n393 & ~new_n501;
  assign new_n503 = ~p_2236_180_ & ~new_n502;
  assign new_n504 = p_2236_180_ & new_n502;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = p_18_5_ & p_160_83_;
  assign new_n507 = ~p_18_5_ & p_138_69_;
  assign new_n508 = ~new_n506 & ~new_n507;
  assign new_n509 = ~p_2218_177_ & new_n508;
  assign new_n510 = p_2218_177_ & ~new_n508;
  assign new_n511 = ~new_n509 & ~new_n510;
  assign new_n512 = p_18_5_ & p_151_74_;
  assign new_n513 = ~p_18_5_ & p_147_72_;
  assign new_n514 = ~new_n512 & ~new_n513;
  assign new_n515 = ~p_2211_176_ & new_n514;
  assign new_n516 = p_2211_176_ & ~new_n514;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = p_159_82_ & p_18_5_;
  assign new_n519 = ~p_18_5_ & p_144_71_;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = ~p_2224_178_ & new_n520;
  assign new_n522 = p_2224_178_ & ~new_n520;
  assign new_n523 = ~new_n521 & ~new_n522;
  assign new_n524 = p_18_5_ & p_158_81_;
  assign new_n525 = ~p_18_5_ & p_135_68_;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = ~p_2230_179_ & new_n526;
  assign new_n528 = p_2230_179_ & ~new_n526;
  assign new_n529 = ~new_n527 & ~new_n528;
  assign new_n530 = ~new_n505 & ~new_n511;
  assign new_n531 = ~new_n517 & new_n530;
  assign new_n532 = ~new_n523 & new_n531;
  assign new_n533 = ~new_n529 & new_n532;
  assign new_n534 = p_153_76_ & p_18_5_;
  assign new_n535 = p_18_5_ & ~new_n534;
  assign new_n536 = ~new_n393 & ~new_n535;
  assign new_n537 = ~p_2256_184_ & ~new_n536;
  assign new_n538 = p_2256_184_ & new_n536;
  assign new_n539 = ~new_n537 & ~new_n538;
  assign new_n540 = p_18_5_ & p_156_79_;
  assign new_n541 = p_18_5_ & ~new_n540;
  assign new_n542 = ~new_n393 & ~new_n541;
  assign new_n543 = ~p_2239_181_ & ~new_n542;
  assign new_n544 = p_2239_181_ & new_n542;
  assign new_n545 = ~new_n543 & ~new_n544;
  assign new_n546 = p_18_5_ & p_155_78_;
  assign new_n547 = p_18_5_ & ~new_n546;
  assign new_n548 = ~new_n393 & ~new_n547;
  assign new_n549 = ~p_2247_182_ & ~new_n548;
  assign new_n550 = p_2247_182_ & new_n548;
  assign new_n551 = ~new_n549 & ~new_n550;
  assign new_n552 = p_18_5_ & p_154_77_;
  assign new_n553 = p_18_5_ & ~new_n552;
  assign new_n554 = ~new_n393 & ~new_n553;
  assign new_n555 = ~p_2253_183_ & ~new_n554;
  assign new_n556 = p_2253_183_ & new_n554;
  assign new_n557 = ~new_n555 & ~new_n556;
  assign new_n558 = ~new_n539 & ~new_n545;
  assign new_n559 = ~new_n551 & new_n558;
  assign new_n560 = ~new_n557 & new_n559;
  assign new_n561 = new_n533 & new_n560;
  assign new_n562 = ~p_18_5_ & p_100_51_;
  assign new_n563 = p_18_5_ & p_231_154_;
  assign new_n564 = ~new_n562 & ~new_n563;
  assign new_n565 = ~p_3749_194_ & new_n564;
  assign new_n566 = p_3749_194_ & ~new_n564;
  assign new_n567 = ~new_n565 & ~new_n566;
  assign new_n568 = ~p_3729_191_ & new_n323;
  assign new_n569 = p_3729_191_ & ~new_n323;
  assign new_n570 = ~new_n568 & ~new_n569;
  assign new_n571 = ~p_18_5_ & p_124_63_;
  assign new_n572 = p_232_155_ & p_18_5_;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = ~p_3743_193_ & new_n573;
  assign new_n575 = p_3743_193_ & ~new_n573;
  assign new_n576 = ~new_n574 & ~new_n575;
  assign new_n577 = ~new_n567 & ~new_n570;
  assign new_n578 = ~new_n320 & new_n577;
  assign new_n579 = ~new_n576 & new_n578;
  assign new_n580 = ~new_n384 & new_n579;
  assign new_n581 = ~new_n567 & ~new_n576;
  assign new_n582 = new_n387 & new_n581;
  assign new_n583 = ~new_n320 & new_n582;
  assign new_n584 = ~p_3743_193_ & ~new_n573;
  assign new_n585 = ~new_n567 & new_n584;
  assign new_n586 = ~p_3737_192_ & ~new_n317;
  assign new_n587 = ~new_n567 & new_n586;
  assign new_n588 = ~new_n576 & new_n587;
  assign new_n589 = ~p_3749_194_ & ~new_n564;
  assign new_n590 = ~new_n583 & ~new_n585;
  assign new_n591 = ~new_n588 & new_n590;
  assign new_n592 = ~new_n589 & new_n591;
  assign new_n593 = ~new_n580 & new_n592;
  assign new_n594 = new_n437 & new_n499;
  assign new_n595 = new_n561 & new_n594;
  assign new_n596 = ~new_n593 & new_n595;
  assign new_n597 = new_n364 & new_n579;
  assign new_n598 = new_n437 & new_n561;
  assign new_n599 = new_n597 & new_n598;
  assign new_n600 = new_n499 & new_n599;
  assign new_n601 = p_4526_205_ & new_n600;
  assign new_n602 = ~p_2218_177_ & ~new_n508;
  assign new_n603 = ~new_n505 & ~new_n529;
  assign new_n604 = new_n602 & new_n603;
  assign new_n605 = ~new_n523 & new_n604;
  assign new_n606 = ~p_2211_176_ & ~new_n514;
  assign new_n607 = ~new_n529 & new_n606;
  assign new_n608 = ~new_n523 & new_n607;
  assign new_n609 = ~new_n505 & new_n608;
  assign new_n610 = ~new_n511 & new_n609;
  assign new_n611 = ~p_2230_179_ & ~new_n526;
  assign new_n612 = ~new_n505 & new_n611;
  assign new_n613 = ~p_2224_178_ & ~new_n520;
  assign new_n614 = ~new_n505 & new_n613;
  assign new_n615 = ~new_n529 & new_n614;
  assign new_n616 = ~p_2236_180_ & new_n502;
  assign new_n617 = ~new_n605 & ~new_n610;
  assign new_n618 = ~new_n612 & new_n617;
  assign new_n619 = ~new_n615 & new_n618;
  assign new_n620 = ~new_n616 & new_n619;
  assign new_n621 = new_n560 & ~new_n620;
  assign new_n622 = ~p_2239_181_ & new_n542;
  assign new_n623 = ~new_n539 & ~new_n557;
  assign new_n624 = new_n622 & new_n623;
  assign new_n625 = ~new_n551 & new_n624;
  assign new_n626 = ~p_2253_183_ & new_n554;
  assign new_n627 = ~new_n539 & new_n626;
  assign new_n628 = ~p_2247_182_ & new_n548;
  assign new_n629 = ~new_n539 & new_n628;
  assign new_n630 = ~new_n557 & new_n629;
  assign new_n631 = ~p_2256_184_ & new_n536;
  assign new_n632 = ~new_n625 & ~new_n627;
  assign new_n633 = ~new_n630 & new_n632;
  assign new_n634 = ~new_n631 & new_n633;
  assign new_n635 = ~new_n621 & new_n634;
  assign new_n636 = new_n437 & ~new_n635;
  assign new_n637 = ~p_4400_197_ & ~new_n446;
  assign new_n638 = ~new_n443 & ~new_n467;
  assign new_n639 = new_n637 & new_n638;
  assign new_n640 = ~new_n461 & new_n639;
  assign new_n641 = ~p_4394_196_ & ~new_n452;
  assign new_n642 = ~new_n467 & new_n641;
  assign new_n643 = ~new_n461 & new_n642;
  assign new_n644 = ~new_n443 & new_n643;
  assign new_n645 = ~new_n449 & new_n644;
  assign new_n646 = ~p_4410_199_ & ~new_n464;
  assign new_n647 = ~new_n443 & new_n646;
  assign new_n648 = ~p_4405_198_ & ~new_n458;
  assign new_n649 = ~new_n443 & new_n648;
  assign new_n650 = ~new_n467 & new_n649;
  assign new_n651 = ~p_4415_200_ & ~new_n440;
  assign new_n652 = ~new_n640 & ~new_n645;
  assign new_n653 = ~new_n647 & new_n652;
  assign new_n654 = ~new_n650 & new_n653;
  assign new_n655 = ~new_n651 & new_n654;
  assign new_n656 = new_n498 & ~new_n655;
  assign new_n657 = ~p_4420_201_ & ~new_n480;
  assign new_n658 = ~new_n477 & ~new_n495;
  assign new_n659 = new_n657 & new_n658;
  assign new_n660 = ~new_n489 & new_n659;
  assign new_n661 = ~p_4432_203_ & ~new_n492;
  assign new_n662 = ~new_n477 & new_n661;
  assign new_n663 = ~p_4427_202_ & ~new_n486;
  assign new_n664 = ~new_n477 & new_n663;
  assign new_n665 = ~new_n495 & new_n664;
  assign new_n666 = ~p_4437_204_ & ~new_n474;
  assign new_n667 = ~new_n660 & ~new_n662;
  assign new_n668 = ~new_n665 & new_n667;
  assign new_n669 = ~new_n666 & new_n668;
  assign new_n670 = ~new_n656 & new_n669;
  assign new_n671 = new_n598 & ~new_n670;
  assign new_n672 = ~p_1469_169_ & new_n402;
  assign new_n673 = ~new_n399 & ~new_n423;
  assign new_n674 = new_n672 & new_n673;
  assign new_n675 = ~new_n417 & new_n674;
  assign new_n676 = ~p_1462_168_ & new_n408;
  assign new_n677 = ~new_n423 & new_n676;
  assign new_n678 = ~new_n417 & new_n677;
  assign new_n679 = ~new_n399 & new_n678;
  assign new_n680 = ~new_n405 & new_n679;
  assign new_n681 = ~p_1480_170_ & new_n420;
  assign new_n682 = ~new_n399 & new_n681;
  assign new_n683 = ~p_106_53_ & new_n414;
  assign new_n684 = ~new_n399 & new_n683;
  assign new_n685 = ~new_n423 & new_n684;
  assign new_n686 = ~p_1486_171_ & new_n396;
  assign new_n687 = ~new_n675 & ~new_n680;
  assign new_n688 = ~new_n682 & new_n687;
  assign new_n689 = ~new_n685 & new_n688;
  assign new_n690 = ~new_n686 & new_n689;
  assign new_n691 = new_n436 & ~new_n690;
  assign new_n692 = p_38_11_ & ~new_n432;
  assign new_n693 = ~new_n431 & new_n692;
  assign new_n694 = p_38_11_ & ~new_n428;
  assign new_n695 = ~new_n693 & ~new_n694;
  assign new_n696 = ~new_n691 & new_n695;
  assign new_n697 = ~new_n596 & ~new_n601;
  assign new_n698 = ~new_n636 & new_n697;
  assign new_n699 = ~new_n671 & new_n698;
  assign p_246_3110_ = ~new_n696 | ~new_n699;
  assign new_n701 = p_4526_205_ & new_n348;
  assign new_n702 = ~p_4526_205_ & ~new_n348;
  assign p_373_2994_ = new_n701 | new_n702;
  assign new_n704 = ~new_n320 & ~new_n576;
  assign new_n705 = ~new_n570 & new_n704;
  assign new_n706 = ~new_n576 & new_n586;
  assign new_n707 = new_n387 & ~new_n576;
  assign new_n708 = ~new_n320 & new_n707;
  assign new_n709 = ~new_n705 & ~new_n706;
  assign new_n710 = ~new_n708 & new_n709;
  assign new_n711 = ~new_n584 & new_n710;
  assign new_n712 = new_n567 & ~new_n711;
  assign new_n713 = ~new_n567 & new_n711;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = ~new_n385 & ~new_n714;
  assign new_n716 = new_n387 & new_n704;
  assign new_n717 = ~new_n706 & ~new_n716;
  assign new_n718 = ~new_n584 & new_n717;
  assign new_n719 = new_n567 & new_n718;
  assign new_n720 = ~new_n567 & ~new_n718;
  assign new_n721 = ~new_n719 & ~new_n720;
  assign new_n722 = new_n385 & new_n721;
  assign p_376_3206_ = new_n715 | new_n722;
  assign new_n724 = ~new_n511 & new_n606;
  assign new_n725 = new_n499 & ~new_n593;
  assign new_n726 = new_n499 & new_n597;
  assign new_n727 = p_4526_205_ & new_n726;
  assign new_n728 = ~new_n725 & ~new_n727;
  assign new_n729 = new_n670 & new_n728;
  assign new_n730 = ~new_n511 & ~new_n517;
  assign new_n731 = ~new_n729 & new_n730;
  assign new_n732 = ~new_n724 & ~new_n731;
  assign new_n733 = ~new_n602 & new_n732;
  assign new_n734 = new_n523 & ~new_n733;
  assign new_n735 = ~new_n523 & new_n733;
  assign p_316_3397_ = new_n734 | new_n735;
  assign p_278_536_ = p_163_86_ & p_1_0_;
  assign new_n738 = ~new_n461 & ~new_n467;
  assign new_n739 = new_n641 & new_n738;
  assign new_n740 = ~new_n449 & new_n739;
  assign new_n741 = ~new_n449 & ~new_n461;
  assign new_n742 = ~new_n467 & new_n741;
  assign new_n743 = ~new_n455 & new_n742;
  assign new_n744 = ~new_n467 & new_n648;
  assign new_n745 = ~new_n467 & new_n637;
  assign new_n746 = ~new_n461 & new_n745;
  assign new_n747 = ~new_n740 & ~new_n743;
  assign new_n748 = ~new_n744 & new_n747;
  assign new_n749 = ~new_n746 & new_n748;
  assign new_n750 = ~new_n646 & new_n749;
  assign new_n751 = ~new_n449 & ~new_n455;
  assign new_n752 = ~new_n449 & new_n641;
  assign new_n753 = ~new_n637 & ~new_n752;
  assign new_n754 = ~new_n751 & new_n753;
  assign new_n755 = ~new_n455 & new_n741;
  assign new_n756 = ~new_n461 & new_n637;
  assign new_n757 = ~new_n461 & new_n641;
  assign new_n758 = ~new_n449 & new_n757;
  assign new_n759 = ~new_n755 & ~new_n756;
  assign new_n760 = ~new_n758 & new_n759;
  assign new_n761 = ~new_n648 & new_n760;
  assign new_n762 = p_4394_196_ & new_n452;
  assign new_n763 = new_n761 & new_n762;
  assign new_n764 = ~new_n761 & ~new_n762;
  assign new_n765 = ~new_n763 & ~new_n764;
  assign new_n766 = new_n754 & ~new_n765;
  assign new_n767 = ~new_n754 & new_n765;
  assign new_n768 = ~new_n766 & ~new_n767;
  assign new_n769 = new_n750 & ~new_n768;
  assign new_n770 = ~new_n750 & new_n768;
  assign new_n771 = ~new_n769 & ~new_n770;
  assign new_n772 = new_n455 & ~new_n771;
  assign new_n773 = ~new_n455 & new_n771;
  assign new_n774 = ~new_n772 & ~new_n773;
  assign new_n775 = new_n449 & ~new_n774;
  assign new_n776 = ~new_n449 & new_n774;
  assign new_n777 = ~new_n775 & ~new_n776;
  assign new_n778 = new_n443 & ~new_n777;
  assign new_n779 = ~new_n443 & new_n777;
  assign new_n780 = ~new_n778 & ~new_n779;
  assign new_n781 = new_n461 & ~new_n780;
  assign new_n782 = ~new_n461 & new_n780;
  assign new_n783 = ~new_n781 & ~new_n782;
  assign new_n784 = new_n467 & ~new_n783;
  assign new_n785 = ~new_n467 & new_n783;
  assign new_n786 = ~new_n784 & ~new_n785;
  assign new_n787 = ~new_n339 & new_n367;
  assign new_n788 = ~new_n354 & new_n787;
  assign new_n789 = ~new_n348 & new_n788;
  assign new_n790 = p_4526_205_ & new_n789;
  assign new_n791 = new_n384 & ~new_n790;
  assign new_n792 = ~new_n592 & new_n791;
  assign new_n793 = ~new_n320 & ~new_n567;
  assign new_n794 = ~new_n576 & new_n793;
  assign new_n795 = ~new_n570 & new_n794;
  assign new_n796 = new_n592 & ~new_n795;
  assign new_n797 = ~new_n791 & ~new_n796;
  assign new_n798 = ~new_n792 & ~new_n797;
  assign new_n799 = ~new_n786 & ~new_n798;
  assign new_n800 = ~new_n740 & ~new_n744;
  assign new_n801 = ~new_n746 & new_n800;
  assign new_n802 = ~new_n646 & new_n801;
  assign new_n803 = ~new_n756 & ~new_n758;
  assign new_n804 = ~new_n648 & new_n803;
  assign new_n805 = new_n641 & ~new_n804;
  assign new_n806 = ~new_n641 & new_n804;
  assign new_n807 = ~new_n805 & ~new_n806;
  assign new_n808 = ~new_n753 & ~new_n807;
  assign new_n809 = new_n753 & new_n807;
  assign new_n810 = ~new_n808 & ~new_n809;
  assign new_n811 = ~new_n802 & ~new_n810;
  assign new_n812 = new_n802 & new_n810;
  assign new_n813 = ~new_n811 & ~new_n812;
  assign new_n814 = new_n455 & ~new_n813;
  assign new_n815 = ~new_n455 & new_n813;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817 = new_n449 & ~new_n816;
  assign new_n818 = ~new_n449 & new_n816;
  assign new_n819 = ~new_n817 & ~new_n818;
  assign new_n820 = new_n443 & ~new_n819;
  assign new_n821 = ~new_n443 & new_n819;
  assign new_n822 = ~new_n820 & ~new_n821;
  assign new_n823 = new_n461 & ~new_n822;
  assign new_n824 = ~new_n461 & new_n822;
  assign new_n825 = ~new_n823 & ~new_n824;
  assign new_n826 = new_n467 & ~new_n825;
  assign new_n827 = ~new_n467 & new_n825;
  assign new_n828 = ~new_n826 & ~new_n827;
  assign new_n829 = new_n798 & new_n828;
  assign new_n830 = ~new_n799 & ~new_n829;
  assign new_n831 = ~new_n449 & new_n638;
  assign new_n832 = ~new_n461 & new_n831;
  assign new_n833 = ~new_n455 & new_n832;
  assign new_n834 = new_n655 & ~new_n833;
  assign new_n835 = ~new_n489 & ~new_n495;
  assign new_n836 = ~new_n483 & new_n835;
  assign new_n837 = ~new_n495 & new_n663;
  assign new_n838 = ~new_n495 & new_n657;
  assign new_n839 = ~new_n489 & new_n838;
  assign new_n840 = ~new_n836 & ~new_n837;
  assign new_n841 = ~new_n839 & new_n840;
  assign new_n842 = ~new_n661 & new_n841;
  assign new_n843 = ~new_n483 & ~new_n489;
  assign new_n844 = ~new_n489 & new_n657;
  assign new_n845 = ~new_n663 & ~new_n844;
  assign new_n846 = ~new_n843 & new_n845;
  assign new_n847 = p_4420_201_ & new_n480;
  assign new_n848 = new_n846 & new_n847;
  assign new_n849 = ~new_n846 & ~new_n847;
  assign new_n850 = ~new_n848 & ~new_n849;
  assign new_n851 = new_n842 & ~new_n850;
  assign new_n852 = ~new_n842 & new_n850;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = new_n483 & ~new_n853;
  assign new_n855 = ~new_n483 & new_n853;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = new_n489 & ~new_n856;
  assign new_n858 = ~new_n489 & new_n856;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = new_n477 & ~new_n859;
  assign new_n861 = ~new_n477 & new_n859;
  assign new_n862 = ~new_n860 & ~new_n861;
  assign new_n863 = new_n495 & ~new_n862;
  assign new_n864 = ~new_n495 & new_n862;
  assign new_n865 = ~new_n863 & ~new_n864;
  assign new_n866 = ~new_n798 & ~new_n834;
  assign new_n867 = ~new_n865 & new_n866;
  assign new_n868 = ~new_n655 & new_n798;
  assign new_n869 = ~new_n865 & new_n868;
  assign new_n870 = ~new_n837 & ~new_n839;
  assign new_n871 = ~new_n661 & new_n870;
  assign new_n872 = new_n657 & ~new_n845;
  assign new_n873 = ~new_n657 & new_n845;
  assign new_n874 = ~new_n872 & ~new_n873;
  assign new_n875 = ~new_n871 & ~new_n874;
  assign new_n876 = new_n871 & new_n874;
  assign new_n877 = ~new_n875 & ~new_n876;
  assign new_n878 = new_n483 & ~new_n877;
  assign new_n879 = ~new_n483 & new_n877;
  assign new_n880 = ~new_n878 & ~new_n879;
  assign new_n881 = new_n489 & ~new_n880;
  assign new_n882 = ~new_n489 & new_n880;
  assign new_n883 = ~new_n881 & ~new_n882;
  assign new_n884 = new_n477 & ~new_n883;
  assign new_n885 = ~new_n477 & new_n883;
  assign new_n886 = ~new_n884 & ~new_n885;
  assign new_n887 = new_n495 & ~new_n886;
  assign new_n888 = ~new_n495 & new_n886;
  assign new_n889 = ~new_n887 & ~new_n888;
  assign new_n890 = ~new_n798 & new_n834;
  assign new_n891 = ~new_n889 & new_n890;
  assign new_n892 = new_n655 & new_n798;
  assign new_n893 = ~new_n889 & new_n892;
  assign new_n894 = ~new_n867 & ~new_n869;
  assign new_n895 = ~new_n891 & new_n894;
  assign new_n896 = ~new_n893 & new_n895;
  assign new_n897 = new_n830 & ~new_n896;
  assign new_n898 = ~new_n830 & new_n896;
  assign p_370_3718_ = ~new_n897 & ~new_n898;
  assign new_n900 = p_18_5_ & p_190_113_;
  assign new_n901 = ~new_n490 & ~new_n900;
  assign new_n902 = p_61_24_ & ~p_18_5_;
  assign new_n903 = ~p_4432_203_ & p_18_5_;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = new_n901 & ~new_n904;
  assign new_n906 = ~new_n901 & new_n904;
  assign new_n907 = ~new_n905 & ~new_n906;
  assign new_n908 = p_189_112_ & p_18_5_;
  assign new_n909 = ~new_n472 & ~new_n908;
  assign new_n910 = ~p_18_5_ & p_62_25_;
  assign new_n911 = p_18_5_ & ~p_4437_204_;
  assign new_n912 = ~new_n910 & ~new_n911;
  assign new_n913 = new_n909 & ~new_n912;
  assign new_n914 = ~new_n909 & new_n912;
  assign new_n915 = ~new_n913 & ~new_n914;
  assign new_n916 = p_192_115_ & p_18_5_;
  assign new_n917 = ~new_n478 & ~new_n916;
  assign new_n918 = ~p_18_5_ & p_79_38_;
  assign new_n919 = p_18_5_ & ~p_4420_201_;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = ~new_n917 & ~new_n920;
  assign new_n922 = p_18_5_ & p_191_114_;
  assign new_n923 = ~new_n484 & ~new_n922;
  assign new_n924 = p_60_23_ & ~p_18_5_;
  assign new_n925 = p_18_5_ & ~p_4427_202_;
  assign new_n926 = ~new_n924 & ~new_n925;
  assign new_n927 = new_n923 & ~new_n926;
  assign new_n928 = ~new_n923 & new_n926;
  assign new_n929 = ~new_n927 & ~new_n928;
  assign new_n930 = ~new_n907 & ~new_n915;
  assign new_n931 = new_n921 & new_n930;
  assign new_n932 = ~new_n929 & new_n931;
  assign new_n933 = ~new_n901 & ~new_n904;
  assign new_n934 = ~new_n915 & new_n933;
  assign new_n935 = ~new_n923 & ~new_n926;
  assign new_n936 = ~new_n915 & new_n935;
  assign new_n937 = ~new_n907 & new_n936;
  assign new_n938 = ~new_n909 & ~new_n912;
  assign new_n939 = ~new_n932 & ~new_n934;
  assign new_n940 = ~new_n937 & new_n939;
  assign new_n941 = ~new_n938 & new_n940;
  assign new_n942 = p_18_5_ & p_201_124_;
  assign new_n943 = ~new_n571 & ~new_n942;
  assign new_n944 = p_55_18_ & ~p_18_5_;
  assign new_n945 = p_18_5_ & ~p_3743_193_;
  assign new_n946 = ~new_n944 & ~new_n945;
  assign new_n947 = new_n943 & ~new_n946;
  assign new_n948 = ~new_n943 & new_n946;
  assign new_n949 = ~new_n947 & ~new_n948;
  assign new_n950 = p_18_5_ & p_200_123_;
  assign new_n951 = ~new_n562 & ~new_n950;
  assign new_n952 = p_56_19_ & ~p_18_5_;
  assign new_n953 = ~p_3749_194_ & p_18_5_;
  assign new_n954 = ~new_n952 & ~new_n953;
  assign new_n955 = new_n951 & ~new_n954;
  assign new_n956 = ~new_n951 & new_n954;
  assign new_n957 = ~new_n955 & ~new_n956;
  assign new_n958 = p_18_5_ & p_203_126_;
  assign new_n959 = ~new_n321 & ~new_n958;
  assign new_n960 = p_53_16_ & ~p_18_5_;
  assign new_n961 = p_18_5_ & ~p_3729_191_;
  assign new_n962 = ~new_n960 & ~new_n961;
  assign new_n963 = ~new_n959 & ~new_n962;
  assign new_n964 = p_18_5_ & p_202_125_;
  assign new_n965 = ~new_n315 & ~new_n964;
  assign new_n966 = p_54_17_ & ~p_18_5_;
  assign new_n967 = ~p_3737_192_ & p_18_5_;
  assign new_n968 = ~new_n966 & ~new_n967;
  assign new_n969 = new_n965 & ~new_n968;
  assign new_n970 = ~new_n965 & new_n968;
  assign new_n971 = ~new_n969 & ~new_n970;
  assign new_n972 = ~new_n949 & ~new_n957;
  assign new_n973 = new_n963 & new_n972;
  assign new_n974 = ~new_n971 & new_n973;
  assign new_n975 = ~new_n943 & ~new_n946;
  assign new_n976 = ~new_n957 & new_n975;
  assign new_n977 = ~new_n965 & ~new_n968;
  assign new_n978 = ~new_n957 & new_n977;
  assign new_n979 = ~new_n949 & new_n978;
  assign new_n980 = ~new_n951 & ~new_n954;
  assign new_n981 = ~new_n974 & ~new_n976;
  assign new_n982 = ~new_n979 & new_n981;
  assign new_n983 = ~new_n980 & new_n982;
  assign new_n984 = p_205_128_ & p_18_5_;
  assign new_n985 = ~new_n355 & ~new_n984;
  assign new_n986 = ~p_18_5_ & p_75_34_;
  assign new_n987 = p_18_5_ & ~p_3717_189_;
  assign new_n988 = ~new_n986 & ~new_n987;
  assign new_n989 = new_n985 & ~new_n988;
  assign new_n990 = ~new_n985 & new_n988;
  assign new_n991 = ~new_n989 & ~new_n990;
  assign new_n992 = p_18_5_ & p_204_127_;
  assign new_n993 = ~new_n328 & ~new_n992;
  assign new_n994 = ~p_18_5_ & p_73_32_;
  assign new_n995 = p_18_5_ & ~p_3723_190_;
  assign new_n996 = ~new_n994 & ~new_n995;
  assign new_n997 = new_n993 & ~new_n996;
  assign new_n998 = ~new_n993 & new_n996;
  assign new_n999 = ~new_n997 & ~new_n998;
  assign new_n1000 = p_207_130_ & p_18_5_;
  assign new_n1001 = ~new_n334 & ~new_n1000;
  assign new_n1002 = ~p_18_5_ & p_74_33_;
  assign new_n1003 = p_18_5_ & ~p_3705_187_;
  assign new_n1004 = ~new_n1002 & ~new_n1003;
  assign new_n1005 = new_n1001 & ~new_n1004;
  assign new_n1006 = ~new_n1001 & new_n1004;
  assign new_n1007 = ~new_n1005 & ~new_n1006;
  assign new_n1008 = p_18_5_ & p_206_129_;
  assign new_n1009 = ~new_n349 & ~new_n1008;
  assign new_n1010 = ~p_18_5_ & p_76_35_;
  assign new_n1011 = p_18_5_ & ~p_3711_188_;
  assign new_n1012 = ~new_n1010 & ~new_n1011;
  assign new_n1013 = new_n1009 & ~new_n1012;
  assign new_n1014 = ~new_n1009 & new_n1012;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = p_18_5_ & p_198_121_;
  assign new_n1017 = ~new_n340 & ~new_n1016;
  assign new_n1018 = ~p_18_5_ & ~new_n1017;
  assign new_n1019 = ~p_18_5_ & p_70_31_;
  assign new_n1020 = ~p_18_5_ & ~new_n1019;
  assign new_n1021 = ~new_n1018 & ~new_n1020;
  assign new_n1022 = new_n1018 & new_n1020;
  assign new_n1023 = ~new_n1021 & ~new_n1022;
  assign new_n1024 = ~new_n991 & ~new_n999;
  assign new_n1025 = ~new_n1007 & new_n1024;
  assign new_n1026 = ~new_n1015 & new_n1025;
  assign new_n1027 = ~new_n1023 & new_n1026;
  assign new_n1028 = p_89_48_ & new_n1027;
  assign new_n1029 = ~new_n1001 & ~new_n1004;
  assign new_n1030 = new_n1024 & new_n1029;
  assign new_n1031 = ~new_n1015 & new_n1030;
  assign new_n1032 = new_n1018 & ~new_n1020;
  assign new_n1033 = ~new_n991 & new_n1032;
  assign new_n1034 = ~new_n1015 & new_n1033;
  assign new_n1035 = ~new_n999 & new_n1034;
  assign new_n1036 = ~new_n1007 & new_n1035;
  assign new_n1037 = ~new_n985 & ~new_n988;
  assign new_n1038 = ~new_n999 & new_n1037;
  assign new_n1039 = ~new_n1009 & ~new_n1012;
  assign new_n1040 = ~new_n999 & new_n1039;
  assign new_n1041 = ~new_n991 & new_n1040;
  assign new_n1042 = ~new_n993 & ~new_n996;
  assign new_n1043 = ~new_n1031 & ~new_n1036;
  assign new_n1044 = ~new_n1038 & new_n1043;
  assign new_n1045 = ~new_n1041 & new_n1044;
  assign new_n1046 = ~new_n1042 & new_n1045;
  assign new_n1047 = ~new_n1028 & new_n1046;
  assign new_n1048 = ~new_n983 & new_n1047;
  assign new_n1049 = new_n959 & ~new_n962;
  assign new_n1050 = ~new_n959 & new_n962;
  assign new_n1051 = ~new_n1049 & ~new_n1050;
  assign new_n1052 = ~new_n957 & ~new_n971;
  assign new_n1053 = ~new_n949 & new_n1052;
  assign new_n1054 = ~new_n1051 & new_n1053;
  assign new_n1055 = new_n983 & ~new_n1054;
  assign new_n1056 = ~new_n1047 & ~new_n1055;
  assign new_n1057 = ~new_n1048 & ~new_n1056;
  assign new_n1058 = p_18_5_ & p_194_117_;
  assign new_n1059 = ~new_n462 & ~new_n1058;
  assign new_n1060 = ~p_18_5_ & p_81_40_;
  assign new_n1061 = p_18_5_ & ~p_4410_199_;
  assign new_n1062 = ~new_n1060 & ~new_n1061;
  assign new_n1063 = new_n1059 & ~new_n1062;
  assign new_n1064 = ~new_n1059 & new_n1062;
  assign new_n1065 = ~new_n1063 & ~new_n1064;
  assign new_n1066 = p_193_116_ & p_18_5_;
  assign new_n1067 = ~new_n438 & ~new_n1066;
  assign new_n1068 = ~p_18_5_ & p_80_39_;
  assign new_n1069 = p_18_5_ & ~p_4415_200_;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = new_n1067 & ~new_n1070;
  assign new_n1072 = ~new_n1067 & new_n1070;
  assign new_n1073 = ~new_n1071 & ~new_n1072;
  assign new_n1074 = p_18_5_ & p_196_119_;
  assign new_n1075 = ~new_n444 & ~new_n1074;
  assign new_n1076 = ~p_18_5_ & p_78_37_;
  assign new_n1077 = p_18_5_ & ~p_4400_197_;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = new_n1075 & ~new_n1078;
  assign new_n1080 = ~new_n1075 & new_n1078;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign new_n1082 = p_195_118_ & p_18_5_;
  assign new_n1083 = ~new_n456 & ~new_n1082;
  assign new_n1084 = ~p_18_5_ & p_59_22_;
  assign new_n1085 = ~p_4405_198_ & p_18_5_;
  assign new_n1086 = ~new_n1084 & ~new_n1085;
  assign new_n1087 = new_n1083 & ~new_n1086;
  assign new_n1088 = ~new_n1083 & new_n1086;
  assign new_n1089 = ~new_n1087 & ~new_n1088;
  assign new_n1090 = p_18_5_ & p_187_110_;
  assign new_n1091 = ~new_n450 & ~new_n1090;
  assign new_n1092 = ~p_18_5_ & p_77_36_;
  assign new_n1093 = ~p_4394_196_ & p_18_5_;
  assign new_n1094 = ~new_n1092 & ~new_n1093;
  assign new_n1095 = new_n1091 & ~new_n1094;
  assign new_n1096 = ~new_n1091 & new_n1094;
  assign new_n1097 = ~new_n1095 & ~new_n1096;
  assign new_n1098 = ~new_n1065 & ~new_n1073;
  assign new_n1099 = ~new_n1081 & new_n1098;
  assign new_n1100 = ~new_n1089 & new_n1099;
  assign new_n1101 = ~new_n1097 & new_n1100;
  assign new_n1102 = ~new_n1057 & new_n1101;
  assign new_n1103 = ~new_n1075 & ~new_n1078;
  assign new_n1104 = new_n1098 & new_n1103;
  assign new_n1105 = ~new_n1089 & new_n1104;
  assign new_n1106 = ~new_n1091 & ~new_n1094;
  assign new_n1107 = ~new_n1065 & new_n1106;
  assign new_n1108 = ~new_n1089 & new_n1107;
  assign new_n1109 = ~new_n1073 & new_n1108;
  assign new_n1110 = ~new_n1081 & new_n1109;
  assign new_n1111 = ~new_n1059 & ~new_n1062;
  assign new_n1112 = ~new_n1073 & new_n1111;
  assign new_n1113 = ~new_n1083 & ~new_n1086;
  assign new_n1114 = ~new_n1073 & new_n1113;
  assign new_n1115 = ~new_n1065 & new_n1114;
  assign new_n1116 = ~new_n1067 & ~new_n1070;
  assign new_n1117 = ~new_n1105 & ~new_n1110;
  assign new_n1118 = ~new_n1112 & new_n1117;
  assign new_n1119 = ~new_n1115 & new_n1118;
  assign new_n1120 = ~new_n1116 & new_n1119;
  assign new_n1121 = ~new_n1102 & new_n1120;
  assign new_n1122 = ~new_n941 & new_n1121;
  assign new_n1123 = new_n917 & ~new_n920;
  assign new_n1124 = ~new_n917 & new_n920;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = ~new_n915 & ~new_n929;
  assign new_n1127 = ~new_n907 & new_n1126;
  assign new_n1128 = ~new_n1125 & new_n1127;
  assign new_n1129 = new_n941 & ~new_n1128;
  assign new_n1130 = ~new_n1121 & ~new_n1129;
  assign p_252_3450_ = new_n1122 | new_n1130;
  assign new_n1132 = new_n561 & new_n597;
  assign new_n1133 = new_n499 & new_n1132;
  assign new_n1134 = p_4526_205_ & new_n1133;
  assign new_n1135 = new_n561 & ~new_n670;
  assign new_n1136 = new_n499 & new_n561;
  assign new_n1137 = ~new_n593 & new_n1136;
  assign new_n1138 = ~new_n1134 & ~new_n1135;
  assign new_n1139 = ~new_n1137 & new_n1138;
  assign new_n1140 = new_n635 & new_n1139;
  assign new_n1141 = new_n427 & ~new_n1140;
  assign new_n1142 = new_n690 & ~new_n1141;
  assign new_n1143 = ~new_n436 & new_n695;
  assign new_n1144 = ~new_n1142 & ~new_n1143;
  assign new_n1145 = ~new_n695 & new_n1142;
  assign p_273_3402_ = new_n1144 | new_n1145;
  assign new_n1147 = ~new_n417 & ~new_n423;
  assign new_n1148 = new_n676 & new_n1147;
  assign new_n1149 = ~new_n405 & new_n1148;
  assign new_n1150 = ~new_n405 & ~new_n423;
  assign new_n1151 = ~new_n411 & new_n1150;
  assign new_n1152 = ~new_n417 & new_n1151;
  assign new_n1153 = ~new_n1140 & new_n1152;
  assign new_n1154 = ~new_n423 & new_n683;
  assign new_n1155 = ~new_n423 & new_n672;
  assign new_n1156 = ~new_n417 & new_n1155;
  assign new_n1157 = ~new_n1149 & ~new_n1153;
  assign new_n1158 = ~new_n1154 & new_n1157;
  assign new_n1159 = ~new_n1156 & new_n1158;
  assign new_n1160 = ~new_n681 & new_n1159;
  assign new_n1161 = new_n399 & ~new_n1160;
  assign new_n1162 = ~new_n399 & new_n1160;
  assign p_327_3408_ = new_n1161 | new_n1162;
  assign new_n1164 = ~new_n405 & ~new_n417;
  assign new_n1165 = ~new_n423 & new_n1164;
  assign new_n1166 = ~new_n411 & new_n1165;
  assign new_n1167 = ~new_n1149 & ~new_n1166;
  assign new_n1168 = ~new_n1154 & new_n1167;
  assign new_n1169 = ~new_n1156 & new_n1168;
  assign new_n1170 = ~new_n681 & new_n1169;
  assign new_n1171 = ~new_n405 & ~new_n411;
  assign new_n1172 = ~new_n405 & new_n676;
  assign new_n1173 = ~new_n672 & ~new_n1172;
  assign new_n1174 = ~new_n1171 & new_n1173;
  assign new_n1175 = ~new_n411 & new_n1164;
  assign new_n1176 = ~new_n417 & new_n672;
  assign new_n1177 = ~new_n417 & new_n676;
  assign new_n1178 = ~new_n405 & new_n1177;
  assign new_n1179 = ~new_n1175 & ~new_n1176;
  assign new_n1180 = ~new_n1178 & new_n1179;
  assign new_n1181 = ~new_n683 & new_n1180;
  assign new_n1182 = p_1462_168_ & ~new_n408;
  assign new_n1183 = new_n1181 & new_n1182;
  assign new_n1184 = ~new_n1181 & ~new_n1182;
  assign new_n1185 = ~new_n1183 & ~new_n1184;
  assign new_n1186 = new_n1174 & ~new_n1185;
  assign new_n1187 = ~new_n1174 & new_n1185;
  assign new_n1188 = ~new_n1186 & ~new_n1187;
  assign new_n1189 = new_n1170 & ~new_n1188;
  assign new_n1190 = ~new_n1170 & new_n1188;
  assign new_n1191 = ~new_n1189 & ~new_n1190;
  assign new_n1192 = new_n411 & ~new_n1191;
  assign new_n1193 = ~new_n411 & new_n1191;
  assign new_n1194 = ~new_n1192 & ~new_n1193;
  assign new_n1195 = new_n405 & ~new_n1194;
  assign new_n1196 = ~new_n405 & new_n1194;
  assign new_n1197 = ~new_n1195 & ~new_n1196;
  assign new_n1198 = new_n399 & ~new_n1197;
  assign new_n1199 = ~new_n399 & new_n1197;
  assign new_n1200 = ~new_n1198 & ~new_n1199;
  assign new_n1201 = new_n417 & ~new_n1200;
  assign new_n1202 = ~new_n417 & new_n1200;
  assign new_n1203 = ~new_n1201 & ~new_n1202;
  assign new_n1204 = new_n423 & ~new_n1203;
  assign new_n1205 = ~new_n423 & new_n1203;
  assign new_n1206 = ~new_n1204 & ~new_n1205;
  assign new_n1207 = ~new_n511 & new_n603;
  assign new_n1208 = ~new_n523 & new_n1207;
  assign new_n1209 = ~new_n517 & new_n1208;
  assign new_n1210 = ~new_n539 & ~new_n551;
  assign new_n1211 = ~new_n557 & new_n1210;
  assign new_n1212 = ~new_n545 & new_n1211;
  assign new_n1213 = new_n1209 & new_n1212;
  assign new_n1214 = new_n789 & new_n795;
  assign new_n1215 = ~new_n477 & ~new_n489;
  assign new_n1216 = ~new_n495 & new_n1215;
  assign new_n1217 = ~new_n483 & new_n1216;
  assign new_n1218 = new_n833 & new_n1217;
  assign new_n1219 = new_n1213 & new_n1214;
  assign new_n1220 = new_n1218 & new_n1219;
  assign new_n1221 = p_4526_205_ & new_n1220;
  assign new_n1222 = ~new_n655 & new_n1217;
  assign new_n1223 = new_n669 & ~new_n1222;
  assign new_n1224 = new_n1213 & ~new_n1223;
  assign new_n1225 = ~new_n384 & new_n795;
  assign new_n1226 = new_n592 & ~new_n1225;
  assign new_n1227 = new_n1213 & new_n1218;
  assign new_n1228 = ~new_n1226 & new_n1227;
  assign new_n1229 = ~new_n620 & new_n1212;
  assign new_n1230 = new_n634 & ~new_n1229;
  assign new_n1231 = ~new_n1221 & ~new_n1224;
  assign new_n1232 = ~new_n1228 & new_n1231;
  assign new_n1233 = new_n1230 & new_n1232;
  assign new_n1234 = ~new_n1206 & ~new_n1233;
  assign new_n1235 = ~new_n1149 & ~new_n1154;
  assign new_n1236 = ~new_n1156 & new_n1235;
  assign new_n1237 = ~new_n681 & new_n1236;
  assign new_n1238 = ~new_n1176 & ~new_n1178;
  assign new_n1239 = ~new_n683 & new_n1238;
  assign new_n1240 = new_n676 & ~new_n1239;
  assign new_n1241 = ~new_n676 & new_n1239;
  assign new_n1242 = ~new_n1240 & ~new_n1241;
  assign new_n1243 = ~new_n1173 & ~new_n1242;
  assign new_n1244 = new_n1173 & new_n1242;
  assign new_n1245 = ~new_n1243 & ~new_n1244;
  assign new_n1246 = ~new_n1237 & ~new_n1245;
  assign new_n1247 = new_n1237 & new_n1245;
  assign new_n1248 = ~new_n1246 & ~new_n1247;
  assign new_n1249 = new_n411 & ~new_n1248;
  assign new_n1250 = ~new_n411 & new_n1248;
  assign new_n1251 = ~new_n1249 & ~new_n1250;
  assign new_n1252 = new_n405 & ~new_n1251;
  assign new_n1253 = ~new_n405 & new_n1251;
  assign new_n1254 = ~new_n1252 & ~new_n1253;
  assign new_n1255 = new_n399 & ~new_n1254;
  assign new_n1256 = ~new_n399 & new_n1254;
  assign new_n1257 = ~new_n1255 & ~new_n1256;
  assign new_n1258 = new_n417 & ~new_n1257;
  assign new_n1259 = ~new_n417 & new_n1257;
  assign new_n1260 = ~new_n1258 & ~new_n1259;
  assign new_n1261 = new_n423 & ~new_n1260;
  assign new_n1262 = ~new_n423 & new_n1260;
  assign new_n1263 = ~new_n1261 & ~new_n1262;
  assign new_n1264 = new_n1233 & new_n1263;
  assign new_n1265 = ~new_n1234 & ~new_n1264;
  assign new_n1266 = ~new_n405 & new_n673;
  assign new_n1267 = ~new_n417 & new_n1266;
  assign new_n1268 = ~new_n411 & new_n1267;
  assign new_n1269 = new_n690 & ~new_n1268;
  assign new_n1270 = ~new_n436 & ~new_n693;
  assign new_n1271 = ~new_n694 & new_n1270;
  assign new_n1272 = ~p_38_11_ & new_n432;
  assign new_n1273 = new_n1143 & new_n1272;
  assign new_n1274 = ~new_n1143 & ~new_n1272;
  assign new_n1275 = ~new_n1273 & ~new_n1274;
  assign new_n1276 = new_n1271 & ~new_n1275;
  assign new_n1277 = ~new_n1271 & new_n1275;
  assign new_n1278 = ~new_n1276 & ~new_n1277;
  assign new_n1279 = new_n435 & ~new_n1278;
  assign new_n1280 = ~new_n435 & new_n1278;
  assign new_n1281 = ~new_n1279 & ~new_n1280;
  assign new_n1282 = new_n431 & ~new_n1281;
  assign new_n1283 = ~new_n431 & new_n1281;
  assign new_n1284 = ~new_n1282 & ~new_n1283;
  assign new_n1285 = ~new_n1233 & ~new_n1269;
  assign new_n1286 = ~new_n1284 & new_n1285;
  assign new_n1287 = ~new_n690 & new_n1233;
  assign new_n1288 = ~new_n1284 & new_n1287;
  assign new_n1289 = new_n692 & ~new_n695;
  assign new_n1290 = ~new_n692 & new_n695;
  assign new_n1291 = ~new_n1289 & ~new_n1290;
  assign new_n1292 = ~new_n695 & ~new_n1291;
  assign new_n1293 = new_n695 & new_n1291;
  assign new_n1294 = ~new_n1292 & ~new_n1293;
  assign new_n1295 = new_n435 & ~new_n1294;
  assign new_n1296 = ~new_n435 & new_n1294;
  assign new_n1297 = ~new_n1295 & ~new_n1296;
  assign new_n1298 = new_n431 & ~new_n1297;
  assign new_n1299 = ~new_n431 & new_n1297;
  assign new_n1300 = ~new_n1298 & ~new_n1299;
  assign new_n1301 = ~new_n1233 & new_n1269;
  assign new_n1302 = ~new_n1300 & new_n1301;
  assign new_n1303 = new_n690 & new_n1233;
  assign new_n1304 = ~new_n1300 & new_n1303;
  assign new_n1305 = ~new_n1286 & ~new_n1288;
  assign new_n1306 = ~new_n1302 & new_n1305;
  assign new_n1307 = ~new_n1304 & new_n1306;
  assign new_n1308 = new_n1265 & ~new_n1307;
  assign new_n1309 = ~new_n1265 & new_n1307;
  assign p_338_3716_ = ~new_n1308 & ~new_n1309;
  assign new_n1311 = p_152_75_ & p_230_153_;
  assign new_n1312 = p_218_141_ & new_n1311;
  assign p_406_388_ = ~p_210_133_ | ~new_n1312;
  assign new_n1314 = new_n431 & new_n1272;
  assign new_n1315 = ~new_n431 & ~new_n1272;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = ~new_n1142 & new_n1316;
  assign new_n1318 = new_n431 & new_n692;
  assign new_n1319 = ~new_n431 & ~new_n692;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = new_n1142 & ~new_n1320;
  assign p_422_3451_ = new_n1317 | new_n1321;
  assign new_n1323 = ~new_n523 & ~new_n529;
  assign new_n1324 = new_n606 & new_n1323;
  assign new_n1325 = ~new_n511 & new_n1324;
  assign new_n1326 = ~new_n511 & ~new_n523;
  assign new_n1327 = ~new_n529 & new_n1326;
  assign new_n1328 = ~new_n517 & new_n1327;
  assign new_n1329 = ~new_n529 & new_n613;
  assign new_n1330 = ~new_n529 & new_n602;
  assign new_n1331 = ~new_n523 & new_n1330;
  assign new_n1332 = ~new_n1325 & ~new_n1328;
  assign new_n1333 = ~new_n1329 & new_n1332;
  assign new_n1334 = ~new_n1331 & new_n1333;
  assign new_n1335 = ~new_n611 & new_n1334;
  assign new_n1336 = ~new_n602 & ~new_n724;
  assign new_n1337 = ~new_n730 & new_n1336;
  assign new_n1338 = ~new_n517 & new_n1326;
  assign new_n1339 = ~new_n523 & new_n602;
  assign new_n1340 = ~new_n523 & new_n606;
  assign new_n1341 = ~new_n511 & new_n1340;
  assign new_n1342 = ~new_n1338 & ~new_n1339;
  assign new_n1343 = ~new_n1341 & new_n1342;
  assign new_n1344 = ~new_n613 & new_n1343;
  assign new_n1345 = p_2211_176_ & new_n514;
  assign new_n1346 = new_n1344 & new_n1345;
  assign new_n1347 = ~new_n1344 & ~new_n1345;
  assign new_n1348 = ~new_n1346 & ~new_n1347;
  assign new_n1349 = new_n1337 & ~new_n1348;
  assign new_n1350 = ~new_n1337 & new_n1348;
  assign new_n1351 = ~new_n1349 & ~new_n1350;
  assign new_n1352 = new_n1335 & ~new_n1351;
  assign new_n1353 = ~new_n1335 & new_n1351;
  assign new_n1354 = ~new_n1352 & ~new_n1353;
  assign new_n1355 = new_n517 & ~new_n1354;
  assign new_n1356 = ~new_n517 & new_n1354;
  assign new_n1357 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = new_n511 & ~new_n1357;
  assign new_n1359 = ~new_n511 & new_n1357;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = new_n505 & ~new_n1360;
  assign new_n1362 = ~new_n505 & new_n1360;
  assign new_n1363 = ~new_n1361 & ~new_n1362;
  assign new_n1364 = new_n523 & ~new_n1363;
  assign new_n1365 = ~new_n523 & new_n1363;
  assign new_n1366 = ~new_n1364 & ~new_n1365;
  assign new_n1367 = new_n529 & ~new_n1366;
  assign new_n1368 = ~new_n529 & new_n1366;
  assign new_n1369 = ~new_n1367 & ~new_n1368;
  assign new_n1370 = new_n1218 & ~new_n1226;
  assign new_n1371 = new_n1214 & new_n1218;
  assign new_n1372 = p_4526_205_ & new_n1371;
  assign new_n1373 = ~new_n1370 & ~new_n1372;
  assign new_n1374 = new_n1223 & new_n1373;
  assign new_n1375 = ~new_n1369 & ~new_n1374;
  assign new_n1376 = ~new_n1325 & ~new_n1329;
  assign new_n1377 = ~new_n1331 & new_n1376;
  assign new_n1378 = ~new_n611 & new_n1377;
  assign new_n1379 = ~new_n1339 & ~new_n1341;
  assign new_n1380 = ~new_n613 & new_n1379;
  assign new_n1381 = new_n606 & ~new_n1380;
  assign new_n1382 = ~new_n606 & new_n1380;
  assign new_n1383 = ~new_n1381 & ~new_n1382;
  assign new_n1384 = ~new_n1336 & ~new_n1383;
  assign new_n1385 = new_n1336 & new_n1383;
  assign new_n1386 = ~new_n1384 & ~new_n1385;
  assign new_n1387 = ~new_n1378 & ~new_n1386;
  assign new_n1388 = new_n1378 & new_n1386;
  assign new_n1389 = ~new_n1387 & ~new_n1388;
  assign new_n1390 = new_n517 & ~new_n1389;
  assign new_n1391 = ~new_n517 & new_n1389;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = new_n511 & ~new_n1392;
  assign new_n1394 = ~new_n511 & new_n1392;
  assign new_n1395 = ~new_n1393 & ~new_n1394;
  assign new_n1396 = new_n505 & ~new_n1395;
  assign new_n1397 = ~new_n505 & new_n1395;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = new_n523 & ~new_n1398;
  assign new_n1400 = ~new_n523 & new_n1398;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = new_n529 & ~new_n1401;
  assign new_n1403 = ~new_n529 & new_n1401;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = new_n1374 & new_n1404;
  assign new_n1406 = ~new_n1375 & ~new_n1405;
  assign new_n1407 = new_n620 & ~new_n1209;
  assign new_n1408 = ~new_n551 & ~new_n557;
  assign new_n1409 = ~new_n545 & new_n1408;
  assign new_n1410 = ~new_n557 & new_n628;
  assign new_n1411 = ~new_n557 & new_n622;
  assign new_n1412 = ~new_n551 & new_n1411;
  assign new_n1413 = ~new_n1409 & ~new_n1410;
  assign new_n1414 = ~new_n1412 & new_n1413;
  assign new_n1415 = ~new_n626 & new_n1414;
  assign new_n1416 = ~new_n545 & ~new_n551;
  assign new_n1417 = ~new_n551 & new_n622;
  assign new_n1418 = ~new_n628 & ~new_n1417;
  assign new_n1419 = ~new_n1416 & new_n1418;
  assign new_n1420 = p_2239_181_ & ~new_n542;
  assign new_n1421 = new_n1419 & new_n1420;
  assign new_n1422 = ~new_n1419 & ~new_n1420;
  assign new_n1423 = ~new_n1421 & ~new_n1422;
  assign new_n1424 = new_n1415 & ~new_n1423;
  assign new_n1425 = ~new_n1415 & new_n1423;
  assign new_n1426 = ~new_n1424 & ~new_n1425;
  assign new_n1427 = new_n545 & ~new_n1426;
  assign new_n1428 = ~new_n545 & new_n1426;
  assign new_n1429 = ~new_n1427 & ~new_n1428;
  assign new_n1430 = new_n551 & ~new_n1429;
  assign new_n1431 = ~new_n551 & new_n1429;
  assign new_n1432 = ~new_n1430 & ~new_n1431;
  assign new_n1433 = new_n539 & ~new_n1432;
  assign new_n1434 = ~new_n539 & new_n1432;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = new_n557 & ~new_n1435;
  assign new_n1437 = ~new_n557 & new_n1435;
  assign new_n1438 = ~new_n1436 & ~new_n1437;
  assign new_n1439 = ~new_n1374 & ~new_n1407;
  assign new_n1440 = ~new_n1438 & new_n1439;
  assign new_n1441 = ~new_n620 & new_n1374;
  assign new_n1442 = ~new_n1438 & new_n1441;
  assign new_n1443 = ~new_n1410 & ~new_n1412;
  assign new_n1444 = ~new_n626 & new_n1443;
  assign new_n1445 = new_n622 & ~new_n1418;
  assign new_n1446 = ~new_n622 & new_n1418;
  assign new_n1447 = ~new_n1445 & ~new_n1446;
  assign new_n1448 = ~new_n1444 & ~new_n1447;
  assign new_n1449 = new_n1444 & new_n1447;
  assign new_n1450 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = new_n545 & ~new_n1450;
  assign new_n1452 = ~new_n545 & new_n1450;
  assign new_n1453 = ~new_n1451 & ~new_n1452;
  assign new_n1454 = new_n551 & ~new_n1453;
  assign new_n1455 = ~new_n551 & new_n1453;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = new_n539 & ~new_n1456;
  assign new_n1458 = ~new_n539 & new_n1456;
  assign new_n1459 = ~new_n1457 & ~new_n1458;
  assign new_n1460 = new_n557 & ~new_n1459;
  assign new_n1461 = ~new_n557 & new_n1459;
  assign new_n1462 = ~new_n1460 & ~new_n1461;
  assign new_n1463 = ~new_n1374 & new_n1407;
  assign new_n1464 = ~new_n1462 & new_n1463;
  assign new_n1465 = new_n620 & new_n1374;
  assign new_n1466 = ~new_n1462 & new_n1465;
  assign new_n1467 = ~new_n1440 & ~new_n1442;
  assign new_n1468 = ~new_n1464 & new_n1467;
  assign new_n1469 = ~new_n1466 & new_n1468;
  assign new_n1470 = new_n1406 & ~new_n1469;
  assign new_n1471 = ~new_n1406 & new_n1469;
  assign p_321_3715_ = ~new_n1470 & ~new_n1471;
  assign new_n1473 = ~new_n579 & new_n592;
  assign new_n1474 = ~new_n385 & ~new_n1473;
  assign new_n1475 = new_n385 & ~new_n592;
  assign new_n1476 = ~new_n1474 & ~new_n1475;
  assign new_n1477 = ~new_n455 & ~new_n1476;
  assign new_n1478 = ~new_n641 & ~new_n1477;
  assign new_n1479 = new_n449 & ~new_n1478;
  assign new_n1480 = ~new_n449 & new_n1478;
  assign p_368_3431_ = new_n1479 | new_n1480;
  assign new_n1482 = p_18_5_ & p_167_90_;
  assign new_n1483 = p_18_5_ & ~new_n1482;
  assign new_n1484 = ~new_n393 & ~new_n1483;
  assign new_n1485 = p_18_5_ & ~p_1480_170_;
  assign new_n1486 = ~p_18_5_ & p_112_57_;
  assign new_n1487 = ~new_n1485 & ~new_n1486;
  assign new_n1488 = ~new_n1484 & ~new_n1487;
  assign new_n1489 = new_n1484 & new_n1487;
  assign new_n1490 = ~new_n1488 & ~new_n1489;
  assign new_n1491 = p_166_89_ & p_18_5_;
  assign new_n1492 = p_18_5_ & ~new_n1491;
  assign new_n1493 = ~new_n393 & ~new_n1492;
  assign new_n1494 = p_18_5_ & ~p_1486_171_;
  assign new_n1495 = ~p_18_5_ & p_88_47_;
  assign new_n1496 = ~new_n1494 & ~new_n1495;
  assign new_n1497 = ~new_n1493 & ~new_n1496;
  assign new_n1498 = new_n1493 & new_n1496;
  assign new_n1499 = ~new_n1497 & ~new_n1498;
  assign new_n1500 = p_169_92_ & p_18_5_;
  assign new_n1501 = p_18_5_ & ~new_n1500;
  assign new_n1502 = ~new_n393 & ~new_n1501;
  assign new_n1503 = p_18_5_ & ~p_1469_169_;
  assign new_n1504 = ~p_18_5_ & p_111_56_;
  assign new_n1505 = ~new_n1503 & ~new_n1504;
  assign new_n1506 = ~new_n1502 & ~new_n1505;
  assign new_n1507 = new_n1502 & new_n1505;
  assign new_n1508 = ~new_n1506 & ~new_n1507;
  assign new_n1509 = p_18_5_ & p_168_91_;
  assign new_n1510 = p_18_5_ & ~new_n1509;
  assign new_n1511 = ~new_n393 & ~new_n1510;
  assign new_n1512 = p_18_5_ & ~p_106_53_;
  assign new_n1513 = ~p_18_5_ & p_87_46_;
  assign new_n1514 = ~new_n1512 & ~new_n1513;
  assign new_n1515 = ~new_n1511 & ~new_n1514;
  assign new_n1516 = new_n1511 & new_n1514;
  assign new_n1517 = ~new_n1515 & ~new_n1516;
  assign new_n1518 = p_18_5_ & ~p_1462_168_;
  assign new_n1519 = p_113_58_ & ~p_18_5_;
  assign new_n1520 = ~new_n1518 & ~new_n1519;
  assign new_n1521 = new_n393 & ~new_n1520;
  assign new_n1522 = ~new_n393 & new_n1520;
  assign new_n1523 = ~new_n1521 & ~new_n1522;
  assign new_n1524 = ~new_n1490 & ~new_n1499;
  assign new_n1525 = ~new_n1508 & new_n1524;
  assign new_n1526 = ~new_n1517 & new_n1525;
  assign new_n1527 = ~new_n1523 & new_n1526;
  assign new_n1528 = p_4528_206_ & ~p_2204_174_;
  assign new_n1529 = ~p_38_11_ & ~new_n1528;
  assign new_n1530 = p_38_11_ & new_n1528;
  assign new_n1531 = ~new_n1529 & ~new_n1530;
  assign new_n1532 = p_4528_206_ & ~p_1455_166_;
  assign new_n1533 = ~p_38_11_ & ~new_n1532;
  assign new_n1534 = p_38_11_ & new_n1532;
  assign new_n1535 = ~new_n1533 & ~new_n1534;
  assign new_n1536 = ~new_n1531 & ~new_n1535;
  assign new_n1537 = new_n1527 & new_n1536;
  assign new_n1538 = new_n1101 & new_n1128;
  assign new_n1539 = p_18_5_ & p_178_101_;
  assign new_n1540 = ~new_n525 & ~new_n1539;
  assign new_n1541 = p_18_5_ & ~p_2230_179_;
  assign new_n1542 = ~p_18_5_ & p_85_44_;
  assign new_n1543 = ~new_n1541 & ~new_n1542;
  assign new_n1544 = new_n1540 & ~new_n1543;
  assign new_n1545 = ~new_n1540 & new_n1543;
  assign new_n1546 = ~new_n1544 & ~new_n1545;
  assign new_n1547 = p_18_5_ & p_177_100_;
  assign new_n1548 = p_18_5_ & ~new_n1547;
  assign new_n1549 = ~new_n393 & ~new_n1548;
  assign new_n1550 = p_18_5_ & ~p_2236_180_;
  assign new_n1551 = ~p_18_5_ & p_64_27_;
  assign new_n1552 = ~new_n1550 & ~new_n1551;
  assign new_n1553 = ~new_n1549 & ~new_n1552;
  assign new_n1554 = new_n1549 & new_n1552;
  assign new_n1555 = ~new_n1553 & ~new_n1554;
  assign new_n1556 = p_18_5_ & p_180_103_;
  assign new_n1557 = ~new_n507 & ~new_n1556;
  assign new_n1558 = p_18_5_ & ~p_2218_177_;
  assign new_n1559 = ~p_18_5_ & p_83_42_;
  assign new_n1560 = ~new_n1558 & ~new_n1559;
  assign new_n1561 = new_n1557 & ~new_n1560;
  assign new_n1562 = ~new_n1557 & new_n1560;
  assign new_n1563 = ~new_n1561 & ~new_n1562;
  assign new_n1564 = p_179_102_ & p_18_5_;
  assign new_n1565 = ~new_n519 & ~new_n1564;
  assign new_n1566 = p_18_5_ & ~p_2224_178_;
  assign new_n1567 = ~p_18_5_ & p_84_43_;
  assign new_n1568 = ~new_n1566 & ~new_n1567;
  assign new_n1569 = new_n1565 & ~new_n1568;
  assign new_n1570 = ~new_n1565 & new_n1568;
  assign new_n1571 = ~new_n1569 & ~new_n1570;
  assign new_n1572 = p_18_5_ & p_171_94_;
  assign new_n1573 = ~new_n513 & ~new_n1572;
  assign new_n1574 = ~p_2211_176_ & p_18_5_;
  assign new_n1575 = ~p_18_5_ & p_65_28_;
  assign new_n1576 = ~new_n1574 & ~new_n1575;
  assign new_n1577 = new_n1573 & ~new_n1576;
  assign new_n1578 = ~new_n1573 & new_n1576;
  assign new_n1579 = ~new_n1577 & ~new_n1578;
  assign new_n1580 = ~new_n1546 & ~new_n1555;
  assign new_n1581 = ~new_n1563 & new_n1580;
  assign new_n1582 = ~new_n1571 & new_n1581;
  assign new_n1583 = ~new_n1579 & new_n1582;
  assign new_n1584 = p_18_5_ & p_173_96_;
  assign new_n1585 = p_18_5_ & ~new_n1584;
  assign new_n1586 = ~new_n393 & ~new_n1585;
  assign new_n1587 = p_18_5_ & ~p_2256_184_;
  assign new_n1588 = ~p_18_5_ & p_110_55_;
  assign new_n1589 = ~new_n1587 & ~new_n1588;
  assign new_n1590 = ~new_n1586 & ~new_n1589;
  assign new_n1591 = new_n1586 & new_n1589;
  assign new_n1592 = ~new_n1590 & ~new_n1591;
  assign new_n1593 = p_18_5_ & p_175_98_;
  assign new_n1594 = p_18_5_ & ~new_n1593;
  assign new_n1595 = ~new_n393 & ~new_n1594;
  assign new_n1596 = p_18_5_ & ~p_2247_182_;
  assign new_n1597 = ~p_18_5_ & p_86_45_;
  assign new_n1598 = ~new_n1596 & ~new_n1597;
  assign new_n1599 = ~new_n1595 & ~new_n1598;
  assign new_n1600 = new_n1595 & new_n1598;
  assign new_n1601 = ~new_n1599 & ~new_n1600;
  assign new_n1602 = p_18_5_ & p_174_97_;
  assign new_n1603 = p_18_5_ & ~new_n1602;
  assign new_n1604 = ~new_n393 & ~new_n1603;
  assign new_n1605 = p_18_5_ & ~p_2253_183_;
  assign new_n1606 = ~p_18_5_ & p_109_54_;
  assign new_n1607 = ~new_n1605 & ~new_n1606;
  assign new_n1608 = ~new_n1604 & ~new_n1607;
  assign new_n1609 = new_n1604 & new_n1607;
  assign new_n1610 = ~new_n1608 & ~new_n1609;
  assign new_n1611 = p_176_99_ & p_18_5_;
  assign new_n1612 = p_18_5_ & ~new_n1611;
  assign new_n1613 = ~new_n393 & ~new_n1612;
  assign new_n1614 = p_18_5_ & ~p_2239_181_;
  assign new_n1615 = ~p_18_5_ & p_63_26_;
  assign new_n1616 = ~new_n1614 & ~new_n1615;
  assign new_n1617 = ~new_n1613 & ~new_n1616;
  assign new_n1618 = new_n1613 & new_n1616;
  assign new_n1619 = ~new_n1617 & ~new_n1618;
  assign new_n1620 = ~new_n1592 & ~new_n1601;
  assign new_n1621 = ~new_n1610 & new_n1620;
  assign new_n1622 = ~new_n1619 & new_n1621;
  assign new_n1623 = new_n1583 & new_n1622;
  assign new_n1624 = ~new_n1046 & new_n1054;
  assign new_n1625 = new_n983 & ~new_n1624;
  assign new_n1626 = new_n1537 & new_n1538;
  assign new_n1627 = new_n1623 & new_n1626;
  assign new_n1628 = ~new_n1625 & new_n1627;
  assign new_n1629 = new_n1027 & new_n1054;
  assign new_n1630 = new_n1537 & new_n1623;
  assign new_n1631 = new_n1629 & new_n1630;
  assign new_n1632 = new_n1538 & new_n1631;
  assign new_n1633 = p_89_48_ & new_n1632;
  assign new_n1634 = ~new_n1557 & ~new_n1560;
  assign new_n1635 = new_n1580 & new_n1634;
  assign new_n1636 = ~new_n1571 & new_n1635;
  assign new_n1637 = ~new_n1573 & ~new_n1576;
  assign new_n1638 = ~new_n1546 & new_n1637;
  assign new_n1639 = ~new_n1571 & new_n1638;
  assign new_n1640 = ~new_n1555 & new_n1639;
  assign new_n1641 = ~new_n1563 & new_n1640;
  assign new_n1642 = ~new_n1540 & ~new_n1543;
  assign new_n1643 = ~new_n1555 & new_n1642;
  assign new_n1644 = ~new_n1565 & ~new_n1568;
  assign new_n1645 = ~new_n1555 & new_n1644;
  assign new_n1646 = ~new_n1546 & new_n1645;
  assign new_n1647 = new_n1549 & ~new_n1552;
  assign new_n1648 = ~new_n1636 & ~new_n1641;
  assign new_n1649 = ~new_n1643 & new_n1648;
  assign new_n1650 = ~new_n1646 & new_n1649;
  assign new_n1651 = ~new_n1647 & new_n1650;
  assign new_n1652 = new_n1622 & ~new_n1651;
  assign new_n1653 = new_n1613 & ~new_n1616;
  assign new_n1654 = ~new_n1592 & ~new_n1610;
  assign new_n1655 = new_n1653 & new_n1654;
  assign new_n1656 = ~new_n1601 & new_n1655;
  assign new_n1657 = new_n1604 & ~new_n1607;
  assign new_n1658 = ~new_n1592 & new_n1657;
  assign new_n1659 = new_n1595 & ~new_n1598;
  assign new_n1660 = ~new_n1592 & new_n1659;
  assign new_n1661 = ~new_n1610 & new_n1660;
  assign new_n1662 = new_n1586 & ~new_n1589;
  assign new_n1663 = ~new_n1656 & ~new_n1658;
  assign new_n1664 = ~new_n1661 & new_n1663;
  assign new_n1665 = ~new_n1662 & new_n1664;
  assign new_n1666 = ~new_n1652 & new_n1665;
  assign new_n1667 = new_n1537 & ~new_n1666;
  assign new_n1668 = ~new_n1120 & new_n1128;
  assign new_n1669 = new_n941 & ~new_n1668;
  assign new_n1670 = new_n1630 & ~new_n1669;
  assign new_n1671 = new_n1502 & ~new_n1505;
  assign new_n1672 = new_n1524 & new_n1671;
  assign new_n1673 = ~new_n1517 & new_n1672;
  assign new_n1674 = ~new_n393 & ~new_n1520;
  assign new_n1675 = ~new_n1490 & new_n1674;
  assign new_n1676 = ~new_n1517 & new_n1675;
  assign new_n1677 = ~new_n1499 & new_n1676;
  assign new_n1678 = ~new_n1508 & new_n1677;
  assign new_n1679 = new_n1484 & ~new_n1487;
  assign new_n1680 = ~new_n1499 & new_n1679;
  assign new_n1681 = new_n1511 & ~new_n1514;
  assign new_n1682 = ~new_n1499 & new_n1681;
  assign new_n1683 = ~new_n1490 & new_n1682;
  assign new_n1684 = new_n1493 & ~new_n1496;
  assign new_n1685 = ~new_n1673 & ~new_n1678;
  assign new_n1686 = ~new_n1680 & new_n1685;
  assign new_n1687 = ~new_n1683 & new_n1686;
  assign new_n1688 = ~new_n1684 & new_n1687;
  assign new_n1689 = new_n1536 & ~new_n1688;
  assign new_n1690 = p_38_11_ & ~new_n1532;
  assign new_n1691 = ~new_n1531 & new_n1690;
  assign new_n1692 = p_38_11_ & ~new_n1528;
  assign new_n1693 = ~new_n1691 & ~new_n1692;
  assign new_n1694 = ~new_n1689 & new_n1693;
  assign new_n1695 = ~new_n1628 & ~new_n1633;
  assign new_n1696 = ~new_n1667 & new_n1695;
  assign new_n1697 = ~new_n1670 & new_n1696;
  assign p_264_3121_ = ~new_n1694 | ~new_n1697;
  assign new_n1699 = new_n533 & ~new_n729;
  assign new_n1700 = new_n620 & ~new_n1699;
  assign new_n1701 = new_n545 & ~new_n1700;
  assign new_n1702 = ~new_n545 & new_n1700;
  assign p_307_3389_ = new_n1701 | new_n1702;
  assign new_n1704 = new_n489 & new_n847;
  assign new_n1705 = ~new_n489 & ~new_n847;
  assign new_n1706 = ~new_n1704 & ~new_n1705;
  assign new_n1707 = new_n471 & ~new_n1476;
  assign new_n1708 = new_n655 & ~new_n1707;
  assign new_n1709 = new_n1706 & ~new_n1708;
  assign new_n1710 = new_n489 & new_n657;
  assign new_n1711 = ~new_n489 & ~new_n657;
  assign new_n1712 = ~new_n1710 & ~new_n1711;
  assign new_n1713 = new_n1708 & ~new_n1712;
  assign p_353_3425_ = new_n1709 | new_n1713;
  assign new_n1715 = ~new_n339 & ~new_n348;
  assign new_n1716 = ~new_n354 & new_n1715;
  assign new_n1717 = p_4526_205_ & new_n1716;
  assign new_n1718 = ~new_n354 & new_n366;
  assign new_n1719 = ~new_n354 & new_n370;
  assign new_n1720 = ~new_n339 & new_n1719;
  assign new_n1721 = ~new_n1717 & ~new_n1718;
  assign new_n1722 = ~new_n1720 & new_n1721;
  assign new_n1723 = ~new_n377 & new_n1722;
  assign new_n1724 = new_n360 & ~new_n1723;
  assign new_n1725 = ~new_n360 & new_n1723;
  assign p_391_3094_ = new_n1724 | new_n1725;
  assign new_n1727 = ~new_n1416 & ~new_n1417;
  assign new_n1728 = ~new_n628 & new_n1727;
  assign new_n1729 = new_n557 & ~new_n1728;
  assign new_n1730 = ~new_n557 & new_n1728;
  assign new_n1731 = ~new_n1729 & ~new_n1730;
  assign new_n1732 = ~new_n1700 & ~new_n1731;
  assign new_n1733 = new_n557 & new_n1418;
  assign new_n1734 = ~new_n557 & ~new_n1418;
  assign new_n1735 = ~new_n1733 & ~new_n1734;
  assign new_n1736 = new_n1700 & new_n1735;
  assign p_301_3388_ = new_n1732 | new_n1736;
  assign new_n1738 = ~new_n354 & ~new_n360;
  assign new_n1739 = new_n370 & new_n1738;
  assign new_n1740 = ~new_n339 & new_n1739;
  assign new_n1741 = ~new_n339 & ~new_n360;
  assign new_n1742 = ~new_n348 & new_n1741;
  assign new_n1743 = ~new_n354 & new_n1742;
  assign new_n1744 = p_4526_205_ & new_n1743;
  assign new_n1745 = ~new_n360 & new_n377;
  assign new_n1746 = ~new_n360 & new_n366;
  assign new_n1747 = ~new_n354 & new_n1746;
  assign new_n1748 = ~new_n1740 & ~new_n1744;
  assign new_n1749 = ~new_n1745 & new_n1748;
  assign new_n1750 = ~new_n1747 & new_n1749;
  assign new_n1751 = ~new_n375 & new_n1750;
  assign new_n1752 = new_n333 & ~new_n1751;
  assign new_n1753 = ~new_n333 & new_n1751;
  assign p_388_3093_ = new_n1752 | new_n1753;
  assign new_n1755 = ~new_n1140 & new_n1171;
  assign new_n1756 = ~new_n1172 & ~new_n1755;
  assign new_n1757 = ~new_n672 & new_n1756;
  assign new_n1758 = new_n417 & ~new_n1757;
  assign new_n1759 = ~new_n417 & new_n1757;
  assign p_333_3416_ = new_n1758 | new_n1759;
  assign new_n1761 = p_199_122_ & p_172_95_;
  assign new_n1762 = p_188_111_ & new_n1761;
  assign p_410_387_ = ~p_162_85_ | ~new_n1762;
  assign new_n1764 = ~new_n449 & ~new_n467;
  assign new_n1765 = ~new_n455 & new_n1764;
  assign new_n1766 = ~new_n461 & new_n1765;
  assign new_n1767 = ~new_n1476 & new_n1766;
  assign new_n1768 = ~new_n740 & ~new_n1767;
  assign new_n1769 = ~new_n744 & new_n1768;
  assign new_n1770 = ~new_n746 & new_n1769;
  assign new_n1771 = ~new_n646 & new_n1770;
  assign new_n1772 = new_n443 & ~new_n1771;
  assign new_n1773 = ~new_n443 & new_n1771;
  assign p_359_3426_ = new_n1772 | new_n1773;
  assign new_n1775 = ~new_n385 & new_n570;
  assign new_n1776 = new_n385 & ~new_n570;
  assign p_385_3151_ = new_n1775 | new_n1776;
  assign new_n1778 = p_4526_205_ & ~new_n348;
  assign new_n1779 = ~new_n370 & ~new_n1778;
  assign new_n1780 = new_n339 & ~new_n1779;
  assign new_n1781 = ~new_n339 & new_n1779;
  assign p_397_3097_ = new_n1780 | new_n1781;
  assign new_n1783 = new_n435 & ~new_n1142;
  assign new_n1784 = ~new_n435 & new_n1142;
  assign p_471_3445_ = new_n1783 | new_n1784;
  assign new_n1786 = p_133_66_ & p_134_67_;
  assign p_281_547_ = p_5_1_ | ~new_n1786;
  assign new_n1788 = ~new_n511 & ~new_n529;
  assign new_n1789 = ~new_n517 & new_n1788;
  assign new_n1790 = ~new_n523 & new_n1789;
  assign new_n1791 = ~new_n729 & new_n1790;
  assign new_n1792 = ~new_n1325 & ~new_n1791;
  assign new_n1793 = ~new_n1329 & new_n1792;
  assign new_n1794 = ~new_n1331 & new_n1793;
  assign new_n1795 = ~new_n611 & new_n1794;
  assign new_n1796 = new_n505 & ~new_n1795;
  assign new_n1797 = ~new_n505 & new_n1795;
  assign p_310_3393_ = new_n1796 | new_n1797;
  assign new_n1799 = new_n411 & ~new_n1140;
  assign new_n1800 = ~new_n411 & new_n1140;
  assign p_324_3363_ = new_n1799 | new_n1800;
  assign new_n1802 = ~new_n317 & new_n323;
  assign new_n1803 = new_n317 & ~new_n323;
  assign new_n1804 = ~new_n1802 & ~new_n1803;
  assign new_n1805 = ~new_n564 & new_n573;
  assign new_n1806 = new_n564 & ~new_n573;
  assign new_n1807 = ~new_n1805 & ~new_n1806;
  assign new_n1808 = new_n1804 & ~new_n1807;
  assign new_n1809 = ~new_n1804 & new_n1807;
  assign new_n1810 = ~new_n1808 & ~new_n1809;
  assign new_n1811 = ~p_18_5_ & p_44_13_;
  assign new_n1812 = p_18_5_ & p_239_162_;
  assign new_n1813 = ~new_n1811 & ~new_n1812;
  assign new_n1814 = ~new_n342 & new_n1813;
  assign new_n1815 = new_n342 & ~new_n1813;
  assign new_n1816 = ~new_n1814 & ~new_n1815;
  assign new_n1817 = ~new_n330 & new_n357;
  assign new_n1818 = new_n330 & ~new_n357;
  assign new_n1819 = ~new_n1817 & ~new_n1818;
  assign new_n1820 = new_n336 & ~new_n351;
  assign new_n1821 = ~new_n336 & new_n351;
  assign new_n1822 = ~new_n1820 & ~new_n1821;
  assign new_n1823 = ~new_n1816 & ~new_n1819;
  assign new_n1824 = ~new_n1822 & new_n1823;
  assign new_n1825 = new_n1819 & ~new_n1822;
  assign new_n1826 = new_n1816 & new_n1825;
  assign new_n1827 = ~new_n1824 & ~new_n1826;
  assign new_n1828 = new_n1816 & ~new_n1819;
  assign new_n1829 = new_n1822 & new_n1828;
  assign new_n1830 = new_n1819 & new_n1822;
  assign new_n1831 = ~new_n1816 & new_n1830;
  assign new_n1832 = ~new_n1829 & ~new_n1831;
  assign new_n1833 = new_n1827 & new_n1832;
  assign new_n1834 = new_n1810 & ~new_n1833;
  assign new_n1835 = ~new_n1810 & new_n1833;
  assign new_n1836 = ~new_n1834 & ~new_n1835;
  assign new_n1837 = ~new_n542 & new_n548;
  assign new_n1838 = new_n542 & ~new_n548;
  assign new_n1839 = ~new_n1837 & ~new_n1838;
  assign new_n1840 = new_n536 & ~new_n554;
  assign new_n1841 = ~new_n536 & new_n554;
  assign new_n1842 = ~new_n1840 & ~new_n1841;
  assign new_n1843 = new_n1839 & ~new_n1842;
  assign new_n1844 = ~new_n1839 & new_n1842;
  assign new_n1845 = ~new_n1843 & ~new_n1844;
  assign new_n1846 = p_18_5_ & p_161_84_;
  assign new_n1847 = ~p_18_5_ & p_141_70_;
  assign new_n1848 = ~new_n1846 & ~new_n1847;
  assign new_n1849 = ~new_n514 & new_n1848;
  assign new_n1850 = new_n514 & ~new_n1848;
  assign new_n1851 = ~new_n1849 & ~new_n1850;
  assign new_n1852 = new_n502 & new_n526;
  assign new_n1853 = ~new_n502 & ~new_n526;
  assign new_n1854 = ~new_n1852 & ~new_n1853;
  assign new_n1855 = new_n508 & ~new_n520;
  assign new_n1856 = ~new_n508 & new_n520;
  assign new_n1857 = ~new_n1855 & ~new_n1856;
  assign new_n1858 = ~new_n1851 & ~new_n1854;
  assign new_n1859 = ~new_n1857 & new_n1858;
  assign new_n1860 = new_n1854 & ~new_n1857;
  assign new_n1861 = new_n1851 & new_n1860;
  assign new_n1862 = ~new_n1859 & ~new_n1861;
  assign new_n1863 = new_n1851 & ~new_n1854;
  assign new_n1864 = new_n1857 & new_n1863;
  assign new_n1865 = new_n1854 & new_n1857;
  assign new_n1866 = ~new_n1851 & new_n1865;
  assign new_n1867 = ~new_n1864 & ~new_n1866;
  assign new_n1868 = new_n1862 & new_n1867;
  assign new_n1869 = new_n1845 & ~new_n1868;
  assign new_n1870 = ~new_n1845 & new_n1868;
  assign new_n1871 = ~new_n1869 & ~new_n1870;
  assign new_n1872 = new_n480 & ~new_n486;
  assign new_n1873 = ~new_n480 & new_n486;
  assign new_n1874 = ~new_n1872 & ~new_n1873;
  assign new_n1875 = ~new_n474 & new_n492;
  assign new_n1876 = new_n474 & ~new_n492;
  assign new_n1877 = ~new_n1875 & ~new_n1876;
  assign new_n1878 = new_n1874 & ~new_n1877;
  assign new_n1879 = ~new_n1874 & new_n1877;
  assign new_n1880 = ~new_n1878 & ~new_n1879;
  assign new_n1881 = p_115_60_ & ~p_18_5_;
  assign new_n1882 = p_18_5_ & p_227_150_;
  assign new_n1883 = ~new_n1881 & ~new_n1882;
  assign new_n1884 = ~new_n452 & new_n1883;
  assign new_n1885 = new_n452 & ~new_n1883;
  assign new_n1886 = ~new_n1884 & ~new_n1885;
  assign new_n1887 = ~new_n440 & new_n464;
  assign new_n1888 = new_n440 & ~new_n464;
  assign new_n1889 = ~new_n1887 & ~new_n1888;
  assign new_n1890 = new_n446 & ~new_n458;
  assign new_n1891 = ~new_n446 & new_n458;
  assign new_n1892 = ~new_n1890 & ~new_n1891;
  assign new_n1893 = ~new_n1886 & ~new_n1889;
  assign new_n1894 = ~new_n1892 & new_n1893;
  assign new_n1895 = new_n1889 & ~new_n1892;
  assign new_n1896 = new_n1886 & new_n1895;
  assign new_n1897 = ~new_n1894 & ~new_n1896;
  assign new_n1898 = new_n1886 & ~new_n1889;
  assign new_n1899 = new_n1892 & new_n1898;
  assign new_n1900 = new_n1889 & new_n1892;
  assign new_n1901 = ~new_n1886 & new_n1900;
  assign new_n1902 = ~new_n1899 & ~new_n1901;
  assign new_n1903 = new_n1897 & new_n1902;
  assign new_n1904 = new_n1880 & ~new_n1903;
  assign new_n1905 = ~new_n1880 & new_n1903;
  assign new_n1906 = ~new_n1904 & ~new_n1905;
  assign new_n1907 = p_212_135_ & p_18_5_;
  assign new_n1908 = p_18_5_ & ~new_n1907;
  assign new_n1909 = ~new_n393 & ~new_n1908;
  assign new_n1910 = p_18_5_ & p_211_134_;
  assign new_n1911 = p_18_5_ & ~new_n1910;
  assign new_n1912 = ~new_n393 & ~new_n1911;
  assign new_n1913 = ~new_n1909 & new_n1912;
  assign new_n1914 = new_n1909 & ~new_n1912;
  assign new_n1915 = ~new_n1913 & ~new_n1914;
  assign new_n1916 = ~new_n393 & new_n408;
  assign new_n1917 = new_n393 & ~new_n408;
  assign new_n1918 = ~new_n1916 & ~new_n1917;
  assign new_n1919 = new_n396 & ~new_n420;
  assign new_n1920 = ~new_n396 & new_n420;
  assign new_n1921 = ~new_n1919 & ~new_n1920;
  assign new_n1922 = ~new_n402 & new_n414;
  assign new_n1923 = new_n402 & ~new_n414;
  assign new_n1924 = ~new_n1922 & ~new_n1923;
  assign new_n1925 = ~new_n1918 & ~new_n1921;
  assign new_n1926 = ~new_n1924 & new_n1925;
  assign new_n1927 = new_n1921 & ~new_n1924;
  assign new_n1928 = new_n1918 & new_n1927;
  assign new_n1929 = ~new_n1926 & ~new_n1928;
  assign new_n1930 = new_n1918 & ~new_n1921;
  assign new_n1931 = new_n1924 & new_n1930;
  assign new_n1932 = new_n1921 & new_n1924;
  assign new_n1933 = ~new_n1918 & new_n1932;
  assign new_n1934 = ~new_n1931 & ~new_n1933;
  assign new_n1935 = new_n1929 & new_n1934;
  assign new_n1936 = new_n1915 & ~new_n1935;
  assign new_n1937 = ~new_n1915 & new_n1935;
  assign new_n1938 = ~new_n1936 & ~new_n1937;
  assign new_n1939 = ~new_n1836 & ~new_n1871;
  assign new_n1940 = ~new_n1906 & new_n1939;
  assign p_412_3369_ = new_n1938 | ~new_n1940;
  assign p_289_383_ = ~p_1197_165_ | p_5_1_;
  assign new_n1943 = ~new_n320 & new_n387;
  assign new_n1944 = ~new_n320 & ~new_n570;
  assign new_n1945 = ~new_n1943 & ~new_n1944;
  assign new_n1946 = ~new_n586 & new_n1945;
  assign new_n1947 = new_n576 & ~new_n1946;
  assign new_n1948 = ~new_n576 & new_n1946;
  assign new_n1949 = ~new_n1947 & ~new_n1948;
  assign new_n1950 = ~new_n385 & ~new_n1949;
  assign new_n1951 = ~new_n586 & ~new_n1943;
  assign new_n1952 = new_n576 & new_n1951;
  assign new_n1953 = ~new_n576 & ~new_n1951;
  assign new_n1954 = ~new_n1952 & ~new_n1953;
  assign new_n1955 = new_n385 & new_n1954;
  assign p_379_3207_ = new_n1950 | new_n1955;
  assign new_n1957 = p_182_105_ & p_186_109_;
  assign new_n1958 = p_185_108_ & new_n1957;
  assign p_408_385_ = ~p_183_106_ | ~new_n1958;
  assign new_n1960 = ~p_410_387_ & ~p_408_385_;
  assign new_n1961 = new_n962 & ~new_n968;
  assign new_n1962 = ~new_n962 & new_n968;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = new_n946 & ~new_n954;
  assign new_n1965 = ~new_n946 & new_n954;
  assign new_n1966 = ~new_n1964 & ~new_n1965;
  assign new_n1967 = new_n1963 & ~new_n1966;
  assign new_n1968 = ~new_n1963 & new_n1966;
  assign new_n1969 = ~new_n1967 & ~new_n1968;
  assign new_n1970 = ~p_18_5_ & p_69_30_;
  assign new_n1971 = ~p_3698_185_ & p_18_5_;
  assign new_n1972 = ~new_n1970 & ~new_n1971;
  assign new_n1973 = p_18_5_ & ~p_3701_186_;
  assign new_n1974 = ~new_n1019 & ~new_n1973;
  assign new_n1975 = new_n1972 & ~new_n1974;
  assign new_n1976 = ~new_n1972 & new_n1974;
  assign new_n1977 = ~new_n1975 & ~new_n1976;
  assign new_n1978 = new_n988 & ~new_n996;
  assign new_n1979 = ~new_n988 & new_n996;
  assign new_n1980 = ~new_n1978 & ~new_n1979;
  assign new_n1981 = new_n1004 & ~new_n1012;
  assign new_n1982 = ~new_n1004 & new_n1012;
  assign new_n1983 = ~new_n1981 & ~new_n1982;
  assign new_n1984 = ~new_n1977 & ~new_n1980;
  assign new_n1985 = ~new_n1983 & new_n1984;
  assign new_n1986 = new_n1980 & ~new_n1983;
  assign new_n1987 = new_n1977 & new_n1986;
  assign new_n1988 = ~new_n1985 & ~new_n1987;
  assign new_n1989 = new_n1977 & ~new_n1980;
  assign new_n1990 = new_n1983 & new_n1989;
  assign new_n1991 = new_n1980 & new_n1983;
  assign new_n1992 = ~new_n1977 & new_n1991;
  assign new_n1993 = ~new_n1990 & ~new_n1992;
  assign new_n1994 = new_n1988 & new_n1993;
  assign new_n1995 = new_n1969 & ~new_n1994;
  assign new_n1996 = ~new_n1969 & new_n1994;
  assign new_n1997 = ~new_n1995 & ~new_n1996;
  assign new_n1998 = ~new_n1598 & new_n1616;
  assign new_n1999 = new_n1598 & ~new_n1616;
  assign new_n2000 = ~new_n1998 & ~new_n1999;
  assign new_n2001 = ~new_n1589 & new_n1607;
  assign new_n2002 = new_n1589 & ~new_n1607;
  assign new_n2003 = ~new_n2001 & ~new_n2002;
  assign new_n2004 = new_n2000 & ~new_n2003;
  assign new_n2005 = ~new_n2000 & new_n2003;
  assign new_n2006 = ~new_n2004 & ~new_n2005;
  assign new_n2007 = ~p_2208_175_ & p_18_5_;
  assign new_n2008 = ~p_18_5_ & p_82_41_;
  assign new_n2009 = ~new_n2007 & ~new_n2008;
  assign new_n2010 = ~new_n1576 & new_n2009;
  assign new_n2011 = new_n1576 & ~new_n2009;
  assign new_n2012 = ~new_n2010 & ~new_n2011;
  assign new_n2013 = new_n1543 & ~new_n1552;
  assign new_n2014 = ~new_n1543 & new_n1552;
  assign new_n2015 = ~new_n2013 & ~new_n2014;
  assign new_n2016 = new_n1560 & ~new_n1568;
  assign new_n2017 = ~new_n1560 & new_n1568;
  assign new_n2018 = ~new_n2016 & ~new_n2017;
  assign new_n2019 = ~new_n2012 & ~new_n2015;
  assign new_n2020 = ~new_n2018 & new_n2019;
  assign new_n2021 = new_n2015 & ~new_n2018;
  assign new_n2022 = new_n2012 & new_n2021;
  assign new_n2023 = ~new_n2020 & ~new_n2022;
  assign new_n2024 = new_n2012 & ~new_n2015;
  assign new_n2025 = new_n2018 & new_n2024;
  assign new_n2026 = new_n2015 & new_n2018;
  assign new_n2027 = ~new_n2012 & new_n2026;
  assign new_n2028 = ~new_n2025 & ~new_n2027;
  assign new_n2029 = new_n2023 & new_n2028;
  assign new_n2030 = new_n2006 & ~new_n2029;
  assign new_n2031 = ~new_n2006 & new_n2029;
  assign new_n2032 = ~new_n2030 & ~new_n2031;
  assign new_n2033 = new_n920 & ~new_n926;
  assign new_n2034 = ~new_n920 & new_n926;
  assign new_n2035 = ~new_n2033 & ~new_n2034;
  assign new_n2036 = new_n904 & ~new_n912;
  assign new_n2037 = ~new_n904 & new_n912;
  assign new_n2038 = ~new_n2036 & ~new_n2037;
  assign new_n2039 = new_n2035 & ~new_n2038;
  assign new_n2040 = ~new_n2035 & new_n2038;
  assign new_n2041 = ~new_n2039 & ~new_n2040;
  assign new_n2042 = ~p_18_5_ & p_58_21_;
  assign new_n2043 = ~p_4393_195_ & p_18_5_;
  assign new_n2044 = ~new_n2042 & ~new_n2043;
  assign new_n2045 = ~new_n1094 & new_n2044;
  assign new_n2046 = new_n1094 & ~new_n2044;
  assign new_n2047 = ~new_n2045 & ~new_n2046;
  assign new_n2048 = new_n1062 & ~new_n1070;
  assign new_n2049 = ~new_n1062 & new_n1070;
  assign new_n2050 = ~new_n2048 & ~new_n2049;
  assign new_n2051 = new_n1078 & ~new_n1086;
  assign new_n2052 = ~new_n1078 & new_n1086;
  assign new_n2053 = ~new_n2051 & ~new_n2052;
  assign new_n2054 = ~new_n2047 & ~new_n2050;
  assign new_n2055 = ~new_n2053 & new_n2054;
  assign new_n2056 = new_n2050 & ~new_n2053;
  assign new_n2057 = new_n2047 & new_n2056;
  assign new_n2058 = ~new_n2055 & ~new_n2057;
  assign new_n2059 = new_n2047 & ~new_n2050;
  assign new_n2060 = new_n2053 & new_n2059;
  assign new_n2061 = new_n2050 & new_n2053;
  assign new_n2062 = ~new_n2047 & new_n2061;
  assign new_n2063 = ~new_n2060 & ~new_n2062;
  assign new_n2064 = new_n2058 & new_n2063;
  assign new_n2065 = new_n2041 & ~new_n2064;
  assign new_n2066 = ~new_n2041 & new_n2064;
  assign new_n2067 = ~new_n2065 & ~new_n2066;
  assign new_n2068 = ~p_1492_172_ & p_18_5_;
  assign new_n2069 = ~p_18_5_ & p_1455_166_;
  assign new_n2070 = ~new_n2068 & ~new_n2069;
  assign new_n2071 = ~p_1496_173_ & p_18_5_;
  assign new_n2072 = p_2204_174_ & ~p_18_5_;
  assign new_n2073 = ~new_n2071 & ~new_n2072;
  assign new_n2074 = new_n2070 & ~new_n2073;
  assign new_n2075 = ~new_n2070 & new_n2073;
  assign new_n2076 = ~new_n2074 & ~new_n2075;
  assign new_n2077 = p_18_5_ & ~p_1459_167_;
  assign new_n2078 = p_114_59_ & ~p_18_5_;
  assign new_n2079 = ~new_n2077 & ~new_n2078;
  assign new_n2080 = ~new_n1520 & new_n2079;
  assign new_n2081 = new_n1520 & ~new_n2079;
  assign new_n2082 = ~new_n2080 & ~new_n2081;
  assign new_n2083 = new_n1487 & ~new_n1496;
  assign new_n2084 = ~new_n1487 & new_n1496;
  assign new_n2085 = ~new_n2083 & ~new_n2084;
  assign new_n2086 = new_n1505 & ~new_n1514;
  assign new_n2087 = ~new_n1505 & new_n1514;
  assign new_n2088 = ~new_n2086 & ~new_n2087;
  assign new_n2089 = ~new_n2082 & ~new_n2085;
  assign new_n2090 = ~new_n2088 & new_n2089;
  assign new_n2091 = new_n2085 & ~new_n2088;
  assign new_n2092 = new_n2082 & new_n2091;
  assign new_n2093 = ~new_n2090 & ~new_n2092;
  assign new_n2094 = new_n2082 & ~new_n2085;
  assign new_n2095 = new_n2088 & new_n2094;
  assign new_n2096 = new_n2085 & new_n2088;
  assign new_n2097 = ~new_n2082 & new_n2096;
  assign new_n2098 = ~new_n2095 & ~new_n2097;
  assign new_n2099 = new_n2093 & new_n2098;
  assign new_n2100 = new_n2076 & ~new_n2099;
  assign new_n2101 = ~new_n2076 & new_n2099;
  assign new_n2102 = ~new_n2100 & ~new_n2101;
  assign new_n2103 = ~new_n1997 & ~new_n2032;
  assign new_n2104 = ~new_n2067 & new_n2103;
  assign p_414_3338_ = new_n2102 | ~new_n2104;
  assign new_n2106 = new_n959 & ~new_n965;
  assign new_n2107 = ~new_n959 & new_n965;
  assign new_n2108 = ~new_n2106 & ~new_n2107;
  assign new_n2109 = new_n943 & ~new_n951;
  assign new_n2110 = ~new_n943 & new_n951;
  assign new_n2111 = ~new_n2109 & ~new_n2110;
  assign new_n2112 = new_n2108 & ~new_n2111;
  assign new_n2113 = ~new_n2108 & new_n2111;
  assign new_n2114 = ~new_n2112 & ~new_n2113;
  assign new_n2115 = p_18_5_ & p_208_131_;
  assign new_n2116 = ~new_n1811 & ~new_n2115;
  assign new_n2117 = ~new_n1017 & new_n2116;
  assign new_n2118 = new_n1017 & ~new_n2116;
  assign new_n2119 = ~new_n2117 & ~new_n2118;
  assign new_n2120 = new_n985 & ~new_n993;
  assign new_n2121 = ~new_n985 & new_n993;
  assign new_n2122 = ~new_n2120 & ~new_n2121;
  assign new_n2123 = new_n1001 & ~new_n1009;
  assign new_n2124 = ~new_n1001 & new_n1009;
  assign new_n2125 = ~new_n2123 & ~new_n2124;
  assign new_n2126 = ~new_n2119 & ~new_n2122;
  assign new_n2127 = ~new_n2125 & new_n2126;
  assign new_n2128 = new_n2122 & ~new_n2125;
  assign new_n2129 = new_n2119 & new_n2128;
  assign new_n2130 = ~new_n2127 & ~new_n2129;
  assign new_n2131 = new_n2119 & ~new_n2122;
  assign new_n2132 = new_n2125 & new_n2131;
  assign new_n2133 = new_n2122 & new_n2125;
  assign new_n2134 = ~new_n2119 & new_n2133;
  assign new_n2135 = ~new_n2132 & ~new_n2134;
  assign new_n2136 = new_n2130 & new_n2135;
  assign new_n2137 = new_n2114 & ~new_n2136;
  assign new_n2138 = ~new_n2114 & new_n2136;
  assign new_n2139 = ~new_n2137 & ~new_n2138;
  assign new_n2140 = new_n1595 & ~new_n1613;
  assign new_n2141 = ~new_n1595 & new_n1613;
  assign new_n2142 = ~new_n2140 & ~new_n2141;
  assign new_n2143 = new_n1586 & ~new_n1604;
  assign new_n2144 = ~new_n1586 & new_n1604;
  assign new_n2145 = ~new_n2143 & ~new_n2144;
  assign new_n2146 = new_n2142 & ~new_n2145;
  assign new_n2147 = ~new_n2142 & new_n2145;
  assign new_n2148 = ~new_n2146 & ~new_n2147;
  assign new_n2149 = p_18_5_ & p_181_104_;
  assign new_n2150 = ~new_n1847 & ~new_n2149;
  assign new_n2151 = ~new_n1573 & new_n2150;
  assign new_n2152 = new_n1573 & ~new_n2150;
  assign new_n2153 = ~new_n2151 & ~new_n2152;
  assign new_n2154 = new_n1540 & new_n1549;
  assign new_n2155 = ~new_n1540 & ~new_n1549;
  assign new_n2156 = ~new_n2154 & ~new_n2155;
  assign new_n2157 = new_n1557 & ~new_n1565;
  assign new_n2158 = ~new_n1557 & new_n1565;
  assign new_n2159 = ~new_n2157 & ~new_n2158;
  assign new_n2160 = ~new_n2153 & ~new_n2156;
  assign new_n2161 = ~new_n2159 & new_n2160;
  assign new_n2162 = new_n2156 & ~new_n2159;
  assign new_n2163 = new_n2153 & new_n2162;
  assign new_n2164 = ~new_n2161 & ~new_n2163;
  assign new_n2165 = new_n2153 & ~new_n2156;
  assign new_n2166 = new_n2159 & new_n2165;
  assign new_n2167 = new_n2156 & new_n2159;
  assign new_n2168 = ~new_n2153 & new_n2167;
  assign new_n2169 = ~new_n2166 & ~new_n2168;
  assign new_n2170 = new_n2164 & new_n2169;
  assign new_n2171 = new_n2148 & ~new_n2170;
  assign new_n2172 = ~new_n2148 & new_n2170;
  assign new_n2173 = ~new_n2171 & ~new_n2172;
  assign new_n2174 = new_n917 & ~new_n923;
  assign new_n2175 = ~new_n917 & new_n923;
  assign new_n2176 = ~new_n2174 & ~new_n2175;
  assign new_n2177 = new_n901 & ~new_n909;
  assign new_n2178 = ~new_n901 & new_n909;
  assign new_n2179 = ~new_n2177 & ~new_n2178;
  assign new_n2180 = new_n2176 & ~new_n2179;
  assign new_n2181 = ~new_n2176 & new_n2179;
  assign new_n2182 = ~new_n2180 & ~new_n2181;
  assign new_n2183 = p_197_120_ & p_18_5_;
  assign new_n2184 = ~new_n1881 & ~new_n2183;
  assign new_n2185 = ~new_n1091 & new_n2184;
  assign new_n2186 = new_n1091 & ~new_n2184;
  assign new_n2187 = ~new_n2185 & ~new_n2186;
  assign new_n2188 = new_n1059 & ~new_n1067;
  assign new_n2189 = ~new_n1059 & new_n1067;
  assign new_n2190 = ~new_n2188 & ~new_n2189;
  assign new_n2191 = new_n1075 & ~new_n1083;
  assign new_n2192 = ~new_n1075 & new_n1083;
  assign new_n2193 = ~new_n2191 & ~new_n2192;
  assign new_n2194 = ~new_n2187 & ~new_n2190;
  assign new_n2195 = ~new_n2193 & new_n2194;
  assign new_n2196 = new_n2190 & ~new_n2193;
  assign new_n2197 = new_n2187 & new_n2196;
  assign new_n2198 = ~new_n2195 & ~new_n2197;
  assign new_n2199 = new_n2187 & ~new_n2190;
  assign new_n2200 = new_n2193 & new_n2199;
  assign new_n2201 = new_n2190 & new_n2193;
  assign new_n2202 = ~new_n2187 & new_n2201;
  assign new_n2203 = ~new_n2200 & ~new_n2202;
  assign new_n2204 = new_n2198 & new_n2203;
  assign new_n2205 = new_n2182 & ~new_n2204;
  assign new_n2206 = ~new_n2182 & new_n2204;
  assign new_n2207 = ~new_n2205 & ~new_n2206;
  assign new_n2208 = p_18_5_ & p_165_88_;
  assign new_n2209 = p_18_5_ & ~new_n2208;
  assign new_n2210 = ~new_n393 & ~new_n2209;
  assign new_n2211 = p_18_5_ & p_164_87_;
  assign new_n2212 = p_18_5_ & ~new_n2211;
  assign new_n2213 = ~new_n393 & ~new_n2212;
  assign new_n2214 = ~new_n2210 & new_n2213;
  assign new_n2215 = new_n2210 & ~new_n2213;
  assign new_n2216 = ~new_n2214 & ~new_n2215;
  assign new_n2217 = p_18_5_ & p_170_93_;
  assign new_n2218 = p_18_5_ & ~new_n2217;
  assign new_n2219 = ~new_n393 & ~new_n2218;
  assign new_n2220 = ~new_n393 & new_n2219;
  assign new_n2221 = new_n393 & ~new_n2219;
  assign new_n2222 = ~new_n2220 & ~new_n2221;
  assign new_n2223 = ~new_n1484 & new_n1493;
  assign new_n2224 = new_n1484 & ~new_n1493;
  assign new_n2225 = ~new_n2223 & ~new_n2224;
  assign new_n2226 = ~new_n1502 & new_n1511;
  assign new_n2227 = new_n1502 & ~new_n1511;
  assign new_n2228 = ~new_n2226 & ~new_n2227;
  assign new_n2229 = ~new_n2222 & ~new_n2225;
  assign new_n2230 = ~new_n2228 & new_n2229;
  assign new_n2231 = new_n2225 & ~new_n2228;
  assign new_n2232 = new_n2222 & new_n2231;
  assign new_n2233 = ~new_n2230 & ~new_n2232;
  assign new_n2234 = new_n2222 & ~new_n2225;
  assign new_n2235 = new_n2228 & new_n2234;
  assign new_n2236 = new_n2225 & new_n2228;
  assign new_n2237 = ~new_n2222 & new_n2236;
  assign new_n2238 = ~new_n2235 & ~new_n2237;
  assign new_n2239 = new_n2233 & new_n2238;
  assign new_n2240 = new_n2216 & ~new_n2239;
  assign new_n2241 = ~new_n2216 & new_n2239;
  assign new_n2242 = ~new_n2240 & ~new_n2241;
  assign new_n2243 = ~new_n2139 & ~new_n2173;
  assign new_n2244 = ~new_n2207 & new_n2243;
  assign p_416_3368_ = new_n2242 | ~new_n2244;
  assign new_n2246 = ~p_414_3338_ & ~p_416_3368_;
  assign new_n2247 = ~p_412_3369_ & new_n2246;
  assign new_n2248 = p_240_163_ & p_184_107_;
  assign new_n2249 = p_228_151_ & new_n2248;
  assign p_404_390_ = ~p_150_73_ | ~new_n2249;
  assign new_n2251 = ~p_406_388_ & ~p_404_390_;
  assign new_n2252 = new_n1960 & new_n2247;
  assign p_418_3449_ = ~new_n2251 | ~new_n2252;
  assign new_n2254 = ~new_n523 & new_n730;
  assign new_n2255 = ~new_n729 & new_n2254;
  assign new_n2256 = ~new_n1339 & ~new_n2255;
  assign new_n2257 = ~new_n1341 & new_n2256;
  assign new_n2258 = ~new_n613 & new_n2257;
  assign new_n2259 = new_n529 & ~new_n2258;
  assign new_n2260 = ~new_n529 & new_n2258;
  assign p_313_3396_ = new_n2259 | new_n2260;
  assign new_n2262 = ~new_n517 & ~new_n729;
  assign new_n2263 = ~new_n606 & ~new_n2262;
  assign new_n2264 = new_n511 & ~new_n2263;
  assign new_n2265 = ~new_n511 & new_n2263;
  assign p_319_3398_ = new_n2264 | new_n2265;
  assign new_n2267 = new_n436 & new_n1268;
  assign new_n2268 = new_n1218 & new_n2267;
  assign new_n2269 = new_n1213 & new_n2268;
  assign new_n2270 = ~new_n1226 & new_n2269;
  assign new_n2271 = new_n1213 & new_n2267;
  assign new_n2272 = new_n1214 & new_n2271;
  assign new_n2273 = new_n1218 & new_n2272;
  assign new_n2274 = p_4526_205_ & new_n2273;
  assign new_n2275 = ~new_n1230 & new_n2267;
  assign new_n2276 = ~new_n1223 & new_n2271;
  assign new_n2277 = ~new_n2270 & ~new_n2274;
  assign new_n2278 = ~new_n2275 & new_n2277;
  assign new_n2279 = ~new_n2276 & new_n2278;
  assign p_270_3109_ = ~new_n696 | ~new_n2279;
  assign new_n2281 = ~new_n1233 & new_n1268;
  assign new_n2282 = new_n690 & ~new_n2281;
  assign new_n2283 = ~new_n695 & new_n2282;
  assign new_n2284 = ~new_n1143 & ~new_n2282;
  assign p_276_3401_ = new_n2283 | new_n2284;
  assign new_n2286 = new_n551 & new_n1420;
  assign new_n2287 = ~new_n551 & ~new_n1420;
  assign new_n2288 = ~new_n2286 & ~new_n2287;
  assign new_n2289 = ~new_n1700 & new_n2288;
  assign new_n2290 = new_n551 & new_n622;
  assign new_n2291 = ~new_n551 & ~new_n622;
  assign new_n2292 = ~new_n2290 & ~new_n2291;
  assign new_n2293 = new_n1700 & ~new_n2292;
  assign p_304_3390_ = new_n2289 | new_n2293;
  assign new_n2295 = ~new_n411 & ~new_n1140;
  assign new_n2296 = ~new_n676 & ~new_n2295;
  assign new_n2297 = new_n405 & ~new_n2296;
  assign new_n2298 = ~new_n405 & new_n2296;
  assign p_336_3412_ = new_n2297 | new_n2298;
  assign new_n2300 = new_n751 & ~new_n1476;
  assign new_n2301 = ~new_n752 & ~new_n2300;
  assign new_n2302 = ~new_n637 & new_n2301;
  assign new_n2303 = new_n461 & ~new_n2302;
  assign new_n2304 = ~new_n461 & new_n2302;
  assign p_365_3430_ = new_n2303 | new_n2304;
  assign new_n2306 = ~new_n417 & new_n1171;
  assign new_n2307 = ~new_n1140 & new_n2306;
  assign new_n2308 = ~new_n1176 & ~new_n2307;
  assign new_n2309 = ~new_n1178 & new_n2308;
  assign new_n2310 = ~new_n683 & new_n2309;
  assign new_n2311 = new_n423 & ~new_n2310;
  assign new_n2312 = ~new_n423 & new_n2310;
  assign p_330_3411_ = new_n2311 | new_n2312;
  assign new_n2314 = new_n455 & ~new_n1476;
  assign new_n2315 = ~new_n455 & new_n1476;
  assign p_344_3382_ = new_n2314 | new_n2315;
  assign new_n2317 = new_n477 & ~new_n842;
  assign new_n2318 = ~new_n477 & new_n842;
  assign new_n2319 = ~new_n2317 & ~new_n2318;
  assign new_n2320 = ~new_n1708 & ~new_n2319;
  assign new_n2321 = new_n657 & new_n835;
  assign new_n2322 = ~new_n837 & ~new_n2321;
  assign new_n2323 = ~new_n661 & new_n2322;
  assign new_n2324 = new_n477 & new_n2323;
  assign new_n2325 = ~new_n477 & ~new_n2323;
  assign new_n2326 = ~new_n2324 & ~new_n2325;
  assign new_n2327 = new_n1708 & new_n2326;
  assign p_347_3420_ = new_n2320 | new_n2327;
  assign new_n2329 = ~new_n339 & ~new_n354;
  assign new_n2330 = ~new_n360 & new_n2329;
  assign new_n2331 = ~new_n348 & new_n2330;
  assign new_n2332 = ~new_n1740 & ~new_n2331;
  assign new_n2333 = ~new_n1745 & new_n2332;
  assign new_n2334 = ~new_n1747 & new_n2333;
  assign new_n2335 = ~new_n375 & new_n2334;
  assign new_n2336 = ~new_n339 & new_n370;
  assign new_n2337 = ~new_n366 & ~new_n2336;
  assign new_n2338 = ~new_n1715 & new_n2337;
  assign new_n2339 = ~new_n348 & new_n2329;
  assign new_n2340 = ~new_n1718 & ~new_n2339;
  assign new_n2341 = ~new_n1720 & new_n2340;
  assign new_n2342 = ~new_n377 & new_n2341;
  assign new_n2343 = ~new_n343 & new_n345;
  assign new_n2344 = new_n2342 & new_n2343;
  assign new_n2345 = ~new_n2342 & ~new_n2343;
  assign new_n2346 = ~new_n2344 & ~new_n2345;
  assign new_n2347 = new_n2338 & ~new_n2346;
  assign new_n2348 = ~new_n2338 & new_n2346;
  assign new_n2349 = ~new_n2347 & ~new_n2348;
  assign new_n2350 = new_n2335 & ~new_n2349;
  assign new_n2351 = ~new_n2335 & new_n2349;
  assign new_n2352 = ~new_n2350 & ~new_n2351;
  assign new_n2353 = new_n348 & ~new_n2352;
  assign new_n2354 = ~new_n348 & new_n2352;
  assign new_n2355 = ~new_n2353 & ~new_n2354;
  assign new_n2356 = new_n339 & ~new_n2355;
  assign new_n2357 = ~new_n339 & new_n2355;
  assign new_n2358 = ~new_n2356 & ~new_n2357;
  assign new_n2359 = new_n333 & ~new_n2358;
  assign new_n2360 = ~new_n333 & new_n2358;
  assign new_n2361 = ~new_n2359 & ~new_n2360;
  assign new_n2362 = new_n354 & ~new_n2361;
  assign new_n2363 = ~new_n354 & new_n2361;
  assign new_n2364 = ~new_n2362 & ~new_n2363;
  assign new_n2365 = new_n360 & ~new_n2364;
  assign new_n2366 = ~new_n360 & new_n2364;
  assign new_n2367 = ~new_n2365 & ~new_n2366;
  assign new_n2368 = p_4526_205_ & ~new_n2367;
  assign new_n2369 = ~new_n1740 & ~new_n1745;
  assign new_n2370 = ~new_n1747 & new_n2369;
  assign new_n2371 = ~new_n375 & new_n2370;
  assign new_n2372 = ~new_n1718 & ~new_n1720;
  assign new_n2373 = ~new_n377 & new_n2372;
  assign new_n2374 = new_n370 & ~new_n2373;
  assign new_n2375 = ~new_n370 & new_n2373;
  assign new_n2376 = ~new_n2374 & ~new_n2375;
  assign new_n2377 = ~new_n2337 & ~new_n2376;
  assign new_n2378 = new_n2337 & new_n2376;
  assign new_n2379 = ~new_n2377 & ~new_n2378;
  assign new_n2380 = ~new_n2371 & ~new_n2379;
  assign new_n2381 = new_n2371 & new_n2379;
  assign new_n2382 = ~new_n2380 & ~new_n2381;
  assign new_n2383 = new_n348 & ~new_n2382;
  assign new_n2384 = ~new_n348 & new_n2382;
  assign new_n2385 = ~new_n2383 & ~new_n2384;
  assign new_n2386 = new_n339 & ~new_n2385;
  assign new_n2387 = ~new_n339 & new_n2385;
  assign new_n2388 = ~new_n2386 & ~new_n2387;
  assign new_n2389 = new_n333 & ~new_n2388;
  assign new_n2390 = ~new_n333 & new_n2388;
  assign new_n2391 = ~new_n2389 & ~new_n2390;
  assign new_n2392 = new_n354 & ~new_n2391;
  assign new_n2393 = ~new_n354 & new_n2391;
  assign new_n2394 = ~new_n2392 & ~new_n2393;
  assign new_n2395 = new_n360 & ~new_n2394;
  assign new_n2396 = ~new_n360 & new_n2394;
  assign new_n2397 = ~new_n2395 & ~new_n2396;
  assign new_n2398 = ~p_4526_205_ & new_n2397;
  assign new_n2399 = ~new_n2368 & ~new_n2398;
  assign new_n2400 = new_n384 & ~new_n789;
  assign new_n2401 = ~new_n1944 & new_n1951;
  assign new_n2402 = new_n324 & new_n2401;
  assign new_n2403 = ~new_n324 & ~new_n2401;
  assign new_n2404 = ~new_n2402 & ~new_n2403;
  assign new_n2405 = new_n711 & ~new_n2404;
  assign new_n2406 = ~new_n711 & new_n2404;
  assign new_n2407 = ~new_n2405 & ~new_n2406;
  assign new_n2408 = new_n570 & ~new_n2407;
  assign new_n2409 = ~new_n570 & new_n2407;
  assign new_n2410 = ~new_n2408 & ~new_n2409;
  assign new_n2411 = new_n320 & ~new_n2410;
  assign new_n2412 = ~new_n320 & new_n2410;
  assign new_n2413 = ~new_n2411 & ~new_n2412;
  assign new_n2414 = new_n567 & ~new_n2413;
  assign new_n2415 = ~new_n567 & new_n2413;
  assign new_n2416 = ~new_n2414 & ~new_n2415;
  assign new_n2417 = new_n576 & ~new_n2416;
  assign new_n2418 = ~new_n576 & new_n2416;
  assign new_n2419 = ~new_n2417 & ~new_n2418;
  assign new_n2420 = p_4526_205_ & ~new_n2400;
  assign new_n2421 = ~new_n2419 & new_n2420;
  assign new_n2422 = ~p_4526_205_ & ~new_n384;
  assign new_n2423 = ~new_n2419 & new_n2422;
  assign new_n2424 = ~new_n706 & ~new_n708;
  assign new_n2425 = ~new_n584 & new_n2424;
  assign new_n2426 = new_n387 & ~new_n1951;
  assign new_n2427 = ~new_n387 & new_n1951;
  assign new_n2428 = ~new_n2426 & ~new_n2427;
  assign new_n2429 = ~new_n2425 & ~new_n2428;
  assign new_n2430 = new_n2425 & new_n2428;
  assign new_n2431 = ~new_n2429 & ~new_n2430;
  assign new_n2432 = new_n570 & ~new_n2431;
  assign new_n2433 = ~new_n570 & new_n2431;
  assign new_n2434 = ~new_n2432 & ~new_n2433;
  assign new_n2435 = new_n320 & ~new_n2434;
  assign new_n2436 = ~new_n320 & new_n2434;
  assign new_n2437 = ~new_n2435 & ~new_n2436;
  assign new_n2438 = new_n567 & ~new_n2437;
  assign new_n2439 = ~new_n567 & new_n2437;
  assign new_n2440 = ~new_n2438 & ~new_n2439;
  assign new_n2441 = new_n576 & ~new_n2440;
  assign new_n2442 = ~new_n576 & new_n2440;
  assign new_n2443 = ~new_n2441 & ~new_n2442;
  assign new_n2444 = p_4526_205_ & new_n2400;
  assign new_n2445 = ~new_n2443 & new_n2444;
  assign new_n2446 = ~p_4526_205_ & new_n384;
  assign new_n2447 = ~new_n2443 & new_n2446;
  assign new_n2448 = ~new_n2421 & ~new_n2423;
  assign new_n2449 = ~new_n2445 & new_n2448;
  assign new_n2450 = ~new_n2447 & new_n2449;
  assign new_n2451 = new_n2399 & ~new_n2450;
  assign new_n2452 = ~new_n2399 & new_n2450;
  assign p_399_3717_ = ~new_n2451 & ~new_n2452;
  assign new_n2454 = ~new_n461 & new_n751;
  assign new_n2455 = ~new_n1476 & new_n2454;
  assign new_n2456 = ~new_n756 & ~new_n2455;
  assign new_n2457 = ~new_n758 & new_n2456;
  assign new_n2458 = ~new_n648 & new_n2457;
  assign new_n2459 = new_n467 & ~new_n2458;
  assign new_n2460 = ~new_n467 & new_n2458;
  assign p_362_3429_ = new_n2459 | new_n2460;
  assign new_n2462 = p_4526_205_ & new_n1715;
  assign new_n2463 = ~new_n2336 & ~new_n2462;
  assign new_n2464 = ~new_n366 & new_n2463;
  assign new_n2465 = new_n354 & ~new_n2464;
  assign new_n2466 = ~new_n354 & new_n2464;
  assign p_394_3095_ = new_n2465 | new_n2466;
  assign p_402_395_ = p_5_1_ | p_57_20_;
  assign new_n2469 = ~new_n843 & ~new_n844;
  assign new_n2470 = ~new_n663 & new_n2469;
  assign new_n2471 = new_n495 & ~new_n2470;
  assign new_n2472 = ~new_n495 & new_n2470;
  assign new_n2473 = ~new_n2471 & ~new_n2472;
  assign new_n2474 = ~new_n1708 & ~new_n2473;
  assign new_n2475 = new_n495 & new_n845;
  assign new_n2476 = ~new_n495 & ~new_n845;
  assign new_n2477 = ~new_n2475 & ~new_n2476;
  assign new_n2478 = new_n1708 & new_n2477;
  assign p_350_3421_ = new_n2474 | new_n2478;
  assign new_n2480 = new_n1623 & new_n1629;
  assign new_n2481 = new_n1538 & new_n2480;
  assign new_n2482 = p_89_48_ & new_n2481;
  assign new_n2483 = new_n1623 & ~new_n1669;
  assign new_n2484 = new_n1538 & new_n1623;
  assign new_n2485 = ~new_n1625 & new_n2484;
  assign new_n2486 = ~new_n2482 & ~new_n2483;
  assign new_n2487 = ~new_n2485 & new_n2486;
  assign new_n2488 = new_n1666 & new_n2487;
  assign new_n2489 = new_n1527 & ~new_n2488;
  assign new_n2490 = new_n1688 & ~new_n2489;
  assign new_n2491 = ~new_n1693 & new_n2490;
  assign new_n2492 = ~new_n1536 & new_n1693;
  assign new_n2493 = ~new_n2490 & ~new_n2492;
  assign p_249_3418_ = new_n2491 | new_n2493;
  assign new_n2495 = new_n539 & ~new_n1415;
  assign new_n2496 = ~new_n539 & new_n1415;
  assign new_n2497 = ~new_n2495 & ~new_n2496;
  assign new_n2498 = ~new_n1700 & ~new_n2497;
  assign new_n2499 = new_n622 & new_n1408;
  assign new_n2500 = ~new_n1410 & ~new_n2499;
  assign new_n2501 = ~new_n626 & new_n2500;
  assign new_n2502 = new_n539 & new_n2501;
  assign new_n2503 = ~new_n539 & ~new_n2501;
  assign new_n2504 = ~new_n2502 & ~new_n2503;
  assign new_n2505 = new_n1700 & new_n2504;
  assign p_298_3387_ = new_n2498 | new_n2505;
  assign new_n2507 = new_n517 & ~new_n729;
  assign new_n2508 = ~new_n517 & new_n729;
  assign p_295_3352_ = new_n2507 | new_n2508;
  assign new_n2510 = new_n483 & ~new_n1708;
  assign new_n2511 = ~new_n483 & new_n1708;
  assign p_356_3424_ = new_n2510 | new_n2511;
  assign p_279_304_ = ~p_15_4_;
  assign p_432_428_ = p_1_0_;
  assign p_450_288_ = p_1459_167_;
  assign p_440_277_ = p_1492_172_;
  assign p_444_282_ = p_1480_170_;
  assign p_488_260_ = p_2236_180_;
  assign p_494_267_ = p_2218_177_;
  assign p_524_210_ = p_4437_204_;
  assign p_530_216_ = p_4420_201_;
  assign p_560_248_ = p_3698_185_;
  assign p_534_220_ = p_4410_199_;
  assign p_544_230_ = p_3749_194_;
  assign p_484_256_ = p_2247_182_;
  assign p_550_236_ = p_3729_191_;
  assign p_448_284_ = p_1469_169_;
  assign p_453_596_ = p_1_0_;
  assign p_540_227_ = p_4393_195_;
  assign p_554_240_ = p_3717_189_;
  assign p_3_312_ = p_1_0_;
  assign p_480_250_ = p_2256_184_;
  assign p_438_274_ = p_1496_173_;
  assign p_490_263_ = p_2230_179_;
  assign p_528_214_ = p_4427_202_;
  assign p_469_3452_ = p_422_3451_;
  assign p_486_258_ = p_2239_181_;
  assign p_538_224_ = p_4400_197_;
  assign p_292_392_ = p_281_547_;
  assign p_548_234_ = p_3737_192_;
  assign p_558_244_ = p_3705_187_;
  assign p_2_313_ = p_1_0_;
  assign p_542_246_ = p_3701_186_;
  assign p_546_232_ = p_3743_193_;
  assign p_552_238_ = p_3723_190_;
  assign p_556_242_ = p_3711_188_;
  assign p_446_393_ = p_106_53_;
  assign p_496_271_ = p_2208_175_;
  assign p_522_226_ = p_4394_196_;
  assign p_341_420_ = p_279_304_;
  assign p_492_265_ = p_2224_178_;
  assign p_526_212_ = p_4432_203_;
  assign p_436_286_ = p_1462_168_;
  assign p_532_218_ = p_4415_200_;
  assign p_286_419_ = p_279_304_;
  assign p_536_222_ = p_4405_198_;
  assign p_478_269_ = p_2211_176_;
  assign p_284_384_ = p_289_383_;
  assign p_419_3444_ = p_471_3445_;
  assign p_258_3122_ = p_264_3121_;
  assign p_442_280_ = p_1486_171_;
  assign p_482_253_ = p_2253_183_;
endmodule


