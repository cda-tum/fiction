module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi106, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi122, pi123, pi124, pi125, pi126, pi127, pi129,
    pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141 );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi106,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi122, pi123, pi124, pi125, pi126, pi127,
    pi129, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output  po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n595, n596, n597, n598, n599, n600, n601, n602, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n620, n621, n622, n623, n624, n625, n626, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n685, n686, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n861, n862, n863, n864, n865, n866, n868, n869, n870, n871, n872,
    n873, n875, n876, n877, n878, n879, n880, n882, n883, n884, n885, n886,
    n887, n889, n890, n891, n892, n893, n894, n896, n897, n898, n899, n900,
    n901, n903, n904, n905, n906, n907, n908, n910, n911, n912, n913, n914,
    n915, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n940,
    n941, n942, n943, n944, n945, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1136, n1137, n1138, n1140, n1141, n1142,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1157, n1158, n1159, n1162, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1236, n1237, n1238, n1240, n1241, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263, n1265, n1266,
    n1267, n1268, n1270, n1271, n1272, n1273, n1274, n1276, n1277, n1278,
    n1280, n1281, n1282, n1283, n1285, n1286, n1287, n1288, n1290, n1291,
    n1292, n1293, n1295, n1296, n1297, n1298, n1300, n1301, n1302, n1304,
    n1305, n1306, n1308, n1309, n1310, n1312, n1313, n1314, n1316, n1317,
    n1318, n1320, n1321, n1322, n1324, n1325, n1326, n1327, n1328, n1330,
    n1331, n1332, n1334, n1335, n1336, n1338, n1339, n1340, n1342, n1343,
    n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1365,
    n1366, n1367, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1377,
    n1378, n1379, n1381, n1382, n1383, n1385, n1386, n1387, n1388, n1389,
    n1391, n1392, n1393, n1395, n1396, n1397, n1399, n1400, n1401, n1403,
    n1404, n1405, n1407, n1408, n1409, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1428, n1429, n1430, n1432, n1433, n1434, n1436, n1437, n1438, n1440,
    n1441, n1442, n1444, n1445, n1446, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1529, n1530, n1531, n1532, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1570,
    n1571, n1572, n1573, n1575, n1576, n1577, n1578, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1588, n1589, n1590, n1591, n1592, n1594,
    n1595, n1596, n1597, n1598, n1600, n1601, n1602, n1603, n1604, n1606,
    n1607, n1608, n1609, n1610, n1613, n1614, n1615, n1616, n1619, n1620,
    n1621, n1623, n1628, n1629, n1631;
  assign n291 = ~pi013 & ~pi014;
  assign n292 = ~pi006 & ~pi007;
  assign n293 = n291 & n292;
  assign n294 = ~pi017 & ~pi021;
  assign n295 = ~pi008 & n294;
  assign n296 = ~pi012 & n295;
  assign n297 = n293 & n296;
  assign n298 = ~pi018 & ~pi019;
  assign n299 = ~pi004 & ~pi016;
  assign n300 = n298 & n299;
  assign n301 = ~pi005 & ~pi022;
  assign n302 = ~pi009 & ~pi011;
  assign n303 = n301 & n302;
  assign n304 = n300 & n303;
  assign n305 = n297 & n304;
  assign n306 = pi054 & ~n305;
  assign n307 = ~pi000 & ~n306;
  assign n308 = n301 & ~n302;
  assign n309 = ~pi056 & n308;
  assign n310 = ~pi056 & ~n301;
  assign n311 = ~pi008 & ~pi021;
  assign n312 = ~pi007 & pi013;
  assign n313 = n311 & n312;
  assign n314 = ~pi007 & n311;
  assign n315 = pi007 & ~n311;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi008 & pi021;
  assign n318 = ~pi013 & ~n317;
  assign n319 = n316 & n318;
  assign n320 = ~n313 & ~n319;
  assign n321 = ~pi014 & ~n320;
  assign n322 = ~pi013 & pi014;
  assign n323 = n314 & n322;
  assign n324 = ~n321 & ~n323;
  assign n325 = ~pi010 & ~n324;
  assign n326 = pi010 & n291;
  assign n327 = n314 & n326;
  assign n328 = ~n325 & ~n327;
  assign n329 = n301 & ~n328;
  assign n330 = n300 & n329;
  assign n331 = ~pi017 & n330;
  assign n332 = ~pi006 & ~pi012;
  assign n333 = n331 & n332;
  assign n334 = ~n310 & ~n333;
  assign n335 = n302 & ~n334;
  assign n336 = ~n309 & ~n335;
  assign n337 = pi054 & ~n336;
  assign n338 = ~n307 & ~n337;
  assign n339 = ~pi129 & ~n338;
  assign po015 = pi003 | ~n339;
  assign n341 = ~pi011 & ~pi012;
  assign n342 = n311 & n341;
  assign n343 = n300 & n342;
  assign n344 = ~pi010 & ~pi022;
  assign n345 = ~pi007 & ~pi013;
  assign n346 = ~pi005 & ~pi006;
  assign n347 = n345 & n346;
  assign n348 = ~pi014 & n347;
  assign n349 = n344 & n348;
  assign n350 = n343 & n349;
  assign n351 = ~pi017 & pi054;
  assign n352 = ~n350 & n351;
  assign n353 = ~pi001 & ~n352;
  assign n354 = ~pi014 & pi054;
  assign n355 = ~pi008 & ~pi011;
  assign n356 = n294 & n355;
  assign n357 = ~pi005 & n332;
  assign n358 = pi005 & ~n332;
  assign n359 = ~n357 & ~n358;
  assign n360 = pi006 & pi012;
  assign n361 = ~pi007 & ~n360;
  assign n362 = n359 & n361;
  assign n363 = pi007 & n357;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~pi013 & ~n364;
  assign n366 = n312 & n357;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~pi009 & ~n367;
  assign n369 = n345 & n357;
  assign n370 = pi009 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = n300 & ~n371;
  assign n373 = n356 & n372;
  assign n374 = n354 & n373;
  assign n375 = n344 & n374;
  assign n376 = ~n353 & ~n375;
  assign n377 = ~pi129 & ~n376;
  assign po016 = pi003 | ~n377;
  assign n379 = pi122 & pi127;
  assign n380 = ~pi045 & ~pi048;
  assign n381 = ~pi043 & ~pi047;
  assign n382 = n380 & n381;
  assign n383 = ~pi015 & ~pi020;
  assign n384 = ~pi024 & ~pi049;
  assign n385 = n383 & n384;
  assign n386 = n382 & n385;
  assign n387 = ~pi041 & ~pi046;
  assign n388 = ~pi038 & ~pi050;
  assign n389 = n387 & n388;
  assign n390 = ~pi042 & ~pi044;
  assign n391 = ~pi040 & n390;
  assign n392 = ~pi002 & n391;
  assign n393 = n389 & n392;
  assign n394 = n386 & n393;
  assign n395 = pi082 & ~n394;
  assign n396 = ~n379 & ~n395;
  assign n397 = ~pi065 & n396;
  assign n398 = ~pi024 & ~pi045;
  assign n399 = ~pi047 & ~pi048;
  assign n400 = n398 & n399;
  assign n401 = ~pi049 & n383;
  assign n402 = n400 & n401;
  assign n403 = ~pi038 & ~pi040;
  assign n404 = n390 & n403;
  assign n405 = ~pi046 & ~pi050;
  assign n406 = ~pi041 & n405;
  assign n407 = n404 & n406;
  assign n408 = ~pi043 & n407;
  assign n409 = n402 & n408;
  assign n410 = pi082 & ~n409;
  assign n411 = ~pi082 & n379;
  assign n412 = ~n410 & ~n411;
  assign n413 = pi002 & ~n412;
  assign n414 = ~n397 & ~n413;
  assign po017 = ~pi129 & ~n414;
  assign n416 = ~pi009 & ~pi014;
  assign n417 = n344 & n416;
  assign n418 = n347 & n417;
  assign n419 = ~pi008 & ~pi017;
  assign n420 = n341 & n419;
  assign n421 = ~pi021 & n300;
  assign n422 = n420 & n421;
  assign n423 = n418 & n422;
  assign n424 = ~pi061 & ~pi118;
  assign n425 = ~n423 & n424;
  assign n426 = pi000 & ~pi123;
  assign n427 = ~pi113 & n426;
  assign n428 = ~n425 & ~n427;
  assign po018 = ~pi129 & ~n428;
  assign n430 = pi010 & ~pi022;
  assign n431 = n416 & n430;
  assign n432 = n369 & n431;
  assign n433 = pi054 & n300;
  assign n434 = n356 & n433;
  assign n435 = n432 & n434;
  assign n436 = pi004 & ~pi054;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~pi129 & ~n437;
  assign po019 = ~pi003 & n438;
  assign n440 = pi005 & ~pi054;
  assign n441 = ~pi007 & n332;
  assign n442 = ~pi025 & ~pi029;
  assign n443 = pi028 & n442;
  assign n444 = n441 & n443;
  assign n445 = ~pi013 & n417;
  assign n446 = n444 & n445;
  assign n447 = ~pi059 & n356;
  assign n448 = ~pi016 & pi054;
  assign n449 = ~pi004 & ~pi019;
  assign n450 = ~pi018 & n449;
  assign n451 = ~pi005 & n450;
  assign n452 = n448 & n451;
  assign n453 = n447 & n452;
  assign n454 = n446 & n453;
  assign n455 = ~n440 & ~n454;
  assign n456 = ~pi129 & ~n455;
  assign po020 = ~pi003 & n456;
  assign n458 = pi006 & ~pi054;
  assign n459 = ~pi005 & ~pi007;
  assign n460 = pi025 & ~pi029;
  assign n461 = ~pi028 & n460;
  assign n462 = ~pi012 & n461;
  assign n463 = n459 & n462;
  assign n464 = n445 & n463;
  assign n465 = ~pi006 & n450;
  assign n466 = n448 & n465;
  assign n467 = n447 & n466;
  assign n468 = n464 & n467;
  assign n469 = ~n458 & ~n468;
  assign n470 = ~pi129 & ~n469;
  assign po021 = ~pi003 & n470;
  assign n472 = pi007 & ~pi054;
  assign n473 = ~pi018 & ~pi021;
  assign n474 = pi008 & ~pi017;
  assign n475 = n473 & n474;
  assign n476 = ~pi007 & n449;
  assign n477 = n448 & n476;
  assign n478 = n475 & n477;
  assign n479 = ~pi006 & n341;
  assign n480 = ~pi005 & n479;
  assign n481 = n445 & n480;
  assign n482 = n478 & n481;
  assign n483 = ~n472 & ~n482;
  assign n484 = ~pi129 & ~n483;
  assign po022 = ~pi003 & n484;
  assign n486 = pi008 & ~pi054;
  assign n487 = n369 & n417;
  assign n488 = ~pi017 & ~pi018;
  assign n489 = ~pi011 & pi021;
  assign n490 = n488 & n489;
  assign n491 = ~pi008 & n449;
  assign n492 = n448 & n491;
  assign n493 = n490 & n492;
  assign n494 = n487 & n493;
  assign n495 = ~n486 & ~n494;
  assign n496 = ~pi129 & ~n495;
  assign po023 = ~pi003 & n496;
  assign n498 = pi009 & ~pi054;
  assign n499 = n291 & n344;
  assign n500 = pi011 & n459;
  assign n501 = n332 & n500;
  assign n502 = n499 & n501;
  assign n503 = n419 & n473;
  assign n504 = ~pi009 & n449;
  assign n505 = n448 & n504;
  assign n506 = n503 & n505;
  assign n507 = n502 & n506;
  assign n508 = ~n498 & ~n507;
  assign n509 = ~pi129 & ~n508;
  assign po024 = ~pi003 & n509;
  assign n511 = pi010 & ~pi054;
  assign n512 = ~pi010 & n449;
  assign n513 = n448 & n512;
  assign n514 = n503 & n513;
  assign n515 = n459 & n479;
  assign n516 = ~pi009 & ~pi022;
  assign n517 = n322 & n516;
  assign n518 = n515 & n517;
  assign n519 = n514 & n518;
  assign n520 = ~n511 & ~n519;
  assign n521 = ~pi129 & ~n520;
  assign po025 = ~pi003 & n521;
  assign n523 = pi011 & ~pi054;
  assign n524 = ~pi011 & n449;
  assign n525 = n448 & n524;
  assign n526 = n503 & n525;
  assign n527 = ~pi010 & pi022;
  assign n528 = n416 & n527;
  assign n529 = n369 & n528;
  assign n530 = n526 & n529;
  assign n531 = ~n523 & ~n530;
  assign n532 = ~pi129 & ~n531;
  assign po026 = ~pi003 & n532;
  assign n534 = pi012 & ~pi054;
  assign n535 = ~pi012 & n449;
  assign n536 = n448 & n535;
  assign n537 = pi018 & n295;
  assign n538 = n536 & n537;
  assign n539 = ~pi011 & n418;
  assign n540 = n538 & n539;
  assign n541 = ~n534 & ~n540;
  assign n542 = ~pi129 & ~n541;
  assign po027 = ~pi003 & n542;
  assign n544 = pi013 & ~pi054;
  assign n545 = ~pi013 & n450;
  assign n546 = n448 & n545;
  assign n547 = n447 & n546;
  assign n548 = ~pi025 & pi029;
  assign n549 = ~pi028 & n548;
  assign n550 = n357 & n549;
  assign n551 = ~pi007 & n417;
  assign n552 = n550 & n551;
  assign n553 = n547 & n552;
  assign n554 = ~n544 & ~n553;
  assign n555 = ~pi129 & ~n554;
  assign po028 = ~pi003 & n555;
  assign n557 = pi014 & ~pi054;
  assign n558 = ~pi016 & n354;
  assign n559 = n449 & n558;
  assign n560 = n503 & n559;
  assign n561 = ~pi009 & pi013;
  assign n562 = n344 & n561;
  assign n563 = n515 & n562;
  assign n564 = n560 & n563;
  assign n565 = ~n557 & ~n564;
  assign n566 = ~pi129 & ~n565;
  assign po029 = ~pi003 & n566;
  assign n568 = ~pi041 & ~pi043;
  assign n569 = n399 & n568;
  assign n570 = ~pi045 & n384;
  assign n571 = n569 & n570;
  assign n572 = ~pi046 & n388;
  assign n573 = n391 & n572;
  assign n574 = ~pi015 & n573;
  assign n575 = n571 & n574;
  assign n576 = pi082 & ~n575;
  assign n577 = ~n379 & ~n576;
  assign n578 = ~pi070 & n577;
  assign n579 = ~pi048 & n381;
  assign n580 = n570 & n579;
  assign n581 = n407 & n580;
  assign n582 = pi015 & ~n581;
  assign n583 = ~pi045 & n399;
  assign n584 = ~pi002 & ~pi020;
  assign n585 = ~pi015 & ~n584;
  assign n586 = n408 & n585;
  assign n587 = n384 & n586;
  assign n588 = n583 & n587;
  assign n589 = ~n582 & ~n588;
  assign n590 = pi082 & ~n589;
  assign n591 = pi015 & n411;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n578 & n592;
  assign po030 = ~pi129 & ~n593;
  assign n595 = pi016 & ~pi054;
  assign n596 = pi006 & ~pi012;
  assign n597 = ~pi005 & n596;
  assign n598 = n345 & n597;
  assign n599 = n417 & n598;
  assign n600 = n434 & n599;
  assign n601 = ~n595 & ~n600;
  assign n602 = ~pi129 & ~n601;
  assign po031 = ~pi003 & n602;
  assign n604 = pi017 & ~pi054;
  assign n605 = ~pi007 & n346;
  assign n606 = ~pi025 & ~pi028;
  assign n607 = ~pi012 & n606;
  assign n608 = n605 & n607;
  assign n609 = n445 & n608;
  assign n610 = ~pi016 & n351;
  assign n611 = n450 & n610;
  assign n612 = ~pi011 & n311;
  assign n613 = ~pi029 & pi059;
  assign n614 = n612 & n613;
  assign n615 = n611 & n614;
  assign n616 = n609 & n615;
  assign n617 = ~n604 & ~n616;
  assign n618 = ~pi129 & ~n617;
  assign po032 = ~pi003 & n618;
  assign n620 = pi018 & ~pi054;
  assign n621 = pi016 & pi054;
  assign n622 = n450 & n621;
  assign n623 = n356 & n622;
  assign n624 = n487 & n623;
  assign n625 = ~n620 & ~n624;
  assign n626 = ~pi129 & ~n625;
  assign po033 = ~pi003 & n626;
  assign n628 = pi019 & ~pi054;
  assign n629 = pi017 & n612;
  assign n630 = ~pi004 & ~pi018;
  assign n631 = ~pi019 & n630;
  assign n632 = n448 & n631;
  assign n633 = n629 & n632;
  assign n634 = n487 & n633;
  assign n635 = ~n628 & ~n634;
  assign n636 = ~pi129 & ~n635;
  assign po034 = ~pi003 & n636;
  assign n638 = n381 & n387;
  assign n639 = ~pi024 & n380;
  assign n640 = n638 & n639;
  assign n641 = ~pi040 & ~pi042;
  assign n642 = n388 & n641;
  assign n643 = ~pi044 & n401;
  assign n644 = n642 & n643;
  assign n645 = n640 & n644;
  assign n646 = pi082 & ~n645;
  assign n647 = ~n379 & ~n646;
  assign n648 = ~pi071 & n647;
  assign n649 = ~pi050 & n403;
  assign n650 = ~pi015 & ~pi049;
  assign n651 = n390 & n650;
  assign n652 = n649 & n651;
  assign n653 = n640 & n652;
  assign n654 = pi020 & ~n653;
  assign n655 = pi002 & n645;
  assign n656 = ~n654 & ~n655;
  assign n657 = pi082 & ~n656;
  assign n658 = pi020 & n411;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~n648 & n659;
  assign po035 = ~pi129 & ~n660;
  assign n662 = pi021 & ~pi054;
  assign n663 = n355 & n488;
  assign n664 = ~pi021 & pi054;
  assign n665 = pi019 & n664;
  assign n666 = n299 & n665;
  assign n667 = n663 & n666;
  assign n668 = n487 & n667;
  assign n669 = ~n662 & ~n668;
  assign n670 = ~pi129 & ~n669;
  assign po036 = ~pi003 & n670;
  assign n672 = pi022 & ~pi054;
  assign n673 = ~pi022 & n449;
  assign n674 = n448 & n673;
  assign n675 = n503 & n674;
  assign n676 = ~pi009 & ~pi010;
  assign n677 = n291 & n676;
  assign n678 = pi005 & ~pi007;
  assign n679 = n479 & n678;
  assign n680 = n677 & n679;
  assign n681 = n675 & n680;
  assign n682 = ~n672 & ~n681;
  assign n683 = ~pi129 & ~n682;
  assign po037 = ~pi003 & n683;
  assign n685 = ~pi023 & pi055;
  assign n686 = ~pi129 & ~n685;
  assign po038 = pi061 & n686;
  assign n688 = ~pi047 & n568;
  assign n689 = n380 & n688;
  assign n690 = n573 & n689;
  assign n691 = pi082 & ~n690;
  assign n692 = n584 & n650;
  assign n693 = pi082 & ~n692;
  assign n694 = n379 & ~n693;
  assign n695 = ~n691 & ~n694;
  assign n696 = ~pi024 & ~n695;
  assign n697 = ~pi002 & ~pi045;
  assign n698 = n399 & n697;
  assign n699 = n401 & n698;
  assign n700 = n408 & n699;
  assign n701 = pi082 & ~n700;
  assign n702 = ~n379 & ~n701;
  assign n703 = pi063 & n702;
  assign n704 = ~pi043 & n387;
  assign n705 = n583 & n704;
  assign n706 = pi024 & pi082;
  assign n707 = n390 & n706;
  assign n708 = n649 & n707;
  assign n709 = n705 & n708;
  assign n710 = ~pi129 & ~n709;
  assign n711 = ~n703 & n710;
  assign po039 = ~n696 & n711;
  assign n713 = pi085 & pi116;
  assign n714 = ~pi085 & ~pi110;
  assign n715 = ~pi096 & n714;
  assign n716 = ~n713 & ~n715;
  assign n717 = pi100 & ~n716;
  assign n718 = pi025 & ~pi116;
  assign n719 = pi085 & n718;
  assign n720 = ~n717 & ~n719;
  assign n721 = ~pi026 & ~n720;
  assign n722 = ~pi051 & ~pi052;
  assign n723 = ~pi039 & n722;
  assign n724 = ~pi095 & ~pi100;
  assign n725 = ~pi097 & n724;
  assign n726 = ~pi110 & ~n725;
  assign n727 = pi025 & ~n726;
  assign n728 = pi026 & pi116;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n723 & ~n729;
  assign n731 = pi026 & n718;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~pi085 & ~n732;
  assign n734 = ~n721 & ~n733;
  assign n735 = ~pi027 & ~n734;
  assign n736 = ~pi039 & ~pi052;
  assign n737 = ~pi051 & n736;
  assign n738 = pi116 & n737;
  assign n739 = ~n718 & ~n738;
  assign n740 = pi027 & ~n739;
  assign n741 = n723 & n727;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~pi026 & ~pi085;
  assign n744 = ~n742 & n743;
  assign n745 = ~n735 & ~n744;
  assign n746 = ~pi053 & ~n745;
  assign n747 = pi025 & ~pi026;
  assign n748 = ~pi116 & n747;
  assign n749 = pi053 & ~pi085;
  assign n750 = ~pi027 & n749;
  assign n751 = n748 & n750;
  assign n752 = ~n746 & ~n751;
  assign n753 = ~pi058 & ~n752;
  assign n754 = ~pi027 & ~pi085;
  assign n755 = ~pi053 & pi058;
  assign n756 = n754 & n755;
  assign n757 = n748 & n756;
  assign n758 = ~n753 & ~n757;
  assign n759 = ~pi129 & ~n758;
  assign po040 = ~pi003 & n759;
  assign n761 = pi085 & ~pi116;
  assign n762 = ~pi110 & ~n761;
  assign n763 = ~n728 & n762;
  assign n764 = ~pi096 & n763;
  assign n765 = ~pi026 & n713;
  assign n766 = ~n764 & ~n765;
  assign n767 = pi100 & ~n766;
  assign n768 = ~pi085 & ~n738;
  assign n769 = pi026 & n768;
  assign n770 = ~n767 & ~n769;
  assign n771 = ~pi129 & ~n770;
  assign n772 = ~pi003 & n771;
  assign n773 = ~pi027 & ~pi053;
  assign n774 = ~pi058 & n773;
  assign po041 = n772 & n774;
  assign n776 = pi095 & ~pi096;
  assign n777 = pi027 & pi116;
  assign n778 = n762 & ~n777;
  assign n779 = n776 & n778;
  assign n780 = ~pi027 & n713;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~pi100 & ~n781;
  assign n783 = pi027 & n768;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~pi129 & ~n784;
  assign n786 = ~pi003 & n785;
  assign n787 = ~pi053 & ~pi058;
  assign n788 = ~pi026 & n787;
  assign po042 = n786 & n788;
  assign n790 = ~pi026 & ~n723;
  assign n791 = ~pi027 & n737;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~n726 & ~n792;
  assign n794 = pi026 & ~pi027;
  assign n795 = ~pi026 & pi027;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~pi116 & ~n796;
  assign n798 = ~n793 & ~n797;
  assign n799 = pi028 & ~n798;
  assign n800 = ~pi026 & ~pi100;
  assign n801 = ~pi110 & n800;
  assign n802 = n776 & n801;
  assign n803 = n728 & n737;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~pi027 & ~n804;
  assign n806 = n777 & n790;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~n799 & n807;
  assign n809 = ~pi085 & ~n808;
  assign n810 = pi028 & ~pi116;
  assign n811 = ~pi100 & pi116;
  assign n812 = ~n810 & ~n811;
  assign n813 = pi085 & ~n812;
  assign n814 = ~pi026 & ~pi027;
  assign n815 = n813 & n814;
  assign n816 = ~n809 & ~n815;
  assign n817 = ~pi053 & ~n816;
  assign n818 = ~pi027 & pi028;
  assign n819 = ~pi116 & n818;
  assign n820 = ~pi026 & n749;
  assign n821 = n819 & n820;
  assign n822 = ~n817 & ~n821;
  assign n823 = ~pi058 & ~n822;
  assign n824 = n743 & n755;
  assign n825 = n819 & n824;
  assign n826 = ~n823 & ~n825;
  assign n827 = ~pi129 & ~n826;
  assign po043 = ~pi003 & n827;
  assign n829 = pi029 & pi110;
  assign n830 = pi097 & ~pi110;
  assign n831 = ~pi096 & n830;
  assign n832 = pi029 & ~pi097;
  assign n833 = ~n831 & ~n832;
  assign n834 = n724 & ~n833;
  assign n835 = ~n829 & ~n834;
  assign n836 = ~pi058 & ~n835;
  assign n837 = pi097 & pi116;
  assign n838 = pi029 & ~pi116;
  assign n839 = ~n837 & ~n838;
  assign n840 = pi058 & ~n839;
  assign n841 = ~n836 & ~n840;
  assign n842 = ~pi053 & ~n841;
  assign n843 = pi053 & ~pi058;
  assign n844 = n838 & n843;
  assign n845 = ~n842 & ~n844;
  assign n846 = ~pi027 & ~n845;
  assign n847 = pi027 & n838;
  assign n848 = n787 & n847;
  assign n849 = ~n846 & ~n848;
  assign n850 = ~pi085 & ~n849;
  assign n851 = pi085 & n774;
  assign n852 = n838 & n851;
  assign n853 = ~n850 & ~n852;
  assign n854 = ~pi026 & ~n853;
  assign n855 = n754 & n787;
  assign n856 = pi026 & n855;
  assign n857 = n838 & n856;
  assign n858 = ~n854 & ~n857;
  assign n859 = ~pi129 & ~n858;
  assign po044 = ~pi003 & n859;
  assign n861 = pi030 & ~pi109;
  assign n862 = pi060 & pi109;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~pi106 & ~n863;
  assign n865 = pi088 & pi106;
  assign n866 = ~n864 & ~n865;
  assign po045 = ~pi129 & ~n866;
  assign n868 = pi089 & pi106;
  assign n869 = pi030 & pi109;
  assign n870 = pi031 & ~pi109;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~pi106 & ~n871;
  assign n873 = ~n868 & ~n872;
  assign po046 = ~pi129 & ~n873;
  assign n875 = pi099 & pi106;
  assign n876 = pi031 & pi109;
  assign n877 = pi032 & ~pi109;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~pi106 & ~n878;
  assign n880 = ~n875 & ~n879;
  assign po047 = ~pi129 & ~n880;
  assign n882 = pi090 & pi106;
  assign n883 = pi032 & pi109;
  assign n884 = pi033 & ~pi109;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~pi106 & ~n885;
  assign n887 = ~n882 & ~n886;
  assign po048 = ~pi129 & ~n887;
  assign n889 = pi091 & pi106;
  assign n890 = pi033 & pi109;
  assign n891 = pi034 & ~pi109;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~pi106 & ~n892;
  assign n894 = ~n889 & ~n893;
  assign po049 = ~pi129 & ~n894;
  assign n896 = pi092 & pi106;
  assign n897 = pi034 & pi109;
  assign n898 = pi035 & ~pi109;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~pi106 & ~n899;
  assign n901 = ~n896 & ~n900;
  assign po050 = ~pi129 & ~n901;
  assign n903 = pi098 & pi106;
  assign n904 = pi035 & pi109;
  assign n905 = pi036 & ~pi109;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~pi106 & ~n906;
  assign n908 = ~n903 & ~n907;
  assign po051 = ~pi129 & ~n908;
  assign n910 = pi093 & pi106;
  assign n911 = pi036 & pi109;
  assign n912 = pi037 & ~pi109;
  assign n913 = ~n911 & ~n912;
  assign n914 = ~pi106 & ~n913;
  assign n915 = ~n910 & ~n914;
  assign po052 = ~pi129 & ~n915;
  assign n917 = pi082 & ~n391;
  assign n918 = n406 & n579;
  assign n919 = n385 & n697;
  assign n920 = n918 & n919;
  assign n921 = pi082 & ~n920;
  assign n922 = n379 & ~n921;
  assign n923 = ~n917 & ~n922;
  assign n924 = ~pi038 & ~n923;
  assign n925 = ~pi002 & ~pi048;
  assign n926 = n398 & n925;
  assign n927 = n401 & n926;
  assign n928 = ~pi050 & n391;
  assign n929 = n638 & n928;
  assign n930 = n927 & n929;
  assign n931 = pi082 & ~n930;
  assign n932 = ~n379 & ~n931;
  assign n933 = pi074 & n932;
  assign n934 = ~pi044 & pi082;
  assign n935 = pi038 & n641;
  assign n936 = n934 & n935;
  assign n937 = ~pi129 & ~n936;
  assign n938 = ~n933 & n937;
  assign po053 = ~n924 & n938;
  assign n940 = ~pi051 & pi109;
  assign n941 = n736 & n940;
  assign n942 = ~pi106 & ~n941;
  assign n943 = pi109 & n722;
  assign n944 = pi039 & ~n943;
  assign n945 = n942 & ~n944;
  assign po054 = ~pi129 & ~n945;
  assign n947 = pi082 & ~n390;
  assign n948 = n579 & n919;
  assign n949 = n389 & n948;
  assign n950 = pi082 & ~n949;
  assign n951 = n379 & ~n950;
  assign n952 = ~n947 & ~n951;
  assign n953 = ~pi040 & ~n952;
  assign n954 = n388 & n390;
  assign n955 = n638 & n954;
  assign n956 = n927 & n955;
  assign n957 = pi082 & ~n956;
  assign n958 = ~n379 & ~n957;
  assign n959 = pi073 & n958;
  assign n960 = pi040 & pi082;
  assign n961 = n390 & n960;
  assign n962 = ~pi129 & ~n961;
  assign n963 = ~n959 & n962;
  assign po055 = ~n953 & n963;
  assign n965 = pi082 & ~n573;
  assign n966 = pi082 & ~n948;
  assign n967 = n379 & ~n966;
  assign n968 = ~n965 & ~n967;
  assign n969 = ~pi041 & ~n968;
  assign n970 = n381 & n405;
  assign n971 = n404 & n970;
  assign n972 = n927 & n971;
  assign n973 = pi082 & ~n972;
  assign n974 = ~n379 & ~n973;
  assign n975 = pi076 & n974;
  assign n976 = n403 & n405;
  assign n977 = pi041 & pi082;
  assign n978 = n390 & n977;
  assign n979 = n976 & n978;
  assign n980 = ~pi129 & ~n979;
  assign n981 = ~n975 & n980;
  assign po056 = ~n969 & n981;
  assign n983 = pi044 & pi082;
  assign n984 = n688 & n976;
  assign n985 = n927 & n984;
  assign n986 = pi082 & ~n985;
  assign n987 = n379 & ~n986;
  assign n988 = ~n983 & ~n987;
  assign n989 = ~pi042 & ~n988;
  assign n990 = ~pi044 & n649;
  assign n991 = n638 & n990;
  assign n992 = n927 & n991;
  assign n993 = pi082 & ~n992;
  assign n994 = ~n379 & ~n993;
  assign n995 = pi072 & n994;
  assign n996 = pi042 & n934;
  assign n997 = ~pi129 & ~n996;
  assign n998 = ~n995 & n997;
  assign po057 = ~n989 & n998;
  assign n1000 = pi082 & ~n407;
  assign n1001 = n385 & n698;
  assign n1002 = pi082 & ~n1001;
  assign n1003 = n379 & ~n1002;
  assign n1004 = ~n1000 & ~n1003;
  assign n1005 = ~pi043 & ~n1004;
  assign n1006 = ~pi047 & n407;
  assign n1007 = n927 & n1006;
  assign n1008 = pi082 & ~n1007;
  assign n1009 = ~n379 & ~n1008;
  assign n1010 = pi077 & n1009;
  assign n1011 = pi043 & n641;
  assign n1012 = n934 & n1011;
  assign n1013 = n389 & n1012;
  assign n1014 = ~pi129 & ~n1013;
  assign n1015 = ~n1010 & n1014;
  assign po058 = ~n1005 & n1015;
  assign n1017 = n638 & n642;
  assign n1018 = n927 & n1017;
  assign n1019 = pi082 & ~n1018;
  assign n1020 = pi067 & ~n379;
  assign n1021 = ~pi044 & n379;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1019 & ~n1022;
  assign n1024 = ~pi129 & ~n983;
  assign po059 = ~n1023 & n1024;
  assign n1026 = n399 & n704;
  assign n1027 = n388 & n391;
  assign n1028 = n1026 & n1027;
  assign n1029 = pi082 & ~n1028;
  assign n1030 = ~pi024 & n692;
  assign n1031 = pi082 & ~n1030;
  assign n1032 = n379 & ~n1031;
  assign n1033 = ~n1029 & ~n1032;
  assign n1034 = ~pi045 & ~n1033;
  assign n1035 = ~pi002 & n399;
  assign n1036 = n385 & n1035;
  assign n1037 = n408 & n1036;
  assign n1038 = pi082 & ~n1037;
  assign n1039 = ~n379 & ~n1038;
  assign n1040 = pi068 & n1039;
  assign n1041 = ~pi038 & n641;
  assign n1042 = pi045 & n1041;
  assign n1043 = n934 & n1042;
  assign n1044 = n918 & n1043;
  assign n1045 = ~pi129 & ~n1044;
  assign n1046 = ~n1040 & n1045;
  assign po060 = ~n1034 & n1046;
  assign n1048 = pi082 & ~n1027;
  assign n1049 = n688 & n927;
  assign n1050 = pi082 & ~n1049;
  assign n1051 = n379 & ~n1050;
  assign n1052 = ~n1048 & ~n1051;
  assign n1053 = ~pi046 & ~n1052;
  assign n1054 = ~pi050 & n404;
  assign n1055 = n1049 & n1054;
  assign n1056 = pi082 & ~n1055;
  assign n1057 = ~n379 & ~n1056;
  assign n1058 = pi075 & n1057;
  assign n1059 = pi046 & pi082;
  assign n1060 = n1054 & n1059;
  assign n1061 = ~pi129 & ~n1060;
  assign n1062 = ~n1058 & n1061;
  assign po061 = ~n1053 & n1062;
  assign n1064 = pi082 & ~n408;
  assign n1065 = pi082 & ~n927;
  assign n1066 = n379 & ~n1065;
  assign n1067 = ~n1064 & ~n1066;
  assign n1068 = ~pi047 & ~n1067;
  assign n1069 = n408 & n927;
  assign n1070 = pi082 & ~n1069;
  assign n1071 = ~n379 & ~n1070;
  assign n1072 = pi064 & n1071;
  assign n1073 = n568 & n572;
  assign n1074 = pi047 & n641;
  assign n1075 = n934 & n1074;
  assign n1076 = n1073 & n1075;
  assign n1077 = ~pi129 & ~n1076;
  assign n1078 = ~n1072 & n1077;
  assign po062 = ~n1068 & n1078;
  assign n1080 = n638 & n1027;
  assign n1081 = pi082 & ~n1080;
  assign n1082 = pi082 & ~n919;
  assign n1083 = n379 & ~n1082;
  assign n1084 = ~n1081 & ~n1083;
  assign n1085 = ~pi048 & ~n1084;
  assign n1086 = ~pi002 & ~pi047;
  assign n1087 = n398 & n401;
  assign n1088 = n1086 & n1087;
  assign n1089 = n408 & n1088;
  assign n1090 = pi082 & ~n1089;
  assign n1091 = ~n379 & ~n1090;
  assign n1092 = pi062 & n1091;
  assign n1093 = n381 & n406;
  assign n1094 = pi048 & n1041;
  assign n1095 = n934 & n1094;
  assign n1096 = n1093 & n1095;
  assign n1097 = ~pi129 & ~n1096;
  assign n1098 = ~n1092 & n1097;
  assign po063 = ~n1085 & n1098;
  assign n1100 = n384 & n1054;
  assign n1101 = n705 & n1100;
  assign n1102 = pi082 & ~n1101;
  assign n1103 = ~n379 & ~n1102;
  assign n1104 = ~pi069 & n1103;
  assign n1105 = ~pi024 & ~pi042;
  assign n1106 = n990 & n1105;
  assign n1107 = n705 & n1106;
  assign n1108 = pi049 & ~n1107;
  assign n1109 = ~pi002 & n383;
  assign n1110 = n1100 & ~n1109;
  assign n1111 = n638 & n1110;
  assign n1112 = n380 & n1111;
  assign n1113 = ~n1108 & ~n1112;
  assign n1114 = pi082 & ~n1113;
  assign n1115 = pi049 & n411;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~n1104 & n1116;
  assign po064 = ~pi129 & ~n1117;
  assign n1119 = pi082 & ~n404;
  assign n1120 = n704 & n1035;
  assign n1121 = n1087 & n1120;
  assign n1122 = pi082 & ~n1121;
  assign n1123 = n379 & ~n1122;
  assign n1124 = ~n1119 & ~n1123;
  assign n1125 = ~pi050 & ~n1124;
  assign n1126 = n404 & n638;
  assign n1127 = n927 & n1126;
  assign n1128 = pi082 & ~n1127;
  assign n1129 = ~n379 & ~n1128;
  assign n1130 = pi066 & n1129;
  assign n1131 = pi050 & n1041;
  assign n1132 = n934 & n1131;
  assign n1133 = ~pi129 & ~n1132;
  assign n1134 = ~n1130 & n1133;
  assign po065 = ~n1125 & n1134;
  assign n1136 = pi051 & ~pi109;
  assign n1137 = ~n940 & ~n1136;
  assign n1138 = ~pi106 & n1137;
  assign po066 = ~pi129 & ~n1138;
  assign n1140 = pi052 & ~n940;
  assign n1141 = ~pi106 & ~n943;
  assign n1142 = ~n1140 & n1141;
  assign po067 = ~pi129 & ~n1142;
  assign n1144 = pi058 & pi116;
  assign n1145 = ~pi058 & ~pi110;
  assign n1146 = ~pi096 & n1145;
  assign n1147 = n724 & n1146;
  assign n1148 = ~n1144 & ~n1147;
  assign n1149 = ~pi053 & ~n1148;
  assign n1150 = pi097 & n1149;
  assign n1151 = ~pi116 & n843;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~pi129 & ~n1152;
  assign n1154 = ~pi003 & n1153;
  assign n1155 = n754 & n1154;
  assign po068 = ~pi026 & n1155;
  assign n1157 = n408 & n1001;
  assign n1158 = pi082 & ~n1157;
  assign n1159 = ~n379 & ~n1158;
  assign po069 = pi129 | n1159;
  assign po129 = pi123 | pi129;
  assign n1162 = pi114 & ~pi122;
  assign po070 = ~po129 & n1162;
  assign n1164 = ~pi026 & pi058;
  assign n1165 = pi026 & ~pi058;
  assign n1166 = pi116 & n1165;
  assign n1167 = ~n1164 & ~n1166;
  assign n1168 = pi094 & ~n1167;
  assign n1169 = pi058 & ~pi116;
  assign n1170 = pi037 & ~pi116;
  assign n1171 = ~n1164 & ~n1170;
  assign n1172 = ~n1169 & ~n1171;
  assign n1173 = ~n1168 & ~n1172;
  assign n1174 = ~pi053 & ~n1173;
  assign n1175 = ~pi026 & pi037;
  assign n1176 = ~pi058 & n1175;
  assign n1177 = ~n1174 & ~n1176;
  assign n1178 = ~pi085 & ~n1177;
  assign n1179 = n787 & n1175;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = ~pi027 & ~n1180;
  assign n1182 = ~pi085 & n787;
  assign n1183 = n1175 & n1182;
  assign n1184 = ~n1181 & ~n1183;
  assign n1185 = ~pi129 & ~n1184;
  assign po071 = ~pi003 & n1185;
  assign n1187 = ~pi026 & ~pi053;
  assign n1188 = pi026 & pi053;
  assign n1189 = ~pi085 & ~n1188;
  assign n1190 = ~n1187 & ~n1189;
  assign n1191 = ~pi058 & ~n1190;
  assign n1192 = ~pi085 & n1187;
  assign n1193 = ~pi116 & n1192;
  assign n1194 = ~n1191 & ~n1193;
  assign n1195 = pi057 & ~n1194;
  assign n1196 = pi060 & n1144;
  assign n1197 = n1192 & n1196;
  assign n1198 = ~n1195 & ~n1197;
  assign n1199 = ~pi027 & ~n1198;
  assign n1200 = pi057 & ~pi058;
  assign n1201 = n1192 & n1200;
  assign n1202 = ~n1199 & ~n1201;
  assign n1203 = ~pi129 & ~n1202;
  assign po072 = ~pi003 & n1203;
  assign n1205 = n814 & n1169;
  assign n1206 = pi116 & ~n796;
  assign n1207 = ~pi058 & n1206;
  assign n1208 = n737 & n1207;
  assign n1209 = ~n1205 & ~n1208;
  assign n1210 = ~pi129 & ~n1209;
  assign n1211 = ~pi003 & n1210;
  assign n1212 = ~pi053 & n1211;
  assign po073 = ~pi085 & n1212;
  assign n1214 = ~n755 & ~n843;
  assign n1215 = ~pi116 & ~n1214;
  assign n1216 = ~n726 & n787;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = pi059 & ~n1217;
  assign n1219 = n726 & n787;
  assign n1220 = pi096 & n1219;
  assign n1221 = ~n1218 & ~n1220;
  assign n1222 = ~pi085 & ~n1221;
  assign n1223 = pi059 & ~pi116;
  assign n1224 = pi085 & n787;
  assign n1225 = n1223 & n1224;
  assign n1226 = ~n1222 & ~n1225;
  assign n1227 = ~pi027 & ~n1226;
  assign n1228 = pi027 & n1182;
  assign n1229 = n1223 & n1228;
  assign n1230 = ~n1227 & ~n1229;
  assign n1231 = ~pi026 & ~n1230;
  assign n1232 = n856 & n1223;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~pi129 & ~n1233;
  assign po074 = ~pi003 & n1234;
  assign n1236 = ~pi117 & ~pi122;
  assign n1237 = pi060 & ~n1236;
  assign n1238 = pi123 & n1236;
  assign po075 = n1237 | n1238;
  assign n1240 = ~pi114 & pi123;
  assign n1241 = ~pi122 & n1240;
  assign po076 = ~pi129 & n1241;
  assign n1243 = ~pi137 & ~pi138;
  assign n1244 = pi136 & n1243;
  assign n1245 = pi132 & pi133;
  assign n1246 = pi131 & n1245;
  assign n1247 = n1244 & n1246;
  assign n1248 = pi062 & ~n1247;
  assign n1249 = pi136 & ~pi137;
  assign n1250 = ~pi140 & n1249;
  assign n1251 = ~pi138 & n1246;
  assign n1252 = n1250 & n1251;
  assign n1253 = ~n1248 & ~n1252;
  assign po077 = pi129 | n1253;
  assign n1255 = pi063 & ~n1247;
  assign n1256 = ~pi142 & n1249;
  assign n1257 = n1251 & n1256;
  assign n1258 = ~n1255 & ~n1257;
  assign po078 = pi129 | n1258;
  assign n1260 = pi064 & ~n1247;
  assign n1261 = ~pi139 & n1249;
  assign n1262 = n1251 & n1261;
  assign n1263 = ~n1260 & ~n1262;
  assign po079 = pi129 | n1263;
  assign n1265 = pi065 & ~n1247;
  assign n1266 = ~pi146 & n1249;
  assign n1267 = n1251 & n1266;
  assign n1268 = ~n1265 & ~n1267;
  assign po080 = pi129 | n1268;
  assign n1270 = ~pi136 & ~pi137;
  assign n1271 = n1251 & n1270;
  assign n1272 = pi066 & ~n1271;
  assign n1273 = ~pi143 & n1271;
  assign n1274 = ~n1272 & ~n1273;
  assign po081 = pi129 | n1274;
  assign n1276 = pi067 & ~n1271;
  assign n1277 = ~pi139 & n1271;
  assign n1278 = ~n1276 & ~n1277;
  assign po082 = pi129 | n1278;
  assign n1280 = pi068 & ~n1247;
  assign n1281 = ~pi141 & n1249;
  assign n1282 = n1251 & n1281;
  assign n1283 = ~n1280 & ~n1282;
  assign po083 = pi129 | n1283;
  assign n1285 = pi069 & ~n1247;
  assign n1286 = ~pi143 & n1249;
  assign n1287 = n1251 & n1286;
  assign n1288 = ~n1285 & ~n1287;
  assign po084 = pi129 | n1288;
  assign n1290 = pi070 & ~n1247;
  assign n1291 = ~pi144 & n1249;
  assign n1292 = n1251 & n1291;
  assign n1293 = ~n1290 & ~n1292;
  assign po085 = pi129 | n1293;
  assign n1295 = pi071 & ~n1247;
  assign n1296 = ~pi145 & n1249;
  assign n1297 = n1251 & n1296;
  assign n1298 = ~n1295 & ~n1297;
  assign po086 = pi129 | n1298;
  assign n1300 = pi072 & ~n1271;
  assign n1301 = ~pi140 & n1271;
  assign n1302 = ~n1300 & ~n1301;
  assign po087 = pi129 | n1302;
  assign n1304 = pi073 & ~n1271;
  assign n1305 = ~pi141 & n1271;
  assign n1306 = ~n1304 & ~n1305;
  assign po088 = pi129 | n1306;
  assign n1308 = pi074 & ~n1271;
  assign n1309 = ~pi142 & n1271;
  assign n1310 = ~n1308 & ~n1309;
  assign po089 = pi129 | n1310;
  assign n1312 = pi075 & ~n1271;
  assign n1313 = ~pi144 & n1271;
  assign n1314 = ~n1312 & ~n1313;
  assign po090 = pi129 | n1314;
  assign n1316 = pi076 & ~n1271;
  assign n1317 = ~pi145 & n1271;
  assign n1318 = ~n1316 & ~n1317;
  assign po091 = pi129 | n1318;
  assign n1320 = pi077 & ~n1271;
  assign n1321 = ~pi146 & n1271;
  assign n1322 = ~n1320 & ~n1321;
  assign po092 = pi129 | n1322;
  assign n1324 = ~pi136 & pi137;
  assign n1325 = n1251 & n1324;
  assign n1326 = pi078 & ~n1325;
  assign n1327 = pi142 & n1325;
  assign n1328 = ~n1326 & ~n1327;
  assign po093 = ~pi129 & ~n1328;
  assign n1330 = pi079 & ~n1325;
  assign n1331 = pi143 & n1325;
  assign n1332 = ~n1330 & ~n1331;
  assign po094 = ~pi129 & ~n1332;
  assign n1334 = pi080 & ~n1325;
  assign n1335 = pi144 & n1325;
  assign n1336 = ~n1334 & ~n1335;
  assign po095 = ~pi129 & ~n1336;
  assign n1338 = pi081 & ~n1325;
  assign n1339 = pi145 & n1325;
  assign n1340 = ~n1338 & ~n1339;
  assign po096 = ~pi129 & ~n1340;
  assign n1342 = pi082 & ~n1325;
  assign n1343 = pi146 & n1325;
  assign n1344 = ~n1342 & ~n1343;
  assign po097 = ~pi129 & ~n1344;
  assign n1346 = pi089 & pi138;
  assign n1347 = ~pi062 & ~pi138;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = pi136 & ~n1348;
  assign n1350 = pi119 & pi138;
  assign n1351 = ~pi072 & ~pi138;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~pi136 & ~n1352;
  assign n1354 = ~n1349 & ~n1353;
  assign n1355 = ~pi137 & ~n1354;
  assign n1356 = ~pi115 & pi138;
  assign n1357 = pi087 & ~pi138;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~pi136 & ~n1358;
  assign n1360 = pi136 & ~pi138;
  assign n1361 = pi031 & n1360;
  assign n1362 = ~n1359 & ~n1361;
  assign n1363 = pi137 & ~n1362;
  assign po098 = n1355 | n1363;
  assign n1365 = pi084 & ~n1325;
  assign n1366 = pi141 & n1325;
  assign n1367 = ~n1365 & ~n1366;
  assign po099 = ~pi129 & ~n1367;
  assign n1369 = ~pi085 & ~n725;
  assign n1370 = ~pi110 & n1369;
  assign n1371 = pi096 & n1370;
  assign n1372 = ~n761 & ~n1371;
  assign n1373 = ~pi129 & ~n1372;
  assign n1374 = ~pi003 & n1373;
  assign n1375 = n774 & n1374;
  assign po100 = ~pi026 & n1375;
  assign n1377 = pi086 & ~n1325;
  assign n1378 = pi139 & n1325;
  assign n1379 = ~n1377 & ~n1378;
  assign po101 = ~pi129 & ~n1379;
  assign n1381 = pi087 & ~n1325;
  assign n1382 = pi140 & n1325;
  assign n1383 = ~n1381 & ~n1382;
  assign po102 = ~pi129 & ~n1383;
  assign n1385 = pi136 & pi137;
  assign n1386 = n1251 & n1385;
  assign n1387 = pi088 & ~n1386;
  assign n1388 = pi139 & n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign po103 = ~pi129 & ~n1389;
  assign n1391 = pi089 & ~n1386;
  assign n1392 = pi140 & n1386;
  assign n1393 = ~n1391 & ~n1392;
  assign po104 = ~pi129 & ~n1393;
  assign n1395 = pi090 & ~n1386;
  assign n1396 = pi142 & n1386;
  assign n1397 = ~n1395 & ~n1396;
  assign po105 = ~pi129 & ~n1397;
  assign n1399 = pi091 & ~n1386;
  assign n1400 = pi143 & n1386;
  assign n1401 = ~n1399 & ~n1400;
  assign po106 = ~pi129 & ~n1401;
  assign n1403 = pi092 & ~n1386;
  assign n1404 = pi144 & n1386;
  assign n1405 = ~n1403 & ~n1404;
  assign po107 = ~pi129 & ~n1405;
  assign n1407 = pi093 & ~n1386;
  assign n1408 = pi146 & n1386;
  assign n1409 = ~n1407 & ~n1408;
  assign po108 = ~pi129 & ~n1409;
  assign n1411 = pi082 & ~pi137;
  assign n1412 = ~pi136 & n1411;
  assign n1413 = pi138 & n1246;
  assign n1414 = n1412 & n1413;
  assign n1415 = pi094 & ~n1414;
  assign n1416 = pi142 & n1414;
  assign n1417 = ~n1415 & ~n1416;
  assign po109 = ~pi129 & ~n1417;
  assign n1419 = ~pi003 & ~n1246;
  assign n1420 = ~pi110 & n1419;
  assign n1421 = pi138 & n1412;
  assign n1422 = n1246 & ~n1421;
  assign n1423 = ~n1420 & ~n1422;
  assign n1424 = pi095 & ~n1423;
  assign n1425 = pi143 & n1414;
  assign n1426 = ~n1424 & ~n1425;
  assign po110 = ~pi129 & ~n1426;
  assign n1428 = pi096 & ~n1423;
  assign n1429 = pi146 & n1414;
  assign n1430 = ~n1428 & ~n1429;
  assign po111 = ~pi129 & ~n1430;
  assign n1432 = pi097 & ~n1423;
  assign n1433 = pi145 & n1414;
  assign n1434 = ~n1432 & ~n1433;
  assign po112 = ~pi129 & ~n1434;
  assign n1436 = pi098 & ~n1386;
  assign n1437 = pi145 & n1386;
  assign n1438 = ~n1436 & ~n1437;
  assign po113 = ~pi129 & ~n1438;
  assign n1440 = pi099 & ~n1386;
  assign n1441 = pi141 & n1386;
  assign n1442 = ~n1440 & ~n1441;
  assign po114 = ~pi129 & ~n1442;
  assign n1444 = pi100 & ~n1423;
  assign n1445 = pi144 & n1414;
  assign n1446 = ~n1444 & ~n1445;
  assign po115 = ~pi129 & ~n1446;
  assign n1448 = pi124 & pi138;
  assign n1449 = ~pi077 & ~pi138;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = ~pi136 & ~n1450;
  assign n1452 = ~pi065 & ~pi138;
  assign n1453 = pi093 & pi138;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = pi136 & ~n1454;
  assign n1456 = ~n1451 & ~n1455;
  assign n1457 = ~pi137 & ~n1456;
  assign n1458 = pi037 & n1360;
  assign n1459 = pi096 & pi138;
  assign n1460 = pi082 & ~pi138;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~pi136 & ~n1461;
  assign n1463 = ~n1458 & ~n1462;
  assign n1464 = pi137 & ~n1463;
  assign po116 = n1457 | n1464;
  assign n1466 = pi091 & n1249;
  assign n1467 = pi095 & n1324;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = pi138 & ~n1468;
  assign n1470 = pi079 & ~pi136;
  assign n1471 = pi034 & pi136;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = pi137 & ~n1472;
  assign n1474 = ~pi069 & pi136;
  assign n1475 = ~pi066 & ~pi136;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~pi137 & ~n1476;
  assign n1478 = ~n1473 & ~n1477;
  assign n1479 = ~pi138 & ~n1478;
  assign po117 = n1469 | n1479;
  assign n1481 = pi090 & n1249;
  assign n1482 = pi094 & n1324;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = pi138 & ~n1483;
  assign n1485 = pi078 & ~pi136;
  assign n1486 = pi033 & pi136;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = pi137 & ~n1487;
  assign n1489 = ~pi063 & pi136;
  assign n1490 = ~pi074 & ~pi136;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~pi137 & ~n1491;
  assign n1493 = ~n1488 & ~n1492;
  assign n1494 = ~pi138 & ~n1493;
  assign po118 = n1484 | n1494;
  assign n1496 = pi099 & n1249;
  assign n1497 = ~pi112 & n1324;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = pi138 & ~n1498;
  assign n1500 = ~pi068 & pi136;
  assign n1501 = ~pi073 & ~pi136;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~pi137 & ~n1502;
  assign n1504 = pi084 & ~pi136;
  assign n1505 = pi032 & pi136;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = pi137 & ~n1506;
  assign n1508 = ~n1503 & ~n1507;
  assign n1509 = ~pi138 & ~n1508;
  assign po119 = n1499 | n1509;
  assign n1511 = pi092 & pi138;
  assign n1512 = ~pi070 & ~pi138;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = pi136 & ~n1513;
  assign n1515 = pi125 & pi138;
  assign n1516 = ~pi075 & ~pi138;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~pi136 & ~n1517;
  assign n1519 = ~n1514 & ~n1518;
  assign n1520 = ~pi137 & ~n1519;
  assign n1521 = pi080 & ~pi138;
  assign n1522 = pi100 & pi138;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~pi136 & ~n1523;
  assign n1525 = pi035 & n1360;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = pi137 & ~n1526;
  assign po120 = n1520 | n1527;
  assign n1529 = n788 & n1370;
  assign n1530 = ~pi027 & n1529;
  assign n1531 = ~n713 & ~n1530;
  assign n1532 = ~pi129 & ~n1531;
  assign po121 = ~pi003 & n1532;
  assign n1534 = pi098 & pi138;
  assign n1535 = ~pi071 & ~pi138;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = pi136 & ~n1536;
  assign n1538 = ~pi076 & ~pi138;
  assign n1539 = pi023 & pi138;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~pi136 & ~n1540;
  assign n1542 = ~n1537 & ~n1541;
  assign n1543 = ~pi137 & ~n1542;
  assign n1544 = pi036 & n1360;
  assign n1545 = pi081 & ~pi138;
  assign n1546 = pi097 & pi138;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~pi136 & ~n1547;
  assign n1549 = ~n1544 & ~n1548;
  assign n1550 = pi137 & ~n1549;
  assign po122 = n1543 | n1550;
  assign n1552 = pi088 & pi138;
  assign n1553 = ~pi064 & ~pi138;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = pi136 & ~n1554;
  assign n1556 = pi120 & pi138;
  assign n1557 = ~pi067 & ~pi138;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~pi136 & ~n1558;
  assign n1560 = ~n1555 & ~n1559;
  assign n1561 = ~pi137 & ~n1560;
  assign n1562 = pi086 & ~pi138;
  assign n1563 = pi111 & pi138;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = ~pi136 & ~n1564;
  assign n1566 = pi030 & n1360;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = pi137 & ~n1567;
  assign po123 = n1561 | n1568;
  assign n1570 = ~n737 & n795;
  assign n1571 = ~n794 & ~n1570;
  assign n1572 = ~pi129 & ~n1571;
  assign n1573 = ~pi003 & n1572;
  assign po124 = pi116 & n1573;
  assign n1575 = ~pi097 & n755;
  assign n1576 = ~n843 & ~n1575;
  assign n1577 = ~pi129 & ~n1576;
  assign n1578 = ~pi003 & n1577;
  assign po125 = pi116 & n1578;
  assign n1580 = pi111 & ~n1421;
  assign n1581 = ~pi136 & pi139;
  assign n1582 = ~pi137 & pi138;
  assign n1583 = pi082 & n1582;
  assign n1584 = n1581 & n1583;
  assign n1585 = ~n1580 & ~n1584;
  assign n1586 = n1246 & ~n1585;
  assign po126 = ~pi129 & n1586;
  assign n1588 = ~pi136 & pi141;
  assign n1589 = n1583 & n1588;
  assign n1590 = ~pi112 & ~n1421;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = n1246 & ~n1591;
  assign po127 = ~pi129 & n1592;
  assign n1594 = ~pi054 & ~pi113;
  assign n1595 = ~pi011 & ~pi022;
  assign n1596 = pi054 & ~n1595;
  assign n1597 = ~n1594 & ~n1596;
  assign n1598 = ~pi129 & ~n1597;
  assign po128 = ~pi003 & n1598;
  assign n1600 = ~pi136 & pi140;
  assign n1601 = n1583 & n1600;
  assign n1602 = ~pi115 & ~n1421;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = n1246 & ~n1603;
  assign po130 = ~pi129 & n1604;
  assign n1606 = ~pi004 & ~pi012;
  assign n1607 = ~pi007 & ~pi009;
  assign n1608 = n1606 & n1607;
  assign n1609 = ~pi129 & ~n1608;
  assign n1610 = ~pi003 & n1609;
  assign po131 = pi054 & n1610;
  assign po132 = ~pi122 | pi129;
  assign n1613 = ~pi054 & pi118;
  assign n1614 = pi054 & ~pi059;
  assign n1615 = n549 & n1614;
  assign n1616 = ~n1613 & ~n1615;
  assign po133 = ~pi129 & ~n1616;
  assign po134 = ~pi129 & ~n724;
  assign n1619 = ~pi110 & ~pi120;
  assign n1620 = ~pi003 & n1619;
  assign n1621 = ~pi129 & ~n1620;
  assign po135 = ~pi111 & n1621;
  assign n1623 = pi081 & pi120;
  assign po136 = ~pi129 & n1623;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi057 & ~pi129;
  assign n1628 = ~pi096 & pi125;
  assign n1629 = ~pi003 & ~n1628;
  assign po140 = ~pi129 & ~n1629;
  assign n1631 = ~pi126 & pi132;
  assign po141 = pi133 & n1631;
endmodule


