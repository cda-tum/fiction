// Benchmark "top" written by ABC on Mon Nov 27 16:54:57 2023

module top ( 
    \1 , \4 , \7 , \10 , \13 , \16 , \19 , \22 , \25 , \28 , \31 , \34 ,
    \37 , \40 , \43 , \46 , \49 , \53 , \56 , \60 , \63 , \66 , \69 , \72 ,
    \76 , \79 , \82 , \85 , \88 , \91 , \94 , \99 , \104 ,
    \2753 , \2754 , \2755 , \2756 , \2762 , \2767 , \2768 , \2779 , \2780 ,
    \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2811 , \2886 ,
    \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2899   );
  input  \1 , \4 , \7 , \10 , \13 , \16 , \19 , \22 , \25 , \28 , \31 ,
    \34 , \37 , \40 , \43 , \46 , \49 , \53 , \56 , \60 , \63 , \66 , \69 ,
    \72 , \76 , \79 , \82 , \85 , \88 , \91 , \94 , \99 , \104 ;
  output \2753 , \2754 , \2755 , \2756 , \2762 , \2767 , \2768 , \2779 ,
    \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2811 ,
    \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2899 ;
  wire new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157, new_n158, new_n159, new_n160,
    new_n161, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n279, new_n280,
    new_n281, new_n283, new_n284, new_n285, new_n286, new_n288, new_n289,
    new_n290, new_n291, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n306,
    new_n307, new_n308, new_n310, new_n311, new_n312, new_n313, new_n315,
    new_n316, new_n317, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n359, new_n360,
    new_n361, new_n362, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n382, new_n383, new_n384,
    new_n385, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n406, new_n407, new_n408,
    new_n409;
  assign new_n59 = ~\28  & ~\43 ;
  assign new_n60 = \28  & \43 ;
  assign new_n61 = ~new_n59 & ~new_n60;
  assign new_n62 = \34  & ~new_n61;
  assign new_n63 = ~\34  & new_n61;
  assign new_n64 = ~new_n62 & ~new_n63;
  assign new_n65 = ~\37  & ~\46 ;
  assign new_n66 = \37  & \46 ;
  assign new_n67 = ~new_n65 & ~new_n66;
  assign new_n68 = \31  & ~new_n67;
  assign new_n69 = ~\31  & new_n67;
  assign new_n70 = ~new_n68 & ~new_n69;
  assign new_n71 = new_n64 & new_n70;
  assign new_n72 = ~new_n64 & ~new_n70;
  assign new_n73 = ~new_n71 & ~new_n72;
  assign new_n74 = \49  & ~\72 ;
  assign new_n75 = ~\104  & new_n74;
  assign new_n76 = ~\1  & ~\13 ;
  assign new_n77 = \1  & \13 ;
  assign new_n78 = ~new_n76 & ~new_n77;
  assign new_n79 = \16  & ~\19 ;
  assign new_n80 = ~\16  & \19 ;
  assign new_n81 = ~new_n79 & ~new_n80;
  assign new_n82 = new_n78 & new_n81;
  assign new_n83 = ~new_n78 & ~new_n81;
  assign new_n84 = ~new_n82 & ~new_n83;
  assign new_n85 = new_n75 & ~new_n84;
  assign new_n86 = ~new_n75 & new_n84;
  assign new_n87 = ~new_n85 & ~new_n86;
  assign new_n88 = new_n73 & new_n87;
  assign new_n89 = ~new_n73 & ~new_n87;
  assign new_n90 = ~new_n88 & ~new_n89;
  assign new_n91 = ~\94  & new_n90;
  assign new_n92 = \79  & ~new_n91;
  assign new_n93 = ~\79  & new_n91;
  assign new_n94 = ~new_n92 & ~new_n93;
  assign new_n95 = \69  & ~\94 ;
  assign new_n96 = \56  & ~new_n95;
  assign new_n97 = \60  & \69 ;
  assign new_n98 = ~\104  & new_n97;
  assign new_n99 = \28  & ~new_n67;
  assign new_n100 = ~\28  & new_n67;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = new_n98 & ~new_n101;
  assign new_n103 = ~new_n98 & new_n101;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = ~\25  & ~\40 ;
  assign new_n106 = \25  & \40 ;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = \10  & ~\19 ;
  assign new_n109 = ~\10  & \19 ;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = new_n107 & ~new_n110;
  assign new_n112 = ~new_n107 & new_n110;
  assign new_n113 = ~new_n111 & ~new_n112;
  assign new_n114 = new_n104 & new_n113;
  assign new_n115 = ~new_n104 & ~new_n113;
  assign new_n116 = ~new_n114 & ~new_n115;
  assign new_n117 = ~\94  & new_n116;
  assign new_n118 = new_n96 & ~new_n117;
  assign new_n119 = ~new_n96 & new_n117;
  assign new_n120 = ~new_n118 & ~new_n119;
  assign new_n121 = ~new_n94 & new_n120;
  assign new_n122 = \53  & ~\72 ;
  assign new_n123 = ~\25  & ~\46 ;
  assign new_n124 = \25  & \46 ;
  assign new_n125 = ~new_n123 & ~new_n124;
  assign new_n126 = ~\4  & ~\13 ;
  assign new_n127 = \4  & \13 ;
  assign new_n128 = ~new_n126 & ~new_n127;
  assign new_n129 = new_n125 & ~new_n128;
  assign new_n130 = ~new_n125 & new_n128;
  assign new_n131 = ~new_n129 & ~new_n130;
  assign new_n132 = ~\40  & ~\43 ;
  assign new_n133 = \40  & \43 ;
  assign new_n134 = ~new_n132 & ~new_n133;
  assign new_n135 = \22  & ~\31 ;
  assign new_n136 = ~\22  & \31 ;
  assign new_n137 = ~new_n135 & ~new_n136;
  assign new_n138 = new_n134 & ~new_n137;
  assign new_n139 = ~new_n134 & new_n137;
  assign new_n140 = ~new_n138 & ~new_n139;
  assign new_n141 = new_n131 & new_n140;
  assign new_n142 = ~new_n131 & ~new_n140;
  assign new_n143 = ~new_n141 & ~new_n142;
  assign new_n144 = ~new_n122 & new_n143;
  assign new_n145 = new_n122 & ~new_n143;
  assign new_n146 = ~new_n144 & ~new_n145;
  assign new_n147 = ~\94  & new_n146;
  assign new_n148 = \82  & ~new_n147;
  assign new_n149 = ~\82  & new_n147;
  assign new_n150 = ~new_n148 & ~new_n149;
  assign new_n151 = \56  & \69 ;
  assign new_n152 = ~\7  & ~\22 ;
  assign new_n153 = \7  & \22 ;
  assign new_n154 = ~new_n152 & ~new_n153;
  assign new_n155 = \16  & ~new_n154;
  assign new_n156 = ~\16  & new_n154;
  assign new_n157 = ~new_n155 & ~new_n156;
  assign new_n158 = new_n64 & new_n157;
  assign new_n159 = ~new_n64 & ~new_n157;
  assign new_n160 = ~new_n158 & ~new_n159;
  assign new_n161 = new_n151 & new_n160;
  assign new_n162 = ~new_n151 & ~new_n160;
  assign new_n163 = ~\94  & ~new_n161;
  assign new_n164 = ~new_n162 & new_n163;
  assign new_n165 = \85  & ~new_n164;
  assign new_n166 = ~\85  & new_n164;
  assign new_n167 = ~new_n165 & ~new_n166;
  assign new_n168 = new_n150 & new_n167;
  assign new_n169 = ~\72  & ~\94 ;
  assign new_n170 = \53  & ~new_n169;
  assign new_n171 = \60  & ~new_n95;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = \49  & ~new_n169;
  assign new_n174 = \63  & ~\104 ;
  assign new_n175 = ~\4  & ~\10 ;
  assign new_n176 = \4  & \10 ;
  assign new_n177 = ~new_n175 & ~new_n176;
  assign new_n178 = new_n154 & ~new_n177;
  assign new_n179 = ~new_n154 & new_n177;
  assign new_n180 = ~new_n178 & ~new_n179;
  assign new_n181 = new_n84 & new_n180;
  assign new_n182 = ~new_n84 & ~new_n180;
  assign new_n183 = ~new_n181 & ~new_n182;
  assign new_n184 = ~new_n125 & ~new_n183;
  assign new_n185 = new_n125 & new_n183;
  assign new_n186 = ~new_n184 & ~new_n185;
  assign new_n187 = new_n61 & ~new_n186;
  assign new_n188 = ~new_n61 & new_n186;
  assign new_n189 = ~new_n187 & ~new_n188;
  assign new_n190 = new_n174 & new_n189;
  assign new_n191 = ~new_n174 & ~new_n189;
  assign new_n192 = ~new_n190 & ~new_n191;
  assign new_n193 = ~\94  & ~new_n192;
  assign new_n194 = new_n173 & ~new_n193;
  assign new_n195 = ~new_n173 & new_n193;
  assign new_n196 = ~new_n194 & ~new_n195;
  assign new_n197 = new_n172 & ~new_n196;
  assign new_n198 = \1  & ~\4 ;
  assign new_n199 = ~\1  & \4 ;
  assign new_n200 = ~new_n198 & ~new_n199;
  assign new_n201 = \66  & ~\104 ;
  assign new_n202 = ~\10  & ~\40 ;
  assign new_n203 = \10  & \40 ;
  assign new_n204 = ~new_n202 & ~new_n203;
  assign new_n205 = \7  & ~new_n204;
  assign new_n206 = ~\7  & new_n204;
  assign new_n207 = ~new_n205 & ~new_n206;
  assign new_n208 = new_n201 & new_n207;
  assign new_n209 = ~new_n201 & ~new_n207;
  assign new_n210 = ~new_n208 & ~new_n209;
  assign new_n211 = new_n73 & ~new_n210;
  assign new_n212 = ~new_n73 & new_n210;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = new_n200 & new_n213;
  assign new_n215 = ~new_n200 & ~new_n213;
  assign new_n216 = ~new_n214 & ~new_n215;
  assign new_n217 = ~\94  & ~new_n216;
  assign new_n218 = \76  & ~new_n217;
  assign new_n219 = ~\76  & new_n217;
  assign new_n220 = ~new_n218 & ~new_n219;
  assign new_n221 = new_n197 & ~new_n220;
  assign new_n222 = \88  & \104 ;
  assign new_n223 = ~\99  & ~\104 ;
  assign new_n224 = \69  & \72 ;
  assign new_n225 = ~\94  & \104 ;
  assign new_n226 = ~new_n223 & ~new_n224;
  assign new_n227 = ~new_n225 & new_n226;
  assign new_n228 = ~new_n222 & new_n227;
  assign new_n229 = new_n221 & new_n228;
  assign new_n230 = new_n168 & new_n229;
  assign new_n231 = new_n121 & new_n230;
  assign new_n232 = ~\1  & ~new_n231;
  assign new_n233 = \1  & new_n231;
  assign \2753  = ~new_n232 & ~new_n233;
  assign new_n235 = new_n94 & new_n120;
  assign new_n236 = new_n229 & new_n235;
  assign new_n237 = ~new_n150 & new_n167;
  assign new_n238 = new_n236 & new_n237;
  assign new_n239 = \4  & ~new_n238;
  assign new_n240 = ~\4  & new_n238;
  assign \2754  = new_n239 | new_n240;
  assign new_n242 = new_n150 & ~new_n167;
  assign new_n243 = new_n236 & new_n242;
  assign new_n244 = \7  & ~new_n243;
  assign new_n245 = ~\7  & new_n243;
  assign \2755  = new_n244 | new_n245;
  assign new_n247 = new_n94 & ~new_n120;
  assign new_n248 = new_n230 & new_n247;
  assign new_n249 = ~\10  & ~new_n248;
  assign new_n250 = \10  & new_n248;
  assign \2756  = ~new_n249 & ~new_n250;
  assign new_n252 = \91  & \104 ;
  assign new_n253 = new_n227 & ~new_n252;
  assign new_n254 = ~new_n94 & ~new_n120;
  assign new_n255 = new_n253 & new_n254;
  assign new_n256 = new_n221 & new_n255;
  assign new_n257 = new_n242 & new_n256;
  assign new_n258 = \28  & ~new_n257;
  assign new_n259 = ~\28  & new_n257;
  assign \2762  = new_n258 | new_n259;
  assign new_n261 = ~new_n150 & ~new_n167;
  assign new_n262 = new_n121 & new_n253;
  assign new_n263 = new_n261 & new_n262;
  assign new_n264 = new_n221 & new_n263;
  assign new_n265 = ~\43  & ~new_n264;
  assign new_n266 = \43  & new_n264;
  assign \2767  = ~new_n265 & ~new_n266;
  assign new_n268 = new_n237 & new_n256;
  assign new_n269 = \46  & ~new_n268;
  assign new_n270 = ~\46  & new_n268;
  assign \2768  = new_n269 | new_n270;
  assign new_n272 = new_n197 & new_n220;
  assign new_n273 = new_n228 & new_n272;
  assign new_n274 = new_n121 & new_n273;
  assign new_n275 = new_n237 & new_n274;
  assign new_n276 = \13  & ~new_n275;
  assign new_n277 = ~\13  & new_n275;
  assign \2779  = new_n276 | new_n277;
  assign new_n279 = new_n242 & new_n274;
  assign new_n280 = \16  & ~new_n279;
  assign new_n281 = ~\16  & new_n279;
  assign \2780  = new_n280 | new_n281;
  assign new_n283 = new_n168 & new_n254;
  assign new_n284 = new_n273 & new_n283;
  assign new_n285 = ~\19  & ~new_n284;
  assign new_n286 = \19  & new_n284;
  assign \2781  = ~new_n285 & ~new_n286;
  assign new_n288 = new_n235 & new_n261;
  assign new_n289 = new_n273 & new_n288;
  assign new_n290 = ~\22  & ~new_n289;
  assign new_n291 = \22  & new_n289;
  assign \2782  = ~new_n290 & ~new_n291;
  assign new_n293 = new_n237 & new_n253;
  assign new_n294 = new_n247 & new_n293;
  assign new_n295 = new_n272 & new_n294;
  assign new_n296 = ~\25  & ~new_n295;
  assign new_n297 = \25  & new_n295;
  assign \2783  = ~new_n296 & ~new_n297;
  assign new_n299 = new_n172 & new_n196;
  assign new_n300 = ~new_n220 & new_n299;
  assign new_n301 = new_n262 & new_n300;
  assign new_n302 = new_n237 & new_n301;
  assign new_n303 = \31  & ~new_n302;
  assign new_n304 = ~\31  & new_n302;
  assign \2784  = new_n303 | new_n304;
  assign new_n306 = new_n242 & new_n301;
  assign new_n307 = \34  & ~new_n306;
  assign new_n308 = ~\34  & new_n306;
  assign \2785  = new_n307 | new_n308;
  assign new_n310 = new_n168 & new_n255;
  assign new_n311 = new_n300 & new_n310;
  assign new_n312 = ~\37  & ~new_n311;
  assign new_n313 = \37  & new_n311;
  assign \2786  = ~new_n312 & ~new_n313;
  assign new_n315 = new_n294 & new_n300;
  assign new_n316 = ~\40  & ~new_n315;
  assign new_n317 = \40  & new_n315;
  assign \2787  = ~new_n316 & ~new_n317;
  assign new_n319 = ~new_n172 & ~new_n196;
  assign new_n320 = new_n168 & new_n235;
  assign new_n321 = \99  & ~new_n224;
  assign new_n322 = ~new_n299 & ~new_n321;
  assign new_n323 = \60  & new_n170;
  assign new_n324 = new_n220 & ~new_n323;
  assign new_n325 = new_n320 & new_n324;
  assign new_n326 = ~new_n319 & new_n325;
  assign new_n327 = ~new_n322 & new_n326;
  assign new_n328 = ~new_n256 & ~new_n301;
  assign new_n329 = ~new_n237 & ~new_n242;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = ~new_n264 & ~new_n295;
  assign new_n332 = ~new_n311 & ~new_n315;
  assign new_n333 = new_n331 & new_n332;
  assign new_n334 = ~new_n330 & new_n333;
  assign new_n335 = ~new_n236 & ~new_n274;
  assign new_n336 = ~new_n329 & ~new_n335;
  assign new_n337 = ~new_n284 & ~new_n289;
  assign new_n338 = ~new_n231 & new_n337;
  assign new_n339 = ~new_n248 & new_n338;
  assign new_n340 = ~new_n336 & new_n339;
  assign new_n341 = new_n334 & new_n340;
  assign new_n342 = ~new_n168 & ~new_n235;
  assign new_n343 = ~new_n254 & ~new_n261;
  assign new_n344 = new_n220 & new_n343;
  assign new_n345 = ~new_n320 & ~new_n344;
  assign new_n346 = new_n321 & ~new_n342;
  assign new_n347 = ~new_n345 & new_n346;
  assign new_n348 = new_n299 & new_n347;
  assign new_n349 = ~\104  & ~new_n348;
  assign new_n350 = ~new_n327 & new_n349;
  assign \2811  = ~new_n341 | ~new_n350;
  assign new_n352 = ~\99  & \104 ;
  assign new_n353 = \94  & ~new_n341;
  assign new_n354 = \49  & new_n353;
  assign new_n355 = ~new_n192 & new_n354;
  assign new_n356 = new_n192 & ~new_n354;
  assign new_n357 = ~new_n352 & ~new_n355;
  assign \2886  = ~new_n356 & new_n357;
  assign new_n359 = \76  & new_n353;
  assign new_n360 = ~new_n216 & new_n359;
  assign new_n361 = new_n216 & ~new_n359;
  assign new_n362 = ~new_n352 & ~new_n360;
  assign \2887  = ~new_n361 & new_n362;
  assign new_n364 = \82  & new_n353;
  assign new_n365 = ~\104  & ~new_n146;
  assign new_n366 = \99  & \104 ;
  assign new_n367 = new_n143 & new_n366;
  assign new_n368 = ~new_n365 & ~new_n367;
  assign new_n369 = ~new_n352 & new_n368;
  assign new_n370 = ~new_n364 & ~new_n369;
  assign new_n371 = new_n364 & new_n368;
  assign \2888  = ~new_n370 & ~new_n371;
  assign new_n373 = ~\104  & new_n151;
  assign new_n374 = \85  & new_n353;
  assign new_n375 = ~new_n160 & new_n374;
  assign new_n376 = new_n160 & ~new_n374;
  assign new_n377 = ~new_n375 & ~new_n376;
  assign new_n378 = new_n373 & new_n377;
  assign new_n379 = ~new_n352 & ~new_n373;
  assign new_n380 = ~new_n377 & new_n379;
  assign \2889  = new_n378 | new_n380;
  assign new_n382 = \56  & new_n353;
  assign new_n383 = new_n116 & new_n382;
  assign new_n384 = ~new_n116 & ~new_n382;
  assign new_n385 = ~new_n352 & ~new_n383;
  assign \2890  = ~new_n384 & new_n385;
  assign new_n387 = ~\88  & \104 ;
  assign new_n388 = ~\63  & \104 ;
  assign new_n389 = new_n340 & ~new_n388;
  assign new_n390 = ~new_n183 & new_n389;
  assign new_n391 = new_n183 & ~new_n389;
  assign new_n392 = ~new_n387 & ~new_n390;
  assign \2891  = new_n391 | ~new_n392;
  assign new_n394 = ~new_n73 & ~new_n107;
  assign new_n395 = new_n73 & new_n107;
  assign new_n396 = ~new_n394 & ~new_n395;
  assign new_n397 = ~new_n334 & new_n396;
  assign new_n398 = new_n334 & ~new_n396;
  assign new_n399 = ~\104  & ~new_n397;
  assign new_n400 = ~new_n398 & new_n399;
  assign new_n401 = \66  & ~new_n396;
  assign new_n402 = ~\66  & new_n396;
  assign new_n403 = new_n252 & ~new_n401;
  assign new_n404 = ~new_n402 & new_n403;
  assign \2892  = ~new_n400 & ~new_n404;
  assign new_n406 = \79  & new_n353;
  assign new_n407 = new_n90 & new_n406;
  assign new_n408 = ~new_n90 & ~new_n406;
  assign new_n409 = ~new_n352 & ~new_n407;
  assign \2899  = ~new_n408 & new_n409;
endmodule


