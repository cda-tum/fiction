// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_,
    i_12_, i_1_, i_11_, i_2_, i_18_, i_17_, i_0_, i_21_, i_16_, i_15_,
    i_19_,
    o_1_, o_19_, o_2_, o_0_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_,
    o_28_, o_13_, o_21_, o_16_, o_22_, o_15_, o_23_, o_18_, o_24_, o_17_,
    o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_  );
  input  i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_,
    i_4_, i_12_, i_1_, i_11_, i_2_, i_18_, i_17_, i_0_, i_21_, i_16_,
    i_15_, i_19_;
  output o_1_, o_19_, o_2_, o_0_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_,
    o_28_, o_13_, o_21_, o_16_, o_22_, o_15_, o_23_, o_18_, o_24_, o_17_,
    o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_;
  wire new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58,
    new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65, new_n66,
    new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73, new_n74,
    new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81, new_n82,
    new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89, new_n90,
    new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97, new_n98,
    new_n99, new_n100, new_n101, new_n102, new_n103, new_n104, new_n105,
    new_n106, new_n107, new_n108, new_n109, new_n110, new_n111, new_n112,
    new_n113, new_n114, new_n115, new_n116, new_n117, new_n118, new_n119,
    new_n120, new_n121, new_n122, new_n123, new_n124, new_n125, new_n126,
    new_n127, new_n128, new_n129, new_n130, new_n131, new_n132, new_n133,
    new_n135, new_n136, new_n137, new_n138, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n280, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n327, new_n329, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n433,
    new_n434, new_n435, new_n436, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n486, new_n487, new_n488, new_n489, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587;
  assign new_n52 = i_18_ & ~i_21_;
  assign new_n53 = ~i_17_ & new_n52;
  assign new_n54 = ~i_14_ & ~i_15_;
  assign new_n55 = i_13_ & new_n54;
  assign new_n56 = new_n53 & new_n55;
  assign new_n57 = ~i_9_ & i_8_;
  assign new_n58 = ~i_7_ & new_n57;
  assign new_n59 = ~i_12_ & i_11_;
  assign new_n60 = i_10_ & new_n59;
  assign new_n61 = ~i_5_ & i_4_;
  assign new_n62 = ~i_2_ & new_n61;
  assign new_n63 = new_n58 & new_n60;
  assign new_n64 = new_n62 & new_n63;
  assign new_n65 = new_n56 & new_n64;
  assign new_n66 = ~i_9_ & ~i_8_;
  assign new_n67 = ~i_7_ & new_n66;
  assign new_n68 = ~i_17_ & ~i_15_;
  assign new_n69 = i_11_ & new_n68;
  assign new_n70 = ~i_5_ & i_6_;
  assign new_n71 = ~i_2_ & new_n70;
  assign new_n72 = new_n67 & new_n69;
  assign new_n73 = new_n71 & new_n72;
  assign new_n74 = new_n52 & new_n73;
  assign new_n75 = ~i_11_ & new_n68;
  assign new_n76 = i_2_ & new_n70;
  assign new_n77 = new_n67 & new_n75;
  assign new_n78 = new_n76 & new_n77;
  assign new_n79 = new_n52 & new_n78;
  assign new_n80 = ~i_9_ & ~i_11_;
  assign new_n81 = i_8_ & new_n80;
  assign new_n82 = i_18_ & ~i_17_;
  assign new_n83 = i_15_ & new_n82;
  assign new_n84 = ~i_7_ & i_5_;
  assign new_n85 = ~i_4_ & new_n84;
  assign new_n86 = new_n81 & new_n83;
  assign new_n87 = new_n85 & new_n86;
  assign new_n88 = ~i_21_ & new_n87;
  assign new_n89 = ~new_n74 & ~new_n79;
  assign new_n90 = ~new_n88 & new_n89;
  assign new_n91 = i_18_ & i_21_;
  assign new_n92 = ~i_17_ & new_n91;
  assign new_n93 = ~i_11_ & new_n54;
  assign new_n94 = new_n67 & new_n93;
  assign new_n95 = new_n76 & new_n94;
  assign new_n96 = new_n92 & new_n95;
  assign new_n97 = ~i_15_ & new_n82;
  assign new_n98 = ~i_21_ & new_n97;
  assign new_n99 = ~i_9_ & ~i_10_;
  assign new_n100 = i_8_ & new_n99;
  assign new_n101 = ~i_14_ & i_13_;
  assign new_n102 = i_11_ & new_n101;
  assign new_n103 = ~i_7_ & ~i_5_;
  assign new_n104 = ~i_2_ & new_n103;
  assign new_n105 = new_n100 & new_n102;
  assign new_n106 = new_n104 & new_n105;
  assign new_n107 = new_n98 & new_n106;
  assign new_n108 = i_11_ & new_n54;
  assign new_n109 = new_n67 & new_n108;
  assign new_n110 = new_n71 & new_n109;
  assign new_n111 = new_n92 & new_n110;
  assign new_n112 = ~new_n96 & ~new_n107;
  assign new_n113 = ~new_n111 & new_n112;
  assign new_n114 = i_9_ & i_11_;
  assign new_n115 = i_8_ & new_n114;
  assign new_n116 = new_n83 & new_n115;
  assign new_n117 = new_n104 & new_n116;
  assign new_n118 = i_11_ & i_15_;
  assign new_n119 = ~i_9_ & new_n118;
  assign new_n120 = ~i_18_ & ~i_17_;
  assign new_n121 = i_7_ & ~i_5_;
  assign new_n122 = i_2_ & new_n121;
  assign new_n123 = new_n119 & new_n120;
  assign new_n124 = new_n122 & new_n123;
  assign new_n125 = ~i_9_ & i_11_;
  assign new_n126 = i_8_ & new_n125;
  assign new_n127 = new_n83 & new_n126;
  assign new_n128 = new_n104 & new_n127;
  assign new_n129 = ~i_21_ & new_n128;
  assign new_n130 = ~new_n117 & ~new_n124;
  assign new_n131 = ~new_n129 & new_n130;
  assign new_n132 = new_n90 & new_n113;
  assign new_n133 = new_n131 & new_n132;
  assign o_1_ = new_n65 | ~new_n133;
  assign new_n135 = ~i_18_ & i_17_;
  assign new_n136 = ~i_15_ & new_n135;
  assign new_n137 = ~i_9_ & ~i_7_;
  assign new_n138 = ~i_5_ & new_n137;
  assign o_19_ = new_n136 & new_n138;
  assign new_n140 = ~i_17_ & i_15_;
  assign new_n141 = ~i_9_ & new_n140;
  assign new_n142 = ~i_7_ & i_8_;
  assign new_n143 = i_5_ & new_n142;
  assign new_n144 = new_n91 & new_n141;
  assign new_n145 = new_n143 & new_n144;
  assign new_n146 = i_18_ & ~i_19_;
  assign new_n147 = ~i_7_ & ~i_8_;
  assign new_n148 = ~i_5_ & new_n147;
  assign new_n149 = new_n141 & new_n146;
  assign new_n150 = new_n148 & new_n149;
  assign new_n151 = ~i_9_ & new_n68;
  assign new_n152 = ~i_7_ & ~i_6_;
  assign new_n153 = ~i_4_ & new_n152;
  assign new_n154 = i_18_ & new_n151;
  assign new_n155 = new_n153 & new_n154;
  assign new_n156 = ~new_n145 & ~new_n150;
  assign new_n157 = ~new_n155 & new_n156;
  assign new_n158 = i_18_ & i_19_;
  assign new_n159 = i_5_ & new_n147;
  assign new_n160 = new_n151 & new_n158;
  assign new_n161 = new_n159 & new_n160;
  assign new_n162 = new_n141 & new_n158;
  assign new_n163 = new_n148 & new_n162;
  assign new_n164 = new_n146 & new_n151;
  assign new_n165 = new_n159 & new_n164;
  assign new_n166 = ~new_n161 & ~new_n163;
  assign new_n167 = ~new_n165 & new_n166;
  assign new_n168 = ~i_12_ & new_n68;
  assign new_n169 = ~i_6_ & new_n137;
  assign new_n170 = i_18_ & new_n168;
  assign new_n171 = new_n169 & new_n170;
  assign new_n172 = i_9_ & new_n68;
  assign new_n173 = i_7_ & i_8_;
  assign new_n174 = i_5_ & new_n173;
  assign new_n175 = i_18_ & new_n172;
  assign new_n176 = new_n174 & new_n175;
  assign new_n177 = ~i_11_ & ~i_17_;
  assign new_n178 = ~i_9_ & new_n177;
  assign new_n179 = ~i_7_ & i_6_;
  assign new_n180 = ~i_5_ & new_n179;
  assign new_n181 = i_18_ & new_n178;
  assign new_n182 = new_n180 & new_n181;
  assign new_n183 = ~new_n171 & ~new_n176;
  assign new_n184 = ~new_n182 & new_n183;
  assign new_n185 = new_n157 & new_n167;
  assign new_n186 = new_n184 & new_n185;
  assign new_n187 = i_9_ & i_12_;
  assign new_n188 = i_8_ & new_n187;
  assign new_n189 = new_n97 & new_n188;
  assign new_n190 = new_n85 & new_n189;
  assign new_n191 = i_16_ & ~i_15_;
  assign new_n192 = ~i_9_ & new_n191;
  assign new_n193 = i_1_ & new_n121;
  assign new_n194 = new_n120 & new_n192;
  assign new_n195 = new_n193 & new_n194;
  assign new_n196 = i_9_ & ~i_11_;
  assign new_n197 = i_8_ & new_n196;
  assign new_n198 = i_2_ & new_n103;
  assign new_n199 = new_n83 & new_n197;
  assign new_n200 = new_n198 & new_n199;
  assign new_n201 = ~new_n190 & ~new_n195;
  assign new_n202 = ~new_n200 & new_n201;
  assign new_n203 = ~i_11_ & i_15_;
  assign new_n204 = i_8_ & new_n203;
  assign new_n205 = new_n53 & new_n204;
  assign new_n206 = new_n198 & new_n205;
  assign new_n207 = i_12_ & ~i_15_;
  assign new_n208 = i_8_ & new_n207;
  assign new_n209 = new_n53 & new_n208;
  assign new_n210 = new_n85 & new_n209;
  assign new_n211 = ~i_9_ & ~i_15_;
  assign new_n212 = i_8_ & new_n211;
  assign new_n213 = new_n120 & new_n212;
  assign new_n214 = new_n193 & new_n213;
  assign new_n215 = ~new_n206 & ~new_n210;
  assign new_n216 = ~new_n214 & new_n215;
  assign new_n217 = ~new_n88 & new_n202;
  assign new_n218 = new_n216 & new_n217;
  assign new_n219 = i_8_ & ~i_12_;
  assign new_n220 = i_5_ & new_n219;
  assign new_n221 = new_n97 & new_n220;
  assign new_n222 = ~i_5_ & new_n57;
  assign new_n223 = i_21_ & new_n83;
  assign new_n224 = new_n222 & new_n223;
  assign new_n225 = new_n154 & new_n174;
  assign new_n226 = ~new_n221 & ~new_n224;
  assign new_n227 = ~new_n225 & new_n226;
  assign new_n228 = ~i_9_ & ~i_17_;
  assign new_n229 = ~i_7_ & new_n228;
  assign new_n230 = i_18_ & new_n229;
  assign new_n231 = new_n71 & new_n230;
  assign new_n232 = i_9_ & new_n140;
  assign new_n233 = ~i_5_ & new_n173;
  assign new_n234 = i_18_ & new_n232;
  assign new_n235 = new_n233 & new_n234;
  assign new_n236 = i_5_ & new_n57;
  assign new_n237 = i_21_ & new_n97;
  assign new_n238 = new_n236 & new_n237;
  assign new_n239 = ~new_n231 & ~new_n235;
  assign new_n240 = ~new_n238 & new_n239;
  assign new_n241 = i_18_ & new_n141;
  assign new_n242 = new_n233 & new_n241;
  assign new_n243 = i_8_ & ~i_5_;
  assign new_n244 = ~i_2_ & new_n243;
  assign new_n245 = new_n83 & new_n244;
  assign new_n246 = ~i_5_ & new_n142;
  assign new_n247 = new_n97 & new_n246;
  assign new_n248 = ~new_n242 & ~new_n245;
  assign new_n249 = ~new_n247 & new_n248;
  assign new_n250 = new_n227 & new_n240;
  assign new_n251 = new_n249 & new_n250;
  assign new_n252 = new_n186 & new_n218;
  assign o_2_ = ~new_n251 | ~new_n252;
  assign new_n254 = i_17_ & i_15_;
  assign new_n255 = ~i_9_ & new_n254;
  assign new_n256 = ~i_0_ & new_n103;
  assign new_n257 = ~i_18_ & new_n255;
  assign new_n258 = new_n256 & new_n257;
  assign new_n259 = ~i_14_ & i_12_;
  assign new_n260 = ~i_9_ & new_n259;
  assign new_n261 = ~i_15_ & new_n120;
  assign new_n262 = i_4_ & new_n103;
  assign new_n263 = new_n260 & new_n261;
  assign new_n264 = new_n262 & new_n263;
  assign new_n265 = ~i_21_ & new_n264;
  assign new_n266 = i_15_ & new_n135;
  assign new_n267 = ~i_9_ & i_7_;
  assign new_n268 = ~i_5_ & new_n267;
  assign new_n269 = new_n266 & new_n268;
  assign new_n270 = ~new_n258 & ~new_n265;
  assign new_n271 = ~new_n269 & new_n270;
  assign new_n272 = i_5_ & new_n137;
  assign new_n273 = new_n135 & new_n272;
  assign new_n274 = i_5_ & new_n211;
  assign new_n275 = new_n135 & new_n274;
  assign new_n276 = ~new_n273 & ~new_n275;
  assign new_n277 = ~o_19_ & new_n276;
  assign o_0_ = ~new_n271 | ~new_n277;
  assign o_23_ = new_n175 & new_n246;
  assign new_n280 = ~new_n150 & ~new_n163;
  assign o_25_ = o_23_ | ~new_n280;
  assign new_n282 = ~i_9_ & i_10_;
  assign new_n283 = i_8_ & new_n282;
  assign new_n284 = ~i_14_ & ~i_13_;
  assign new_n285 = ~i_12_ & new_n284;
  assign new_n286 = new_n283 & new_n285;
  assign new_n287 = new_n262 & new_n286;
  assign new_n288 = new_n98 & new_n287;
  assign new_n289 = ~new_n107 & ~new_n288;
  assign new_n290 = ~new_n79 & new_n289;
  assign new_n291 = ~new_n65 & new_n290;
  assign new_n292 = ~i_10_ & ~i_13_;
  assign new_n293 = ~i_9_ & new_n292;
  assign new_n294 = ~i_14_ & new_n68;
  assign new_n295 = new_n293 & new_n294;
  assign new_n296 = new_n246 & new_n295;
  assign new_n297 = new_n52 & new_n296;
  assign new_n298 = ~i_9_ & ~i_12_;
  assign new_n299 = i_8_ & new_n298;
  assign new_n300 = i_4_ & new_n84;
  assign new_n301 = new_n97 & new_n299;
  assign new_n302 = new_n300 & new_n301;
  assign new_n303 = ~i_21_ & new_n302;
  assign new_n304 = ~new_n88 & ~new_n297;
  assign new_n305 = ~new_n303 & new_n304;
  assign new_n306 = ~i_5_ & ~i_6_;
  assign new_n307 = i_4_ & new_n306;
  assign new_n308 = new_n67 & new_n168;
  assign new_n309 = new_n307 & new_n308;
  assign new_n310 = new_n52 & new_n309;
  assign new_n311 = i_12_ & new_n68;
  assign new_n312 = ~i_4_ & new_n306;
  assign new_n313 = new_n67 & new_n311;
  assign new_n314 = new_n312 & new_n313;
  assign new_n315 = new_n52 & new_n314;
  assign new_n316 = ~new_n310 & ~new_n315;
  assign new_n317 = ~new_n74 & new_n316;
  assign new_n318 = i_0_ & new_n103;
  assign new_n319 = new_n257 & new_n318;
  assign new_n320 = new_n136 & new_n268;
  assign new_n321 = ~new_n129 & ~new_n319;
  assign new_n322 = ~new_n320 & new_n321;
  assign new_n323 = new_n305 & new_n317;
  assign new_n324 = new_n322 & new_n323;
  assign o_12_ = ~new_n291 | ~new_n324;
  assign o_8_ = ~i_20_ & i_14_;
  assign new_n327 = ~i_20_ & i_21_;
  assign o_26_ = o_8_ | new_n327;
  assign new_n329 = ~i_18_ & new_n151;
  assign o_11_ = new_n193 & new_n329;
  assign new_n331 = new_n160 & new_n174;
  assign new_n332 = i_9_ & ~i_15_;
  assign new_n333 = i_8_ & new_n332;
  assign new_n334 = ~i_17_ & new_n158;
  assign new_n335 = i_3_ & new_n103;
  assign new_n336 = new_n333 & new_n334;
  assign new_n337 = new_n335 & new_n336;
  assign new_n338 = new_n162 & new_n233;
  assign new_n339 = ~new_n331 & ~new_n337;
  assign new_n340 = ~new_n338 & new_n339;
  assign new_n341 = ~new_n79 & ~new_n315;
  assign new_n342 = ~new_n88 & new_n341;
  assign new_n343 = ~new_n161 & ~new_n319;
  assign new_n344 = ~new_n320 & new_n343;
  assign new_n345 = new_n340 & new_n342;
  assign o_27_ = ~new_n344 | ~new_n345;
  assign new_n347 = i_9_ & ~i_12_;
  assign new_n348 = i_8_ & new_n347;
  assign new_n349 = new_n97 & new_n348;
  assign new_n350 = new_n300 & new_n349;
  assign new_n351 = ~new_n265 & ~new_n350;
  assign new_n352 = ~new_n124 & new_n351;
  assign new_n353 = ~new_n117 & ~new_n303;
  assign new_n354 = ~new_n129 & new_n353;
  assign new_n355 = new_n352 & new_n354;
  assign new_n356 = ~i_19_ & new_n83;
  assign new_n357 = new_n233 & new_n356;
  assign new_n358 = ~i_2_ & new_n121;
  assign new_n359 = ~i_18_ & new_n141;
  assign new_n360 = new_n358 & new_n359;
  assign new_n361 = ~new_n357 & ~new_n360;
  assign new_n362 = ~new_n269 & new_n361;
  assign new_n363 = ~i_11_ & new_n140;
  assign new_n364 = ~i_18_ & new_n363;
  assign new_n365 = new_n268 & new_n364;
  assign new_n366 = ~i_19_ & new_n97;
  assign new_n367 = new_n174 & new_n366;
  assign new_n368 = ~new_n365 & ~new_n367;
  assign new_n369 = ~new_n258 & new_n368;
  assign new_n370 = ~i_9_ & ~i_18_;
  assign new_n371 = ~i_1_ & new_n121;
  assign new_n372 = new_n370 & new_n371;
  assign new_n373 = ~new_n319 & ~new_n372;
  assign new_n374 = ~new_n320 & new_n373;
  assign new_n375 = new_n362 & new_n369;
  assign new_n376 = new_n374 & new_n375;
  assign o_14_ = ~new_n355 | ~new_n376;
  assign new_n378 = ~new_n200 & ~new_n210;
  assign new_n379 = ~new_n206 & new_n378;
  assign new_n380 = ~i_12_ & new_n54;
  assign new_n381 = new_n67 & new_n380;
  assign new_n382 = new_n307 & new_n381;
  assign new_n383 = new_n92 & new_n382;
  assign new_n384 = ~new_n111 & ~new_n383;
  assign new_n385 = ~new_n190 & new_n384;
  assign new_n386 = ~i_18_ & ~i_19_;
  assign new_n387 = i_17_ & new_n386;
  assign new_n388 = ~i_9_ & i_15_;
  assign new_n389 = ~i_5_ & new_n388;
  assign new_n390 = new_n387 & new_n389;
  assign new_n391 = ~new_n365 & ~new_n390;
  assign new_n392 = ~new_n258 & new_n391;
  assign new_n393 = new_n379 & new_n385;
  assign new_n394 = new_n392 & new_n393;
  assign new_n395 = ~i_17_ & i_16_;
  assign new_n396 = ~i_15_ & new_n395;
  assign new_n397 = new_n52 & new_n396;
  assign new_n398 = i_12_ & new_n284;
  assign new_n399 = ~i_5_ & new_n152;
  assign new_n400 = new_n283 & new_n398;
  assign new_n401 = new_n399 & new_n400;
  assign new_n402 = new_n397 & new_n401;
  assign new_n403 = ~i_17_ & ~i_16_;
  assign new_n404 = ~i_15_ & new_n403;
  assign new_n405 = new_n52 & new_n404;
  assign new_n406 = new_n180 & new_n400;
  assign new_n407 = new_n405 & new_n406;
  assign new_n408 = new_n401 & new_n405;
  assign new_n409 = ~new_n402 & ~new_n407;
  assign new_n410 = ~new_n408 & new_n409;
  assign new_n411 = i_12_ & new_n101;
  assign new_n412 = new_n283 & new_n411;
  assign new_n413 = new_n198 & new_n412;
  assign new_n414 = new_n98 & new_n413;
  assign new_n415 = new_n397 & new_n406;
  assign new_n416 = i_11_ & new_n259;
  assign new_n417 = new_n283 & new_n416;
  assign new_n418 = new_n104 & new_n417;
  assign new_n419 = new_n53 & new_n418;
  assign new_n420 = ~new_n414 & ~new_n415;
  assign new_n421 = ~new_n419 & new_n420;
  assign new_n422 = new_n410 & new_n421;
  assign new_n423 = ~new_n235 & ~new_n319;
  assign new_n424 = ~new_n224 & new_n423;
  assign new_n425 = ~new_n150 & ~new_n360;
  assign new_n426 = ~new_n145 & new_n425;
  assign new_n427 = ~new_n245 & ~new_n273;
  assign new_n428 = ~new_n242 & new_n427;
  assign new_n429 = new_n424 & new_n426;
  assign new_n430 = new_n428 & new_n429;
  assign new_n431 = new_n394 & new_n422;
  assign o_28_ = ~new_n430 | ~new_n431;
  assign new_n433 = ~new_n258 & ~new_n269;
  assign new_n434 = ~new_n319 & new_n433;
  assign new_n435 = ~new_n273 & ~new_n320;
  assign new_n436 = ~o_19_ & new_n435;
  assign o_13_ = ~new_n434 | ~new_n436;
  assign new_n438 = ~i_8_ & new_n211;
  assign new_n439 = i_5_ & new_n179;
  assign new_n440 = new_n82 & new_n438;
  assign new_n441 = new_n439 & new_n440;
  assign new_n442 = new_n82 & new_n333;
  assign new_n443 = new_n180 & new_n442;
  assign new_n444 = ~i_8_ & new_n388;
  assign new_n445 = new_n82 & new_n444;
  assign new_n446 = new_n399 & new_n445;
  assign new_n447 = ~new_n443 & ~new_n446;
  assign new_n448 = ~new_n242 & new_n447;
  assign o_21_ = new_n441 | ~new_n448;
  assign new_n450 = new_n58 & new_n416;
  assign new_n451 = new_n71 & new_n450;
  assign new_n452 = new_n405 & new_n451;
  assign new_n453 = ~i_2_ & new_n306;
  assign new_n454 = new_n450 & new_n453;
  assign new_n455 = new_n397 & new_n454;
  assign new_n456 = ~new_n65 & ~new_n452;
  assign new_n457 = ~new_n455 & new_n456;
  assign new_n458 = i_6_ & new_n142;
  assign new_n459 = ~i_14_ & ~i_12_;
  assign new_n460 = ~i_9_ & new_n459;
  assign new_n461 = i_2_ & new_n61;
  assign new_n462 = new_n458 & new_n460;
  assign new_n463 = new_n461 & new_n462;
  assign new_n464 = new_n98 & new_n463;
  assign new_n465 = new_n409 & ~new_n464;
  assign new_n466 = new_n457 & new_n465;
  assign new_n467 = i_9_ & i_8_;
  assign new_n468 = i_5_ & new_n467;
  assign new_n469 = new_n170 & new_n468;
  assign new_n470 = new_n146 & new_n172;
  assign new_n471 = new_n246 & new_n470;
  assign new_n472 = ~new_n297 & ~new_n469;
  assign new_n473 = ~new_n471 & new_n472;
  assign new_n474 = ~i_10_ & new_n101;
  assign new_n475 = new_n58 & new_n474;
  assign new_n476 = new_n76 & new_n475;
  assign new_n477 = new_n98 & new_n476;
  assign new_n478 = ~new_n107 & ~new_n477;
  assign new_n479 = ~new_n288 & new_n478;
  assign new_n480 = new_n234 & new_n244;
  assign new_n481 = ~new_n176 & ~new_n480;
  assign new_n482 = ~new_n235 & new_n481;
  assign new_n483 = new_n473 & new_n479;
  assign new_n484 = new_n482 & new_n483;
  assign o_16_ = ~new_n466 | ~new_n484;
  assign new_n486 = new_n180 & new_n445;
  assign new_n487 = ~new_n441 & ~new_n486;
  assign new_n488 = ~new_n235 & ~o_23_;
  assign new_n489 = ~new_n242 & new_n488;
  assign o_22_ = ~new_n487 | ~new_n489;
  assign o_15_ = new_n136 & new_n272;
  assign new_n492 = i_2_ & new_n306;
  assign new_n493 = new_n475 & new_n492;
  assign new_n494 = new_n98 & new_n493;
  assign new_n495 = ~new_n408 & ~new_n415;
  assign new_n496 = ~new_n494 & new_n495;
  assign new_n497 = i_12_ & new_n54;
  assign new_n498 = new_n67 & new_n497;
  assign new_n499 = new_n312 & new_n498;
  assign new_n500 = new_n92 & new_n499;
  assign new_n501 = ~new_n96 & ~new_n500;
  assign new_n502 = ~new_n163 & new_n501;
  assign o_18_ = ~new_n496 | ~new_n502;
  assign new_n504 = ~new_n88 & ~new_n265;
  assign new_n505 = ~new_n303 & new_n504;
  assign new_n506 = new_n148 & new_n154;
  assign new_n507 = ~new_n129 & ~new_n214;
  assign new_n508 = ~new_n506 & new_n507;
  assign o_24_ = ~new_n505 | ~new_n508;
  assign new_n510 = ~new_n79 & ~new_n500;
  assign new_n511 = ~new_n315 & new_n510;
  assign new_n512 = ~new_n88 & ~new_n319;
  assign new_n513 = ~new_n320 & new_n512;
  assign new_n514 = ~new_n96 & new_n511;
  assign o_17_ = ~new_n513 | ~new_n514;
  assign new_n516 = ~new_n265 & new_n316;
  assign new_n517 = ~new_n288 & ~new_n500;
  assign new_n518 = ~new_n383 & new_n517;
  assign new_n519 = ~new_n88 & ~new_n350;
  assign new_n520 = ~new_n303 & new_n519;
  assign new_n521 = new_n516 & new_n518;
  assign new_n522 = new_n520 & new_n521;
  assign o_20_ = new_n65 | ~new_n522;
  assign new_n524 = i_5_ & new_n152;
  assign new_n525 = new_n440 & new_n524;
  assign new_n526 = ~new_n446 & ~new_n525;
  assign new_n527 = ~new_n176 & ~new_n320;
  assign new_n528 = ~new_n273 & new_n527;
  assign new_n529 = ~o_19_ & ~o_23_;
  assign new_n530 = ~new_n225 & new_n529;
  assign new_n531 = new_n434 & new_n528;
  assign new_n532 = new_n530 & new_n531;
  assign o_10_ = ~new_n526 | ~new_n532;
  assign new_n534 = ~new_n74 & ~new_n310;
  assign new_n535 = ~new_n265 & new_n534;
  assign new_n536 = ~i_7_ & i_4_;
  assign new_n537 = i_2_ & new_n536;
  assign new_n538 = new_n55 & new_n299;
  assign new_n539 = new_n537 & new_n538;
  assign new_n540 = new_n53 & new_n539;
  assign new_n541 = ~new_n414 & ~new_n494;
  assign new_n542 = ~new_n540 & new_n541;
  assign new_n543 = ~new_n190 & ~new_n200;
  assign new_n544 = ~new_n210 & new_n543;
  assign new_n545 = new_n535 & new_n542;
  assign new_n546 = new_n544 & new_n545;
  assign new_n547 = ~new_n145 & ~new_n176;
  assign new_n548 = ~new_n238 & new_n547;
  assign new_n549 = ~new_n206 & ~o_15_;
  assign new_n550 = ~new_n165 & new_n549;
  assign new_n551 = ~o_19_ & ~new_n221;
  assign new_n552 = ~new_n225 & new_n551;
  assign new_n553 = new_n548 & new_n550;
  assign new_n554 = new_n552 & new_n553;
  assign new_n555 = ~new_n477 & new_n546;
  assign o_9_ = ~new_n554 | ~new_n555;
  assign new_n557 = i_9_ & new_n191;
  assign new_n558 = new_n82 & new_n557;
  assign new_n559 = new_n246 & new_n558;
  assign new_n560 = ~new_n150 & ~new_n225;
  assign new_n561 = ~new_n242 & new_n560;
  assign new_n562 = new_n167 & ~new_n559;
  assign o_7_ = ~new_n561 | ~new_n562;
  assign new_n564 = ~new_n415 & ~new_n494;
  assign new_n565 = ~new_n96 & new_n564;
  assign new_n566 = ~new_n383 & ~new_n500;
  assign new_n567 = ~new_n111 & new_n566;
  assign new_n568 = ~new_n408 & new_n565;
  assign o_5_ = ~new_n567 | ~new_n568;
  assign new_n570 = ~new_n65 & ~new_n408;
  assign new_n571 = ~new_n415 & new_n570;
  assign new_n572 = ~new_n107 & ~new_n494;
  assign new_n573 = ~new_n288 & new_n572;
  assign new_n574 = new_n571 & new_n573;
  assign new_n575 = ~new_n74 & ~new_n297;
  assign new_n576 = ~new_n303 & new_n575;
  assign new_n577 = ~new_n310 & new_n384;
  assign new_n578 = new_n576 & new_n577;
  assign new_n579 = new_n322 & new_n578;
  assign o_6_ = ~new_n574 | ~new_n579;
  assign new_n581 = ~new_n161 & ~new_n258;
  assign new_n582 = ~new_n165 & ~new_n269;
  assign new_n583 = ~new_n319 & new_n582;
  assign new_n584 = ~new_n225 & ~o_23_;
  assign new_n585 = ~new_n242 & new_n584;
  assign new_n586 = new_n436 & new_n583;
  assign new_n587 = new_n585 & new_n586;
  assign o_3_ = ~new_n581 | ~new_n587;
  assign o_4_ = ~i_20_ & ~i_14_;
endmodule


