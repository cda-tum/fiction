// Benchmark "top" written by ABC on Mon Nov 27 16:49:22 2023

module top ( 
    \1 , \5 , \9 , \13 , \17 , \21 , \25 , \29 , \33 , \37 , \41 , \45 ,
    \49 , \53 , \57 , \61 , \65 , \69 , \73 , \77 , \81 , \85 , \89 , \93 ,
    \97 , \101 , \105 , \109 , \113 , \117 , \121 , \125 , \129 , \130 ,
    \131 , \132 , \133 , \134 , \135 , \136 , \137 ,
    \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 ,
    \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 ,
    \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 ,
    \754 , \755   );
  input  \1 , \5 , \9 , \13 , \17 , \21 , \25 , \29 , \33 , \37 , \41 ,
    \45 , \49 , \53 , \57 , \61 , \65 , \69 , \73 , \77 , \81 , \85 , \89 ,
    \93 , \97 , \101 , \105 , \109 , \113 , \117 , \121 , \125 , \129 ,
    \130 , \131 , \132 , \133 , \134 , \135 , \136 , \137 ;
  output \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 ,
    \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 ,
    \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 ,
    \754 , \755 ;
  wire new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n323,
    new_n324, new_n325, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n334, new_n335, new_n336, new_n338, new_n339, new_n340,
    new_n342, new_n343, new_n344, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n352, new_n353, new_n354, new_n356, new_n357, new_n358,
    new_n360, new_n361, new_n362, new_n364, new_n365, new_n366, new_n367,
    new_n369, new_n370, new_n371, new_n373, new_n374, new_n375, new_n377,
    new_n378, new_n379, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n396, new_n397, new_n398, new_n400, new_n401,
    new_n402, new_n404, new_n405, new_n406, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n414, new_n415, new_n416, new_n418, new_n419,
    new_n420, new_n422, new_n423, new_n424, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n433, new_n434, new_n435, new_n437,
    new_n438, new_n439, new_n441, new_n442, new_n443, new_n445, new_n446,
    new_n447, new_n448, new_n450, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n458, new_n459, new_n460;
  assign new_n74 = ~\81  & ~\85 ;
  assign new_n75 = \81  & \85 ;
  assign new_n76 = ~new_n74 & ~new_n75;
  assign new_n77 = \89  & ~\93 ;
  assign new_n78 = ~\89  & \93 ;
  assign new_n79 = ~new_n77 & ~new_n78;
  assign new_n80 = new_n76 & new_n79;
  assign new_n81 = ~new_n76 & ~new_n79;
  assign new_n82 = ~new_n80 & ~new_n81;
  assign new_n83 = ~\1  & ~\33 ;
  assign new_n84 = \1  & \33 ;
  assign new_n85 = ~new_n83 & ~new_n84;
  assign new_n86 = \17  & ~\49 ;
  assign new_n87 = ~\17  & \49 ;
  assign new_n88 = ~new_n86 & ~new_n87;
  assign new_n89 = \129  & \137 ;
  assign new_n90 = ~\65  & ~\69 ;
  assign new_n91 = \65  & \69 ;
  assign new_n92 = ~new_n90 & ~new_n91;
  assign new_n93 = \73  & ~\77 ;
  assign new_n94 = ~\73  & \77 ;
  assign new_n95 = ~new_n93 & ~new_n94;
  assign new_n96 = new_n92 & new_n95;
  assign new_n97 = ~new_n92 & ~new_n95;
  assign new_n98 = ~new_n96 & ~new_n97;
  assign new_n99 = new_n89 & ~new_n98;
  assign new_n100 = ~new_n89 & new_n98;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = new_n88 & new_n101;
  assign new_n103 = ~new_n88 & ~new_n101;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = new_n85 & ~new_n104;
  assign new_n106 = ~new_n85 & new_n104;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = new_n82 & new_n107;
  assign new_n109 = ~new_n82 & ~new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = ~\49  & ~\53 ;
  assign new_n112 = \49  & \53 ;
  assign new_n113 = ~new_n111 & ~new_n112;
  assign new_n114 = \57  & ~\61 ;
  assign new_n115 = ~\57  & \61 ;
  assign new_n116 = ~new_n114 & ~new_n115;
  assign new_n117 = new_n113 & new_n116;
  assign new_n118 = ~new_n113 & ~new_n116;
  assign new_n119 = ~new_n117 & ~new_n118;
  assign new_n120 = \93  & ~new_n119;
  assign new_n121 = ~\93  & new_n119;
  assign new_n122 = ~new_n120 & ~new_n121;
  assign new_n123 = \136  & \137 ;
  assign new_n124 = ~\17  & ~\21 ;
  assign new_n125 = \17  & \21 ;
  assign new_n126 = ~new_n124 & ~new_n125;
  assign new_n127 = \25  & ~\29 ;
  assign new_n128 = ~\25  & \29 ;
  assign new_n129 = ~new_n127 & ~new_n128;
  assign new_n130 = new_n126 & new_n129;
  assign new_n131 = ~new_n126 & ~new_n129;
  assign new_n132 = ~new_n130 & ~new_n131;
  assign new_n133 = ~\77  & ~\109 ;
  assign new_n134 = \77  & \109 ;
  assign new_n135 = ~new_n133 & ~new_n134;
  assign new_n136 = \125  & ~new_n135;
  assign new_n137 = ~\125  & new_n135;
  assign new_n138 = ~new_n136 & ~new_n137;
  assign new_n139 = new_n132 & new_n138;
  assign new_n140 = ~new_n132 & ~new_n138;
  assign new_n141 = ~new_n139 & ~new_n140;
  assign new_n142 = new_n123 & ~new_n141;
  assign new_n143 = ~new_n123 & new_n141;
  assign new_n144 = ~new_n142 & ~new_n143;
  assign new_n145 = new_n122 & new_n144;
  assign new_n146 = ~new_n122 & ~new_n144;
  assign new_n147 = ~new_n145 & ~new_n146;
  assign new_n148 = ~\1  & ~\5 ;
  assign new_n149 = \1  & \5 ;
  assign new_n150 = ~new_n148 & ~new_n149;
  assign new_n151 = \9  & ~\13 ;
  assign new_n152 = ~\9  & \13 ;
  assign new_n153 = ~new_n151 & ~new_n152;
  assign new_n154 = new_n150 & new_n153;
  assign new_n155 = ~new_n150 & ~new_n153;
  assign new_n156 = ~new_n154 & ~new_n155;
  assign new_n157 = \121  & ~new_n156;
  assign new_n158 = ~\121  & new_n156;
  assign new_n159 = ~new_n157 & ~new_n158;
  assign new_n160 = \135  & \137 ;
  assign new_n161 = ~\33  & ~\37 ;
  assign new_n162 = \33  & \37 ;
  assign new_n163 = ~new_n161 & ~new_n162;
  assign new_n164 = \41  & ~\45 ;
  assign new_n165 = ~\41  & \45 ;
  assign new_n166 = ~new_n164 & ~new_n165;
  assign new_n167 = new_n163 & new_n166;
  assign new_n168 = ~new_n163 & ~new_n166;
  assign new_n169 = ~new_n167 & ~new_n168;
  assign new_n170 = ~\89  & ~\105 ;
  assign new_n171 = \89  & \105 ;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = \73  & ~new_n172;
  assign new_n174 = ~\73  & new_n172;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176 = new_n169 & new_n175;
  assign new_n177 = ~new_n169 & ~new_n175;
  assign new_n178 = ~new_n176 & ~new_n177;
  assign new_n179 = new_n160 & ~new_n178;
  assign new_n180 = ~new_n160 & new_n178;
  assign new_n181 = ~new_n179 & ~new_n180;
  assign new_n182 = new_n159 & new_n181;
  assign new_n183 = ~new_n159 & ~new_n181;
  assign new_n184 = ~new_n182 & ~new_n183;
  assign new_n185 = new_n147 & ~new_n184;
  assign new_n186 = ~\97  & ~\101 ;
  assign new_n187 = \97  & \101 ;
  assign new_n188 = ~new_n186 & ~new_n187;
  assign new_n189 = \105  & ~\109 ;
  assign new_n190 = ~\105  & \109 ;
  assign new_n191 = ~new_n189 & ~new_n190;
  assign new_n192 = new_n188 & new_n191;
  assign new_n193 = ~new_n188 & ~new_n191;
  assign new_n194 = ~new_n192 & ~new_n193;
  assign new_n195 = ~\9  & ~\25 ;
  assign new_n196 = \9  & \25 ;
  assign new_n197 = ~new_n195 & ~new_n196;
  assign new_n198 = \41  & ~\57 ;
  assign new_n199 = ~\41  & \57 ;
  assign new_n200 = ~new_n198 & ~new_n199;
  assign new_n201 = \131  & \137 ;
  assign new_n202 = ~new_n98 & new_n201;
  assign new_n203 = new_n98 & ~new_n201;
  assign new_n204 = ~new_n202 & ~new_n203;
  assign new_n205 = new_n200 & new_n204;
  assign new_n206 = ~new_n200 & ~new_n204;
  assign new_n207 = ~new_n205 & ~new_n206;
  assign new_n208 = new_n197 & ~new_n207;
  assign new_n209 = ~new_n197 & new_n207;
  assign new_n210 = ~new_n208 & ~new_n209;
  assign new_n211 = new_n194 & new_n210;
  assign new_n212 = ~new_n194 & ~new_n210;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = new_n110 & new_n213;
  assign new_n215 = \37  & ~\53 ;
  assign new_n216 = ~\37  & \53 ;
  assign new_n217 = ~new_n215 & ~new_n216;
  assign new_n218 = new_n194 & ~new_n217;
  assign new_n219 = ~new_n194 & new_n217;
  assign new_n220 = ~new_n218 & ~new_n219;
  assign new_n221 = ~\113  & ~\117 ;
  assign new_n222 = \113  & \117 ;
  assign new_n223 = ~new_n221 & ~new_n222;
  assign new_n224 = \121  & ~\125 ;
  assign new_n225 = ~\121  & \125 ;
  assign new_n226 = ~new_n224 & ~new_n225;
  assign new_n227 = new_n223 & new_n226;
  assign new_n228 = ~new_n223 & ~new_n226;
  assign new_n229 = ~new_n227 & ~new_n228;
  assign new_n230 = \130  & \137 ;
  assign new_n231 = ~\5  & ~\21 ;
  assign new_n232 = \5  & \21 ;
  assign new_n233 = ~new_n231 & ~new_n232;
  assign new_n234 = new_n230 & ~new_n233;
  assign new_n235 = ~new_n230 & new_n233;
  assign new_n236 = ~new_n234 & ~new_n235;
  assign new_n237 = new_n229 & ~new_n236;
  assign new_n238 = ~new_n229 & new_n236;
  assign new_n239 = ~new_n237 & ~new_n238;
  assign new_n240 = new_n220 & new_n239;
  assign new_n241 = ~new_n220 & ~new_n239;
  assign new_n242 = ~new_n240 & ~new_n241;
  assign new_n243 = \132  & \137 ;
  assign new_n244 = ~new_n82 & new_n243;
  assign new_n245 = new_n82 & ~new_n243;
  assign new_n246 = ~new_n244 & ~new_n245;
  assign new_n247 = ~\13  & ~\61 ;
  assign new_n248 = \13  & \61 ;
  assign new_n249 = ~new_n247 & ~new_n248;
  assign new_n250 = new_n229 & new_n249;
  assign new_n251 = ~new_n229 & ~new_n249;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253 = \29  & ~\45 ;
  assign new_n254 = ~\29  & \45 ;
  assign new_n255 = ~new_n253 & ~new_n254;
  assign new_n256 = new_n252 & ~new_n255;
  assign new_n257 = ~new_n252 & new_n255;
  assign new_n258 = ~new_n256 & ~new_n257;
  assign new_n259 = new_n246 & new_n258;
  assign new_n260 = ~new_n246 & ~new_n258;
  assign new_n261 = ~new_n259 & ~new_n260;
  assign new_n262 = ~new_n242 & new_n261;
  assign new_n263 = ~new_n214 & ~new_n262;
  assign new_n264 = new_n242 & ~new_n261;
  assign new_n265 = ~new_n262 & ~new_n264;
  assign new_n266 = new_n214 & ~new_n265;
  assign new_n267 = ~new_n110 & ~new_n213;
  assign new_n268 = ~new_n263 & ~new_n267;
  assign new_n269 = ~new_n266 & new_n268;
  assign new_n270 = new_n185 & new_n269;
  assign new_n271 = \133  & \137 ;
  assign new_n272 = ~new_n132 & new_n271;
  assign new_n273 = new_n132 & ~new_n271;
  assign new_n274 = ~new_n272 & ~new_n273;
  assign new_n275 = ~\65  & ~\81 ;
  assign new_n276 = \65  & \81 ;
  assign new_n277 = ~new_n275 & ~new_n276;
  assign new_n278 = new_n156 & new_n277;
  assign new_n279 = ~new_n156 & ~new_n277;
  assign new_n280 = ~new_n278 & ~new_n279;
  assign new_n281 = \97  & ~\113 ;
  assign new_n282 = ~\97  & \113 ;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = new_n280 & ~new_n283;
  assign new_n285 = ~new_n280 & new_n283;
  assign new_n286 = ~new_n284 & ~new_n285;
  assign new_n287 = new_n274 & new_n286;
  assign new_n288 = ~new_n274 & ~new_n286;
  assign new_n289 = ~new_n287 & ~new_n288;
  assign new_n290 = \134  & \137 ;
  assign new_n291 = ~new_n119 & new_n290;
  assign new_n292 = new_n119 & ~new_n290;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294 = ~\69  & ~\85 ;
  assign new_n295 = \69  & \85 ;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = new_n169 & new_n296;
  assign new_n298 = ~new_n169 & ~new_n296;
  assign new_n299 = ~new_n297 & ~new_n298;
  assign new_n300 = \101  & ~\117 ;
  assign new_n301 = ~\101  & \117 ;
  assign new_n302 = ~new_n300 & ~new_n301;
  assign new_n303 = new_n299 & ~new_n302;
  assign new_n304 = ~new_n299 & new_n302;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = new_n293 & new_n305;
  assign new_n307 = ~new_n293 & ~new_n305;
  assign new_n308 = ~new_n306 & ~new_n307;
  assign new_n309 = ~new_n289 & new_n308;
  assign new_n310 = new_n270 & new_n309;
  assign new_n311 = ~new_n110 & new_n310;
  assign new_n312 = \1  & ~new_n311;
  assign new_n313 = ~\1  & new_n311;
  assign \724  = new_n312 | new_n313;
  assign new_n315 = new_n242 & new_n310;
  assign new_n316 = \5  & ~new_n315;
  assign new_n317 = ~\5  & new_n315;
  assign \725  = new_n316 | new_n317;
  assign new_n319 = ~new_n213 & new_n310;
  assign new_n320 = \9  & ~new_n319;
  assign new_n321 = ~\9  & new_n319;
  assign \726  = new_n320 | new_n321;
  assign new_n323 = ~new_n261 & new_n310;
  assign new_n324 = \13  & ~new_n323;
  assign new_n325 = ~\13  & new_n323;
  assign \727  = new_n324 | new_n325;
  assign new_n327 = ~new_n147 & new_n184;
  assign new_n328 = new_n269 & new_n327;
  assign new_n329 = new_n309 & new_n328;
  assign new_n330 = ~new_n110 & new_n329;
  assign new_n331 = \17  & ~new_n330;
  assign new_n332 = ~\17  & new_n330;
  assign \728  = new_n331 | new_n332;
  assign new_n334 = new_n242 & new_n329;
  assign new_n335 = \21  & ~new_n334;
  assign new_n336 = ~\21  & new_n334;
  assign \729  = new_n335 | new_n336;
  assign new_n338 = ~new_n213 & new_n329;
  assign new_n339 = \25  & ~new_n338;
  assign new_n340 = ~\25  & new_n338;
  assign \730  = new_n339 | new_n340;
  assign new_n342 = ~new_n261 & new_n329;
  assign new_n343 = \29  & ~new_n342;
  assign new_n344 = ~\29  & new_n342;
  assign \731  = new_n343 | new_n344;
  assign new_n346 = new_n289 & ~new_n308;
  assign new_n347 = new_n270 & new_n346;
  assign new_n348 = ~new_n110 & new_n347;
  assign new_n349 = \33  & ~new_n348;
  assign new_n350 = ~\33  & new_n348;
  assign \732  = new_n349 | new_n350;
  assign new_n352 = new_n242 & new_n347;
  assign new_n353 = \37  & ~new_n352;
  assign new_n354 = ~\37  & new_n352;
  assign \733  = new_n353 | new_n354;
  assign new_n356 = ~new_n213 & new_n347;
  assign new_n357 = \41  & ~new_n356;
  assign new_n358 = ~\41  & new_n356;
  assign \734  = new_n357 | new_n358;
  assign new_n360 = ~new_n261 & new_n347;
  assign new_n361 = \45  & ~new_n360;
  assign new_n362 = ~\45  & new_n360;
  assign \735  = new_n361 | new_n362;
  assign new_n364 = new_n328 & new_n346;
  assign new_n365 = ~new_n110 & new_n364;
  assign new_n366 = \49  & ~new_n365;
  assign new_n367 = ~\49  & new_n365;
  assign \736  = new_n366 | new_n367;
  assign new_n369 = new_n242 & new_n364;
  assign new_n370 = \53  & ~new_n369;
  assign new_n371 = ~\53  & new_n369;
  assign \737  = new_n370 | new_n371;
  assign new_n373 = ~new_n213 & new_n364;
  assign new_n374 = \57  & ~new_n373;
  assign new_n375 = ~\57  & new_n373;
  assign \738  = new_n374 | new_n375;
  assign new_n377 = ~new_n261 & new_n364;
  assign new_n378 = \61  & ~new_n377;
  assign new_n379 = ~\61  & new_n377;
  assign \739  = new_n378 | new_n379;
  assign new_n381 = ~new_n213 & new_n261;
  assign new_n382 = ~new_n185 & ~new_n327;
  assign new_n383 = new_n289 & new_n308;
  assign new_n384 = ~new_n382 & new_n383;
  assign new_n385 = ~new_n309 & ~new_n346;
  assign new_n386 = new_n147 & new_n184;
  assign new_n387 = ~new_n385 & new_n386;
  assign new_n388 = ~new_n384 & ~new_n387;
  assign new_n389 = ~new_n110 & ~new_n242;
  assign new_n390 = ~new_n388 & new_n389;
  assign new_n391 = new_n381 & new_n390;
  assign new_n392 = ~new_n289 & new_n391;
  assign new_n393 = \65  & ~new_n392;
  assign new_n394 = ~\65  & new_n392;
  assign \740  = new_n393 | new_n394;
  assign new_n396 = ~new_n308 & new_n391;
  assign new_n397 = \69  & ~new_n396;
  assign new_n398 = ~\69  & new_n396;
  assign \741  = new_n397 | new_n398;
  assign new_n400 = ~new_n184 & new_n391;
  assign new_n401 = \73  & ~new_n400;
  assign new_n402 = ~\73  & new_n400;
  assign \742  = new_n401 | new_n402;
  assign new_n404 = ~new_n147 & new_n391;
  assign new_n405 = \77  & ~new_n404;
  assign new_n406 = ~\77  & new_n404;
  assign \743  = new_n405 | new_n406;
  assign new_n408 = new_n213 & ~new_n261;
  assign new_n409 = new_n390 & new_n408;
  assign new_n410 = ~new_n289 & new_n409;
  assign new_n411 = \81  & ~new_n410;
  assign new_n412 = ~\81  & new_n410;
  assign \744  = new_n411 | new_n412;
  assign new_n414 = ~new_n308 & new_n409;
  assign new_n415 = \85  & ~new_n414;
  assign new_n416 = ~\85  & new_n414;
  assign \745  = new_n415 | new_n416;
  assign new_n418 = ~new_n184 & new_n409;
  assign new_n419 = \89  & ~new_n418;
  assign new_n420 = ~\89  & new_n418;
  assign \746  = new_n419 | new_n420;
  assign new_n422 = ~new_n147 & new_n409;
  assign new_n423 = \93  & ~new_n422;
  assign new_n424 = ~\93  & new_n422;
  assign \747  = new_n423 | new_n424;
  assign new_n426 = new_n110 & new_n242;
  assign new_n427 = ~new_n388 & new_n426;
  assign new_n428 = new_n381 & new_n427;
  assign new_n429 = ~new_n289 & new_n428;
  assign new_n430 = \97  & ~new_n429;
  assign new_n431 = ~\97  & new_n429;
  assign \748  = new_n430 | new_n431;
  assign new_n433 = ~new_n308 & new_n428;
  assign new_n434 = \101  & ~new_n433;
  assign new_n435 = ~\101  & new_n433;
  assign \749  = new_n434 | new_n435;
  assign new_n437 = ~new_n184 & new_n428;
  assign new_n438 = \105  & ~new_n437;
  assign new_n439 = ~\105  & new_n437;
  assign \750  = new_n438 | new_n439;
  assign new_n441 = ~new_n147 & new_n428;
  assign new_n442 = \109  & ~new_n441;
  assign new_n443 = ~\109  & new_n441;
  assign \751  = new_n442 | new_n443;
  assign new_n445 = new_n408 & new_n427;
  assign new_n446 = ~new_n289 & new_n445;
  assign new_n447 = \113  & ~new_n446;
  assign new_n448 = ~\113  & new_n446;
  assign \752  = new_n447 | new_n448;
  assign new_n450 = ~new_n308 & new_n445;
  assign new_n451 = \117  & ~new_n450;
  assign new_n452 = ~\117  & new_n450;
  assign \753  = new_n451 | new_n452;
  assign new_n454 = ~new_n184 & new_n445;
  assign new_n455 = \121  & ~new_n454;
  assign new_n456 = ~\121  & new_n454;
  assign \754  = new_n455 | new_n456;
  assign new_n458 = ~new_n147 & new_n445;
  assign new_n459 = \125  & ~new_n458;
  assign new_n460 = ~\125  & new_n458;
  assign \755  = new_n459 | new_n460;
endmodule


