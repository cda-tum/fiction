// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pt, pu, pv, pw, px, py, pz, pa, pb, pc,
    pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    pd0, pe0, pf0  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pt, pu, pv, pw, px, py, pz, pa,
    pb, pc, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po;
  output pd0, pe0, pf0;
  wire new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38,
    new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46,
    new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53, new_n54,
    new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61, new_n62,
    new_n63, new_n64, new_n65, new_n66, new_n67, new_n68, new_n69, new_n70,
    new_n71, new_n72, new_n73, new_n74, new_n75, new_n76, new_n77, new_n78,
    new_n79, new_n80, new_n81, new_n82, new_n83, new_n84, new_n85, new_n86,
    new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93, new_n94,
    new_n95, new_n96, new_n97, new_n98, new_n99, new_n100, new_n101,
    new_n102, new_n103, new_n104, new_n105, new_n106, new_n107, new_n108,
    new_n109, new_n110, new_n111, new_n112, new_n113, new_n114, new_n115,
    new_n116, new_n117, new_n118, new_n119, new_n120, new_n121, new_n122,
    new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689;
  assign new_n32 = pe & ~pi;
  assign new_n33 = ~pj & new_n32;
  assign new_n34 = ~pc & new_n33;
  assign new_n35 = ~pi & ~pj;
  assign new_n36 = pa & new_n35;
  assign new_n37 = ~pc & new_n36;
  assign new_n38 = ~pq & ~pv;
  assign new_n39 = pe & new_n38;
  assign new_n40 = ~pr & new_n39;
  assign new_n41 = ~pc & new_n40;
  assign new_n42 = ~pm & new_n41;
  assign new_n43 = ~pu & new_n42;
  assign new_n44 = ~ps & new_n43;
  assign new_n45 = ~pt & new_n44;
  assign new_n46 = ~po & new_n45;
  assign new_n47 = ~pp & new_n46;
  assign new_n48 = pe & ~pg;
  assign new_n49 = ~ph & new_n48;
  assign new_n50 = ~pc & new_n49;
  assign new_n51 = ~pq & pa;
  assign new_n52 = ~pr & new_n51;
  assign new_n53 = ~pv & new_n52;
  assign new_n54 = ~pc & new_n53;
  assign new_n55 = ~pm & new_n54;
  assign new_n56 = ~pu & new_n55;
  assign new_n57 = ~ps & new_n56;
  assign new_n58 = ~pt & new_n57;
  assign new_n59 = ~po & new_n58;
  assign new_n60 = ~pp & new_n59;
  assign new_n61 = pa & ~ph;
  assign new_n62 = ~pg & new_n61;
  assign new_n63 = ~pc & new_n62;
  assign new_n64 = ~pz & ~pk;
  assign new_n65 = pe & new_n64;
  assign new_n66 = ~pr & new_n65;
  assign new_n67 = ~pc & new_n66;
  assign new_n68 = ~px & new_n67;
  assign new_n69 = ~pw & new_n68;
  assign new_n70 = ~po & new_n69;
  assign new_n71 = ~pp & new_n70;
  assign new_n72 = ~pq & new_n71;
  assign new_n73 = ~py & new_n72;
  assign new_n74 = ~pq & ~pk;
  assign new_n75 = ~pr & new_n74;
  assign new_n76 = ~pz & new_n75;
  assign new_n77 = ~pc & new_n76;
  assign new_n78 = ~px & new_n77;
  assign new_n79 = ~pw & new_n78;
  assign new_n80 = ~po & new_n79;
  assign new_n81 = ~pp & new_n80;
  assign new_n82 = ~py & new_n81;
  assign new_n83 = pa & new_n82;
  assign new_n84 = ~pb & pc;
  assign new_n85 = ~pr & ~pv;
  assign new_n86 = pe & new_n85;
  assign new_n87 = ~ph & new_n86;
  assign new_n88 = ~pc & new_n87;
  assign new_n89 = ~px & new_n88;
  assign new_n90 = ~ps & new_n89;
  assign new_n91 = ~pt & new_n90;
  assign new_n92 = ~pz & new_n91;
  assign new_n93 = ~pp & new_n92;
  assign new_n94 = ~pv & ~pz;
  assign new_n95 = ~ph & new_n94;
  assign new_n96 = ~pr & new_n95;
  assign new_n97 = ~pc & new_n96;
  assign new_n98 = ~px & new_n97;
  assign new_n99 = ~ps & new_n98;
  assign new_n100 = ~pt & new_n99;
  assign new_n101 = pa & new_n100;
  assign new_n102 = ~pp & new_n101;
  assign new_n103 = ~pp & ~ps;
  assign new_n104 = pe & new_n103;
  assign new_n105 = ~po & new_n104;
  assign new_n106 = ~pc & new_n105;
  assign new_n107 = ~px & new_n106;
  assign new_n108 = ~pi & new_n107;
  assign new_n109 = ~pt & new_n108;
  assign new_n110 = ~pw & new_n109;
  assign new_n111 = ~pq & ~py;
  assign new_n112 = ~pj & new_n111;
  assign new_n113 = ~pg & new_n112;
  assign new_n114 = ~pc & new_n113;
  assign new_n115 = pa & new_n114;
  assign new_n116 = ~pu & new_n115;
  assign new_n117 = ~px & ~pi;
  assign new_n118 = pe & new_n117;
  assign new_n119 = ~ph & new_n118;
  assign new_n120 = ~pc & new_n119;
  assign new_n121 = ~pn & new_n120;
  assign new_n122 = ~py & ~pz;
  assign new_n123 = pe & new_n122;
  assign new_n124 = ~pj & new_n123;
  assign new_n125 = ~pc & new_n124;
  assign new_n126 = ~pn & new_n125;
  assign new_n127 = ~pw & ~po;
  assign new_n128 = pe & new_n127;
  assign new_n129 = ~pg & new_n128;
  assign new_n130 = ~pc & new_n129;
  assign new_n131 = ~pi & new_n130;
  assign new_n132 = pa & new_n103;
  assign new_n133 = ~po & new_n132;
  assign new_n134 = ~pc & new_n133;
  assign new_n135 = ~px & new_n134;
  assign new_n136 = ~pi & new_n135;
  assign new_n137 = ~pt & new_n136;
  assign new_n138 = ~pw & new_n137;
  assign new_n139 = ~pq & ~pg;
  assign new_n140 = pe & new_n139;
  assign new_n141 = ~pj & new_n140;
  assign new_n142 = ~pc & new_n141;
  assign new_n143 = ~py & new_n142;
  assign new_n144 = ~pu & new_n143;
  assign new_n145 = ~ph & new_n117;
  assign new_n146 = pa & new_n145;
  assign new_n147 = ~pc & new_n146;
  assign new_n148 = ~pn & new_n147;
  assign new_n149 = ~pz & ~pj;
  assign new_n150 = pe & new_n149;
  assign new_n151 = ~ph & new_n150;
  assign new_n152 = ~pc & new_n151;
  assign new_n153 = ~pn & new_n152;
  assign new_n154 = ~pg & new_n127;
  assign new_n155 = pa & new_n154;
  assign new_n156 = ~pc & new_n155;
  assign new_n157 = ~pi & new_n156;
  assign new_n158 = ~pq & ~pz;
  assign new_n159 = ~pr & new_n158;
  assign new_n160 = ~pv & new_n159;
  assign new_n161 = ~pc & new_n160;
  assign new_n162 = ~pw & new_n161;
  assign new_n163 = ~px & new_n162;
  assign new_n164 = ~pt & new_n163;
  assign new_n165 = ~pu & new_n164;
  assign new_n166 = ~ps & new_n165;
  assign new_n167 = ~po & new_n166;
  assign new_n168 = ~pp & new_n167;
  assign new_n169 = ~py & new_n168;
  assign new_n170 = pa & new_n169;
  assign new_n171 = ~pt & new_n88;
  assign new_n172 = ~pm & new_n171;
  assign new_n173 = ~pp & new_n172;
  assign new_n174 = ~ps & new_n173;
  assign new_n175 = ~ph & new_n104;
  assign new_n176 = ~pc & new_n175;
  assign new_n177 = ~pi & new_n176;
  assign new_n178 = ~pt & new_n177;
  assign new_n179 = ~px & new_n178;
  assign new_n180 = ~pj & new_n74;
  assign new_n181 = ~pg & new_n180;
  assign new_n182 = ~pc & new_n181;
  assign new_n183 = ~py & new_n182;
  assign new_n184 = pa & new_n183;
  assign new_n185 = ~pw & ~pi;
  assign new_n186 = pe & new_n185;
  assign new_n187 = ~pg & new_n186;
  assign new_n188 = ~pc & new_n187;
  assign new_n189 = ~pn & new_n188;
  assign new_n190 = ~pz & pa;
  assign new_n191 = ~ph & new_n190;
  assign new_n192 = ~pj & new_n191;
  assign new_n193 = ~pc & new_n192;
  assign new_n194 = ~pn & new_n193;
  assign new_n195 = ~pm & ~po;
  assign new_n196 = pe & new_n195;
  assign new_n197 = ~pg & new_n196;
  assign new_n198 = ~pc & new_n197;
  assign new_n199 = ~pi & new_n198;
  assign new_n200 = pe & new_n94;
  assign new_n201 = ~pr & new_n200;
  assign new_n202 = ~pc & new_n201;
  assign new_n203 = ~pw & new_n202;
  assign new_n204 = ~px & new_n203;
  assign new_n205 = ~pt & new_n204;
  assign new_n206 = ~pu & new_n205;
  assign new_n207 = ~ps & new_n206;
  assign new_n208 = ~po & new_n207;
  assign new_n209 = ~pp & new_n208;
  assign new_n210 = ~pq & new_n209;
  assign new_n211 = ~py & new_n210;
  assign new_n212 = ~pv & pa;
  assign new_n213 = ~ph & new_n212;
  assign new_n214 = ~pr & new_n213;
  assign new_n215 = ~pc & new_n214;
  assign new_n216 = ~pt & new_n215;
  assign new_n217 = ~pm & new_n216;
  assign new_n218 = ~pp & new_n217;
  assign new_n219 = ~ps & new_n218;
  assign new_n220 = ~ph & new_n103;
  assign new_n221 = pa & new_n220;
  assign new_n222 = ~pc & new_n221;
  assign new_n223 = ~pi & new_n222;
  assign new_n224 = ~pt & new_n223;
  assign new_n225 = ~px & new_n224;
  assign new_n226 = ~pr & ~pz;
  assign new_n227 = ~ph & new_n226;
  assign new_n228 = ~pj & new_n227;
  assign new_n229 = ~pc & new_n228;
  assign new_n230 = ~pk & new_n229;
  assign new_n231 = pa & new_n230;
  assign new_n232 = ~pg & new_n185;
  assign new_n233 = pa & new_n232;
  assign new_n234 = ~pc & new_n233;
  assign new_n235 = ~pn & new_n234;
  assign new_n236 = ~py & ~pg;
  assign new_n237 = pe & new_n236;
  assign new_n238 = ~pj & new_n237;
  assign new_n239 = ~pc & new_n238;
  assign new_n240 = ~pn & new_n239;
  assign new_n241 = ~pg & new_n195;
  assign new_n242 = pa & new_n241;
  assign new_n243 = ~pc & new_n242;
  assign new_n244 = ~pi & new_n243;
  assign new_n245 = ~pg & new_n111;
  assign new_n246 = ~pk & new_n245;
  assign new_n247 = ~pc & new_n246;
  assign new_n248 = ~pw & new_n247;
  assign new_n249 = pa & new_n248;
  assign new_n250 = ~po & new_n249;
  assign new_n251 = ~pp & ~po;
  assign new_n252 = pe & new_n251;
  assign new_n253 = ~pk & new_n252;
  assign new_n254 = ~pc & new_n253;
  assign new_n255 = ~pm & new_n254;
  assign new_n256 = ~pi & new_n255;
  assign new_n257 = ~ph & new_n85;
  assign new_n258 = ~pj & new_n257;
  assign new_n259 = ~pc & new_n258;
  assign new_n260 = ~pz & new_n259;
  assign new_n261 = pa & new_n260;
  assign new_n262 = ~px & ~pz;
  assign new_n263 = pe & new_n262;
  assign new_n264 = ~ph & new_n263;
  assign new_n265 = ~pc & new_n264;
  assign new_n266 = ~pn & new_n265;
  assign new_n267 = ~pu & pa;
  assign new_n268 = ~pj & new_n267;
  assign new_n269 = ~pv & new_n268;
  assign new_n270 = ~pc & new_n269;
  assign new_n271 = ~pl & new_n270;
  assign new_n272 = ~pu & ~pl;
  assign new_n273 = pe & new_n272;
  assign new_n274 = ~pg & new_n273;
  assign new_n275 = ~pc & new_n274;
  assign new_n276 = pe & new_n74;
  assign new_n277 = ~pg & new_n276;
  assign new_n278 = ~pc & new_n277;
  assign new_n279 = ~pw & new_n278;
  assign new_n280 = ~py & new_n279;
  assign new_n281 = ~po & new_n280;
  assign new_n282 = ~pk & new_n251;
  assign new_n283 = pa & new_n282;
  assign new_n284 = ~pc & new_n283;
  assign new_n285 = ~pm & new_n284;
  assign new_n286 = ~pi & new_n285;
  assign new_n287 = ~pg & ~pk;
  assign new_n288 = pe & new_n287;
  assign new_n289 = ~pj & new_n288;
  assign new_n290 = ~pc & new_n289;
  assign new_n291 = ~pq & new_n290;
  assign new_n292 = ~py & new_n291;
  assign new_n293 = ~px & pa;
  assign new_n294 = ~ph & new_n293;
  assign new_n295 = ~pz & new_n294;
  assign new_n296 = ~pc & new_n295;
  assign new_n297 = ~pn & new_n296;
  assign new_n298 = ~pu & ~pv;
  assign new_n299 = pe & new_n298;
  assign new_n300 = ~pj & new_n299;
  assign new_n301 = ~pc & new_n300;
  assign new_n302 = ~pl & new_n301;
  assign new_n303 = ~pg & new_n272;
  assign new_n304 = pa & new_n303;
  assign new_n305 = ~pc & new_n304;
  assign new_n306 = pa & ~pk;
  assign new_n307 = ~ph & new_n306;
  assign new_n308 = ~pr & new_n307;
  assign new_n309 = ~pc & new_n308;
  assign new_n310 = ~pp & new_n309;
  assign new_n311 = ~pm & new_n310;
  assign new_n312 = ~pr & ~pj;
  assign new_n313 = pe & new_n312;
  assign new_n314 = ~ph & new_n313;
  assign new_n315 = ~pc & new_n314;
  assign new_n316 = ~pv & new_n315;
  assign new_n317 = ~pm & new_n316;
  assign new_n318 = ~pz & new_n315;
  assign new_n319 = ~pk & new_n318;
  assign new_n320 = ~pw & ~py;
  assign new_n321 = pe & new_n320;
  assign new_n322 = ~pg & new_n321;
  assign new_n323 = ~pc & new_n322;
  assign new_n324 = ~pn & new_n323;
  assign new_n325 = ~pt & ~pi;
  assign new_n326 = pa & new_n325;
  assign new_n327 = ~ps & new_n326;
  assign new_n328 = ~pc & new_n327;
  assign new_n329 = ~pl & new_n328;
  assign new_n330 = ~pi & ~pl;
  assign new_n331 = pe & new_n330;
  assign new_n332 = ~pg & new_n331;
  assign new_n333 = ~pc & new_n332;
  assign new_n334 = ~pr & ~pk;
  assign new_n335 = pe & new_n334;
  assign new_n336 = ~ph & new_n335;
  assign new_n337 = ~pc & new_n336;
  assign new_n338 = ~pp & new_n337;
  assign new_n339 = ~pm & new_n338;
  assign new_n340 = ~pk & new_n315;
  assign new_n341 = ~pm & new_n340;
  assign new_n342 = ~pz & new_n316;
  assign new_n343 = ~pw & pa;
  assign new_n344 = ~pg & new_n343;
  assign new_n345 = ~py & new_n344;
  assign new_n346 = ~pc & new_n345;
  assign new_n347 = ~pn & new_n346;
  assign new_n348 = pe & new_n325;
  assign new_n349 = ~ps & new_n348;
  assign new_n350 = ~pc & new_n349;
  assign new_n351 = ~pl & new_n350;
  assign new_n352 = ~pg & new_n330;
  assign new_n353 = pa & new_n352;
  assign new_n354 = ~pc & new_n353;
  assign new_n355 = ~pi & new_n106;
  assign new_n356 = ~pt & new_n355;
  assign new_n357 = ~pm & new_n356;
  assign new_n358 = ~ph & new_n64;
  assign new_n359 = ~pr & new_n358;
  assign new_n360 = ~pc & new_n359;
  assign new_n361 = ~px & new_n360;
  assign new_n362 = pa & new_n361;
  assign new_n363 = ~pp & new_n362;
  assign new_n364 = ~ps & ~pt;
  assign new_n365 = pe & new_n364;
  assign new_n366 = ~pv & new_n365;
  assign new_n367 = ~pc & new_n366;
  assign new_n368 = ~pu & new_n367;
  assign new_n369 = ~pl & new_n368;
  assign new_n370 = ~pj & new_n51;
  assign new_n371 = ~pg & new_n370;
  assign new_n372 = ~pc & new_n371;
  assign new_n373 = ~pu & new_n372;
  assign new_n374 = ~pm & new_n373;
  assign new_n375 = ~pj & new_n335;
  assign new_n376 = ~pc & new_n375;
  assign new_n377 = ~pq & new_n376;
  assign new_n378 = ~pm & new_n377;
  assign new_n379 = pa & new_n117;
  assign new_n380 = ~pw & new_n379;
  assign new_n381 = ~pc & new_n380;
  assign new_n382 = ~pn & new_n381;
  assign new_n383 = ~py & pa;
  assign new_n384 = ~pj & new_n383;
  assign new_n385 = ~pz & new_n384;
  assign new_n386 = ~pc & new_n385;
  assign new_n387 = ~pn & new_n386;
  assign new_n388 = ~pi & new_n134;
  assign new_n389 = ~pt & new_n388;
  assign new_n390 = ~pm & new_n389;
  assign new_n391 = pe & new_n226;
  assign new_n392 = ~ph & new_n391;
  assign new_n393 = ~pc & new_n392;
  assign new_n394 = ~px & new_n393;
  assign new_n395 = ~pk & new_n394;
  assign new_n396 = ~pp & new_n395;
  assign new_n397 = ~pv & new_n364;
  assign new_n398 = pa & new_n397;
  assign new_n399 = ~pc & new_n398;
  assign new_n400 = ~pu & new_n399;
  assign new_n401 = ~pl & new_n400;
  assign new_n402 = ~pu & new_n142;
  assign new_n403 = ~pm & new_n402;
  assign new_n404 = ~pm & new_n291;
  assign new_n405 = ~pw & new_n118;
  assign new_n406 = ~pc & new_n405;
  assign new_n407 = ~pn & new_n406;
  assign new_n408 = ~pg & new_n384;
  assign new_n409 = ~pc & new_n408;
  assign new_n410 = ~pn & new_n409;
  assign new_n411 = ~pj & new_n86;
  assign new_n412 = ~pc & new_n411;
  assign new_n413 = ~py & new_n412;
  assign new_n414 = ~pu & new_n413;
  assign new_n415 = ~pz & new_n414;
  assign new_n416 = ~pq & new_n415;
  assign new_n417 = ~pg & new_n383;
  assign new_n418 = ~pq & new_n417;
  assign new_n419 = ~pc & new_n418;
  assign new_n420 = ~pw & new_n419;
  assign new_n421 = ~po & new_n420;
  assign new_n422 = ~pu & new_n421;
  assign new_n423 = ~ps & ~pv;
  assign new_n424 = pe & new_n423;
  assign new_n425 = ~ph & new_n424;
  assign new_n426 = ~pc & new_n425;
  assign new_n427 = ~pt & new_n426;
  assign new_n428 = ~pl & new_n427;
  assign new_n429 = pa & ~po;
  assign new_n430 = ~pg & new_n429;
  assign new_n431 = ~pq & new_n430;
  assign new_n432 = ~pc & new_n431;
  assign new_n433 = ~pu & new_n432;
  assign new_n434 = ~pm & new_n433;
  assign new_n435 = pa & new_n259;
  assign new_n436 = ~pm & new_n435;
  assign new_n437 = ~pj & new_n213;
  assign new_n438 = ~pc & new_n437;
  assign new_n439 = ~pl & new_n438;
  assign new_n440 = pa & ~pn;
  assign new_n441 = ~pl & new_n440;
  assign new_n442 = ~pc & new_n441;
  assign new_n443 = ~pj & new_n94;
  assign new_n444 = ~pr & new_n443;
  assign new_n445 = ~pc & new_n444;
  assign new_n446 = pa & new_n445;
  assign new_n447 = ~pu & new_n446;
  assign new_n448 = ~pq & new_n447;
  assign new_n449 = ~py & new_n448;
  assign new_n450 = pe & new_n111;
  assign new_n451 = ~pg & new_n450;
  assign new_n452 = ~pc & new_n451;
  assign new_n453 = ~pw & new_n452;
  assign new_n454 = ~po & new_n453;
  assign new_n455 = ~pu & new_n454;
  assign new_n456 = ~ps & pa;
  assign new_n457 = ~ph & new_n456;
  assign new_n458 = ~pv & new_n457;
  assign new_n459 = ~pc & new_n458;
  assign new_n460 = ~pt & new_n459;
  assign new_n461 = ~pl & new_n460;
  assign new_n462 = ~pq & ~po;
  assign new_n463 = pe & new_n462;
  assign new_n464 = ~pg & new_n463;
  assign new_n465 = ~pc & new_n464;
  assign new_n466 = ~pu & new_n465;
  assign new_n467 = ~pm & new_n466;
  assign new_n468 = ~ph & new_n334;
  assign new_n469 = ~pj & new_n468;
  assign new_n470 = ~pc & new_n469;
  assign new_n471 = pa & new_n470;
  assign new_n472 = ~pm & new_n471;
  assign new_n473 = ~pv & ~pj;
  assign new_n474 = pe & new_n473;
  assign new_n475 = ~ph & new_n474;
  assign new_n476 = ~pc & new_n475;
  assign new_n477 = ~pl & new_n476;
  assign new_n478 = ~pc0 & ~pe;
  assign new_n479 = ~pa & new_n478;
  assign new_n480 = ~pc & new_n479;
  assign new_n481 = ~pi & new_n254;
  assign new_n482 = ~pw & new_n481;
  assign new_n483 = ~px & new_n482;
  assign new_n484 = ~pj & new_n38;
  assign new_n485 = ~pr & new_n484;
  assign new_n486 = ~pc & new_n485;
  assign new_n487 = ~pm & new_n486;
  assign new_n488 = pa & new_n487;
  assign new_n489 = ~pu & new_n488;
  assign new_n490 = ~pj & new_n391;
  assign new_n491 = ~pc & new_n490;
  assign new_n492 = ~py & new_n491;
  assign new_n493 = ~pk & new_n492;
  assign new_n494 = ~pq & new_n493;
  assign new_n495 = ~pp & pa;
  assign new_n496 = ~ph & new_n495;
  assign new_n497 = ~pk & new_n496;
  assign new_n498 = ~pc & new_n497;
  assign new_n499 = ~px & new_n498;
  assign new_n500 = ~pi & new_n499;
  assign new_n501 = ~pr & new_n180;
  assign new_n502 = ~pc & new_n501;
  assign new_n503 = pa & new_n502;
  assign new_n504 = ~pm & new_n503;
  assign new_n505 = ~pi & new_n284;
  assign new_n506 = ~pw & new_n505;
  assign new_n507 = ~px & new_n506;
  assign new_n508 = ~pm & new_n412;
  assign new_n509 = ~pq & new_n508;
  assign new_n510 = ~pu & new_n509;
  assign new_n511 = ~pj & new_n64;
  assign new_n512 = ~pr & new_n511;
  assign new_n513 = ~pc & new_n512;
  assign new_n514 = pa & new_n513;
  assign new_n515 = ~pq & new_n514;
  assign new_n516 = ~py & new_n515;
  assign new_n517 = ~pp & ~pk;
  assign new_n518 = pe & new_n517;
  assign new_n519 = ~ph & new_n518;
  assign new_n520 = ~pc & new_n519;
  assign new_n521 = ~px & new_n520;
  assign new_n522 = ~pi & new_n521;
  assign new_n523 = pa & new_n182;
  assign new_n524 = ~pm & new_n523;
  assign new_n525 = ~pm & new_n178;
  assign new_n526 = ~pk & new_n52;
  assign new_n527 = ~pc & new_n526;
  assign new_n528 = ~pm & new_n527;
  assign new_n529 = ~po & new_n528;
  assign new_n530 = ~pp & new_n529;
  assign new_n531 = ~pz & new_n321;
  assign new_n532 = ~pc & new_n531;
  assign new_n533 = ~px & new_n532;
  assign new_n534 = ~pn & new_n533;
  assign new_n535 = ~pm & new_n498;
  assign new_n536 = ~pi & new_n535;
  assign new_n537 = ~po & new_n278;
  assign new_n538 = ~pm & new_n537;
  assign new_n539 = ~pm & new_n224;
  assign new_n540 = ~pr & new_n276;
  assign new_n541 = ~pc & new_n540;
  assign new_n542 = ~pm & new_n541;
  assign new_n543 = ~po & new_n542;
  assign new_n544 = ~pp & new_n543;
  assign new_n545 = ~pz & new_n343;
  assign new_n546 = ~py & new_n545;
  assign new_n547 = ~pc & new_n546;
  assign new_n548 = ~px & new_n547;
  assign new_n549 = ~pn & new_n548;
  assign new_n550 = ~pm & new_n520;
  assign new_n551 = ~pi & new_n550;
  assign new_n552 = ~pg & new_n51;
  assign new_n553 = ~pk & new_n552;
  assign new_n554 = ~pc & new_n553;
  assign new_n555 = ~po & new_n554;
  assign new_n556 = ~pm & new_n555;
  assign new_n557 = pe & ~pn;
  assign new_n558 = ~pl & new_n557;
  assign new_n559 = ~pc & new_n558;
  assign new_n560 = ~pm & new_n557;
  assign new_n561 = ~pc & new_n560;
  assign new_n562 = ~pm & new_n440;
  assign new_n563 = ~pc & new_n562;
  assign new_n564 = pe & ~pl;
  assign new_n565 = ~pk & new_n564;
  assign new_n566 = ~pc & new_n565;
  assign new_n567 = ~pk & ~pl;
  assign new_n568 = pa & new_n567;
  assign new_n569 = ~pc & new_n568;
  assign new_n570 = ~new_n563 & ~new_n566;
  assign new_n571 = ~new_n569 & new_n570;
  assign new_n572 = ~new_n559 & ~new_n561;
  assign new_n573 = ~new_n551 & ~new_n556;
  assign new_n574 = new_n572 & new_n573;
  assign new_n575 = new_n571 & new_n574;
  assign new_n576 = ~new_n539 & ~new_n544;
  assign new_n577 = ~new_n549 & new_n576;
  assign new_n578 = ~new_n536 & ~new_n538;
  assign new_n579 = ~new_n530 & ~new_n534;
  assign new_n580 = new_n578 & new_n579;
  assign new_n581 = new_n577 & new_n580;
  assign new_n582 = new_n575 & new_n581;
  assign new_n583 = ~new_n522 & ~new_n524;
  assign new_n584 = ~new_n525 & new_n583;
  assign new_n585 = ~new_n510 & ~new_n516;
  assign new_n586 = ~new_n504 & ~new_n507;
  assign new_n587 = new_n585 & new_n586;
  assign new_n588 = new_n584 & new_n587;
  assign new_n589 = ~new_n489 & ~new_n494;
  assign new_n590 = ~new_n500 & new_n589;
  assign new_n591 = ~new_n480 & ~new_n483;
  assign new_n592 = ~new_n472 & ~new_n477;
  assign new_n593 = new_n591 & new_n592;
  assign new_n594 = new_n590 & new_n593;
  assign new_n595 = new_n588 & new_n594;
  assign new_n596 = new_n582 & new_n595;
  assign new_n597 = ~new_n455 & ~new_n461;
  assign new_n598 = ~new_n467 & new_n597;
  assign new_n599 = ~new_n442 & ~new_n449;
  assign new_n600 = ~new_n436 & ~new_n439;
  assign new_n601 = new_n599 & new_n600;
  assign new_n602 = new_n598 & new_n601;
  assign new_n603 = ~new_n422 & ~new_n428;
  assign new_n604 = ~new_n434 & new_n603;
  assign new_n605 = ~new_n410 & ~new_n416;
  assign new_n606 = ~new_n404 & ~new_n407;
  assign new_n607 = new_n605 & new_n606;
  assign new_n608 = new_n604 & new_n607;
  assign new_n609 = new_n602 & new_n608;
  assign new_n610 = ~new_n396 & ~new_n401;
  assign new_n611 = ~new_n403 & new_n610;
  assign new_n612 = ~new_n387 & ~new_n390;
  assign new_n613 = ~new_n378 & ~new_n382;
  assign new_n614 = new_n612 & new_n613;
  assign new_n615 = new_n611 & new_n614;
  assign new_n616 = ~new_n363 & ~new_n369;
  assign new_n617 = ~new_n374 & new_n616;
  assign new_n618 = ~new_n354 & ~new_n357;
  assign new_n619 = ~new_n347 & ~new_n351;
  assign new_n620 = new_n618 & new_n619;
  assign new_n621 = new_n617 & new_n620;
  assign new_n622 = new_n615 & new_n621;
  assign new_n623 = new_n609 & new_n622;
  assign new_n624 = new_n596 & new_n623;
  assign new_n625 = ~new_n339 & ~new_n341;
  assign new_n626 = ~new_n342 & new_n625;
  assign new_n627 = ~new_n329 & ~new_n333;
  assign new_n628 = ~new_n319 & ~new_n324;
  assign new_n629 = new_n627 & new_n628;
  assign new_n630 = new_n626 & new_n629;
  assign new_n631 = ~new_n305 & ~new_n311;
  assign new_n632 = ~new_n317 & new_n631;
  assign new_n633 = ~new_n297 & ~new_n302;
  assign new_n634 = ~new_n286 & ~new_n292;
  assign new_n635 = new_n633 & new_n634;
  assign new_n636 = new_n632 & new_n635;
  assign new_n637 = new_n630 & new_n636;
  assign new_n638 = ~new_n271 & ~new_n275;
  assign new_n639 = ~new_n281 & new_n638;
  assign new_n640 = ~new_n261 & ~new_n266;
  assign new_n641 = ~new_n250 & ~new_n256;
  assign new_n642 = new_n640 & new_n641;
  assign new_n643 = new_n639 & new_n642;
  assign new_n644 = ~new_n235 & ~new_n240;
  assign new_n645 = ~new_n244 & new_n644;
  assign new_n646 = ~new_n225 & ~new_n231;
  assign new_n647 = ~new_n211 & ~new_n219;
  assign new_n648 = new_n646 & new_n647;
  assign new_n649 = new_n645 & new_n648;
  assign new_n650 = new_n643 & new_n649;
  assign new_n651 = new_n637 & new_n650;
  assign new_n652 = ~new_n189 & ~new_n194;
  assign new_n653 = ~new_n199 & new_n652;
  assign new_n654 = ~new_n179 & ~new_n184;
  assign new_n655 = ~new_n170 & ~new_n174;
  assign new_n656 = new_n654 & new_n655;
  assign new_n657 = new_n653 & new_n656;
  assign new_n658 = ~new_n148 & ~new_n153;
  assign new_n659 = ~new_n157 & new_n658;
  assign new_n660 = ~new_n138 & ~new_n144;
  assign new_n661 = ~new_n126 & ~new_n131;
  assign new_n662 = new_n660 & new_n661;
  assign new_n663 = new_n659 & new_n662;
  assign new_n664 = new_n657 & new_n663;
  assign new_n665 = ~new_n110 & ~new_n116;
  assign new_n666 = ~new_n121 & new_n665;
  assign new_n667 = ~new_n93 & ~new_n102;
  assign new_n668 = ~new_n83 & ~new_n84;
  assign new_n669 = new_n667 & new_n668;
  assign new_n670 = new_n666 & new_n669;
  assign new_n671 = ~new_n60 & ~new_n63;
  assign new_n672 = ~new_n73 & new_n671;
  assign new_n673 = ~new_n47 & ~new_n50;
  assign new_n674 = ~new_n34 & ~new_n37;
  assign new_n675 = new_n673 & new_n674;
  assign new_n676 = new_n672 & new_n675;
  assign new_n677 = new_n670 & new_n676;
  assign new_n678 = new_n664 & new_n677;
  assign new_n679 = new_n651 & new_n678;
  assign pd0 = ~new_n624 | ~new_n679;
  assign new_n681 = pe & pf;
  assign new_n682 = ~pa0 & pf;
  assign new_n683 = ~pa & ~new_n682;
  assign new_n684 = ~pc & ~new_n681;
  assign pe0 = ~new_n683 | ~new_n684;
  assign new_n686 = ~pb0 & ~pe;
  assign new_n687 = pc & ~pe;
  assign new_n688 = pa & ~pe;
  assign new_n689 = ~new_n686 & ~new_n687;
  assign pf0 = new_n688 | ~new_n689;
endmodule


