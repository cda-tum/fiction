// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3, pb0,
    pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1, pf2,
    pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0, pg1, pv,
    pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4, pm5, ph1,
    pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5, pz, ph3,
    pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5, pi4, pl1,
    pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3, pm2, pn1,
    po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4, pb, pp2,
    pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5, pt0,
    pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2, pu3,
    pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1,
    py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4, pn,
    pz4, po,
    pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8, pk9,
    ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7, pc6,
    pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9, pn6,
    po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7, pm6,
    pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9, pg8,
    ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8, pc10,
    pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7, pd10,
    pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9, ph10,
    pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5, pz6,
    pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9, pw8,
    px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pe5, pp, pa0, pb3, pc2, pd5, pe4, pq, pa3,
    pb0, pc1, pf4, pg5, pr, pa2, pb1, pc0, pf5, pg4, ps, pa5, pd0, pe1,
    pf2, pg3, pt, pa4, pd1, pe0, pf3, pg2, pu, pb4, pc5, pd2, pe3, pf0,
    pg1, pv, pb5, pc4, pd3, pe2, pf1, pg0, pw, ph0, pi1, pj2, pk3, pl4,
    pm5, ph1, pi0, pj3, pk2, pl5, pm4, py, ph2, pi3, pj0, pk1, pn4, po5,
    pz, ph3, pi2, pj1, pk0, pn5, po4, ph4, pi5, pl0, pm1, pn2, po3, ph5,
    pi4, pl1, pm0, pn3, po2, pj4, pk5, pl2, pm3, pn0, po1, pj5, pk4, pl3,
    pm2, pn1, po0, pp0, pq1, pr2, ps3, pt4, pa, pp1, pq0, pr3, ps2, pu4,
    pb, pp2, pq3, pr0, ps1, pv4, pc, pp3, pq2, pr1, ps0, pw4, pd, pp4, pq5,
    pt0, pu1, pv2, pw3, pe, pp5, pq4, pt1, pu0, pv3, pw2, pf, pr4, pt2,
    pu3, pv0, pw1, pg, pr5, ps4, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi,
    px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, px4, pm, py4,
    pn, pz4, po;
  output pf6, pg7, ph8, pi9, pq10, pf7, pg6, ph9, pi8, pp10, pd6, pe7, pj8,
    pk9, ps10, pd7, pe6, pj9, pk8, pr10, pb6, pc7, pl8, pm9, pu10, pb7,
    pc6, pl9, pm8, pt10, pa7, pn8, po9, pw10, pa6, pn9, po8, pv10, pa9,
    pn6, po7, py10, pa8, pn7, po6, px10, pb8, pc9, pl6, pm7, pb9, pc8, pl7,
    pm6, pd8, pe9, pj6, pk7, pd9, pe8, pj7, pk6, pf8, pg9, ph6, pi7, pf9,
    pg8, ph7, pi6, pa10, pu5, pv6, pw7, px8, py9, pt5, pv7, pw6, px9, py8,
    pc10, pt6, pu7, pw5, pz8, pb10, pt7, pu6, pv5, pz9, pe10, pr6, ps7,
    pd10, pr7, ps6, pg10, pp6, pq7, ps5, pf10, pp7, pq6, pi10, pp8, pq9,
    ph10, pp9, pq8, pk10, pr8, ps9, pj10, pr9, ps8, pm10, pt8, pu9, py5,
    pz6, pl10, pt9, pu8, px5, pz7, po10, pv8, pw9, px6, py7, pn10, pv9,
    pw8, px7, py6, pz5;
  wire new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n334, new_n335, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1395, new_n1396, new_n1397, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1420,
    new_n1421, new_n1422, new_n1423, new_n1424, new_n1425, new_n1426,
    new_n1427, new_n1428, new_n1429, new_n1430, new_n1431, new_n1432,
    new_n1433, new_n1434, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1541, new_n1542, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1634, new_n1635, new_n1636, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1654, new_n1655, new_n1656, new_n1657, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1675, new_n1676, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1719, new_n1720,
    new_n1721, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1728, new_n1729, new_n1730, new_n1731, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1751, new_n1752, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1768, new_n1769,
    new_n1770, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1873, new_n1874, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1879, new_n1880, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1926, new_n1927, new_n1928,
    new_n1929, new_n1930, new_n1931, new_n1932, new_n1933, new_n1934,
    new_n1935, new_n1936, new_n1937, new_n1938, new_n1939, new_n1940,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1951, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1994,
    new_n1995, new_n1996, new_n1997, new_n1998, new_n1999, new_n2000,
    new_n2001, new_n2002, new_n2003, new_n2005, new_n2006, new_n2007,
    new_n2009, new_n2010, new_n2011, new_n2012, new_n2013, new_n2014,
    new_n2015, new_n2016, new_n2017, new_n2018, new_n2019, new_n2020,
    new_n2021, new_n2022, new_n2023, new_n2024, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045;
  assign new_n311 = ~pm1 & ~pb;
  assign new_n312 = pl1 & pn1;
  assign new_n313 = new_n311 & new_n312;
  assign new_n314 = ~pn1 & ~pb;
  assign new_n315 = pm1 & pl1;
  assign new_n316 = new_n314 & new_n315;
  assign new_n317 = pv0 & new_n316;
  assign new_n318 = pr1 & new_n317;
  assign new_n319 = ~pj1 & ~po1;
  assign new_n320 = ~pk1 & po1;
  assign new_n321 = ~new_n319 & ~new_n320;
  assign new_n322 = pj1 & ~new_n321;
  assign new_n323 = pe1 & ~pf1;
  assign new_n324 = new_n322 & ~new_n323;
  assign new_n325 = ~new_n322 & new_n323;
  assign new_n326 = ~new_n324 & ~new_n325;
  assign new_n327 = ~pi1 & ~ph1;
  assign new_n328 = new_n322 & ~new_n326;
  assign new_n329 = new_n327 & new_n328;
  assign new_n330 = ~ph1 & ~new_n329;
  assign new_n331 = ~pm1 & ~pl1;
  assign new_n332 = ~pn1 & new_n331;
  assign pv6 = pb | new_n332;
  assign new_n334 = ~new_n326 & new_n327;
  assign new_n335 = new_n323 & new_n334;
  assign pn6 = pi1 | new_n335;
  assign new_n337 = ~pg1 & ~pn6;
  assign new_n338 = new_n330 & pv6;
  assign new_n339 = new_n337 & new_n338;
  assign new_n340 = ~new_n313 & ~new_n318;
  assign new_n341 = ~pb & ~new_n339;
  assign new_n342 = new_n340 & new_n341;
  assign new_n343 = ~pr1 & new_n337;
  assign new_n344 = ~new_n316 & new_n337;
  assign new_n345 = ~new_n343 & ~new_n344;
  assign new_n346 = new_n330 & ~new_n345;
  assign new_n347 = pw0 & ~new_n346;
  assign new_n348 = px0 & new_n347;
  assign new_n349 = pv0 & new_n348;
  assign new_n350 = ~py0 & ~new_n349;
  assign new_n351 = py0 & new_n349;
  assign new_n352 = ~new_n350 & ~new_n351;
  assign pf6 = new_n342 & new_n352;
  assign new_n354 = ~px0 & ~py0;
  assign new_n355 = ~pz0 & new_n354;
  assign new_n356 = ~pp1 & ~new_n355;
  assign new_n357 = ~pr1 & new_n356;
  assign new_n358 = ~pa1 & ~pc1;
  assign new_n359 = ~pb1 & new_n358;
  assign new_n360 = new_n355 & new_n359;
  assign new_n361 = new_n356 & ~new_n360;
  assign new_n362 = ~new_n354 & ~new_n355;
  assign new_n363 = ~pr1 & new_n362;
  assign new_n364 = ~new_n360 & new_n362;
  assign new_n365 = ~pv0 & pw0;
  assign new_n366 = ~pq1 & ~pp1;
  assign new_n367 = ~pr1 & new_n366;
  assign new_n368 = ~new_n360 & new_n366;
  assign new_n369 = ~pq1 & ~new_n354;
  assign new_n370 = ~pr1 & new_n369;
  assign new_n371 = ~new_n360 & new_n369;
  assign new_n372 = ~new_n370 & ~new_n371;
  assign new_n373 = ~new_n367 & ~new_n368;
  assign new_n374 = new_n372 & new_n373;
  assign new_n375 = ~new_n357 & ~new_n361;
  assign new_n376 = ~new_n363 & new_n375;
  assign new_n377 = ~new_n364 & new_n365;
  assign new_n378 = new_n376 & new_n377;
  assign new_n379 = new_n374 & new_n378;
  assign new_n380 = pv6 & new_n379;
  assign new_n381 = ~ph & ~new_n380;
  assign new_n382 = ps1 & pt1;
  assign new_n383 = pu1 & new_n382;
  assign new_n384 = ~pk & ~new_n383;
  assign new_n385 = pw1 & ~new_n384;
  assign new_n386 = pv1 & new_n385;
  assign new_n387 = px1 & new_n386;
  assign new_n388 = ~pk & ~new_n387;
  assign new_n389 = py1 & ~new_n388;
  assign new_n390 = ~pi & new_n337;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = ~ps1 & ~pt1;
  assign new_n393 = ~pu1 & new_n392;
  assign new_n394 = ~pk & ~new_n393;
  assign new_n395 = ~pw1 & ~new_n394;
  assign new_n396 = ~pv1 & new_n395;
  assign new_n397 = ~px1 & new_n396;
  assign new_n398 = ~pk & ~new_n397;
  assign new_n399 = ~py1 & ~new_n398;
  assign new_n400 = ~new_n389 & ~new_n399;
  assign new_n401 = new_n390 & ~new_n399;
  assign new_n402 = ~new_n391 & ~new_n400;
  assign new_n403 = ~new_n401 & new_n402;
  assign new_n404 = ~new_n381 & new_n403;
  assign new_n405 = ~pz1 & new_n404;
  assign new_n406 = pz1 & ~new_n404;
  assign new_n407 = ~new_n405 & ~new_n406;
  assign new_n408 = ~pd3 & new_n407;
  assign new_n409 = ~pn1 & new_n311;
  assign new_n410 = pl1 & new_n409;
  assign new_n411 = ~pv6 & ~new_n410;
  assign new_n412 = ~pd1 & ~pw0;
  assign new_n413 = new_n360 & new_n412;
  assign new_n414 = pv0 & new_n413;
  assign new_n415 = ~new_n410 & ~new_n414;
  assign new_n416 = ~new_n411 & ~new_n415;
  assign new_n417 = new_n407 & ~new_n416;
  assign new_n418 = ~pd3 & new_n416;
  assign new_n419 = ~new_n408 & ~new_n417;
  assign new_n420 = ~new_n418 & new_n419;
  assign pg7 = pb | new_n420;
  assign new_n422 = pv6 & ~new_n337;
  assign new_n423 = ~pg & ~new_n422;
  assign new_n424 = pm1 & ~pb;
  assign new_n425 = ~pn1 & new_n424;
  assign new_n426 = ~pl1 & new_n425;
  assign new_n427 = ~pb & ~new_n426;
  assign new_n428 = ~new_n423 & ~new_n427;
  assign new_n429 = pr1 & ~pv6;
  assign new_n430 = ~pv0 & new_n429;
  assign new_n431 = ~new_n316 & ~pv6;
  assign new_n432 = new_n330 & new_n337;
  assign new_n433 = ~pv0 & new_n413;
  assign new_n434 = ~new_n432 & new_n433;
  assign new_n435 = pr1 & ~new_n434;
  assign new_n436 = ~pv0 & new_n435;
  assign new_n437 = ~new_n316 & ~new_n434;
  assign new_n438 = ~new_n430 & ~new_n431;
  assign new_n439 = ~new_n436 & ~new_n437;
  assign new_n440 = new_n438 & new_n439;
  assign new_n441 = ~pf & ~new_n440;
  assign new_n442 = pp1 & new_n316;
  assign new_n443 = ~pj & new_n442;
  assign new_n444 = pr2 & pq2;
  assign new_n445 = pq1 & new_n316;
  assign new_n446 = ~pj & new_n445;
  assign new_n447 = ~new_n444 & ~new_n446;
  assign new_n448 = ~new_n443 & new_n447;
  assign new_n449 = ~ps2 & ~new_n443;
  assign new_n450 = ~new_n448 & ~new_n449;
  assign new_n451 = pt2 & new_n450;
  assign new_n452 = ~pj & ~new_n451;
  assign new_n453 = pv2 & ~new_n452;
  assign new_n454 = ~new_n423 & ~new_n453;
  assign new_n455 = ~pr2 & ~pq2;
  assign new_n456 = ~new_n446 & ~new_n455;
  assign new_n457 = ~new_n443 & new_n456;
  assign new_n458 = ps2 & ~new_n443;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = ~pt2 & new_n459;
  assign new_n461 = ~pj & ~new_n460;
  assign new_n462 = pu2 & ~new_n461;
  assign new_n463 = ~new_n453 & ~new_n462;
  assign new_n464 = new_n423 & ~new_n462;
  assign new_n465 = ~new_n454 & ~new_n463;
  assign new_n466 = ~new_n464 & new_n465;
  assign new_n467 = ~new_n441 & new_n466;
  assign new_n468 = ~pa3 & new_n467;
  assign new_n469 = pa3 & ~new_n467;
  assign new_n470 = ~new_n468 & ~new_n469;
  assign new_n471 = new_n427 & ~new_n470;
  assign ph8 = new_n428 | new_n471;
  assign new_n473 = ~pm5 & ~pz;
  assign new_n474 = ~pn5 & new_n473;
  assign new_n475 = pl5 & new_n474;
  assign new_n476 = ~pm5 & ~pl5;
  assign new_n477 = ~pn5 & new_n476;
  assign pv10 = pz | new_n477;
  assign new_n479 = ~new_n475 & ~pv10;
  assign new_n480 = ~pt4 & ~pu4;
  assign new_n481 = ~pv4 & new_n480;
  assign new_n482 = ~pw4 & ~py4;
  assign new_n483 = ~px4 & new_n482;
  assign new_n484 = new_n481 & new_n483;
  assign new_n485 = ~ps4 & ~pz4;
  assign new_n486 = new_n484 & new_n485;
  assign new_n487 = pr4 & new_n486;
  assign new_n488 = ~new_n475 & ~new_n487;
  assign new_n489 = ~new_n479 & ~new_n488;
  assign new_n490 = ~pr5 & ~new_n480;
  assign new_n491 = ~pq5 & new_n490;
  assign new_n492 = ~new_n480 & ~new_n484;
  assign new_n493 = ~pq5 & new_n492;
  assign new_n494 = ~pp5 & ~pr5;
  assign new_n495 = ~pq5 & new_n494;
  assign new_n496 = ~pp5 & ~new_n484;
  assign new_n497 = ~pq5 & new_n496;
  assign new_n498 = ~pr4 & ps4;
  assign new_n499 = ~new_n480 & ~new_n481;
  assign new_n500 = ~pr5 & new_n499;
  assign new_n501 = ~new_n484 & new_n499;
  assign new_n502 = ~pr5 & ~new_n481;
  assign new_n503 = ~pp5 & new_n502;
  assign new_n504 = ~new_n481 & ~new_n484;
  assign new_n505 = ~pp5 & new_n504;
  assign new_n506 = ~new_n503 & ~new_n505;
  assign new_n507 = ~new_n500 & ~new_n501;
  assign new_n508 = new_n506 & new_n507;
  assign new_n509 = ~new_n491 & ~new_n493;
  assign new_n510 = ~new_n495 & new_n509;
  assign new_n511 = ~new_n497 & new_n498;
  assign new_n512 = new_n510 & new_n511;
  assign new_n513 = new_n508 & new_n512;
  assign new_n514 = pv10 & new_n513;
  assign new_n515 = ~pf0 & ~new_n514;
  assign new_n516 = ~pg5 & ~po5;
  assign new_n517 = po5 & ~pi5;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = pg5 & ~new_n518;
  assign new_n520 = pa5 & ~pb5;
  assign new_n521 = new_n519 & ~new_n520;
  assign new_n522 = ~new_n519 & new_n520;
  assign new_n523 = ~new_n521 & ~new_n522;
  assign new_n524 = ~pe5 & ~pd5;
  assign new_n525 = ~new_n523 & new_n524;
  assign new_n526 = new_n520 & new_n525;
  assign pj10 = pe5 | new_n526;
  assign new_n528 = ~pc5 & ~pj10;
  assign new_n529 = ~pg0 & new_n528;
  assign new_n530 = ~pv3 & ~pu3;
  assign new_n531 = ~pw3 & new_n530;
  assign new_n532 = ~pi0 & ~new_n531;
  assign new_n533 = ~py3 & ~new_n532;
  assign new_n534 = ~px3 & new_n533;
  assign new_n535 = ~pz3 & new_n534;
  assign new_n536 = ~pi0 & ~new_n535;
  assign new_n537 = ~pa4 & ~new_n536;
  assign new_n538 = new_n529 & ~new_n537;
  assign new_n539 = pv3 & pu3;
  assign new_n540 = pw3 & new_n539;
  assign new_n541 = ~pi0 & ~new_n540;
  assign new_n542 = py3 & ~new_n541;
  assign new_n543 = px3 & new_n542;
  assign new_n544 = pz3 & new_n543;
  assign new_n545 = ~pi0 & ~new_n544;
  assign new_n546 = pa4 & ~new_n545;
  assign new_n547 = ~new_n529 & ~new_n546;
  assign new_n548 = ~new_n537 & ~new_n546;
  assign new_n549 = ~new_n538 & ~new_n547;
  assign new_n550 = ~new_n548 & new_n549;
  assign new_n551 = ~new_n515 & new_n550;
  assign new_n552 = ~pb4 & new_n551;
  assign new_n553 = pb4 & ~new_n551;
  assign new_n554 = ~new_n552 & ~new_n553;
  assign new_n555 = ~new_n489 & new_n554;
  assign new_n556 = ~ps3 & new_n489;
  assign new_n557 = ~ps3 & new_n554;
  assign new_n558 = ~new_n555 & ~new_n556;
  assign new_n559 = ~new_n557 & new_n558;
  assign pi9 = pz | new_n559;
  assign new_n561 = pk5 & ~pj5;
  assign new_n562 = ~pz & ~new_n561;
  assign new_n563 = ~pz & ~pn5;
  assign new_n564 = pm5 & pl5;
  assign new_n565 = new_n563 & new_n564;
  assign new_n566 = pj5 & new_n565;
  assign new_n567 = ~pj5 & ~new_n565;
  assign new_n568 = ~new_n566 & ~new_n567;
  assign pq10 = new_n562 & new_n568;
  assign new_n570 = new_n388 & ~new_n390;
  assign new_n571 = new_n388 & new_n398;
  assign new_n572 = new_n390 & new_n398;
  assign new_n573 = ~new_n570 & ~new_n571;
  assign new_n574 = ~new_n572 & new_n573;
  assign new_n575 = ~new_n381 & new_n574;
  assign new_n576 = ~py1 & new_n575;
  assign new_n577 = py1 & ~new_n575;
  assign new_n578 = ~new_n576 & ~new_n577;
  assign new_n579 = ~pc3 & new_n578;
  assign new_n580 = ~new_n416 & new_n578;
  assign new_n581 = ~pc3 & new_n416;
  assign new_n582 = ~new_n579 & ~new_n580;
  assign new_n583 = ~new_n581 & new_n582;
  assign pf7 = ~pb & new_n583;
  assign new_n585 = pw0 & py0;
  assign new_n586 = pv0 & px0;
  assign new_n587 = new_n585 & new_n586;
  assign new_n588 = ~new_n346 & new_n587;
  assign new_n589 = ~pz0 & ~new_n588;
  assign new_n590 = pz0 & new_n588;
  assign new_n591 = ~new_n589 & ~new_n590;
  assign pg6 = new_n342 & new_n591;
  assign new_n593 = new_n529 & new_n536;
  assign new_n594 = ~new_n529 & new_n545;
  assign new_n595 = new_n536 & new_n545;
  assign new_n596 = ~new_n593 & ~new_n594;
  assign new_n597 = ~new_n595 & new_n596;
  assign new_n598 = ~new_n515 & new_n597;
  assign new_n599 = ~pa4 & new_n598;
  assign new_n600 = pa4 & ~new_n598;
  assign new_n601 = ~new_n599 & ~new_n600;
  assign new_n602 = ~new_n489 & new_n601;
  assign new_n603 = ~pr3 & new_n489;
  assign new_n604 = ~pr3 & new_n601;
  assign new_n605 = ~new_n602 & ~new_n603;
  assign new_n606 = ~new_n604 & new_n605;
  assign ph9 = ~pz & new_n606;
  assign new_n608 = pa3 & new_n453;
  assign new_n609 = ~pj & ~new_n608;
  assign new_n610 = ~new_n423 & new_n609;
  assign new_n611 = ~pa3 & new_n462;
  assign new_n612 = ~pj & ~new_n611;
  assign new_n613 = new_n609 & new_n612;
  assign new_n614 = new_n423 & new_n612;
  assign new_n615 = ~new_n610 & ~new_n613;
  assign new_n616 = ~new_n614 & new_n615;
  assign new_n617 = ~new_n441 & new_n616;
  assign new_n618 = ~pb3 & new_n617;
  assign new_n619 = pb3 & ~new_n617;
  assign new_n620 = ~new_n618 & ~new_n619;
  assign new_n621 = new_n427 & ~new_n620;
  assign pi8 = new_n428 | new_n621;
  assign new_n623 = pv0 & ~new_n346;
  assign new_n624 = ~pw0 & ~new_n623;
  assign new_n625 = pw0 & new_n623;
  assign new_n626 = ~new_n624 & ~new_n625;
  assign pd6 = new_n342 & new_n626;
  assign new_n628 = pv1 & ~new_n384;
  assign new_n629 = pw1 & new_n628;
  assign new_n630 = ~new_n390 & ~new_n629;
  assign new_n631 = ~pw1 & ~pv1;
  assign new_n632 = ~new_n394 & new_n631;
  assign new_n633 = ~new_n629 & ~new_n632;
  assign new_n634 = new_n390 & ~new_n632;
  assign new_n635 = ~new_n630 & ~new_n633;
  assign new_n636 = ~new_n634 & new_n635;
  assign new_n637 = ~new_n381 & new_n636;
  assign new_n638 = ~px1 & new_n637;
  assign new_n639 = px1 & ~new_n637;
  assign new_n640 = ~new_n638 & ~new_n639;
  assign new_n641 = ~pb3 & new_n640;
  assign new_n642 = ~new_n416 & new_n640;
  assign new_n643 = ~pb3 & new_n416;
  assign new_n644 = ~new_n641 & ~new_n642;
  assign new_n645 = ~new_n643 & new_n644;
  assign pe7 = pb | new_n645;
  assign new_n647 = pb3 & ~new_n609;
  assign new_n648 = ~new_n423 & ~new_n647;
  assign new_n649 = ~pb3 & ~new_n612;
  assign new_n650 = ~new_n647 & ~new_n649;
  assign new_n651 = new_n423 & ~new_n649;
  assign new_n652 = ~new_n648 & ~new_n650;
  assign new_n653 = ~new_n651 & new_n652;
  assign new_n654 = ~new_n441 & new_n653;
  assign new_n655 = ~pc3 & ~new_n654;
  assign new_n656 = pc3 & new_n654;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign pj8 = new_n427 & new_n657;
  assign pk9 = ~pd4 | pz;
  assign new_n660 = pm5 & ~pz;
  assign new_n661 = ~pn5 & new_n660;
  assign new_n662 = ~pl5 & new_n661;
  assign new_n663 = new_n520 & new_n662;
  assign new_n664 = pq3 & pp3;
  assign new_n665 = ps3 & new_n664;
  assign new_n666 = pr3 & new_n665;
  assign new_n667 = pt3 & new_n666;
  assign new_n668 = ~pr3 & ~pt3;
  assign new_n669 = ~ps3 & ~pq3;
  assign new_n670 = new_n668 & new_n669;
  assign new_n671 = ~po3 & ~pp3;
  assign new_n672 = pn3 & new_n671;
  assign new_n673 = new_n670 & new_n672;
  assign new_n674 = new_n520 & new_n667;
  assign new_n675 = ~new_n673 & new_n674;
  assign new_n676 = new_n565 & ~new_n675;
  assign new_n677 = ~new_n475 & ~new_n663;
  assign new_n678 = ~new_n676 & new_n677;
  assign ps10 = ~pz & ~new_n678;
  assign new_n680 = ~new_n390 & ~new_n628;
  assign new_n681 = ~pv1 & ~new_n394;
  assign new_n682 = ~new_n628 & ~new_n681;
  assign new_n683 = new_n390 & ~new_n681;
  assign new_n684 = ~new_n680 & ~new_n682;
  assign new_n685 = ~new_n683 & new_n684;
  assign new_n686 = ~new_n381 & new_n685;
  assign new_n687 = ~pw1 & new_n686;
  assign new_n688 = pw1 & ~new_n686;
  assign new_n689 = ~new_n687 & ~new_n688;
  assign new_n690 = ~pa3 & new_n689;
  assign new_n691 = ~new_n416 & new_n689;
  assign new_n692 = ~pa3 & new_n416;
  assign new_n693 = ~new_n690 & ~new_n691;
  assign new_n694 = ~new_n692 & new_n693;
  assign pd7 = pb | new_n694;
  assign new_n696 = pv0 & new_n347;
  assign new_n697 = ~px0 & ~new_n696;
  assign new_n698 = px0 & new_n696;
  assign new_n699 = ~new_n697 & ~new_n698;
  assign pe6 = new_n342 & new_n699;
  assign new_n701 = ~pa4 & ~pb4;
  assign new_n702 = ~new_n536 & new_n701;
  assign new_n703 = new_n529 & ~new_n702;
  assign new_n704 = pb4 & new_n546;
  assign new_n705 = ~new_n529 & ~new_n704;
  assign new_n706 = ~new_n702 & ~new_n704;
  assign new_n707 = ~new_n703 & ~new_n705;
  assign new_n708 = ~new_n706 & new_n707;
  assign new_n709 = ~new_n515 & new_n708;
  assign new_n710 = ~pc4 & new_n709;
  assign new_n711 = pc4 & ~new_n709;
  assign new_n712 = ~new_n710 & ~new_n711;
  assign new_n713 = ~new_n489 & new_n712;
  assign new_n714 = ~pt3 & new_n489;
  assign new_n715 = ~pt3 & new_n712;
  assign new_n716 = ~new_n713 & ~new_n714;
  assign new_n717 = ~new_n715 & new_n716;
  assign pj9 = pz | new_n717;
  assign new_n719 = pc3 & new_n647;
  assign new_n720 = ~new_n423 & ~new_n719;
  assign new_n721 = ~pc3 & new_n649;
  assign new_n722 = ~new_n719 & ~new_n721;
  assign new_n723 = new_n423 & ~new_n721;
  assign new_n724 = ~new_n720 & ~new_n722;
  assign new_n725 = ~new_n723 & new_n724;
  assign new_n726 = ~new_n441 & new_n725;
  assign new_n727 = ~pd3 & new_n726;
  assign new_n728 = pd3 & ~new_n726;
  assign new_n729 = ~new_n727 & ~new_n728;
  assign new_n730 = new_n427 & ~new_n729;
  assign pk8 = new_n428 | new_n730;
  assign new_n732 = ~pk5 & ~new_n566;
  assign new_n733 = pk5 & new_n566;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign pr10 = new_n562 & new_n734;
  assign new_n736 = pn0 & pq5;
  assign new_n737 = pn5 & pp0;
  assign new_n738 = ~pz & ~new_n662;
  assign new_n739 = po0 & ~new_n738;
  assign new_n740 = ~pj0 & ~pp5;
  assign new_n741 = pd4 & pe4;
  assign new_n742 = pf4 & new_n741;
  assign new_n743 = ~pj0 & pq5;
  assign new_n744 = ~new_n742 & ~new_n743;
  assign new_n745 = pi4 & ~new_n744;
  assign new_n746 = new_n740 & ~new_n745;
  assign new_n747 = pg4 & pp4;
  assign new_n748 = ~new_n746 & new_n747;
  assign new_n749 = pq0 & new_n748;
  assign new_n750 = ~new_n736 & ~new_n737;
  assign new_n751 = ~new_n739 & ~new_n749;
  assign new_n752 = new_n750 & new_n751;
  assign new_n753 = pl0 & pl3;
  assign new_n754 = pk0 & new_n673;
  assign new_n755 = pm0 & new_n667;
  assign new_n756 = ~new_n753 & ~new_n754;
  assign new_n757 = ~new_n755 & new_n756;
  assign new_n758 = pg4 & pr0;
  assign new_n759 = pv4 & pt0;
  assign new_n760 = pr5 & ~pv10;
  assign new_n761 = ~pr4 & new_n760;
  assign new_n762 = ~pv10 & ~new_n561;
  assign new_n763 = new_n519 & ~new_n523;
  assign new_n764 = new_n524 & new_n763;
  assign new_n765 = ~pd5 & ~new_n764;
  assign new_n766 = new_n528 & new_n765;
  assign new_n767 = ~pr4 & new_n486;
  assign new_n768 = ~new_n766 & new_n767;
  assign new_n769 = pr5 & ~new_n768;
  assign new_n770 = ~pr4 & new_n769;
  assign new_n771 = ~new_n561 & ~new_n768;
  assign new_n772 = ~new_n761 & ~new_n762;
  assign new_n773 = ~new_n770 & ~new_n771;
  assign new_n774 = new_n772 & new_n773;
  assign new_n775 = ~pd0 & ~new_n774;
  assign new_n776 = ps0 & new_n775;
  assign new_n777 = pl5 & pu0;
  assign new_n778 = ~new_n758 & ~new_n759;
  assign new_n779 = ~new_n776 & ~new_n777;
  assign new_n780 = new_n778 & new_n779;
  assign new_n781 = new_n752 & new_n757;
  assign pb6 = ~new_n780 | ~new_n781;
  assign new_n783 = new_n384 & ~new_n390;
  assign new_n784 = new_n384 & new_n394;
  assign new_n785 = new_n390 & new_n394;
  assign new_n786 = ~new_n783 & ~new_n784;
  assign new_n787 = ~new_n785 & new_n786;
  assign new_n788 = ~new_n381 & new_n787;
  assign new_n789 = ~pv1 & new_n788;
  assign new_n790 = pv1 & ~new_n788;
  assign new_n791 = ~new_n789 & ~new_n790;
  assign new_n792 = ~pz2 & new_n791;
  assign new_n793 = ~new_n416 & new_n791;
  assign new_n794 = ~pz2 & new_n416;
  assign new_n795 = ~new_n792 & ~new_n793;
  assign new_n796 = ~new_n794 & new_n795;
  assign pc7 = pb | new_n796;
  assign new_n798 = pd3 & new_n719;
  assign new_n799 = ~new_n423 & ~new_n798;
  assign new_n800 = ~pc3 & ~pd3;
  assign new_n801 = new_n649 & new_n800;
  assign new_n802 = ~new_n798 & ~new_n801;
  assign new_n803 = new_n423 & ~new_n801;
  assign new_n804 = ~new_n799 & ~new_n802;
  assign new_n805 = ~new_n803 & new_n804;
  assign new_n806 = ~new_n441 & new_n805;
  assign new_n807 = ~pe3 & new_n806;
  assign new_n808 = pe3 & ~new_n806;
  assign new_n809 = ~new_n807 & ~new_n808;
  assign new_n810 = new_n427 & ~new_n809;
  assign pl8 = new_n428 | new_n810;
  assign new_n812 = ~pf4 & ~new_n741;
  assign new_n813 = ~new_n742 & ~new_n812;
  assign pm9 = pz | new_n813;
  assign new_n815 = pn5 & new_n660;
  assign new_n816 = pl5 & new_n815;
  assign new_n817 = ~new_n667 & ~new_n816;
  assign new_n818 = ~new_n520 & ~new_n816;
  assign new_n819 = new_n673 & ~new_n816;
  assign new_n820 = ~new_n565 & ~new_n816;
  assign new_n821 = ~new_n817 & ~new_n818;
  assign new_n822 = ~new_n819 & ~new_n820;
  assign new_n823 = new_n821 & new_n822;
  assign new_n824 = pn5 & new_n473;
  assign new_n825 = ~pl5 & new_n824;
  assign new_n826 = ~new_n475 & ~new_n825;
  assign new_n827 = ~new_n673 & new_n826;
  assign new_n828 = ~new_n565 & new_n826;
  assign new_n829 = ~new_n827 & ~new_n828;
  assign new_n830 = ~new_n823 & ~new_n829;
  assign pu10 = ~pz & ~new_n830;
  assign new_n832 = ~new_n382 & ~new_n390;
  assign new_n833 = ~new_n382 & ~new_n392;
  assign new_n834 = new_n390 & ~new_n392;
  assign new_n835 = ~new_n832 & ~new_n833;
  assign new_n836 = ~new_n834 & new_n835;
  assign new_n837 = ~new_n381 & new_n836;
  assign new_n838 = ~pu1 & new_n837;
  assign new_n839 = pu1 & ~new_n837;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = ~py2 & new_n840;
  assign new_n842 = ~new_n416 & new_n840;
  assign new_n843 = ~py2 & new_n416;
  assign new_n844 = ~new_n841 & ~new_n842;
  assign new_n845 = ~new_n843 & new_n844;
  assign pb7 = ~pb & new_n845;
  assign new_n847 = ~pv0 & new_n346;
  assign new_n848 = ~new_n623 & ~new_n847;
  assign pc6 = new_n342 & new_n848;
  assign new_n850 = ~pd4 & ~pe4;
  assign new_n851 = ~new_n741 & ~new_n850;
  assign pl9 = pz | new_n851;
  assign new_n853 = ~pf3 & new_n775;
  assign new_n854 = pf3 & ~new_n775;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign pm8 = new_n738 & new_n855;
  assign new_n857 = ~pm5 & ~new_n816;
  assign new_n858 = ~new_n565 & new_n857;
  assign new_n859 = new_n520 & new_n857;
  assign new_n860 = ~pn5 & ~new_n816;
  assign new_n861 = new_n520 & new_n860;
  assign new_n862 = new_n673 & new_n860;
  assign new_n863 = ~new_n565 & new_n860;
  assign new_n864 = new_n673 & new_n857;
  assign new_n865 = ~new_n858 & ~new_n859;
  assign new_n866 = ~new_n861 & new_n865;
  assign new_n867 = ~new_n862 & ~new_n863;
  assign new_n868 = ~new_n864 & new_n867;
  assign new_n869 = new_n866 & new_n868;
  assign new_n870 = new_n565 & new_n673;
  assign new_n871 = ~pr5 & new_n528;
  assign new_n872 = new_n528 & ~new_n565;
  assign new_n873 = ~new_n871 & ~new_n872;
  assign new_n874 = new_n765 & ~new_n873;
  assign new_n875 = py4 & ~new_n874;
  assign new_n876 = pw4 & px4;
  assign new_n877 = pv4 & new_n876;
  assign new_n878 = pu4 & ps4;
  assign new_n879 = pt4 & pr4;
  assign new_n880 = new_n878 & new_n879;
  assign new_n881 = new_n877 & new_n880;
  assign new_n882 = new_n875 & new_n881;
  assign new_n883 = pz4 & new_n882;
  assign new_n884 = ~pz4 & ~new_n883;
  assign new_n885 = ~pa0 & new_n884;
  assign new_n886 = pr5 & ~new_n883;
  assign new_n887 = ~pa0 & new_n886;
  assign new_n888 = ~pr5 & ~pz4;
  assign new_n889 = ~pa0 & new_n888;
  assign new_n890 = ~new_n885 & ~new_n887;
  assign new_n891 = ~new_n889 & new_n890;
  assign new_n892 = pv10 & new_n891;
  assign new_n893 = ~new_n870 & ~new_n892;
  assign new_n894 = ~new_n662 & ~new_n825;
  assign new_n895 = new_n893 & new_n894;
  assign new_n896 = ~new_n869 & new_n895;
  assign pt10 = ~pz & ~new_n896;
  assign new_n898 = ~ps1 & ~new_n390;
  assign new_n899 = ps1 & new_n390;
  assign new_n900 = ~new_n898 & ~new_n899;
  assign new_n901 = ~new_n381 & new_n900;
  assign new_n902 = ~pt1 & new_n901;
  assign new_n903 = pt1 & ~new_n901;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = ~px2 & new_n904;
  assign new_n906 = ~new_n416 & new_n904;
  assign new_n907 = ~px2 & new_n416;
  assign new_n908 = ~new_n905 & ~new_n906;
  assign new_n909 = ~new_n907 & new_n908;
  assign pa7 = ~pb & new_n909;
  assign new_n911 = pv10 & ~new_n528;
  assign new_n912 = ~pe0 & ~new_n911;
  assign new_n913 = ~pf3 & ~new_n912;
  assign new_n914 = pf3 & new_n912;
  assign new_n915 = ~new_n913 & ~new_n914;
  assign new_n916 = ~new_n775 & new_n915;
  assign new_n917 = ~pg3 & ~new_n916;
  assign new_n918 = pg3 & new_n916;
  assign new_n919 = ~new_n917 & ~new_n918;
  assign pn8 = new_n738 & new_n919;
  assign new_n921 = pl5 & pn5;
  assign new_n922 = new_n473 & new_n921;
  assign new_n923 = ~new_n748 & ~new_n922;
  assign new_n924 = ~pv3 & ~new_n923;
  assign new_n925 = pg4 & ~new_n746;
  assign new_n926 = ~ph4 & new_n925;
  assign new_n927 = ph4 & ~new_n925;
  assign new_n928 = ~new_n926 & ~new_n927;
  assign new_n929 = new_n923 & new_n928;
  assign new_n930 = ~pv3 & new_n928;
  assign new_n931 = ~new_n924 & ~new_n929;
  assign new_n932 = ~new_n930 & new_n931;
  assign po9 = pz | new_n932;
  assign new_n934 = ~pb0 & ~new_n825;
  assign new_n935 = ~pr5 & new_n934;
  assign new_n936 = ~pp5 & new_n935;
  assign new_n937 = ~pc0 & ~new_n816;
  assign new_n938 = new_n934 & new_n937;
  assign new_n939 = ~pp5 & new_n938;
  assign new_n940 = ~pq5 & new_n937;
  assign new_n941 = ~pp5 & new_n940;
  assign new_n942 = ~pr5 & ~new_n937;
  assign new_n943 = ~pq5 & new_n942;
  assign new_n944 = ~pq5 & ~pr5;
  assign new_n945 = ~pp5 & new_n944;
  assign new_n946 = ~new_n934 & new_n937;
  assign new_n947 = ~pq5 & new_n946;
  assign new_n948 = new_n934 & ~new_n937;
  assign new_n949 = ~pr5 & new_n948;
  assign new_n950 = ~pr5 & ~new_n934;
  assign new_n951 = ~pq5 & new_n950;
  assign new_n952 = ~new_n936 & ~new_n939;
  assign new_n953 = ~new_n941 & ~new_n943;
  assign new_n954 = new_n952 & new_n953;
  assign new_n955 = ~new_n949 & ~new_n951;
  assign new_n956 = ~new_n945 & ~new_n947;
  assign new_n957 = new_n955 & new_n956;
  assign new_n958 = new_n954 & new_n957;
  assign new_n959 = ~pq5 & ~pp5;
  assign new_n960 = ~new_n494 & ~new_n944;
  assign new_n961 = ~new_n959 & new_n960;
  assign new_n962 = ~pz & ~new_n961;
  assign new_n963 = pr5 & new_n962;
  assign new_n964 = pq5 & new_n962;
  assign new_n965 = pp5 & new_n962;
  assign new_n966 = ~new_n963 & ~new_n964;
  assign new_n967 = ~new_n965 & new_n966;
  assign pw10 = new_n958 | new_n967;
  assign new_n969 = pn0 & pp5;
  assign new_n970 = pm5 & pp0;
  assign new_n971 = po0 & pr5;
  assign new_n972 = pm4 & pq0;
  assign new_n973 = ~new_n969 & ~new_n970;
  assign new_n974 = ~new_n971 & ~new_n972;
  assign new_n975 = new_n973 & new_n974;
  assign new_n976 = pl0 & pm3;
  assign new_n977 = pk0 & pq3;
  assign new_n978 = pf3 & pm0;
  assign new_n979 = ~new_n976 & ~new_n977;
  assign new_n980 = ~new_n978 & new_n979;
  assign new_n981 = ph4 & pr0;
  assign new_n982 = pw4 & pt0;
  assign new_n983 = pd4 & ps0;
  assign new_n984 = pu0 & pr4;
  assign new_n985 = ~new_n981 & ~new_n982;
  assign new_n986 = ~new_n983 & ~new_n984;
  assign new_n987 = new_n985 & new_n986;
  assign new_n988 = new_n975 & new_n980;
  assign pa6 = ~new_n987 | ~new_n988;
  assign new_n990 = ~pu3 & ~new_n923;
  assign new_n991 = ~pg4 & ~new_n746;
  assign new_n992 = pg4 & new_n746;
  assign new_n993 = ~new_n991 & ~new_n992;
  assign new_n994 = new_n923 & new_n993;
  assign new_n995 = ~pu3 & new_n993;
  assign new_n996 = ~new_n990 & ~new_n994;
  assign new_n997 = ~new_n995 & new_n996;
  assign pn9 = pz | new_n997;
  assign new_n999 = ~pg3 & ~pf3;
  assign new_n1000 = pq5 & new_n565;
  assign new_n1001 = ~ph0 & new_n1000;
  assign new_n1002 = ~new_n999 & ~new_n1001;
  assign new_n1003 = new_n912 & new_n1002;
  assign new_n1004 = pg3 & pf3;
  assign new_n1005 = ~new_n1001 & ~new_n1004;
  assign new_n1006 = ~new_n912 & new_n1005;
  assign new_n1007 = new_n1002 & new_n1005;
  assign new_n1008 = ~new_n1003 & ~new_n1006;
  assign new_n1009 = ~new_n1007 & new_n1008;
  assign new_n1010 = ~new_n775 & new_n1009;
  assign new_n1011 = ~ph3 & ~new_n1010;
  assign new_n1012 = ph3 & new_n1010;
  assign new_n1013 = ~new_n1011 & ~new_n1012;
  assign po8 = new_n738 & new_n1013;
  assign new_n1015 = ~new_n738 & ~new_n912;
  assign new_n1016 = pp5 & new_n565;
  assign new_n1017 = ~ph0 & new_n1016;
  assign new_n1018 = new_n1002 & ~new_n1017;
  assign new_n1019 = ph3 & ~new_n1017;
  assign new_n1020 = ~new_n1018 & ~new_n1019;
  assign new_n1021 = ~pi3 & new_n1020;
  assign new_n1022 = ~ph0 & ~new_n1021;
  assign new_n1023 = pj3 & ~new_n1022;
  assign new_n1024 = ~pp3 & new_n1023;
  assign new_n1025 = ~ph0 & ~new_n1024;
  assign new_n1026 = ~pq3 & ~new_n1025;
  assign new_n1027 = ~ps3 & ~pr3;
  assign new_n1028 = new_n1026 & new_n1027;
  assign new_n1029 = new_n912 & ~new_n1028;
  assign new_n1030 = new_n1005 & ~new_n1017;
  assign new_n1031 = ~ph3 & ~new_n1017;
  assign new_n1032 = ~new_n1030 & ~new_n1031;
  assign new_n1033 = pi3 & new_n1032;
  assign new_n1034 = ~ph0 & ~new_n1033;
  assign new_n1035 = pk3 & ~new_n1034;
  assign new_n1036 = pp3 & new_n1035;
  assign new_n1037 = ~ph0 & ~new_n1036;
  assign new_n1038 = pq3 & ~new_n1037;
  assign new_n1039 = pr3 & new_n1038;
  assign new_n1040 = ps3 & new_n1039;
  assign new_n1041 = ~new_n912 & ~new_n1040;
  assign new_n1042 = ~new_n1028 & ~new_n1040;
  assign new_n1043 = ~new_n1029 & ~new_n1041;
  assign new_n1044 = ~new_n1042 & new_n1043;
  assign new_n1045 = ~new_n775 & new_n1044;
  assign new_n1046 = ~pt3 & new_n1045;
  assign new_n1047 = pt3 & ~new_n1045;
  assign new_n1048 = ~new_n1046 & ~new_n1047;
  assign new_n1049 = new_n738 & ~new_n1048;
  assign pa9 = new_n1015 | new_n1049;
  assign new_n1051 = ~pp1 & ~pl;
  assign new_n1052 = pb2 & pc2;
  assign new_n1053 = pd2 & new_n1052;
  assign new_n1054 = pq1 & ~pl;
  assign new_n1055 = ~new_n1053 & ~new_n1054;
  assign new_n1056 = pg2 & ~new_n1055;
  assign new_n1057 = new_n1051 & ~new_n1056;
  assign new_n1058 = pe2 & ~new_n1057;
  assign new_n1059 = pf2 & new_n1058;
  assign new_n1060 = ~ph2 & new_n1059;
  assign new_n1061 = ph2 & ~new_n1059;
  assign new_n1062 = ~new_n1060 & ~new_n1061;
  assign new_n1063 = ~pu1 & new_n1062;
  assign new_n1064 = pe2 & pn2;
  assign new_n1065 = ~new_n1057 & new_n1064;
  assign new_n1066 = ~new_n313 & ~new_n1065;
  assign new_n1067 = new_n1062 & new_n1066;
  assign new_n1068 = ~pu1 & ~new_n1066;
  assign new_n1069 = ~new_n1063 & ~new_n1067;
  assign new_n1070 = ~new_n1068 & new_n1069;
  assign po7 = pb | new_n1070;
  assign new_n1072 = ~pq5 & new_n935;
  assign new_n1073 = ~pr5 & new_n938;
  assign new_n1074 = ~pr5 & new_n937;
  assign new_n1075 = ~pp5 & new_n1074;
  assign new_n1076 = ~pq5 & ~new_n937;
  assign new_n1077 = ~pp5 & new_n1076;
  assign new_n1078 = ~pp5 & new_n946;
  assign new_n1079 = ~pq5 & new_n948;
  assign new_n1080 = ~pq5 & ~new_n934;
  assign new_n1081 = ~pp5 & new_n1080;
  assign new_n1082 = ~new_n1072 & ~new_n1073;
  assign new_n1083 = ~new_n1075 & ~new_n1077;
  assign new_n1084 = new_n1082 & new_n1083;
  assign new_n1085 = ~new_n1079 & ~new_n1081;
  assign new_n1086 = ~new_n945 & ~new_n1078;
  assign new_n1087 = new_n1085 & new_n1086;
  assign new_n1088 = new_n1084 & new_n1087;
  assign py10 = ~new_n967 & new_n1088;
  assign new_n1090 = ~new_n423 & new_n450;
  assign new_n1091 = new_n423 & new_n459;
  assign new_n1092 = ~new_n1090 & ~new_n1091;
  assign new_n1093 = ~new_n441 & ~new_n1092;
  assign new_n1094 = ~pt2 & new_n1093;
  assign new_n1095 = pt2 & ~new_n1093;
  assign new_n1096 = ~new_n1094 & ~new_n1095;
  assign new_n1097 = new_n427 & ~new_n1096;
  assign pa8 = new_n428 | new_n1097;
  assign new_n1099 = ~pg2 & new_n1055;
  assign new_n1100 = ~new_n1056 & ~new_n1099;
  assign pn7 = pb | new_n1100;
  assign new_n1102 = ~pb & ~new_n313;
  assign new_n1103 = ~new_n323 & new_n1102;
  assign new_n1104 = ~ph1 & new_n1102;
  assign new_n1105 = ~new_n1103 & ~new_n1104;
  assign new_n1106 = ph1 & ~new_n1105;
  assign po6 = new_n329 | new_n1106;
  assign new_n1108 = ~pq5 & new_n934;
  assign new_n1109 = ~pp5 & new_n1108;
  assign new_n1110 = ~pq5 & new_n938;
  assign new_n1111 = ~pq5 & new_n1074;
  assign new_n1112 = ~pp5 & new_n942;
  assign new_n1113 = ~pr5 & new_n946;
  assign new_n1114 = ~pp5 & new_n948;
  assign new_n1115 = ~pp5 & new_n950;
  assign new_n1116 = ~new_n1109 & ~new_n1110;
  assign new_n1117 = ~new_n1111 & ~new_n1112;
  assign new_n1118 = new_n1116 & new_n1117;
  assign new_n1119 = ~new_n1114 & ~new_n1115;
  assign new_n1120 = ~new_n945 & ~new_n1113;
  assign new_n1121 = new_n1119 & new_n1120;
  assign new_n1122 = new_n1118 & new_n1121;
  assign px10 = ~new_n967 & new_n1122;
  assign new_n1124 = ~pz2 & ~px2;
  assign new_n1125 = ~pw2 & ~py2;
  assign new_n1126 = new_n1124 & new_n1125;
  assign new_n1127 = new_n423 & new_n1126;
  assign new_n1128 = new_n427 & new_n1126;
  assign new_n1129 = new_n423 & ~new_n427;
  assign new_n1130 = ~new_n1127 & ~new_n1128;
  assign pb8 = new_n1129 | ~new_n1130;
  assign new_n1132 = ~pu3 & ~new_n529;
  assign new_n1133 = pu3 & new_n529;
  assign new_n1134 = ~new_n1132 & ~new_n1133;
  assign new_n1135 = ~new_n515 & new_n1134;
  assign new_n1136 = ~pv3 & new_n1135;
  assign new_n1137 = pv3 & ~new_n1135;
  assign new_n1138 = ~new_n1136 & ~new_n1137;
  assign new_n1139 = ~new_n489 & new_n1138;
  assign new_n1140 = ~pm3 & new_n489;
  assign new_n1141 = ~pm3 & new_n1138;
  assign new_n1142 = ~new_n1139 & ~new_n1140;
  assign new_n1143 = ~new_n1141 & new_n1142;
  assign pc9 = ~pz & new_n1143;
  assign new_n1145 = ~pf2 & new_n1058;
  assign new_n1146 = pf2 & ~new_n1058;
  assign new_n1147 = ~new_n1145 & ~new_n1146;
  assign new_n1148 = ~pt1 & new_n1147;
  assign new_n1149 = new_n1066 & new_n1147;
  assign new_n1150 = ~pt1 & ~new_n1066;
  assign new_n1151 = ~new_n1148 & ~new_n1149;
  assign new_n1152 = ~new_n1150 & new_n1151;
  assign pm7 = pb | new_n1152;
  assign new_n1154 = ~pu3 & ~new_n515;
  assign new_n1155 = pu3 & new_n515;
  assign new_n1156 = ~new_n1154 & ~new_n1155;
  assign new_n1157 = ~new_n489 & new_n1156;
  assign new_n1158 = ~pl3 & new_n489;
  assign new_n1159 = ~pl3 & new_n1156;
  assign new_n1160 = ~new_n1157 & ~new_n1158;
  assign new_n1161 = ~new_n1159 & new_n1160;
  assign pb9 = ~pz & new_n1161;
  assign new_n1163 = pz2 & px2;
  assign new_n1164 = pw2 & py2;
  assign new_n1165 = new_n1163 & new_n1164;
  assign pc8 = new_n427 & new_n1165;
  assign new_n1167 = ~pe2 & ~new_n1057;
  assign new_n1168 = pe2 & new_n1057;
  assign new_n1169 = ~new_n1167 & ~new_n1168;
  assign new_n1170 = ~ps1 & new_n1169;
  assign new_n1171 = new_n1066 & new_n1169;
  assign new_n1172 = ~ps1 & ~new_n1066;
  assign new_n1173 = ~new_n1170 & ~new_n1171;
  assign new_n1174 = ~new_n1172 & new_n1173;
  assign pl7 = pb | new_n1174;
  assign new_n1176 = ~new_n423 & new_n452;
  assign new_n1177 = new_n452 & new_n461;
  assign new_n1178 = new_n423 & new_n461;
  assign new_n1179 = ~new_n1176 & ~new_n1177;
  assign new_n1180 = ~new_n1178 & new_n1179;
  assign new_n1181 = ~new_n441 & new_n1180;
  assign new_n1182 = ~pw2 & ~new_n1181;
  assign new_n1183 = pw2 & new_n1181;
  assign new_n1184 = ~new_n1182 & ~new_n1183;
  assign pd8 = new_n427 & new_n1184;
  assign new_n1186 = new_n529 & new_n532;
  assign new_n1187 = ~new_n529 & new_n541;
  assign new_n1188 = new_n532 & new_n541;
  assign new_n1189 = ~new_n1186 & ~new_n1187;
  assign new_n1190 = ~new_n1188 & new_n1189;
  assign new_n1191 = ~new_n515 & new_n1190;
  assign new_n1192 = ~px3 & new_n1191;
  assign new_n1193 = px3 & ~new_n1191;
  assign new_n1194 = ~new_n1192 & ~new_n1193;
  assign new_n1195 = ~new_n489 & new_n1194;
  assign new_n1196 = ~po3 & new_n489;
  assign new_n1197 = ~po3 & new_n1194;
  assign new_n1198 = ~new_n1195 & ~new_n1196;
  assign new_n1199 = ~new_n1197 & new_n1198;
  assign pe9 = pz | new_n1199;
  assign new_n1201 = pa1 & pb1;
  assign new_n1202 = pz0 & new_n1201;
  assign new_n1203 = ~new_n346 & new_n1202;
  assign new_n1204 = new_n587 & new_n1203;
  assign new_n1205 = ~pc1 & ~new_n1204;
  assign new_n1206 = pc1 & new_n1204;
  assign new_n1207 = ~new_n1205 & ~new_n1206;
  assign pj6 = new_n342 & new_n1207;
  assign new_n1209 = ~pd2 & ~new_n1052;
  assign new_n1210 = ~new_n1053 & ~new_n1209;
  assign pk7 = pb | new_n1210;
  assign new_n1212 = new_n529 & ~new_n530;
  assign new_n1213 = ~new_n529 & ~new_n539;
  assign new_n1214 = ~new_n530 & ~new_n539;
  assign new_n1215 = ~new_n1212 & ~new_n1213;
  assign new_n1216 = ~new_n1214 & new_n1215;
  assign new_n1217 = ~new_n515 & new_n1216;
  assign new_n1218 = ~pw3 & new_n1217;
  assign new_n1219 = pw3 & ~new_n1217;
  assign new_n1220 = ~new_n1218 & ~new_n1219;
  assign new_n1221 = ~new_n489 & new_n1220;
  assign new_n1222 = ~pn3 & new_n489;
  assign new_n1223 = ~pn3 & new_n1220;
  assign new_n1224 = ~new_n1221 & ~new_n1222;
  assign new_n1225 = ~new_n1223 & new_n1224;
  assign pd9 = ~pz & new_n1225;
  assign new_n1227 = pw2 & ~new_n452;
  assign new_n1228 = ~new_n423 & ~new_n1227;
  assign new_n1229 = ~pw2 & ~new_n461;
  assign new_n1230 = ~new_n1227 & ~new_n1229;
  assign new_n1231 = new_n423 & ~new_n1229;
  assign new_n1232 = ~new_n1228 & ~new_n1230;
  assign new_n1233 = ~new_n1231 & new_n1232;
  assign new_n1234 = ~new_n441 & new_n1233;
  assign new_n1235 = ~px2 & ~new_n1234;
  assign new_n1236 = px2 & new_n1234;
  assign new_n1237 = ~new_n1235 & ~new_n1236;
  assign pe8 = new_n427 & new_n1237;
  assign new_n1239 = ~pb2 & ~pc2;
  assign new_n1240 = ~new_n1052 & ~new_n1239;
  assign pj7 = pb | new_n1240;
  assign new_n1242 = pc1 & ~new_n346;
  assign new_n1243 = new_n587 & new_n1202;
  assign new_n1244 = new_n1242 & new_n1243;
  assign new_n1245 = pd1 & new_n1244;
  assign new_n1246 = ~pd1 & ~new_n1244;
  assign new_n1247 = ~new_n1245 & ~new_n1246;
  assign pk6 = new_n342 & new_n1247;
  assign new_n1249 = px2 & new_n1227;
  assign new_n1250 = ~new_n423 & ~new_n1249;
  assign new_n1251 = ~pw2 & ~px2;
  assign new_n1252 = ~new_n461 & new_n1251;
  assign new_n1253 = ~new_n1249 & ~new_n1252;
  assign new_n1254 = new_n423 & ~new_n1252;
  assign new_n1255 = ~new_n1250 & ~new_n1253;
  assign new_n1256 = ~new_n1254 & new_n1255;
  assign new_n1257 = ~new_n441 & new_n1256;
  assign new_n1258 = ~py2 & ~new_n1257;
  assign new_n1259 = py2 & new_n1257;
  assign new_n1260 = ~new_n1258 & ~new_n1259;
  assign pf8 = new_n427 & new_n1260;
  assign new_n1262 = ~py3 & ~px3;
  assign new_n1263 = ~new_n532 & new_n1262;
  assign new_n1264 = new_n529 & ~new_n1263;
  assign new_n1265 = px3 & ~new_n541;
  assign new_n1266 = py3 & new_n1265;
  assign new_n1267 = ~new_n529 & ~new_n1266;
  assign new_n1268 = ~new_n1263 & ~new_n1266;
  assign new_n1269 = ~new_n1264 & ~new_n1267;
  assign new_n1270 = ~new_n1268 & new_n1269;
  assign new_n1271 = ~new_n515 & new_n1270;
  assign new_n1272 = ~pz3 & new_n1271;
  assign new_n1273 = pz3 & ~new_n1271;
  assign new_n1274 = ~new_n1272 & ~new_n1273;
  assign new_n1275 = ~new_n489 & new_n1274;
  assign new_n1276 = ~pq3 & new_n489;
  assign new_n1277 = ~pq3 & new_n1274;
  assign new_n1278 = ~new_n1275 & ~new_n1276;
  assign new_n1279 = ~new_n1277 & new_n1278;
  assign pg9 = pz | new_n1279;
  assign new_n1281 = pz0 & ~new_n346;
  assign new_n1282 = new_n587 & new_n1281;
  assign new_n1283 = ~pa1 & ~new_n1282;
  assign new_n1284 = pa1 & new_n1282;
  assign new_n1285 = ~new_n1283 & ~new_n1284;
  assign ph6 = new_n342 & new_n1285;
  assign pi7 = ~pb2 | pb;
  assign new_n1288 = ~px3 & ~new_n532;
  assign new_n1289 = new_n529 & ~new_n1288;
  assign new_n1290 = ~new_n529 & ~new_n1265;
  assign new_n1291 = ~new_n1265 & ~new_n1288;
  assign new_n1292 = ~new_n1289 & ~new_n1290;
  assign new_n1293 = ~new_n1291 & new_n1292;
  assign new_n1294 = ~new_n515 & new_n1293;
  assign new_n1295 = ~py3 & new_n1294;
  assign new_n1296 = py3 & ~new_n1294;
  assign new_n1297 = ~new_n1295 & ~new_n1296;
  assign new_n1298 = ~new_n489 & new_n1297;
  assign new_n1299 = ~pp3 & new_n489;
  assign new_n1300 = ~pp3 & new_n1297;
  assign new_n1301 = ~new_n1298 & ~new_n1299;
  assign new_n1302 = ~new_n1300 & new_n1301;
  assign pf9 = pz | new_n1302;
  assign new_n1304 = px2 & ~new_n452;
  assign new_n1305 = pw2 & new_n1304;
  assign new_n1306 = py2 & new_n1305;
  assign new_n1307 = ~new_n423 & ~new_n1306;
  assign new_n1308 = ~px2 & new_n1125;
  assign new_n1309 = ~new_n461 & new_n1308;
  assign new_n1310 = ~new_n1306 & ~new_n1309;
  assign new_n1311 = new_n423 & ~new_n1309;
  assign new_n1312 = ~new_n1307 & ~new_n1310;
  assign new_n1313 = ~new_n1311 & new_n1312;
  assign new_n1314 = ~new_n441 & new_n1313;
  assign new_n1315 = ~pz2 & new_n1314;
  assign new_n1316 = pz2 & ~new_n1314;
  assign new_n1317 = ~new_n1315 & ~new_n1316;
  assign new_n1318 = new_n427 & ~new_n1317;
  assign pg8 = new_n428 | new_n1318;
  assign new_n1320 = pz1 & new_n389;
  assign new_n1321 = ~new_n390 & ~new_n1320;
  assign new_n1322 = ~py1 & ~pz1;
  assign new_n1323 = ~new_n398 & new_n1322;
  assign new_n1324 = ~new_n1320 & ~new_n1323;
  assign new_n1325 = new_n390 & ~new_n1323;
  assign new_n1326 = ~new_n1321 & ~new_n1324;
  assign new_n1327 = ~new_n1325 & new_n1326;
  assign new_n1328 = ~new_n381 & new_n1327;
  assign new_n1329 = ~pa2 & new_n1328;
  assign new_n1330 = pa2 & ~new_n1328;
  assign new_n1331 = ~new_n1329 & ~new_n1330;
  assign new_n1332 = ~pe3 & new_n1331;
  assign new_n1333 = ~new_n416 & new_n1331;
  assign new_n1334 = ~pe3 & new_n416;
  assign new_n1335 = ~new_n1332 & ~new_n1333;
  assign new_n1336 = ~new_n1334 & new_n1335;
  assign ph7 = pb | new_n1336;
  assign new_n1338 = pa1 & new_n1281;
  assign new_n1339 = new_n587 & new_n1338;
  assign new_n1340 = ~pb1 & ~new_n1339;
  assign new_n1341 = pb1 & new_n1339;
  assign new_n1342 = ~new_n1340 & ~new_n1341;
  assign pi6 = new_n342 & new_n1342;
  assign new_n1344 = pr4 & new_n565;
  assign new_n1345 = pr5 & new_n1344;
  assign new_n1346 = pv10 & new_n765;
  assign new_n1347 = new_n528 & new_n1346;
  assign new_n1348 = ~new_n922 & ~new_n1345;
  assign new_n1349 = ~pz & ~new_n1347;
  assign new_n1350 = new_n1348 & new_n1349;
  assign new_n1351 = ps4 & ~new_n874;
  assign new_n1352 = pr4 & new_n1351;
  assign new_n1353 = ~pt4 & ~new_n1352;
  assign new_n1354 = pt4 & new_n1352;
  assign new_n1355 = ~new_n1353 & ~new_n1354;
  assign pa10 = new_n1350 & new_n1355;
  assign new_n1357 = pp & py1;
  assign new_n1358 = pr & ps1;
  assign new_n1359 = pq & pv1;
  assign new_n1360 = ps & pl2;
  assign new_n1361 = ~new_n1357 & ~new_n1358;
  assign new_n1362 = ~new_n1359 & ~new_n1360;
  assign new_n1363 = new_n1361 & new_n1362;
  assign new_n1364 = py2 & pn;
  assign new_n1365 = pc3 & pm;
  assign new_n1366 = pr2 & po;
  assign new_n1367 = ~new_n1364 & ~new_n1365;
  assign new_n1368 = ~new_n1366 & new_n1367;
  assign new_n1369 = pt & ph2;
  assign new_n1370 = pb1 & pv;
  assign new_n1371 = pc2 & pu;
  assign new_n1372 = pw & pw0;
  assign new_n1373 = ~new_n1369 & ~new_n1370;
  assign new_n1374 = ~new_n1371 & ~new_n1372;
  assign new_n1375 = new_n1373 & new_n1374;
  assign new_n1376 = new_n1363 & new_n1368;
  assign pu5 = ~new_n1375 | ~new_n1376;
  assign new_n1378 = pj1 & new_n1065;
  assign new_n1379 = pp2 & ~new_n1378;
  assign new_n1380 = ~pa & new_n1378;
  assign new_n1381 = ~pa & pp2;
  assign new_n1382 = ~new_n1379 & ~new_n1380;
  assign pw7 = new_n1381 | ~new_n1382;
  assign new_n1384 = new_n912 & new_n1025;
  assign new_n1385 = ~new_n912 & new_n1037;
  assign new_n1386 = new_n1025 & new_n1037;
  assign new_n1387 = ~new_n1384 & ~new_n1385;
  assign new_n1388 = ~new_n1386 & new_n1387;
  assign new_n1389 = ~new_n775 & new_n1388;
  assign new_n1390 = ~pq3 & new_n1389;
  assign new_n1391 = pq3 & ~new_n1389;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = new_n738 & ~new_n1392;
  assign px8 = new_n1015 | new_n1393;
  assign new_n1395 = ~pr4 & new_n874;
  assign new_n1396 = pr4 & ~new_n874;
  assign new_n1397 = ~new_n1395 & ~new_n1396;
  assign py9 = new_n1350 & new_n1397;
  assign new_n1399 = pp & pz1;
  assign new_n1400 = pr & pt1;
  assign new_n1401 = pq & pw1;
  assign new_n1402 = ps & pm2;
  assign new_n1403 = ~new_n1399 & ~new_n1400;
  assign new_n1404 = ~new_n1401 & ~new_n1402;
  assign new_n1405 = new_n1403 & new_n1404;
  assign new_n1406 = pz2 & pn;
  assign new_n1407 = pd3 & pm;
  assign new_n1408 = ps2 & po;
  assign new_n1409 = ~new_n1406 & ~new_n1407;
  assign new_n1410 = ~new_n1408 & new_n1409;
  assign new_n1411 = pt & pi2;
  assign new_n1412 = pc1 & pv;
  assign new_n1413 = pu & pd2;
  assign new_n1414 = pw & px0;
  assign new_n1415 = ~new_n1411 & ~new_n1412;
  assign new_n1416 = ~new_n1413 & ~new_n1414;
  assign new_n1417 = new_n1415 & new_n1416;
  assign new_n1418 = new_n1405 & new_n1410;
  assign pt5 = ~new_n1417 | ~new_n1418;
  assign new_n1420 = ph2 & new_n1059;
  assign new_n1421 = pi2 & new_n1420;
  assign new_n1422 = pj2 & new_n1421;
  assign new_n1423 = ~pl & ~new_n1422;
  assign new_n1424 = pk2 & ~new_n1423;
  assign new_n1425 = pl2 & new_n1424;
  assign new_n1426 = pm2 & new_n1425;
  assign new_n1427 = ~po2 & new_n1426;
  assign new_n1428 = po2 & ~new_n1426;
  assign new_n1429 = ~new_n1427 & ~new_n1428;
  assign new_n1430 = ~pa2 & new_n1429;
  assign new_n1431 = new_n1066 & new_n1429;
  assign new_n1432 = ~pa2 & ~new_n1066;
  assign new_n1433 = ~new_n1430 & ~new_n1431;
  assign new_n1434 = ~new_n1432 & new_n1433;
  assign pv7 = pb | new_n1434;
  assign new_n1436 = pn1 & new_n311;
  assign new_n1437 = ~pl1 & new_n1436;
  assign new_n1438 = ~pd & ~new_n1437;
  assign new_n1439 = ~pr1 & new_n1438;
  assign new_n1440 = ~pp1 & new_n1439;
  assign new_n1441 = pn1 & new_n424;
  assign new_n1442 = pl1 & new_n1441;
  assign new_n1443 = ~pe & ~new_n1442;
  assign new_n1444 = new_n1438 & new_n1443;
  assign new_n1445 = ~pp1 & new_n1444;
  assign new_n1446 = ~pq1 & new_n1443;
  assign new_n1447 = ~pp1 & new_n1446;
  assign new_n1448 = ~pr1 & ~new_n1443;
  assign new_n1449 = ~pq1 & new_n1448;
  assign new_n1450 = ~pq1 & ~pr1;
  assign new_n1451 = ~pp1 & new_n1450;
  assign new_n1452 = ~new_n1438 & new_n1443;
  assign new_n1453 = ~pq1 & new_n1452;
  assign new_n1454 = new_n1438 & ~new_n1443;
  assign new_n1455 = ~pr1 & new_n1454;
  assign new_n1456 = ~pr1 & ~new_n1438;
  assign new_n1457 = ~pq1 & new_n1456;
  assign new_n1458 = ~new_n1440 & ~new_n1445;
  assign new_n1459 = ~new_n1447 & ~new_n1449;
  assign new_n1460 = new_n1458 & new_n1459;
  assign new_n1461 = ~new_n1455 & ~new_n1457;
  assign new_n1462 = ~new_n1451 & ~new_n1453;
  assign new_n1463 = new_n1461 & new_n1462;
  assign new_n1464 = new_n1460 & new_n1463;
  assign new_n1465 = ~pp1 & ~pr1;
  assign new_n1466 = ~new_n1450 & ~new_n1465;
  assign new_n1467 = ~new_n366 & new_n1466;
  assign new_n1468 = ~pb & ~new_n1467;
  assign new_n1469 = pr1 & new_n1468;
  assign new_n1470 = pq1 & new_n1468;
  assign new_n1471 = pp1 & new_n1468;
  assign new_n1472 = ~new_n1469 & ~new_n1470;
  assign new_n1473 = ~new_n1471 & new_n1472;
  assign pw6 = new_n1464 | new_n1473;
  assign new_n1475 = ~pc4 & ~new_n923;
  assign new_n1476 = ph4 & new_n925;
  assign new_n1477 = pj4 & new_n1476;
  assign new_n1478 = pk4 & new_n1477;
  assign new_n1479 = pl4 & new_n1478;
  assign new_n1480 = ~pj0 & ~new_n1479;
  assign new_n1481 = pm4 & ~new_n1480;
  assign new_n1482 = pn4 & new_n1481;
  assign new_n1483 = po4 & new_n1482;
  assign new_n1484 = ~pq4 & new_n1483;
  assign new_n1485 = pq4 & ~new_n1483;
  assign new_n1486 = ~new_n1484 & ~new_n1485;
  assign new_n1487 = new_n923 & new_n1486;
  assign new_n1488 = ~pc4 & new_n1486;
  assign new_n1489 = ~new_n1475 & ~new_n1487;
  assign new_n1490 = ~new_n1488 & new_n1489;
  assign px9 = pz | new_n1490;
  assign new_n1492 = new_n912 & ~new_n1026;
  assign new_n1493 = ~new_n912 & ~new_n1038;
  assign new_n1494 = ~new_n1026 & ~new_n1038;
  assign new_n1495 = ~new_n1492 & ~new_n1493;
  assign new_n1496 = ~new_n1494 & new_n1495;
  assign new_n1497 = ~new_n775 & new_n1496;
  assign new_n1498 = ~pr3 & ~new_n1497;
  assign new_n1499 = pr3 & new_n1497;
  assign new_n1500 = ~new_n1498 & ~new_n1499;
  assign py8 = new_n738 & new_n1500;
  assign new_n1502 = ~new_n874 & new_n880;
  assign new_n1503 = ~pv4 & ~new_n1502;
  assign new_n1504 = pv4 & new_n1502;
  assign new_n1505 = ~new_n1503 & ~new_n1504;
  assign pc10 = new_n1350 & new_n1505;
  assign new_n1507 = ~pm1 & ~new_n1442;
  assign new_n1508 = ~new_n316 & new_n1507;
  assign new_n1509 = new_n323 & new_n1507;
  assign new_n1510 = ~pn1 & ~new_n1442;
  assign new_n1511 = new_n323 & new_n1510;
  assign new_n1512 = ~pc3 & ~pe3;
  assign new_n1513 = ~pb3 & ~pd3;
  assign new_n1514 = new_n1512 & new_n1513;
  assign new_n1515 = ~pa3 & ~pz2;
  assign new_n1516 = py2 & new_n1515;
  assign new_n1517 = new_n1514 & new_n1516;
  assign new_n1518 = new_n1510 & new_n1517;
  assign new_n1519 = ~new_n316 & new_n1510;
  assign new_n1520 = new_n1507 & new_n1517;
  assign new_n1521 = ~new_n1508 & ~new_n1509;
  assign new_n1522 = ~new_n1511 & new_n1521;
  assign new_n1523 = ~new_n1518 & ~new_n1519;
  assign new_n1524 = ~new_n1520 & new_n1523;
  assign new_n1525 = new_n1522 & new_n1524;
  assign new_n1526 = new_n316 & new_n1517;
  assign new_n1527 = ~pd1 & ~new_n1245;
  assign new_n1528 = ~pc & new_n1527;
  assign new_n1529 = pr1 & ~new_n1245;
  assign new_n1530 = ~pc & new_n1529;
  assign new_n1531 = ~pd1 & ~pr1;
  assign new_n1532 = ~pc & new_n1531;
  assign new_n1533 = ~new_n1528 & ~new_n1530;
  assign new_n1534 = ~new_n1532 & new_n1533;
  assign new_n1535 = pv6 & new_n1534;
  assign new_n1536 = ~new_n1526 & ~new_n1535;
  assign new_n1537 = ~new_n426 & ~new_n1437;
  assign new_n1538 = new_n1536 & new_n1537;
  assign new_n1539 = ~new_n1525 & new_n1538;
  assign pt6 = ~pb & ~new_n1539;
  assign new_n1541 = ~pb & ~new_n1066;
  assign new_n1542 = pj2 & pi2;
  assign new_n1543 = pk2 & new_n1542;
  assign new_n1544 = pf2 & ph2;
  assign new_n1545 = pl2 & pm2;
  assign new_n1546 = po2 & new_n1545;
  assign new_n1547 = ~new_n1541 & new_n1543;
  assign new_n1548 = new_n1544 & new_n1547;
  assign pu7 = new_n1546 & new_n1548;
  assign new_n1550 = pp & pq1;
  assign new_n1551 = pr & pn1;
  assign new_n1552 = pq & ~new_n427;
  assign new_n1553 = ps & new_n1065;
  assign new_n1554 = ~new_n1550 & ~new_n1551;
  assign new_n1555 = ~new_n1552 & ~new_n1553;
  assign new_n1556 = new_n1554 & new_n1555;
  assign new_n1557 = pw2 & pn;
  assign new_n1558 = pm & new_n1517;
  assign new_n1559 = pc3 & pd3;
  assign new_n1560 = pe3 & new_n1559;
  assign new_n1561 = po & new_n1560;
  assign new_n1562 = ~new_n1557 & ~new_n1558;
  assign new_n1563 = ~new_n1561 & new_n1562;
  assign new_n1564 = pt & pe2;
  assign new_n1565 = pv & pz0;
  assign new_n1566 = pu & new_n441;
  assign new_n1567 = pw & pl1;
  assign new_n1568 = ~new_n1564 & ~new_n1565;
  assign new_n1569 = ~new_n1566 & ~new_n1567;
  assign new_n1570 = new_n1568 & new_n1569;
  assign new_n1571 = new_n1556 & new_n1563;
  assign pw5 = ~new_n1570 | ~new_n1571;
  assign new_n1573 = ~pr3 & new_n1026;
  assign new_n1574 = new_n912 & ~new_n1573;
  assign new_n1575 = ~new_n912 & ~new_n1039;
  assign new_n1576 = ~new_n1039 & ~new_n1573;
  assign new_n1577 = ~new_n1574 & ~new_n1575;
  assign new_n1578 = ~new_n1576 & new_n1577;
  assign new_n1579 = ~new_n775 & new_n1578;
  assign new_n1580 = ~ps3 & new_n1579;
  assign new_n1581 = ps3 & ~new_n1579;
  assign new_n1582 = ~new_n1580 & ~new_n1581;
  assign new_n1583 = new_n738 & ~new_n1582;
  assign pz8 = new_n1015 | new_n1583;
  assign new_n1585 = pt4 & new_n1351;
  assign new_n1586 = pr4 & new_n1585;
  assign new_n1587 = ~pu4 & ~new_n1586;
  assign new_n1588 = pu4 & new_n1586;
  assign new_n1589 = ~new_n1587 & ~new_n1588;
  assign pb10 = new_n1350 & new_n1589;
  assign new_n1591 = ~pm2 & new_n1425;
  assign new_n1592 = pm2 & ~new_n1425;
  assign new_n1593 = ~new_n1591 & ~new_n1592;
  assign new_n1594 = ~pz1 & new_n1593;
  assign new_n1595 = new_n1066 & new_n1593;
  assign new_n1596 = ~pz1 & ~new_n1066;
  assign new_n1597 = ~new_n1594 & ~new_n1595;
  assign new_n1598 = ~new_n1596 & new_n1597;
  assign pt7 = pb | new_n1598;
  assign new_n1600 = ~new_n1442 & ~new_n1560;
  assign new_n1601 = ~new_n323 & ~new_n1442;
  assign new_n1602 = ~new_n1442 & new_n1517;
  assign new_n1603 = ~new_n316 & ~new_n1442;
  assign new_n1604 = ~new_n1600 & ~new_n1601;
  assign new_n1605 = ~new_n1602 & ~new_n1603;
  assign new_n1606 = new_n1604 & new_n1605;
  assign new_n1607 = ~new_n410 & ~new_n1437;
  assign new_n1608 = ~new_n1517 & new_n1607;
  assign new_n1609 = ~new_n316 & new_n1607;
  assign new_n1610 = ~new_n1608 & ~new_n1609;
  assign new_n1611 = ~new_n1606 & ~new_n1610;
  assign pu6 = ~pb & ~new_n1611;
  assign new_n1613 = pp & pp1;
  assign new_n1614 = pr & pm1;
  assign new_n1615 = pq & pr1;
  assign new_n1616 = ps & pk2;
  assign new_n1617 = ~new_n1613 & ~new_n1614;
  assign new_n1618 = ~new_n1615 & ~new_n1616;
  assign new_n1619 = new_n1617 & new_n1618;
  assign new_n1620 = px2 & pn;
  assign new_n1621 = pb3 & pm;
  assign new_n1622 = pq2 & po;
  assign new_n1623 = ~new_n1620 & ~new_n1621;
  assign new_n1624 = ~new_n1622 & new_n1623;
  assign new_n1625 = pf2 & pt;
  assign new_n1626 = pa1 & pv;
  assign new_n1627 = pb2 & pu;
  assign new_n1628 = pw & pv0;
  assign new_n1629 = ~new_n1625 & ~new_n1626;
  assign new_n1630 = ~new_n1627 & ~new_n1628;
  assign new_n1631 = new_n1629 & new_n1630;
  assign new_n1632 = new_n1619 & new_n1624;
  assign pv5 = ~new_n1631 | ~new_n1632;
  assign new_n1634 = ~ps4 & ~new_n1396;
  assign new_n1635 = ps4 & new_n1396;
  assign new_n1636 = ~new_n1634 & ~new_n1635;
  assign pz9 = new_n1350 & new_n1636;
  assign new_n1638 = pv4 & ~new_n874;
  assign new_n1639 = pw4 & new_n1638;
  assign new_n1640 = new_n880 & new_n1639;
  assign new_n1641 = ~px4 & ~new_n1640;
  assign new_n1642 = px4 & new_n1640;
  assign new_n1643 = ~new_n1641 & ~new_n1642;
  assign pe10 = new_n1350 & new_n1643;
  assign new_n1645 = ~pl2 & new_n1424;
  assign new_n1646 = pl2 & ~new_n1424;
  assign new_n1647 = ~new_n1645 & ~new_n1646;
  assign new_n1648 = ~py1 & new_n1647;
  assign new_n1649 = new_n1066 & new_n1647;
  assign new_n1650 = ~py1 & ~new_n1066;
  assign new_n1651 = ~new_n1648 & ~new_n1649;
  assign new_n1652 = ~new_n1650 & new_n1651;
  assign ps7 = pb | new_n1652;
  assign new_n1654 = new_n880 & new_n1638;
  assign new_n1655 = ~pw4 & ~new_n1654;
  assign new_n1656 = pw4 & new_n1654;
  assign new_n1657 = ~new_n1655 & ~new_n1656;
  assign pd10 = new_n1350 & new_n1657;
  assign new_n1659 = ~pk2 & ~new_n1423;
  assign new_n1660 = pk2 & new_n1423;
  assign new_n1661 = ~new_n1659 & ~new_n1660;
  assign new_n1662 = ~px1 & new_n1661;
  assign new_n1663 = new_n1066 & new_n1661;
  assign new_n1664 = ~px1 & ~new_n1066;
  assign new_n1665 = ~new_n1662 & ~new_n1663;
  assign new_n1666 = ~new_n1664 & new_n1665;
  assign pr7 = pb | new_n1666;
  assign new_n1668 = new_n323 & new_n426;
  assign new_n1669 = new_n323 & new_n1560;
  assign new_n1670 = ~new_n1517 & new_n1669;
  assign new_n1671 = new_n316 & ~new_n1670;
  assign new_n1672 = ~new_n410 & ~new_n1668;
  assign new_n1673 = ~new_n1671 & new_n1672;
  assign ps6 = ~pb & ~new_n1673;
  assign new_n1675 = ~pz4 & ~new_n882;
  assign new_n1676 = ~new_n883 & ~new_n1675;
  assign pg10 = new_n1350 & new_n1676;
  assign new_n1678 = ~pi1 & new_n1102;
  assign new_n1679 = ~new_n322 & new_n1102;
  assign new_n1680 = ~new_n1678 & ~new_n1679;
  assign new_n1681 = pi1 & ~new_n1680;
  assign pp6 = new_n335 | new_n1681;
  assign new_n1683 = ~pj2 & new_n1421;
  assign new_n1684 = pj2 & ~new_n1421;
  assign new_n1685 = ~new_n1683 & ~new_n1684;
  assign new_n1686 = ~pw1 & new_n1685;
  assign new_n1687 = new_n1066 & new_n1685;
  assign new_n1688 = ~pw1 & ~new_n1066;
  assign new_n1689 = ~new_n1686 & ~new_n1687;
  assign new_n1690 = ~new_n1688 & new_n1689;
  assign pq7 = pb | new_n1690;
  assign new_n1692 = pp & pa2;
  assign new_n1693 = pr & pu1;
  assign new_n1694 = pq & px1;
  assign new_n1695 = ps & po2;
  assign new_n1696 = ~new_n1692 & ~new_n1693;
  assign new_n1697 = ~new_n1694 & ~new_n1695;
  assign new_n1698 = new_n1696 & new_n1697;
  assign new_n1699 = pa3 & pn;
  assign new_n1700 = pe3 & pm;
  assign new_n1701 = pt2 & po;
  assign new_n1702 = ~new_n1699 & ~new_n1700;
  assign new_n1703 = ~new_n1701 & new_n1702;
  assign new_n1704 = pt & pj2;
  assign new_n1705 = pd1 & pv;
  assign new_n1706 = pg2 & pu;
  assign new_n1707 = pw & py0;
  assign new_n1708 = ~new_n1704 & ~new_n1705;
  assign new_n1709 = ~new_n1706 & ~new_n1707;
  assign new_n1710 = new_n1708 & new_n1709;
  assign new_n1711 = new_n1698 & new_n1703;
  assign ps5 = ~new_n1710 | ~new_n1711;
  assign new_n1713 = ~new_n874 & new_n877;
  assign new_n1714 = new_n880 & new_n1713;
  assign new_n1715 = ~py4 & ~new_n1714;
  assign new_n1716 = py4 & new_n1714;
  assign new_n1717 = ~new_n1715 & ~new_n1716;
  assign pf10 = new_n1350 & new_n1717;
  assign new_n1719 = ~pi2 & new_n1420;
  assign new_n1720 = pi2 & ~new_n1420;
  assign new_n1721 = ~new_n1719 & ~new_n1720;
  assign new_n1722 = ~pv1 & new_n1721;
  assign new_n1723 = new_n1066 & new_n1721;
  assign new_n1724 = ~pv1 & ~new_n1066;
  assign new_n1725 = ~new_n1722 & ~new_n1723;
  assign new_n1726 = ~new_n1724 & new_n1725;
  assign pp7 = pb | new_n1726;
  assign new_n1728 = ~new_n313 & ~new_n410;
  assign new_n1729 = ~pj1 & ~new_n1065;
  assign new_n1730 = ~new_n1378 & ~new_n1729;
  assign new_n1731 = ~pb & new_n1730;
  assign pq6 = ~new_n1728 | new_n1731;
  assign new_n1733 = ~new_n912 & new_n1032;
  assign new_n1734 = new_n912 & new_n1020;
  assign new_n1735 = ~new_n1733 & ~new_n1734;
  assign new_n1736 = ~new_n775 & ~new_n1735;
  assign new_n1737 = ~pi3 & new_n1736;
  assign new_n1738 = pi3 & ~new_n1736;
  assign new_n1739 = ~new_n1737 & ~new_n1738;
  assign new_n1740 = new_n738 & ~new_n1739;
  assign pp8 = new_n1015 | new_n1740;
  assign new_n1742 = ~pw3 & ~new_n923;
  assign new_n1743 = ~pj4 & new_n1476;
  assign new_n1744 = pj4 & ~new_n1476;
  assign new_n1745 = ~new_n1743 & ~new_n1744;
  assign new_n1746 = new_n923 & new_n1745;
  assign new_n1747 = ~pw3 & new_n1745;
  assign new_n1748 = ~new_n1742 & ~new_n1746;
  assign new_n1749 = ~new_n1747 & new_n1748;
  assign pq9 = pz | new_n1749;
  assign new_n1751 = ~pi4 & new_n744;
  assign new_n1752 = ~new_n745 & ~new_n1751;
  assign pp9 = pz | new_n1752;
  assign new_n1754 = ~po3 & ~pm3;
  assign new_n1755 = ~pn3 & ~pl3;
  assign new_n1756 = new_n1754 & new_n1755;
  assign new_n1757 = new_n738 & new_n1756;
  assign new_n1758 = ~new_n738 & new_n912;
  assign new_n1759 = new_n912 & new_n1756;
  assign new_n1760 = ~new_n1757 & ~new_n1758;
  assign pq8 = new_n1759 | ~new_n1760;
  assign new_n1762 = ~pz & ~new_n922;
  assign new_n1763 = ~new_n520 & new_n1762;
  assign new_n1764 = ~pd5 & new_n1762;
  assign new_n1765 = ~new_n1763 & ~new_n1764;
  assign new_n1766 = pd5 & ~new_n1765;
  assign pk10 = new_n764 | new_n1766;
  assign new_n1768 = po3 & pm3;
  assign new_n1769 = pn3 & pl3;
  assign new_n1770 = new_n1768 & new_n1769;
  assign pr8 = new_n738 & new_n1770;
  assign new_n1772 = ~py3 & ~new_n923;
  assign new_n1773 = ~pl4 & new_n1478;
  assign new_n1774 = pl4 & ~new_n1478;
  assign new_n1775 = ~new_n1773 & ~new_n1774;
  assign new_n1776 = new_n923 & new_n1775;
  assign new_n1777 = ~py3 & new_n1775;
  assign new_n1778 = ~new_n1772 & ~new_n1776;
  assign new_n1779 = ~new_n1777 & new_n1778;
  assign ps9 = pz | new_n1779;
  assign new_n1781 = ~px3 & ~new_n923;
  assign new_n1782 = ~pk4 & new_n1477;
  assign new_n1783 = pk4 & ~new_n1477;
  assign new_n1784 = ~new_n1782 & ~new_n1783;
  assign new_n1785 = new_n923 & new_n1784;
  assign new_n1786 = ~px3 & new_n1784;
  assign new_n1787 = ~new_n1781 & ~new_n1785;
  assign new_n1788 = ~new_n1786 & new_n1787;
  assign pr9 = pz | new_n1788;
  assign new_n1790 = new_n912 & new_n1022;
  assign new_n1791 = ~new_n912 & new_n1034;
  assign new_n1792 = new_n1022 & new_n1034;
  assign new_n1793 = ~new_n1790 & ~new_n1791;
  assign new_n1794 = ~new_n1792 & new_n1793;
  assign new_n1795 = ~new_n775 & new_n1794;
  assign new_n1796 = ~pl3 & ~new_n1795;
  assign new_n1797 = pl3 & new_n1795;
  assign new_n1798 = ~new_n1796 & ~new_n1797;
  assign ps8 = new_n738 & new_n1798;
  assign new_n1800 = ~new_n475 & ~new_n922;
  assign new_n1801 = ~pg5 & ~pf5;
  assign new_n1802 = ~pf5 & ~new_n1801;
  assign new_n1803 = ~pz & new_n1802;
  assign new_n1804 = ~ph5 & ~new_n748;
  assign new_n1805 = ph5 & new_n748;
  assign new_n1806 = ~new_n1804 & ~new_n1805;
  assign new_n1807 = ~pz & new_n1806;
  assign po10 = ~new_n1800 | new_n1807;
  assign new_n1809 = ~ph5 & po10;
  assign new_n1810 = ~new_n1801 & new_n1809;
  assign new_n1811 = ~pz & new_n1810;
  assign new_n1812 = ~pf5 & ~new_n1809;
  assign new_n1813 = ~pz & new_n1812;
  assign new_n1814 = ~new_n1803 & ~new_n1811;
  assign new_n1815 = ~new_n1813 & new_n1814;
  assign pm10 = new_n1800 & new_n1815;
  assign new_n1817 = ~pl3 & ~new_n1022;
  assign new_n1818 = new_n912 & ~new_n1817;
  assign new_n1819 = pl3 & ~new_n1034;
  assign new_n1820 = ~new_n912 & ~new_n1819;
  assign new_n1821 = ~new_n1817 & ~new_n1819;
  assign new_n1822 = ~new_n1818 & ~new_n1820;
  assign new_n1823 = ~new_n1821 & new_n1822;
  assign new_n1824 = ~new_n775 & new_n1823;
  assign new_n1825 = ~pm3 & ~new_n1824;
  assign new_n1826 = pm3 & new_n1824;
  assign new_n1827 = ~new_n1825 & ~new_n1826;
  assign pt8 = new_n738 & new_n1827;
  assign new_n1829 = ~pa4 & ~new_n923;
  assign new_n1830 = ~pn4 & new_n1481;
  assign new_n1831 = pn4 & ~new_n1481;
  assign new_n1832 = ~new_n1830 & ~new_n1831;
  assign new_n1833 = new_n923 & new_n1832;
  assign new_n1834 = ~pa4 & new_n1832;
  assign new_n1835 = ~new_n1829 & ~new_n1833;
  assign new_n1836 = ~new_n1834 & new_n1835;
  assign pu9 = pz | new_n1836;
  assign new_n1838 = pb4 & pn0;
  assign new_n1839 = pp0 & pv3;
  assign new_n1840 = po0 & py3;
  assign new_n1841 = po4 & pq0;
  assign new_n1842 = ~new_n1838 & ~new_n1839;
  assign new_n1843 = ~new_n1840 & ~new_n1841;
  assign new_n1844 = new_n1842 & new_n1843;
  assign new_n1845 = pl0 & po3;
  assign new_n1846 = pk0 & ps3;
  assign new_n1847 = ph3 & pm0;
  assign new_n1848 = ~new_n1845 & ~new_n1846;
  assign new_n1849 = ~new_n1847 & new_n1848;
  assign new_n1850 = pk4 & pr0;
  assign new_n1851 = pt0 & py4;
  assign new_n1852 = pf4 & ps0;
  assign new_n1853 = pt4 & pu0;
  assign new_n1854 = ~new_n1850 & ~new_n1851;
  assign new_n1855 = ~new_n1852 & ~new_n1853;
  assign new_n1856 = new_n1854 & new_n1855;
  assign new_n1857 = new_n1844 & new_n1849;
  assign py5 = ~new_n1856 | ~new_n1857;
  assign new_n1859 = ~ps1 & ~new_n381;
  assign new_n1860 = ps1 & new_n381;
  assign new_n1861 = ~new_n1859 & ~new_n1860;
  assign new_n1862 = ~pw2 & new_n1861;
  assign new_n1863 = ~new_n416 & new_n1861;
  assign new_n1864 = ~pw2 & new_n416;
  assign new_n1865 = ~new_n1862 & ~new_n1863;
  assign new_n1866 = ~new_n1864 & new_n1865;
  assign pz6 = ~pb & new_n1866;
  assign new_n1868 = ~pe5 & new_n1762;
  assign new_n1869 = ~new_n519 & new_n1762;
  assign new_n1870 = ~new_n1868 & ~new_n1869;
  assign new_n1871 = pe5 & ~new_n1870;
  assign pl10 = new_n526 | new_n1871;
  assign new_n1873 = ~pz3 & ~new_n923;
  assign new_n1874 = ~pm4 & ~new_n1480;
  assign new_n1875 = pm4 & new_n1480;
  assign new_n1876 = ~new_n1874 & ~new_n1875;
  assign new_n1877 = new_n923 & new_n1876;
  assign new_n1878 = ~pz3 & new_n1876;
  assign new_n1879 = ~new_n1873 & ~new_n1877;
  assign new_n1880 = ~new_n1878 & new_n1879;
  assign pt9 = pz | new_n1880;
  assign new_n1882 = ~pm3 & ~pl3;
  assign new_n1883 = ~new_n1022 & new_n1882;
  assign new_n1884 = new_n912 & ~new_n1883;
  assign new_n1885 = pm3 & new_n1819;
  assign new_n1886 = ~new_n912 & ~new_n1885;
  assign new_n1887 = ~new_n1883 & ~new_n1885;
  assign new_n1888 = ~new_n1884 & ~new_n1886;
  assign new_n1889 = ~new_n1887 & new_n1888;
  assign new_n1890 = ~new_n775 & new_n1889;
  assign new_n1891 = ~pn3 & ~new_n1890;
  assign new_n1892 = pn3 & new_n1890;
  assign new_n1893 = ~new_n1891 & ~new_n1892;
  assign pu8 = new_n738 & new_n1893;
  assign new_n1895 = pc4 & pn0;
  assign new_n1896 = pp0 & pw3;
  assign new_n1897 = po0 & pz3;
  assign new_n1898 = pq0 & pq4;
  assign new_n1899 = ~new_n1895 & ~new_n1896;
  assign new_n1900 = ~new_n1897 & ~new_n1898;
  assign new_n1901 = new_n1899 & new_n1900;
  assign new_n1902 = pl0 & pp3;
  assign new_n1903 = pk0 & pt3;
  assign new_n1904 = pi3 & pm0;
  assign new_n1905 = ~new_n1902 & ~new_n1903;
  assign new_n1906 = ~new_n1904 & new_n1905;
  assign new_n1907 = pl4 & pr0;
  assign new_n1908 = pt0 & pz4;
  assign new_n1909 = pi4 & ps0;
  assign new_n1910 = pu4 & pu0;
  assign new_n1911 = ~new_n1907 & ~new_n1908;
  assign new_n1912 = ~new_n1909 & ~new_n1910;
  assign new_n1913 = new_n1911 & new_n1912;
  assign new_n1914 = new_n1901 & new_n1906;
  assign px5 = ~new_n1913 | ~new_n1914;
  assign new_n1916 = ~new_n423 & new_n447;
  assign new_n1917 = new_n447 & new_n456;
  assign new_n1918 = new_n423 & new_n456;
  assign new_n1919 = ~new_n1916 & ~new_n1917;
  assign new_n1920 = ~new_n1918 & new_n1919;
  assign new_n1921 = ~new_n441 & new_n1920;
  assign new_n1922 = ~ps2 & ~new_n1921;
  assign new_n1923 = ps2 & new_n1921;
  assign new_n1924 = ~new_n1922 & ~new_n1923;
  assign pz7 = new_n427 & new_n1924;
  assign new_n1926 = ~pm3 & new_n1755;
  assign new_n1927 = ~new_n1022 & new_n1926;
  assign new_n1928 = new_n912 & ~new_n1927;
  assign new_n1929 = pm3 & ~new_n1034;
  assign new_n1930 = pl3 & new_n1929;
  assign new_n1931 = pn3 & new_n1930;
  assign new_n1932 = ~new_n912 & ~new_n1931;
  assign new_n1933 = ~new_n1927 & ~new_n1931;
  assign new_n1934 = ~new_n1928 & ~new_n1932;
  assign new_n1935 = ~new_n1933 & new_n1934;
  assign new_n1936 = ~new_n775 & new_n1935;
  assign new_n1937 = ~po3 & new_n1936;
  assign new_n1938 = po3 & ~new_n1936;
  assign new_n1939 = ~new_n1937 & ~new_n1938;
  assign new_n1940 = new_n738 & ~new_n1939;
  assign pv8 = new_n1015 | new_n1940;
  assign new_n1942 = ~pz & ~new_n923;
  assign new_n1943 = pl4 & pk4;
  assign new_n1944 = pm4 & new_n1943;
  assign new_n1945 = ph4 & pj4;
  assign new_n1946 = pn4 & po4;
  assign new_n1947 = pq4 & new_n1946;
  assign new_n1948 = ~new_n1942 & new_n1944;
  assign new_n1949 = new_n1945 & new_n1948;
  assign pw9 = new_n1947 & new_n1949;
  assign new_n1951 = ~pq1 & new_n1438;
  assign new_n1952 = ~pp1 & new_n1951;
  assign new_n1953 = ~pq1 & new_n1444;
  assign new_n1954 = ~pr1 & new_n1443;
  assign new_n1955 = ~pq1 & new_n1954;
  assign new_n1956 = ~pp1 & new_n1448;
  assign new_n1957 = ~pr1 & new_n1452;
  assign new_n1958 = ~pp1 & new_n1454;
  assign new_n1959 = ~pp1 & new_n1456;
  assign new_n1960 = ~new_n1952 & ~new_n1953;
  assign new_n1961 = ~new_n1955 & ~new_n1956;
  assign new_n1962 = new_n1960 & new_n1961;
  assign new_n1963 = ~new_n1958 & ~new_n1959;
  assign new_n1964 = ~new_n1451 & ~new_n1957;
  assign new_n1965 = new_n1963 & new_n1964;
  assign new_n1966 = new_n1962 & new_n1965;
  assign px6 = ~new_n1473 & new_n1966;
  assign new_n1968 = ~pq2 & ~new_n423;
  assign new_n1969 = pq2 & new_n423;
  assign new_n1970 = ~new_n1968 & ~new_n1969;
  assign new_n1971 = ~new_n441 & new_n1970;
  assign new_n1972 = ~pr2 & ~new_n1971;
  assign new_n1973 = pr2 & new_n1971;
  assign new_n1974 = ~new_n1972 & ~new_n1973;
  assign py7 = new_n427 & new_n1974;
  assign new_n1976 = new_n1800 & ~new_n1809;
  assign new_n1977 = ~pg5 & new_n1976;
  assign new_n1978 = new_n1800 & new_n1809;
  assign new_n1979 = ~pf5 & new_n1978;
  assign new_n1980 = ~pg5 & new_n1800;
  assign new_n1981 = ~pf5 & new_n1980;
  assign new_n1982 = ~new_n1977 & ~new_n1979;
  assign new_n1983 = ~new_n1981 & new_n1982;
  assign pn10 = ~pz & new_n1983;
  assign new_n1985 = ~pb4 & ~new_n923;
  assign new_n1986 = ~po4 & new_n1482;
  assign new_n1987 = po4 & ~new_n1482;
  assign new_n1988 = ~new_n1986 & ~new_n1987;
  assign new_n1989 = new_n923 & new_n1988;
  assign new_n1990 = ~pb4 & new_n1988;
  assign new_n1991 = ~new_n1985 & ~new_n1989;
  assign new_n1992 = ~new_n1990 & new_n1991;
  assign pv9 = pz | new_n1992;
  assign new_n1994 = new_n912 & ~new_n1023;
  assign new_n1995 = ~new_n912 & ~new_n1035;
  assign new_n1996 = ~new_n1023 & ~new_n1035;
  assign new_n1997 = ~new_n1994 & ~new_n1995;
  assign new_n1998 = ~new_n1996 & new_n1997;
  assign new_n1999 = ~new_n775 & new_n1998;
  assign new_n2000 = ~pp3 & new_n1999;
  assign new_n2001 = pp3 & ~new_n1999;
  assign new_n2002 = ~new_n2000 & ~new_n2001;
  assign new_n2003 = new_n738 & ~new_n2002;
  assign pw8 = new_n1015 | new_n2003;
  assign new_n2005 = ~pq2 & new_n441;
  assign new_n2006 = pq2 & ~new_n441;
  assign new_n2007 = ~new_n2005 & ~new_n2006;
  assign px7 = new_n427 & new_n2007;
  assign new_n2009 = ~pq1 & new_n1439;
  assign new_n2010 = ~pr1 & new_n1444;
  assign new_n2011 = ~pp1 & new_n1954;
  assign new_n2012 = ~pq1 & ~new_n1443;
  assign new_n2013 = ~pp1 & new_n2012;
  assign new_n2014 = ~pp1 & new_n1452;
  assign new_n2015 = ~pq1 & new_n1454;
  assign new_n2016 = ~pq1 & ~new_n1438;
  assign new_n2017 = ~pp1 & new_n2016;
  assign new_n2018 = ~new_n2009 & ~new_n2010;
  assign new_n2019 = ~new_n2011 & ~new_n2013;
  assign new_n2020 = new_n2018 & new_n2019;
  assign new_n2021 = ~new_n2015 & ~new_n2017;
  assign new_n2022 = ~new_n1451 & ~new_n2014;
  assign new_n2023 = new_n2021 & new_n2022;
  assign new_n2024 = new_n2020 & new_n2023;
  assign py6 = ~new_n1473 & new_n2024;
  assign new_n2026 = pa4 & pn0;
  assign new_n2027 = pp0 & pu3;
  assign new_n2028 = po0 & px3;
  assign new_n2029 = pn4 & pq0;
  assign new_n2030 = ~new_n2026 & ~new_n2027;
  assign new_n2031 = ~new_n2028 & ~new_n2029;
  assign new_n2032 = new_n2030 & new_n2031;
  assign new_n2033 = pl0 & pn3;
  assign new_n2034 = pk0 & pr3;
  assign new_n2035 = pg3 & pm0;
  assign new_n2036 = ~new_n2033 & ~new_n2034;
  assign new_n2037 = ~new_n2035 & new_n2036;
  assign new_n2038 = pj4 & pr0;
  assign new_n2039 = pt0 & px4;
  assign new_n2040 = pe4 & ps0;
  assign new_n2041 = pu0 & ps4;
  assign new_n2042 = ~new_n2038 & ~new_n2039;
  assign new_n2043 = ~new_n2040 & ~new_n2041;
  assign new_n2044 = new_n2042 & new_n2043;
  assign new_n2045 = new_n2032 & new_n2037;
  assign pz5 = ~new_n2044 | ~new_n2045;
  assign pp10 = pg5;
  assign pl6 = pa;
  assign pm6 = pe1;
  assign pr6 = pj1;
  assign pi10 = pa5;
  assign ph10 = py;
endmodule


