// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_, o_3_  );
  input  i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_, o_3_;
  wire new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21,
    new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29,
    new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37,
    new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45,
    new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53,
    new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61,
    new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68, new_n69,
    new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76, new_n77,
    new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84, new_n85,
    new_n86, new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n101, new_n102, new_n103, new_n104, new_n105, new_n106, new_n107,
    new_n108, new_n109, new_n110, new_n111, new_n112, new_n113, new_n115,
    new_n116, new_n117, new_n118, new_n119, new_n120, new_n121, new_n122,
    new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277;
  assign new_n15 = ~i_5_ & i_4_;
  assign new_n16 = i_3_ & new_n15;
  assign new_n17 = i_7_ & ~i_8_;
  assign new_n18 = i_6_ & new_n17;
  assign new_n19 = i_1_ & i_2_;
  assign new_n20 = i_0_ & new_n19;
  assign new_n21 = new_n16 & new_n18;
  assign new_n22 = new_n20 & new_n21;
  assign new_n23 = ~i_9_ & new_n22;
  assign new_n24 = ~i_5_ & ~i_4_;
  assign new_n25 = i_3_ & new_n24;
  assign new_n26 = i_7_ & i_8_;
  assign new_n27 = i_6_ & new_n26;
  assign new_n28 = new_n25 & new_n27;
  assign new_n29 = new_n20 & new_n28;
  assign new_n30 = ~i_9_ & new_n29;
  assign new_n31 = i_1_ & ~i_2_;
  assign new_n32 = i_0_ & new_n31;
  assign new_n33 = new_n16 & new_n27;
  assign new_n34 = new_n32 & new_n33;
  assign new_n35 = ~i_9_ & new_n34;
  assign new_n36 = ~new_n23 & ~new_n30;
  assign new_n37 = ~new_n35 & new_n36;
  assign new_n38 = ~i_0_ & new_n31;
  assign new_n39 = new_n28 & new_n38;
  assign new_n40 = ~i_9_ & new_n39;
  assign new_n41 = ~i_6_ & new_n17;
  assign new_n42 = ~i_1_ & i_2_;
  assign new_n43 = i_0_ & new_n42;
  assign new_n44 = new_n16 & new_n41;
  assign new_n45 = new_n43 & new_n44;
  assign new_n46 = ~i_9_ & new_n45;
  assign new_n47 = ~i_6_ & new_n26;
  assign new_n48 = new_n16 & new_n47;
  assign new_n49 = new_n20 & new_n48;
  assign new_n50 = ~i_9_ & new_n49;
  assign new_n51 = ~new_n40 & ~new_n46;
  assign new_n52 = ~new_n50 & new_n51;
  assign new_n53 = ~i_3_ & new_n24;
  assign new_n54 = new_n41 & new_n53;
  assign new_n55 = new_n43 & new_n54;
  assign new_n56 = ~i_9_ & new_n55;
  assign new_n57 = new_n33 & new_n43;
  assign new_n58 = ~i_9_ & new_n57;
  assign new_n59 = ~i_0_ & new_n19;
  assign new_n60 = new_n33 & new_n59;
  assign new_n61 = ~i_9_ & new_n60;
  assign new_n62 = ~new_n56 & ~new_n58;
  assign new_n63 = ~new_n61 & new_n62;
  assign new_n64 = new_n37 & new_n52;
  assign new_n65 = new_n63 & new_n64;
  assign new_n66 = new_n25 & new_n41;
  assign new_n67 = new_n20 & new_n66;
  assign new_n68 = ~i_9_ & new_n67;
  assign new_n69 = new_n25 & new_n47;
  assign new_n70 = new_n32 & new_n69;
  assign new_n71 = ~i_9_ & new_n70;
  assign new_n72 = ~new_n68 & ~new_n71;
  assign new_n73 = ~i_1_ & ~i_2_;
  assign new_n74 = i_0_ & new_n73;
  assign new_n75 = new_n66 & new_n74;
  assign new_n76 = ~i_9_ & new_n75;
  assign new_n77 = ~i_3_ & new_n15;
  assign new_n78 = new_n27 & new_n77;
  assign new_n79 = new_n20 & new_n78;
  assign new_n80 = ~i_9_ & new_n79;
  assign new_n81 = new_n38 & new_n66;
  assign new_n82 = ~i_9_ & new_n81;
  assign new_n83 = ~new_n76 & ~new_n80;
  assign new_n84 = ~new_n82 & new_n83;
  assign new_n85 = ~i_7_ & i_8_;
  assign new_n86 = i_6_ & new_n85;
  assign new_n87 = new_n16 & new_n86;
  assign new_n88 = new_n20 & new_n87;
  assign new_n89 = ~i_9_ & new_n88;
  assign new_n90 = new_n38 & new_n87;
  assign new_n91 = ~i_9_ & new_n90;
  assign new_n92 = new_n18 & new_n77;
  assign new_n93 = new_n43 & new_n92;
  assign new_n94 = ~i_9_ & new_n93;
  assign new_n95 = ~new_n89 & ~new_n91;
  assign new_n96 = ~new_n94 & new_n95;
  assign new_n97 = ~i_7_ & ~i_8_;
  assign new_n98 = ~i_6_ & new_n97;
  assign new_n99 = ~i_0_ & new_n73;
  assign new_n100 = new_n25 & new_n98;
  assign new_n101 = new_n99 & new_n100;
  assign new_n102 = ~i_9_ & new_n101;
  assign new_n103 = ~i_6_ & new_n85;
  assign new_n104 = new_n25 & new_n103;
  assign new_n105 = new_n38 & new_n104;
  assign new_n106 = ~i_9_ & new_n105;
  assign new_n107 = new_n54 & new_n99;
  assign new_n108 = ~i_9_ & new_n107;
  assign new_n109 = ~new_n102 & ~new_n106;
  assign new_n110 = ~new_n108 & new_n109;
  assign new_n111 = new_n84 & new_n96;
  assign new_n112 = new_n110 & new_n111;
  assign new_n113 = new_n65 & new_n72;
  assign o_1_ = ~new_n112 | ~new_n113;
  assign new_n115 = ~i_9_ & ~i_7_;
  assign new_n116 = i_2_ & new_n24;
  assign new_n117 = new_n115 & new_n116;
  assign new_n118 = ~i_9_ & i_5_;
  assign new_n119 = ~i_6_ & i_4_;
  assign new_n120 = ~i_0_ & new_n119;
  assign new_n121 = ~i_9_ & new_n120;
  assign new_n122 = ~new_n117 & ~new_n118;
  assign new_n123 = ~new_n121 & new_n122;
  assign new_n124 = ~i_5_ & ~i_2_;
  assign new_n125 = i_0_ & new_n124;
  assign new_n126 = new_n115 & new_n125;
  assign new_n127 = ~i_9_ & ~i_8_;
  assign new_n128 = ~i_5_ & ~i_3_;
  assign new_n129 = i_1_ & new_n128;
  assign new_n130 = new_n127 & new_n129;
  assign new_n131 = ~i_3_ & new_n115;
  assign new_n132 = ~new_n126 & ~new_n130;
  assign new_n133 = ~new_n131 & new_n132;
  assign new_n134 = ~i_9_ & ~i_5_;
  assign new_n135 = ~i_3_ & i_1_;
  assign new_n136 = ~i_0_ & new_n135;
  assign new_n137 = new_n134 & new_n136;
  assign new_n138 = ~i_9_ & i_8_;
  assign new_n139 = ~i_7_ & ~i_5_;
  assign new_n140 = ~i_1_ & new_n139;
  assign new_n141 = new_n138 & new_n140;
  assign new_n142 = ~i_5_ & i_6_;
  assign new_n143 = ~i_2_ & new_n142;
  assign new_n144 = new_n127 & new_n143;
  assign new_n145 = ~new_n137 & ~new_n141;
  assign new_n146 = ~new_n144 & new_n145;
  assign new_n147 = new_n123 & new_n133;
  assign new_n148 = new_n146 & new_n147;
  assign new_n149 = ~i_9_ & ~i_6_;
  assign new_n150 = ~i_2_ & new_n15;
  assign new_n151 = new_n149 & new_n150;
  assign new_n152 = ~i_5_ & ~i_6_;
  assign new_n153 = ~i_1_ & new_n152;
  assign new_n154 = new_n138 & new_n153;
  assign new_n155 = ~i_4_ & new_n142;
  assign new_n156 = new_n127 & new_n155;
  assign new_n157 = ~i_4_ & i_2_;
  assign new_n158 = ~i_0_ & new_n157;
  assign new_n159 = new_n134 & new_n158;
  assign new_n160 = ~new_n154 & ~new_n156;
  assign new_n161 = ~new_n159 & new_n160;
  assign new_n162 = ~new_n151 & new_n161;
  assign new_n163 = i_4_ & new_n152;
  assign new_n164 = new_n115 & new_n163;
  assign new_n165 = ~i_1_ & new_n24;
  assign new_n166 = new_n138 & new_n165;
  assign new_n167 = ~i_1_ & new_n124;
  assign new_n168 = new_n138 & new_n167;
  assign new_n169 = ~new_n164 & ~new_n166;
  assign new_n170 = ~new_n168 & new_n169;
  assign new_n171 = ~i_3_ & ~i_2_;
  assign new_n172 = i_1_ & new_n171;
  assign new_n173 = new_n134 & new_n172;
  assign new_n174 = ~i_7_ & i_6_;
  assign new_n175 = ~i_5_ & new_n174;
  assign new_n176 = new_n127 & new_n175;
  assign new_n177 = ~i_5_ & ~i_1_;
  assign new_n178 = ~i_0_ & new_n177;
  assign new_n179 = new_n138 & new_n178;
  assign new_n180 = ~new_n173 & ~new_n176;
  assign new_n181 = ~new_n179 & new_n180;
  assign new_n182 = ~i_3_ & ~i_4_;
  assign new_n183 = i_1_ & new_n182;
  assign new_n184 = new_n134 & new_n183;
  assign new_n185 = ~i_0_ & new_n142;
  assign new_n186 = new_n127 & new_n185;
  assign new_n187 = ~i_6_ & ~i_3_;
  assign new_n188 = i_1_ & new_n187;
  assign new_n189 = ~i_9_ & new_n188;
  assign new_n190 = ~new_n184 & ~new_n186;
  assign new_n191 = ~new_n189 & new_n190;
  assign new_n192 = new_n170 & new_n181;
  assign new_n193 = new_n191 & new_n192;
  assign new_n194 = new_n148 & new_n162;
  assign o_2_ = ~new_n193 | ~new_n194;
  assign new_n196 = ~i_4_ & new_n152;
  assign new_n197 = i_7_ & new_n127;
  assign new_n198 = ~i_1_ & new_n171;
  assign new_n199 = new_n196 & new_n197;
  assign new_n200 = new_n198 & new_n199;
  assign new_n201 = new_n16 & new_n197;
  assign new_n202 = new_n43 & new_n201;
  assign new_n203 = ~i_6_ & new_n127;
  assign new_n204 = new_n25 & new_n203;
  assign new_n205 = new_n99 & new_n204;
  assign new_n206 = i_3_ & new_n152;
  assign new_n207 = new_n197 & new_n206;
  assign new_n208 = new_n20 & new_n207;
  assign new_n209 = ~new_n202 & ~new_n205;
  assign new_n210 = ~new_n208 & new_n209;
  assign new_n211 = ~i_9_ & i_7_;
  assign new_n212 = i_6_ & new_n211;
  assign new_n213 = new_n77 & new_n212;
  assign new_n214 = new_n43 & new_n213;
  assign new_n215 = i_4_ & new_n142;
  assign new_n216 = ~i_7_ & new_n138;
  assign new_n217 = i_3_ & i_1_;
  assign new_n218 = ~i_0_ & new_n217;
  assign new_n219 = new_n215 & new_n216;
  assign new_n220 = new_n218 & new_n219;
  assign new_n221 = ~i_7_ & new_n127;
  assign new_n222 = i_3_ & ~i_2_;
  assign new_n223 = ~i_0_ & new_n222;
  assign new_n224 = new_n196 & new_n221;
  assign new_n225 = new_n223 & new_n224;
  assign new_n226 = ~new_n214 & ~new_n220;
  assign new_n227 = ~new_n225 & new_n226;
  assign new_n228 = i_7_ & new_n138;
  assign new_n229 = i_1_ & new_n222;
  assign new_n230 = new_n155 & new_n228;
  assign new_n231 = new_n229 & new_n230;
  assign new_n232 = i_6_ & new_n138;
  assign new_n233 = new_n16 & new_n232;
  assign new_n234 = new_n38 & new_n233;
  assign new_n235 = i_0_ & new_n217;
  assign new_n236 = new_n196 & new_n228;
  assign new_n237 = new_n235 & new_n236;
  assign new_n238 = ~new_n231 & ~new_n234;
  assign new_n239 = ~new_n237 & new_n238;
  assign new_n240 = new_n210 & new_n227;
  assign new_n241 = new_n239 & new_n240;
  assign o_0_ = new_n200 | ~new_n241;
  assign new_n243 = new_n115 & new_n129;
  assign new_n244 = ~i_5_ & i_3_;
  assign new_n245 = ~i_0_ & new_n244;
  assign new_n246 = new_n149 & new_n245;
  assign new_n247 = i_3_ & ~i_4_;
  assign new_n248 = ~i_1_ & new_n247;
  assign new_n249 = new_n134 & new_n248;
  assign new_n250 = ~new_n243 & ~new_n246;
  assign new_n251 = ~new_n249 & new_n250;
  assign new_n252 = ~i_2_ & new_n244;
  assign new_n253 = new_n127 & new_n252;
  assign new_n254 = new_n77 & new_n149;
  assign new_n255 = new_n25 & new_n115;
  assign new_n256 = ~new_n253 & ~new_n254;
  assign new_n257 = ~new_n255 & new_n256;
  assign new_n258 = ~new_n117 & ~new_n141;
  assign new_n259 = ~new_n137 & new_n258;
  assign new_n260 = new_n251 & new_n257;
  assign new_n261 = new_n259 & new_n260;
  assign new_n262 = ~new_n154 & ~new_n159;
  assign new_n263 = ~new_n130 & new_n262;
  assign new_n264 = ~new_n151 & ~new_n156;
  assign new_n265 = ~new_n126 & ~new_n200;
  assign new_n266 = ~new_n56 & new_n265;
  assign new_n267 = new_n263 & new_n264;
  assign new_n268 = new_n266 & new_n267;
  assign new_n269 = ~new_n166 & ~new_n179;
  assign new_n270 = ~new_n164 & new_n269;
  assign new_n271 = ~new_n144 & ~new_n176;
  assign new_n272 = ~new_n173 & new_n271;
  assign new_n273 = ~new_n168 & ~new_n186;
  assign new_n274 = ~new_n184 & new_n273;
  assign new_n275 = new_n270 & new_n272;
  assign new_n276 = new_n274 & new_n275;
  assign new_n277 = new_n261 & new_n268;
  assign o_3_ = ~new_n276 | ~new_n277;
endmodule


