// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_,
    pv202_0_  );
  input  pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_;
  output pv202_0_;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378, new_n379, new_n380, new_n381, new_n382, new_n383, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433;
  assign new_n203 = ~pv190_1_ & ~pv188_30_;
  assign new_n204 = ~pv190_0_ & ~pv188_31_;
  assign new_n205 = new_n203 & new_n204;
  assign new_n206 = pv201_4_ & ~new_n205;
  assign new_n207 = pv201_5_ & new_n206;
  assign new_n208 = pv193_1_ & pv201_6_;
  assign new_n209 = pv201_7_ & new_n208;
  assign new_n210 = pv191_31_ & pv201_6_;
  assign new_n211 = pv201_7_ & new_n210;
  assign new_n212 = ~pv176_3_ & ~pv176_2_;
  assign new_n213 = ~pv176_6_ & ~pv176_4_;
  assign new_n214 = new_n212 & new_n213;
  assign new_n215 = ~pv176_5_ & ~pv176_9_;
  assign new_n216 = ~pv176_7_ & ~pv176_17_;
  assign new_n217 = new_n215 & new_n216;
  assign new_n218 = new_n214 & new_n217;
  assign new_n219 = ~pv176_13_ & ~pv176_15_;
  assign new_n220 = ~pv176_11_ & ~pv176_16_;
  assign new_n221 = new_n219 & new_n220;
  assign new_n222 = ~pv176_8_ & ~pv176_10_;
  assign new_n223 = ~pv176_12_ & ~pv176_14_;
  assign new_n224 = new_n222 & new_n223;
  assign new_n225 = new_n221 & new_n224;
  assign new_n226 = new_n218 & new_n225;
  assign new_n227 = pv201_2_ & ~new_n226;
  assign new_n228 = ~pv176_19_ & ~pv176_18_;
  assign new_n229 = ~pv176_22_ & ~pv176_20_;
  assign new_n230 = new_n228 & new_n229;
  assign new_n231 = ~pv176_21_ & ~pv176_25_;
  assign new_n232 = ~pv176_23_ & ~pv178_1_;
  assign new_n233 = new_n231 & new_n232;
  assign new_n234 = new_n230 & new_n233;
  assign new_n235 = ~pv176_31_ & ~pv176_29_;
  assign new_n236 = ~pv178_0_ & ~pv176_27_;
  assign new_n237 = new_n235 & new_n236;
  assign new_n238 = ~pv176_26_ & ~pv176_24_;
  assign new_n239 = ~pv176_30_ & ~pv176_28_;
  assign new_n240 = new_n238 & new_n239;
  assign new_n241 = new_n237 & new_n240;
  assign new_n242 = new_n234 & new_n241;
  assign new_n243 = pv201_3_ & ~new_n242;
  assign new_n244 = ~pv188_26_ & ~pv188_29_;
  assign new_n245 = ~pv188_27_ & ~pv188_28_;
  assign new_n246 = new_n244 & new_n245;
  assign new_n247 = pv201_4_ & ~new_n246;
  assign new_n248 = pv201_5_ & new_n247;
  assign new_n249 = pv201_7_ & pv193_1_;
  assign new_n250 = ~pv30_22_ & ~pv30_20_;
  assign new_n251 = ~pv30_18_ & ~pv30_16_;
  assign new_n252 = new_n250 & new_n251;
  assign new_n253 = ~pv30_14_ & ~pv30_10_;
  assign new_n254 = ~pv30_12_ & ~pv30_11_;
  assign new_n255 = new_n253 & new_n254;
  assign new_n256 = new_n252 & new_n255;
  assign new_n257 = ~pv62_1_ & ~pv30_13_;
  assign new_n258 = ~pv30_2_ & ~pv30_31_;
  assign new_n259 = new_n257 & new_n258;
  assign new_n260 = ~pv30_19_ & ~pv30_4_;
  assign new_n261 = ~pv30_6_ & ~pv30_21_;
  assign new_n262 = new_n260 & new_n261;
  assign new_n263 = new_n259 & new_n262;
  assign new_n264 = new_n256 & new_n263;
  assign new_n265 = ~pv30_9_ & ~pv30_17_;
  assign new_n266 = ~pv30_8_ & ~pv30_15_;
  assign new_n267 = new_n265 & new_n266;
  assign new_n268 = ~pv30_7_ & ~pv30_27_;
  assign new_n269 = ~pv30_29_ & ~pv30_5_;
  assign new_n270 = new_n268 & new_n269;
  assign new_n271 = new_n267 & new_n270;
  assign new_n272 = ~pv30_3_ & ~pv30_23_;
  assign new_n273 = ~pv62_0_ & ~pv30_25_;
  assign new_n274 = new_n272 & new_n273;
  assign new_n275 = ~pv30_26_ & ~pv30_24_;
  assign new_n276 = ~pv30_28_ & ~pv30_30_;
  assign new_n277 = new_n275 & new_n276;
  assign new_n278 = new_n274 & new_n277;
  assign new_n279 = new_n271 & new_n278;
  assign new_n280 = new_n264 & new_n279;
  assign new_n281 = ~pv201_0_ & ~new_n280;
  assign new_n282 = pv201_1_ & new_n281;
  assign new_n283 = pv193_0_ & pv201_6_;
  assign new_n284 = pv130_0_ & pv201_0_;
  assign new_n285 = ~pv126_20_ & ~pv126_22_;
  assign new_n286 = ~pv126_18_ & ~pv126_16_;
  assign new_n287 = new_n285 & new_n286;
  assign new_n288 = ~pv126_10_ & ~pv126_14_;
  assign new_n289 = ~pv126_12_ & ~pv126_11_;
  assign new_n290 = new_n288 & new_n289;
  assign new_n291 = new_n287 & new_n290;
  assign new_n292 = ~pv128_0_ & ~pv126_13_;
  assign new_n293 = ~pv126_31_ & ~pv126_2_;
  assign new_n294 = new_n292 & new_n293;
  assign new_n295 = ~pv126_19_ & ~pv126_4_;
  assign new_n296 = ~pv126_6_ & ~pv126_21_;
  assign new_n297 = new_n295 & new_n296;
  assign new_n298 = new_n294 & new_n297;
  assign new_n299 = new_n291 & new_n298;
  assign new_n300 = ~pv126_9_ & ~pv126_17_;
  assign new_n301 = ~pv126_8_ & ~pv126_15_;
  assign new_n302 = new_n300 & new_n301;
  assign new_n303 = ~pv126_7_ & ~pv126_27_;
  assign new_n304 = ~pv126_5_ & ~pv126_29_;
  assign new_n305 = new_n303 & new_n304;
  assign new_n306 = new_n302 & new_n305;
  assign new_n307 = ~pv126_23_ & ~pv126_3_;
  assign new_n308 = ~pv126_25_ & ~pv127_0_;
  assign new_n309 = new_n307 & new_n308;
  assign new_n310 = ~pv126_26_ & ~pv126_24_;
  assign new_n311 = ~pv126_28_ & ~pv126_30_;
  assign new_n312 = new_n310 & new_n311;
  assign new_n313 = new_n309 & new_n312;
  assign new_n314 = new_n306 & new_n313;
  assign new_n315 = new_n299 & new_n314;
  assign new_n316 = pv201_0_ & ~new_n315;
  assign new_n317 = pv201_1_ & new_n316;
  assign new_n318 = pv201_3_ & new_n227;
  assign new_n319 = pv201_7_ & new_n283;
  assign new_n320 = ~pv62_20_ & ~pv62_22_;
  assign new_n321 = ~pv62_16_ & ~pv62_18_;
  assign new_n322 = new_n320 & new_n321;
  assign new_n323 = ~pv62_10_ & ~pv62_14_;
  assign new_n324 = ~pv62_11_ & ~pv62_12_;
  assign new_n325 = new_n323 & new_n324;
  assign new_n326 = new_n322 & new_n325;
  assign new_n327 = ~pv64_0_ & ~pv62_13_;
  assign new_n328 = ~pv62_2_ & ~pv62_31_;
  assign new_n329 = new_n327 & new_n328;
  assign new_n330 = ~pv62_4_ & ~pv62_19_;
  assign new_n331 = ~pv62_6_ & ~pv62_21_;
  assign new_n332 = new_n330 & new_n331;
  assign new_n333 = new_n329 & new_n332;
  assign new_n334 = new_n326 & new_n333;
  assign new_n335 = ~pv62_17_ & ~pv62_9_;
  assign new_n336 = ~pv62_15_ & ~pv62_8_;
  assign new_n337 = new_n335 & new_n336;
  assign new_n338 = ~pv62_7_ & ~pv62_27_;
  assign new_n339 = ~pv62_5_ & ~pv62_29_;
  assign new_n340 = new_n338 & new_n339;
  assign new_n341 = new_n337 & new_n340;
  assign new_n342 = ~pv62_3_ & ~pv62_23_;
  assign new_n343 = ~pv63_0_ & ~pv62_25_;
  assign new_n344 = new_n342 & new_n343;
  assign new_n345 = ~pv62_26_ & ~pv62_24_;
  assign new_n346 = ~pv62_28_ & ~pv62_30_;
  assign new_n347 = new_n345 & new_n346;
  assign new_n348 = new_n344 & new_n347;
  assign new_n349 = new_n341 & new_n348;
  assign new_n350 = new_n334 & new_n349;
  assign new_n351 = ~pv201_0_ & ~new_n350;
  assign new_n352 = pv201_1_ & new_n351;
  assign new_n353 = pv201_5_ & ~new_n205;
  assign new_n354 = pv129_0_ & ~pv201_0_;
  assign new_n355 = ~pv94_20_ & ~pv94_22_;
  assign new_n356 = ~pv94_18_ & ~pv94_16_;
  assign new_n357 = new_n355 & new_n356;
  assign new_n358 = ~pv94_10_ & ~pv94_14_;
  assign new_n359 = ~pv94_11_ & ~pv94_12_;
  assign new_n360 = new_n358 & new_n359;
  assign new_n361 = new_n357 & new_n360;
  assign new_n362 = ~pv126_1_ & ~pv94_13_;
  assign new_n363 = ~pv94_31_ & ~pv94_2_;
  assign new_n364 = new_n362 & new_n363;
  assign new_n365 = ~pv94_4_ & ~pv94_19_;
  assign new_n366 = ~pv94_21_ & ~pv94_6_;
  assign new_n367 = new_n365 & new_n366;
  assign new_n368 = new_n364 & new_n367;
  assign new_n369 = new_n361 & new_n368;
  assign new_n370 = ~pv94_9_ & ~pv94_17_;
  assign new_n371 = ~pv94_8_ & ~pv94_15_;
  assign new_n372 = new_n370 & new_n371;
  assign new_n373 = ~pv94_7_ & ~pv94_27_;
  assign new_n374 = ~pv94_5_ & ~pv94_29_;
  assign new_n375 = new_n373 & new_n374;
  assign new_n376 = new_n372 & new_n375;
  assign new_n377 = ~pv94_3_ & ~pv94_23_;
  assign new_n378 = ~pv94_25_ & ~pv126_0_;
  assign new_n379 = new_n377 & new_n378;
  assign new_n380 = ~pv94_24_ & ~pv94_26_;
  assign new_n381 = ~pv94_30_ & ~pv94_28_;
  assign new_n382 = new_n380 & new_n381;
  assign new_n383 = new_n379 & new_n382;
  assign new_n384 = new_n376 & new_n383;
  assign new_n385 = new_n369 & new_n384;
  assign new_n386 = pv201_0_ & ~new_n385;
  assign new_n387 = pv201_1_ & new_n386;
  assign new_n388 = pv201_2_ & ~new_n242;
  assign new_n389 = pv201_3_ & new_n388;
  assign new_n390 = ~pv144_18_ & ~pv144_19_;
  assign new_n391 = ~pv144_20_ & ~pv144_22_;
  assign new_n392 = new_n390 & new_n391;
  assign new_n393 = ~pv144_25_ & ~pv144_21_;
  assign new_n394 = ~pv176_1_ & ~pv144_23_;
  assign new_n395 = new_n393 & new_n394;
  assign new_n396 = new_n392 & new_n395;
  assign new_n397 = ~pv144_29_ & ~pv144_31_;
  assign new_n398 = ~pv144_27_ & ~pv176_0_;
  assign new_n399 = new_n397 & new_n398;
  assign new_n400 = ~pv144_24_ & ~pv144_26_;
  assign new_n401 = ~pv144_28_ & ~pv144_30_;
  assign new_n402 = new_n400 & new_n401;
  assign new_n403 = new_n399 & new_n402;
  assign new_n404 = new_n396 & new_n403;
  assign new_n405 = pv201_2_ & ~new_n404;
  assign new_n406 = pv201_3_ & new_n405;
  assign new_n407 = ~pv188_25_ & ~pv188_22_;
  assign new_n408 = ~pv188_23_ & ~pv188_24_;
  assign new_n409 = new_n407 & new_n408;
  assign new_n410 = pv201_4_ & ~new_n409;
  assign new_n411 = pv201_5_ & new_n410;
  assign new_n412 = ~new_n406 & ~new_n411;
  assign new_n413 = ~new_n388 & new_n412;
  assign new_n414 = ~new_n354 & ~new_n387;
  assign new_n415 = ~new_n389 & new_n414;
  assign new_n416 = new_n413 & new_n415;
  assign new_n417 = ~new_n319 & ~new_n352;
  assign new_n418 = ~new_n353 & new_n417;
  assign new_n419 = ~new_n284 & ~new_n317;
  assign new_n420 = ~new_n318 & new_n419;
  assign new_n421 = new_n418 & new_n420;
  assign new_n422 = new_n416 & new_n421;
  assign new_n423 = ~new_n249 & ~new_n282;
  assign new_n424 = ~new_n283 & new_n423;
  assign new_n425 = ~new_n243 & ~new_n248;
  assign new_n426 = ~new_n247 & new_n425;
  assign new_n427 = new_n424 & new_n426;
  assign new_n428 = ~new_n208 & ~new_n211;
  assign new_n429 = ~new_n227 & new_n428;
  assign new_n430 = ~new_n206 & ~new_n207;
  assign new_n431 = ~new_n209 & new_n430;
  assign new_n432 = new_n429 & new_n431;
  assign new_n433 = new_n427 & new_n432;
  assign pv202_0_ = ~new_n422 | ~new_n433;
endmodule


