// Benchmark "top" written by ABC on Mon Nov 27 17:39:42 2023

module top ( 
    A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15,
    A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28, A29,
    A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42, A43,
    A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56, A57,
    A58, A59, A60, A61, A62, A63, A64, A65, A66, A67, A68, A69, A70, A71,
    A72, A73, A74, A75, A76, A77, A78, A79, A80, A81, A82, A83, A84, A85,
    A86, A87, A88, A89, A90, A91, A92, A93, A94, A95, A96, A97, A98, A99,
    A100, A101, A102, A103, A104, A105, A106, A107, A108, A109, A110, A111,
    A112, A113, A114, A115, A116, A117, A118, A119, A120, A121, A122, A123,
    A124, A125, A126, A127, A128, A129, A130, A131, A132, A133, A134, A135,
    A136, A137, A138, A139, A140, A141, A142, A143, A144, A145, A146, A147,
    A148, A149, A150, A151, A152, A153, A154, A155, A156, A157, A158, A159,
    A160, A161, A162, A163, A164, A165, A166, A167, A168, A169, A170, A171,
    A172, A173, A174, A175, A176, A177, A178, A179, A180, A181, A182, A183,
    A184, A185, A186, A187, A188, A189, A190, A191, A192, A193, A194, A195,
    A196, A197, A198, A199, A200, A201, A202, A203, A204, A205, A206, A207,
    A208, A209, A210, A211, A212, A213, A214, A215, A216, A217, A218, A219,
    A220, A221, A222, A223, A224, A225, A226, A227, A228, A229, A230, A231,
    A232, A233, A234, A235, A236, A237, A238, A239, A240, A241, A242, A243,
    A244, A245, A246, A247, A248, A249, A250, A251, A252, A253, A254, A255,
    A256, A257, A258, A259, A260, A261, A262, A263, A264, A265, A266, A267,
    A268, A269, A270, A271, A272, A273, A274, A275, A276, A277, A278, A279,
    A280, A281, A282, A283, A284, A285, A286, A287, A288, A289, A290, A291,
    A292, A293, A294, A295, A296, A297, A298, A299, A300, A301, A302, A303,
    A304, A305, A306, A307, A308, A309, A310, A311, A312, A313, A314, A315,
    A316, A317, A318, A319, A320, A321, A322, A323, A324, A325, A326, A327,
    A328, A329, A330, A331, A332, A333, A334, A335, A336, A337, A338, A339,
    A340, A341, A342, A343, A344, A345, A346, A347, A348, A349, A350, A351,
    A352, A353, A354, A355, A356, A357, A358, A359, A360, A361, A362, A363,
    A364, A365, A366, A367, A368, A369, A370, A371, A372, A373, A374, A375,
    A376, A377, A378, A379, A380, A381, A382, A383, A384, A385, A386, A387,
    A388, A389, A390, A391, A392, A393, A394, A395, A396, A397, A398, A399,
    A400, A401, A402, A403, A404, A405, A406, A407, A408, A409, A410, A411,
    A412, A413, A414, A415, A416, A417, A418, A419, A420, A421, A422, A423,
    A424, A425, A426, A427, A428, A429, A430, A431, A432, A433, A434, A435,
    A436, A437, A438, A439, A440, A441, A442, A443, A444, A445, A446, A447,
    A448, A449, A450, A451, A452, A453, A454, A455, A456, A457, A458, A459,
    A460, A461, A462, A463, A464, A465, A466, A467, A468, A469, A470, A471,
    A472, A473, A474, A475, A476, A477, A478, A479, A480, A481, A482, A483,
    A484, A485, A486, A487, A488, A489, A490, A491, A492, A493, A494, A495,
    A496, A497, A498, A499, A500, A501, A502, A503, A504, A505, A506, A507,
    A508, A509, A510, A511, A512, A513, A514, A515, A516, A517, A518, A519,
    A520, A521, A522, A523, A524, A525, A526, A527, A528, A529, A530, A531,
    A532, A533, A534, A535, A536, A537, A538, A539, A540, A541, A542, A543,
    A544, A545, A546, A547, A548, A549, A550, A551, A552, A553, A554, A555,
    A556, A557, A558, A559, A560, A561, A562, A563, A564, A565, A566, A567,
    A568, A569, A570, A571, A572, A573, A574, A575, A576, A577, A578, A579,
    A580, A581, A582, A583, A584, A585, A586, A587, A588, A589, A590, A591,
    A592, A593, A594, A595, A596, A597, A598, A599, A600, A601, A602, A603,
    A604, A605, A606, A607, A608, A609, A610, A611, A612, A613, A614, A615,
    A616, A617, A618, A619, A620, A621, A622, A623, A624, A625, A626, A627,
    A628, A629, A630, A631, A632, A633, A634, A635, A636, A637, A638, A639,
    A640, A641, A642, A643, A644, A645, A646, A647, A648, A649, A650, A651,
    A652, A653, A654, A655, A656, A657, A658, A659, A660, A661, A662, A663,
    A664, A665, A666, A667, A668, A669, A670, A671, A672, A673, A674, A675,
    A676, A677, A678, A679, A680, A681, A682, A683, A684, A685, A686, A687,
    A688, A689, A690, A691, A692, A693, A694, A695, A696, A697, A698, A699,
    A700, A701, A702, A703, A704, A705, A706, A707, A708, A709, A710, A711,
    A712, A713, A714, A715, A716, A717, A718, A719, A720, A721, A722, A723,
    A724, A725, A726, A727, A728, A729, A730, A731, A732, A733, A734, A735,
    A736, A737, A738, A739, A740, A741, A742, A743, A744, A745, A746, A747,
    A748, A749, A750, A751, A752, A753, A754, A755, A756, A757, A758, A759,
    A760, A761, A762, A763, A764, A765, A766, A767, A768, A769, A770, A771,
    A772, A773, A774, A775, A776, A777, A778, A779, A780, A781, A782, A783,
    A784, A785, A786, A787, A788, A789, A790, A791, A792, A793, A794, A795,
    A796, A797, A798, A799, A800, A801, A802, A803, A804, A805, A806, A807,
    A808, A809, A810, A811, A812, A813, A814, A815, A816, A817, A818, A819,
    A820, A821, A822, A823, A824, A825, A826, A827, A828, A829, A830, A831,
    A832, A833, A834, A835, A836, A837, A838, A839, A840, A841, A842, A843,
    A844, A845, A846, A847, A848, A849, A850, A851, A852, A853, A854, A855,
    A856, A857, A858, A859, A860, A861, A862, A863, A864, A865, A866, A867,
    A868, A869, A870, A871, A872, A873, A874, A875, A876, A877, A878, A879,
    A880, A881, A882, A883, A884, A885, A886, A887, A888, A889, A890, A891,
    A892, A893, A894, A895, A896, A897, A898, A899, A900, A901, A902, A903,
    A904, A905, A906, A907, A908, A909, A910, A911, A912, A913, A914, A915,
    A916, A917, A918, A919, A920, A921, A922, A923, A924, A925, A926, A927,
    A928, A929, A930, A931, A932, A933, A934, A935, A936, A937, A938, A939,
    A940, A941, A942, A943, A944, A945, A946, A947, A948, A949, A950, A951,
    A952, A953, A954, A955, A956, A957, A958, A959, A960, A961, A962, A963,
    A964, A965, A966, A967, A968, A969, A970, A971, A972, A973, A974, A975,
    A976, A977, A978, A979, A980, A981, A982, A983, A984, A985, A986, A987,
    A988, A989, A990, A991, A992, A993, A994, A995, A996, A997, A998, A999,
    A1000,
    maj  );
  input  A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14,
    A15, A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28,
    A29, A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42,
    A43, A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56,
    A57, A58, A59, A60, A61, A62, A63, A64, A65, A66, A67, A68, A69, A70,
    A71, A72, A73, A74, A75, A76, A77, A78, A79, A80, A81, A82, A83, A84,
    A85, A86, A87, A88, A89, A90, A91, A92, A93, A94, A95, A96, A97, A98,
    A99, A100, A101, A102, A103, A104, A105, A106, A107, A108, A109, A110,
    A111, A112, A113, A114, A115, A116, A117, A118, A119, A120, A121, A122,
    A123, A124, A125, A126, A127, A128, A129, A130, A131, A132, A133, A134,
    A135, A136, A137, A138, A139, A140, A141, A142, A143, A144, A145, A146,
    A147, A148, A149, A150, A151, A152, A153, A154, A155, A156, A157, A158,
    A159, A160, A161, A162, A163, A164, A165, A166, A167, A168, A169, A170,
    A171, A172, A173, A174, A175, A176, A177, A178, A179, A180, A181, A182,
    A183, A184, A185, A186, A187, A188, A189, A190, A191, A192, A193, A194,
    A195, A196, A197, A198, A199, A200, A201, A202, A203, A204, A205, A206,
    A207, A208, A209, A210, A211, A212, A213, A214, A215, A216, A217, A218,
    A219, A220, A221, A222, A223, A224, A225, A226, A227, A228, A229, A230,
    A231, A232, A233, A234, A235, A236, A237, A238, A239, A240, A241, A242,
    A243, A244, A245, A246, A247, A248, A249, A250, A251, A252, A253, A254,
    A255, A256, A257, A258, A259, A260, A261, A262, A263, A264, A265, A266,
    A267, A268, A269, A270, A271, A272, A273, A274, A275, A276, A277, A278,
    A279, A280, A281, A282, A283, A284, A285, A286, A287, A288, A289, A290,
    A291, A292, A293, A294, A295, A296, A297, A298, A299, A300, A301, A302,
    A303, A304, A305, A306, A307, A308, A309, A310, A311, A312, A313, A314,
    A315, A316, A317, A318, A319, A320, A321, A322, A323, A324, A325, A326,
    A327, A328, A329, A330, A331, A332, A333, A334, A335, A336, A337, A338,
    A339, A340, A341, A342, A343, A344, A345, A346, A347, A348, A349, A350,
    A351, A352, A353, A354, A355, A356, A357, A358, A359, A360, A361, A362,
    A363, A364, A365, A366, A367, A368, A369, A370, A371, A372, A373, A374,
    A375, A376, A377, A378, A379, A380, A381, A382, A383, A384, A385, A386,
    A387, A388, A389, A390, A391, A392, A393, A394, A395, A396, A397, A398,
    A399, A400, A401, A402, A403, A404, A405, A406, A407, A408, A409, A410,
    A411, A412, A413, A414, A415, A416, A417, A418, A419, A420, A421, A422,
    A423, A424, A425, A426, A427, A428, A429, A430, A431, A432, A433, A434,
    A435, A436, A437, A438, A439, A440, A441, A442, A443, A444, A445, A446,
    A447, A448, A449, A450, A451, A452, A453, A454, A455, A456, A457, A458,
    A459, A460, A461, A462, A463, A464, A465, A466, A467, A468, A469, A470,
    A471, A472, A473, A474, A475, A476, A477, A478, A479, A480, A481, A482,
    A483, A484, A485, A486, A487, A488, A489, A490, A491, A492, A493, A494,
    A495, A496, A497, A498, A499, A500, A501, A502, A503, A504, A505, A506,
    A507, A508, A509, A510, A511, A512, A513, A514, A515, A516, A517, A518,
    A519, A520, A521, A522, A523, A524, A525, A526, A527, A528, A529, A530,
    A531, A532, A533, A534, A535, A536, A537, A538, A539, A540, A541, A542,
    A543, A544, A545, A546, A547, A548, A549, A550, A551, A552, A553, A554,
    A555, A556, A557, A558, A559, A560, A561, A562, A563, A564, A565, A566,
    A567, A568, A569, A570, A571, A572, A573, A574, A575, A576, A577, A578,
    A579, A580, A581, A582, A583, A584, A585, A586, A587, A588, A589, A590,
    A591, A592, A593, A594, A595, A596, A597, A598, A599, A600, A601, A602,
    A603, A604, A605, A606, A607, A608, A609, A610, A611, A612, A613, A614,
    A615, A616, A617, A618, A619, A620, A621, A622, A623, A624, A625, A626,
    A627, A628, A629, A630, A631, A632, A633, A634, A635, A636, A637, A638,
    A639, A640, A641, A642, A643, A644, A645, A646, A647, A648, A649, A650,
    A651, A652, A653, A654, A655, A656, A657, A658, A659, A660, A661, A662,
    A663, A664, A665, A666, A667, A668, A669, A670, A671, A672, A673, A674,
    A675, A676, A677, A678, A679, A680, A681, A682, A683, A684, A685, A686,
    A687, A688, A689, A690, A691, A692, A693, A694, A695, A696, A697, A698,
    A699, A700, A701, A702, A703, A704, A705, A706, A707, A708, A709, A710,
    A711, A712, A713, A714, A715, A716, A717, A718, A719, A720, A721, A722,
    A723, A724, A725, A726, A727, A728, A729, A730, A731, A732, A733, A734,
    A735, A736, A737, A738, A739, A740, A741, A742, A743, A744, A745, A746,
    A747, A748, A749, A750, A751, A752, A753, A754, A755, A756, A757, A758,
    A759, A760, A761, A762, A763, A764, A765, A766, A767, A768, A769, A770,
    A771, A772, A773, A774, A775, A776, A777, A778, A779, A780, A781, A782,
    A783, A784, A785, A786, A787, A788, A789, A790, A791, A792, A793, A794,
    A795, A796, A797, A798, A799, A800, A801, A802, A803, A804, A805, A806,
    A807, A808, A809, A810, A811, A812, A813, A814, A815, A816, A817, A818,
    A819, A820, A821, A822, A823, A824, A825, A826, A827, A828, A829, A830,
    A831, A832, A833, A834, A835, A836, A837, A838, A839, A840, A841, A842,
    A843, A844, A845, A846, A847, A848, A849, A850, A851, A852, A853, A854,
    A855, A856, A857, A858, A859, A860, A861, A862, A863, A864, A865, A866,
    A867, A868, A869, A870, A871, A872, A873, A874, A875, A876, A877, A878,
    A879, A880, A881, A882, A883, A884, A885, A886, A887, A888, A889, A890,
    A891, A892, A893, A894, A895, A896, A897, A898, A899, A900, A901, A902,
    A903, A904, A905, A906, A907, A908, A909, A910, A911, A912, A913, A914,
    A915, A916, A917, A918, A919, A920, A921, A922, A923, A924, A925, A926,
    A927, A928, A929, A930, A931, A932, A933, A934, A935, A936, A937, A938,
    A939, A940, A941, A942, A943, A944, A945, A946, A947, A948, A949, A950,
    A951, A952, A953, A954, A955, A956, A957, A958, A959, A960, A961, A962,
    A963, A964, A965, A966, A967, A968, A969, A970, A971, A972, A973, A974,
    A975, A976, A977, A978, A979, A980, A981, A982, A983, A984, A985, A986,
    A987, A988, A989, A990, A991, A992, A993, A994, A995, A996, A997, A998,
    A999, A1000;
  output maj;
  wire new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1824,
    new_n1825, new_n1826, new_n1827, new_n1828, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1866,
    new_n1867, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436,
    new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604,
    new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610,
    new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628,
    new_n2629, new_n2630, new_n2631, new_n2632, new_n2633, new_n2634,
    new_n2635, new_n2636, new_n2637, new_n2638, new_n2639, new_n2640,
    new_n2641, new_n2642, new_n2643, new_n2644, new_n2645, new_n2646,
    new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658,
    new_n2659, new_n2660, new_n2661, new_n2662, new_n2663, new_n2664,
    new_n2665, new_n2666, new_n2667, new_n2668, new_n2669, new_n2670,
    new_n2671, new_n2672, new_n2673, new_n2674, new_n2675, new_n2676,
    new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682,
    new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694,
    new_n2695, new_n2696, new_n2697, new_n2698, new_n2699, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712,
    new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774, new_n2775, new_n2776, new_n2777, new_n2778,
    new_n2779, new_n2780, new_n2781, new_n2782, new_n2783, new_n2784,
    new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790,
    new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808,
    new_n2809, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570,
    new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576,
    new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582,
    new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588,
    new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594,
    new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600,
    new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606,
    new_n3607, new_n3608, new_n3609, new_n3610, new_n3611, new_n3612,
    new_n3613, new_n3614, new_n3615, new_n3616, new_n3617, new_n3618,
    new_n3619, new_n3620, new_n3621, new_n3622, new_n3623, new_n3624,
    new_n3625, new_n3626, new_n3627, new_n3628, new_n3629, new_n3630,
    new_n3631, new_n3632, new_n3633, new_n3634, new_n3635, new_n3636,
    new_n3637, new_n3638, new_n3639, new_n3640, new_n3641, new_n3642,
    new_n3643, new_n3644, new_n3645, new_n3646, new_n3647, new_n3648,
    new_n3649, new_n3650, new_n3651, new_n3652, new_n3653, new_n3654,
    new_n3655, new_n3656, new_n3657, new_n3658, new_n3659, new_n3660,
    new_n3661, new_n3662, new_n3663, new_n3664, new_n3665, new_n3666,
    new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672,
    new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684,
    new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690,
    new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696,
    new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702,
    new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708,
    new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726,
    new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732,
    new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738,
    new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744,
    new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750,
    new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756,
    new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774,
    new_n3775, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780,
    new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786,
    new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804,
    new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810,
    new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3816,
    new_n3817, new_n3818, new_n3819, new_n3820, new_n3821, new_n3822,
    new_n3823, new_n3824, new_n3825, new_n3826, new_n3827, new_n3828,
    new_n3829, new_n3830, new_n3831, new_n3832, new_n3833, new_n3834,
    new_n3835, new_n3836, new_n3837, new_n3838, new_n3839, new_n3840,
    new_n3841, new_n3842, new_n3843, new_n3844, new_n3845, new_n3846,
    new_n3847, new_n3848, new_n3849, new_n3850, new_n3851, new_n3852,
    new_n3853, new_n3854, new_n3855, new_n3856, new_n3857, new_n3858,
    new_n3859, new_n3860, new_n3861, new_n3862, new_n3863, new_n3864,
    new_n3865, new_n3866, new_n3867, new_n3868, new_n3869, new_n3870,
    new_n3871, new_n3872, new_n3873, new_n3874, new_n3875, new_n3876,
    new_n3877, new_n3878, new_n3879, new_n3880, new_n3881, new_n3882,
    new_n3883, new_n3884, new_n3885, new_n3886, new_n3887, new_n3888,
    new_n3889, new_n3890, new_n3891, new_n3892, new_n3893, new_n3894,
    new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900,
    new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906,
    new_n3907, new_n3908, new_n3909, new_n3910, new_n3911, new_n3912,
    new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918,
    new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924,
    new_n3925, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960,
    new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3979, new_n3980, new_n3981, new_n3982, new_n3983, new_n3984,
    new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964, new_n4965, new_n4966, new_n4967, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022,
    new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202,
    new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208,
    new_n5209, new_n5210, new_n5211, new_n5212, new_n5213, new_n5214,
    new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226,
    new_n5227, new_n5228, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255, new_n5256,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273, new_n5274,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300, new_n5301, new_n5302, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351, new_n5352,
    new_n5353, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630,
    new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726,
    new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732,
    new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738,
    new_n6739, new_n6740, new_n6741, new_n6742, new_n6743, new_n6744,
    new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750,
    new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756,
    new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762,
    new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768,
    new_n6769, new_n6770, new_n6771, new_n6772, new_n6773, new_n6774,
    new_n6775, new_n6776, new_n6777, new_n6778, new_n6779, new_n6780,
    new_n6781, new_n6782, new_n6783, new_n6784, new_n6785, new_n6786,
    new_n6787, new_n6788, new_n6789, new_n6790, new_n6791, new_n6792,
    new_n6793, new_n6794, new_n6795, new_n6796, new_n6797, new_n6798,
    new_n6799, new_n6800, new_n6801, new_n6802, new_n6803, new_n6804,
    new_n6805, new_n6806, new_n6807, new_n6808, new_n6809, new_n6810,
    new_n6811, new_n6812, new_n6813, new_n6814, new_n6815, new_n6816,
    new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822,
    new_n6823, new_n6824, new_n6825, new_n6826, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134,
    new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140,
    new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146,
    new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152,
    new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158,
    new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148,
    new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154,
    new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160,
    new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166,
    new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172,
    new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178,
    new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184,
    new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190,
    new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196,
    new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448,
    new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454,
    new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8460,
    new_n8461, new_n8462, new_n8463, new_n8464, new_n8465, new_n8466,
    new_n8467, new_n8468, new_n8469, new_n8470, new_n8471, new_n8472,
    new_n8473, new_n8474, new_n8475, new_n8476, new_n8477, new_n8478,
    new_n8479, new_n8480, new_n8481, new_n8482, new_n8483, new_n8484,
    new_n8485, new_n8486, new_n8487, new_n8488, new_n8489, new_n8490,
    new_n8491, new_n8492, new_n8493, new_n8494, new_n8495, new_n8496,
    new_n8497, new_n8498, new_n8499, new_n8500, new_n8501, new_n8502,
    new_n8503, new_n8504, new_n8505, new_n8506, new_n8507, new_n8508,
    new_n8509, new_n8510, new_n8511, new_n8512, new_n8513, new_n8514,
    new_n8515, new_n8516, new_n8517, new_n8518, new_n8519, new_n8520,
    new_n8521, new_n8522, new_n8523, new_n8524, new_n8525, new_n8526,
    new_n8527, new_n8528, new_n8529, new_n8530, new_n8531, new_n8532,
    new_n8533, new_n8534, new_n8535, new_n8536, new_n8537, new_n8538,
    new_n8539, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544,
    new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550,
    new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556,
    new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562,
    new_n8563, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568,
    new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574,
    new_n8575, new_n8576, new_n8577, new_n8578, new_n8579, new_n8580,
    new_n8581, new_n8582, new_n8583, new_n8584, new_n8585, new_n8586,
    new_n8587, new_n8588, new_n8589, new_n8590, new_n8591, new_n8592,
    new_n8593, new_n8594, new_n8595, new_n8596, new_n8597, new_n8598,
    new_n8599, new_n8600, new_n8601, new_n8602, new_n8603, new_n8604,
    new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610,
    new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616,
    new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622,
    new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628,
    new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634,
    new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552,
    new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558,
    new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564,
    new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570,
    new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576,
    new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582,
    new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912,
    new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9918,
    new_n9919, new_n9920, new_n9921, new_n9922, new_n9923, new_n9924,
    new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930,
    new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936,
    new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942,
    new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948,
    new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954,
    new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960,
    new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966,
    new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972,
    new_n9973, new_n9974, new_n9975, new_n9976, new_n9977, new_n9978,
    new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984,
    new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990,
    new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996,
    new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020,
    new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218,
    new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578,
    new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584,
    new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644,
    new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650,
    new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656,
    new_n10657, new_n10658, new_n10659, new_n10660, new_n10661, new_n10662,
    new_n10663, new_n10664, new_n10665, new_n10666, new_n10667, new_n10668,
    new_n10669, new_n10670, new_n10671, new_n10672, new_n10673, new_n10674,
    new_n10675, new_n10676, new_n10677, new_n10678, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685, new_n10686,
    new_n10687, new_n10688, new_n10689, new_n10690, new_n10691, new_n10692,
    new_n10693, new_n10694, new_n10695, new_n10696, new_n10697, new_n10698,
    new_n10699, new_n10700, new_n10701, new_n10702, new_n10703, new_n10704,
    new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710,
    new_n10711, new_n10712, new_n10713, new_n10714, new_n10715;
  assign new_n1003 = ~A961 & ~A962;
  assign new_n1004 = A961 & A962;
  assign new_n1005 = ~A963 & ~new_n1004;
  assign new_n1006 = ~new_n1003 & ~new_n1005;
  assign new_n1007 = A965 & A966;
  assign new_n1008 = new_n1006 & new_n1007;
  assign new_n1009 = A963 & new_n1004;
  assign new_n1010 = ~A964 & ~new_n1009;
  assign new_n1011 = new_n1006 & ~new_n1010;
  assign new_n1012 = A965 & new_n1011;
  assign new_n1013 = A963 & A964;
  assign new_n1014 = new_n1004 & new_n1013;
  assign new_n1015 = ~new_n1012 & ~new_n1014;
  assign new_n1016 = ~A966 & ~new_n1015;
  assign new_n1017 = ~A965 & ~A966;
  assign new_n1018 = ~new_n1003 & ~new_n1017;
  assign new_n1019 = new_n1005 & ~new_n1007;
  assign new_n1020 = ~new_n1018 & new_n1019;
  assign new_n1021 = ~new_n1008 & ~new_n1020;
  assign new_n1022 = ~A964 & ~new_n1021;
  assign new_n1023 = ~A965 & A966;
  assign new_n1024 = new_n1011 & new_n1023;
  assign new_n1025 = new_n1003 & ~new_n1013;
  assign new_n1026 = A964 & new_n1007;
  assign new_n1027 = ~new_n1009 & new_n1026;
  assign new_n1028 = ~new_n1025 & new_n1027;
  assign new_n1029 = ~new_n1024 & ~new_n1028;
  assign new_n1030 = ~new_n1022 & new_n1029;
  assign new_n1031 = ~new_n1016 & new_n1030;
  assign new_n1032 = ~new_n1010 & ~new_n1031;
  assign new_n1033 = ~new_n1008 & ~new_n1032;
  assign new_n1034 = A957 & A960;
  assign new_n1035 = A958 & A959;
  assign new_n1036 = A955 & A956;
  assign new_n1037 = ~new_n1035 & ~new_n1036;
  assign new_n1038 = new_n1034 & ~new_n1037;
  assign new_n1039 = ~A955 & ~A956;
  assign new_n1040 = ~A957 & A960;
  assign new_n1041 = new_n1035 & new_n1040;
  assign new_n1042 = ~A957 & ~new_n1036;
  assign new_n1043 = ~A958 & ~A959;
  assign new_n1044 = ~new_n1035 & ~new_n1043;
  assign new_n1045 = A960 & ~new_n1044;
  assign new_n1046 = ~A960 & ~new_n1035;
  assign new_n1047 = ~new_n1042 & ~new_n1046;
  assign new_n1048 = ~new_n1045 & new_n1047;
  assign new_n1049 = ~new_n1041 & ~new_n1048;
  assign new_n1050 = ~new_n1039 & ~new_n1049;
  assign new_n1051 = A959 & new_n1036;
  assign new_n1052 = new_n1038 & ~new_n1051;
  assign new_n1053 = ~new_n1034 & new_n1039;
  assign new_n1054 = new_n1043 & new_n1053;
  assign new_n1055 = A957 & ~A960;
  assign new_n1056 = new_n1036 & ~new_n1043;
  assign new_n1057 = new_n1055 & new_n1056;
  assign new_n1058 = ~new_n1054 & ~new_n1057;
  assign new_n1059 = ~new_n1052 & new_n1058;
  assign new_n1060 = ~new_n1050 & new_n1059;
  assign new_n1061 = ~new_n1039 & ~new_n1060;
  assign new_n1062 = ~new_n1038 & ~new_n1061;
  assign new_n1063 = new_n1033 & new_n1062;
  assign new_n1064 = ~new_n1036 & ~new_n1039;
  assign new_n1065 = ~new_n1040 & ~new_n1055;
  assign new_n1066 = new_n1064 & ~new_n1065;
  assign new_n1067 = ~new_n1064 & new_n1065;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n1044 & new_n1068;
  assign new_n1070 = ~new_n1044 & ~new_n1068;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = A964 & ~A966;
  assign new_n1073 = ~A964 & A966;
  assign new_n1074 = ~new_n1072 & ~new_n1073;
  assign new_n1075 = ~new_n1003 & ~new_n1004;
  assign new_n1076 = ~A963 & ~A965;
  assign new_n1077 = A963 & A965;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = new_n1075 & ~new_n1078;
  assign new_n1080 = ~new_n1075 & new_n1078;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign new_n1082 = new_n1074 & new_n1081;
  assign new_n1083 = ~new_n1074 & ~new_n1081;
  assign new_n1084 = ~new_n1082 & ~new_n1083;
  assign new_n1085 = new_n1071 & new_n1084;
  assign new_n1086 = new_n1042 & new_n1046;
  assign new_n1087 = ~new_n1069 & new_n1086;
  assign new_n1088 = new_n1060 & ~new_n1087;
  assign new_n1089 = ~new_n1085 & ~new_n1088;
  assign new_n1090 = new_n1017 & new_n1025;
  assign new_n1091 = new_n1031 & ~new_n1090;
  assign new_n1092 = new_n1085 & new_n1088;
  assign new_n1093 = ~new_n1089 & ~new_n1092;
  assign new_n1094 = ~new_n1091 & new_n1093;
  assign new_n1095 = ~new_n1089 & ~new_n1094;
  assign new_n1096 = ~new_n1033 & ~new_n1062;
  assign new_n1097 = ~new_n1063 & ~new_n1096;
  assign new_n1098 = ~new_n1095 & new_n1097;
  assign new_n1099 = ~new_n1063 & ~new_n1098;
  assign new_n1100 = A945 & A948;
  assign new_n1101 = A946 & A947;
  assign new_n1102 = A943 & A944;
  assign new_n1103 = ~new_n1101 & ~new_n1102;
  assign new_n1104 = new_n1100 & ~new_n1103;
  assign new_n1105 = ~A943 & ~A944;
  assign new_n1106 = ~A945 & A948;
  assign new_n1107 = new_n1101 & new_n1106;
  assign new_n1108 = ~A945 & ~new_n1102;
  assign new_n1109 = ~A946 & ~A947;
  assign new_n1110 = ~new_n1101 & ~new_n1109;
  assign new_n1111 = A948 & ~new_n1110;
  assign new_n1112 = ~A948 & ~new_n1101;
  assign new_n1113 = ~new_n1108 & ~new_n1112;
  assign new_n1114 = ~new_n1111 & new_n1113;
  assign new_n1115 = ~new_n1107 & ~new_n1114;
  assign new_n1116 = ~new_n1105 & ~new_n1115;
  assign new_n1117 = A947 & new_n1102;
  assign new_n1118 = new_n1104 & ~new_n1117;
  assign new_n1119 = ~new_n1100 & new_n1105;
  assign new_n1120 = new_n1109 & new_n1119;
  assign new_n1121 = A945 & ~A948;
  assign new_n1122 = new_n1102 & ~new_n1109;
  assign new_n1123 = new_n1121 & new_n1122;
  assign new_n1124 = ~new_n1120 & ~new_n1123;
  assign new_n1125 = ~new_n1118 & new_n1124;
  assign new_n1126 = ~new_n1116 & new_n1125;
  assign new_n1127 = ~new_n1105 & ~new_n1126;
  assign new_n1128 = ~new_n1104 & ~new_n1127;
  assign new_n1129 = A951 & A954;
  assign new_n1130 = A952 & A953;
  assign new_n1131 = A949 & A950;
  assign new_n1132 = ~new_n1130 & ~new_n1131;
  assign new_n1133 = new_n1129 & ~new_n1132;
  assign new_n1134 = ~A949 & ~A950;
  assign new_n1135 = ~A951 & A954;
  assign new_n1136 = new_n1130 & new_n1135;
  assign new_n1137 = ~A951 & ~new_n1131;
  assign new_n1138 = ~A952 & ~A953;
  assign new_n1139 = ~new_n1130 & ~new_n1138;
  assign new_n1140 = A954 & ~new_n1139;
  assign new_n1141 = ~A954 & ~new_n1130;
  assign new_n1142 = ~new_n1137 & ~new_n1141;
  assign new_n1143 = ~new_n1140 & new_n1142;
  assign new_n1144 = ~new_n1136 & ~new_n1143;
  assign new_n1145 = ~new_n1134 & ~new_n1144;
  assign new_n1146 = A953 & new_n1131;
  assign new_n1147 = new_n1133 & ~new_n1146;
  assign new_n1148 = ~new_n1129 & new_n1134;
  assign new_n1149 = new_n1138 & new_n1148;
  assign new_n1150 = A951 & ~A954;
  assign new_n1151 = new_n1131 & ~new_n1138;
  assign new_n1152 = new_n1150 & new_n1151;
  assign new_n1153 = ~new_n1149 & ~new_n1152;
  assign new_n1154 = ~new_n1147 & new_n1153;
  assign new_n1155 = ~new_n1145 & new_n1154;
  assign new_n1156 = ~new_n1134 & ~new_n1155;
  assign new_n1157 = ~new_n1133 & ~new_n1156;
  assign new_n1158 = new_n1128 & new_n1157;
  assign new_n1159 = ~new_n1102 & ~new_n1105;
  assign new_n1160 = ~new_n1106 & ~new_n1121;
  assign new_n1161 = new_n1159 & ~new_n1160;
  assign new_n1162 = ~new_n1159 & new_n1160;
  assign new_n1163 = ~new_n1161 & ~new_n1162;
  assign new_n1164 = new_n1110 & new_n1163;
  assign new_n1165 = ~new_n1110 & ~new_n1163;
  assign new_n1166 = ~new_n1164 & ~new_n1165;
  assign new_n1167 = ~new_n1131 & ~new_n1134;
  assign new_n1168 = ~new_n1135 & ~new_n1150;
  assign new_n1169 = new_n1167 & ~new_n1168;
  assign new_n1170 = ~new_n1167 & new_n1168;
  assign new_n1171 = ~new_n1169 & ~new_n1170;
  assign new_n1172 = new_n1139 & new_n1171;
  assign new_n1173 = ~new_n1139 & ~new_n1171;
  assign new_n1174 = ~new_n1172 & ~new_n1173;
  assign new_n1175 = new_n1166 & new_n1174;
  assign new_n1176 = new_n1137 & new_n1141;
  assign new_n1177 = ~new_n1172 & new_n1176;
  assign new_n1178 = new_n1155 & ~new_n1177;
  assign new_n1179 = ~new_n1175 & ~new_n1178;
  assign new_n1180 = new_n1175 & new_n1178;
  assign new_n1181 = ~new_n1179 & ~new_n1180;
  assign new_n1182 = new_n1108 & new_n1112;
  assign new_n1183 = ~new_n1164 & new_n1182;
  assign new_n1184 = new_n1126 & ~new_n1183;
  assign new_n1185 = new_n1181 & ~new_n1184;
  assign new_n1186 = ~new_n1179 & ~new_n1185;
  assign new_n1187 = ~new_n1128 & ~new_n1157;
  assign new_n1188 = ~new_n1158 & ~new_n1187;
  assign new_n1189 = ~new_n1186 & new_n1188;
  assign new_n1190 = ~new_n1158 & ~new_n1189;
  assign new_n1191 = new_n1099 & new_n1190;
  assign new_n1192 = ~new_n1099 & ~new_n1190;
  assign new_n1193 = ~new_n1191 & ~new_n1192;
  assign new_n1194 = new_n1186 & ~new_n1188;
  assign new_n1195 = ~new_n1189 & ~new_n1194;
  assign new_n1196 = new_n1091 & ~new_n1093;
  assign new_n1197 = ~new_n1094 & ~new_n1196;
  assign new_n1198 = ~new_n1181 & new_n1184;
  assign new_n1199 = ~new_n1185 & ~new_n1198;
  assign new_n1200 = new_n1197 & new_n1199;
  assign new_n1201 = ~new_n1166 & ~new_n1174;
  assign new_n1202 = ~new_n1175 & ~new_n1201;
  assign new_n1203 = ~new_n1071 & ~new_n1084;
  assign new_n1204 = ~new_n1085 & ~new_n1203;
  assign new_n1205 = new_n1202 & new_n1204;
  assign new_n1206 = ~new_n1197 & ~new_n1199;
  assign new_n1207 = ~new_n1200 & ~new_n1206;
  assign new_n1208 = ~new_n1205 & new_n1207;
  assign new_n1209 = ~new_n1200 & ~new_n1208;
  assign new_n1210 = ~new_n1195 & new_n1209;
  assign new_n1211 = new_n1095 & ~new_n1097;
  assign new_n1212 = ~new_n1098 & ~new_n1211;
  assign new_n1213 = new_n1195 & ~new_n1209;
  assign new_n1214 = ~new_n1210 & ~new_n1213;
  assign new_n1215 = ~new_n1212 & new_n1214;
  assign new_n1216 = ~new_n1210 & ~new_n1215;
  assign new_n1217 = new_n1193 & ~new_n1216;
  assign new_n1218 = ~new_n1191 & ~new_n1217;
  assign new_n1219 = A981 & A984;
  assign new_n1220 = A982 & A983;
  assign new_n1221 = A979 & A980;
  assign new_n1222 = ~new_n1220 & ~new_n1221;
  assign new_n1223 = new_n1219 & ~new_n1222;
  assign new_n1224 = ~A979 & ~A980;
  assign new_n1225 = ~A981 & A984;
  assign new_n1226 = new_n1220 & new_n1225;
  assign new_n1227 = ~A981 & ~new_n1221;
  assign new_n1228 = ~A982 & ~A983;
  assign new_n1229 = ~new_n1220 & ~new_n1228;
  assign new_n1230 = A984 & ~new_n1229;
  assign new_n1231 = ~A984 & ~new_n1220;
  assign new_n1232 = ~new_n1227 & ~new_n1231;
  assign new_n1233 = ~new_n1230 & new_n1232;
  assign new_n1234 = ~new_n1226 & ~new_n1233;
  assign new_n1235 = ~new_n1224 & ~new_n1234;
  assign new_n1236 = A983 & new_n1221;
  assign new_n1237 = new_n1223 & ~new_n1236;
  assign new_n1238 = ~new_n1219 & new_n1224;
  assign new_n1239 = new_n1228 & new_n1238;
  assign new_n1240 = A981 & ~A984;
  assign new_n1241 = new_n1221 & ~new_n1228;
  assign new_n1242 = new_n1240 & new_n1241;
  assign new_n1243 = ~new_n1239 & ~new_n1242;
  assign new_n1244 = ~new_n1237 & new_n1243;
  assign new_n1245 = ~new_n1235 & new_n1244;
  assign new_n1246 = ~new_n1224 & ~new_n1245;
  assign new_n1247 = ~new_n1223 & ~new_n1246;
  assign new_n1248 = ~A989 & ~A990;
  assign new_n1249 = A989 & A990;
  assign new_n1250 = ~new_n1248 & ~new_n1249;
  assign new_n1251 = ~A988 & new_n1250;
  assign new_n1252 = ~new_n1248 & ~new_n1251;
  assign new_n1253 = ~A986 & ~A987;
  assign new_n1254 = A986 & A987;
  assign new_n1255 = ~new_n1253 & ~new_n1254;
  assign new_n1256 = ~A985 & new_n1255;
  assign new_n1257 = ~new_n1253 & ~new_n1256;
  assign new_n1258 = ~new_n1252 & ~new_n1257;
  assign new_n1259 = A985 & ~new_n1255;
  assign new_n1260 = ~new_n1256 & ~new_n1259;
  assign new_n1261 = A988 & ~new_n1250;
  assign new_n1262 = ~new_n1251 & ~new_n1261;
  assign new_n1263 = ~new_n1260 & ~new_n1262;
  assign new_n1264 = new_n1252 & new_n1257;
  assign new_n1265 = ~new_n1258 & ~new_n1264;
  assign new_n1266 = ~new_n1263 & new_n1265;
  assign new_n1267 = ~new_n1258 & ~new_n1266;
  assign new_n1268 = ~new_n1247 & new_n1267;
  assign new_n1269 = new_n1263 & ~new_n1265;
  assign new_n1270 = ~new_n1266 & ~new_n1269;
  assign new_n1271 = ~new_n1221 & ~new_n1224;
  assign new_n1272 = ~new_n1225 & ~new_n1240;
  assign new_n1273 = new_n1271 & ~new_n1272;
  assign new_n1274 = ~new_n1271 & new_n1272;
  assign new_n1275 = ~new_n1273 & ~new_n1274;
  assign new_n1276 = new_n1229 & new_n1275;
  assign new_n1277 = new_n1227 & new_n1231;
  assign new_n1278 = ~new_n1276 & new_n1277;
  assign new_n1279 = new_n1245 & ~new_n1278;
  assign new_n1280 = ~new_n1270 & new_n1279;
  assign new_n1281 = ~new_n1229 & ~new_n1275;
  assign new_n1282 = ~new_n1276 & ~new_n1281;
  assign new_n1283 = new_n1260 & new_n1262;
  assign new_n1284 = ~new_n1263 & ~new_n1283;
  assign new_n1285 = new_n1282 & new_n1284;
  assign new_n1286 = ~new_n1265 & ~new_n1279;
  assign new_n1287 = new_n1285 & ~new_n1286;
  assign new_n1288 = ~new_n1280 & ~new_n1287;
  assign new_n1289 = new_n1247 & ~new_n1267;
  assign new_n1290 = ~new_n1268 & ~new_n1289;
  assign new_n1291 = ~new_n1288 & new_n1290;
  assign new_n1292 = ~new_n1268 & ~new_n1291;
  assign new_n1293 = ~A968 & ~A969;
  assign new_n1294 = A968 & A969;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = ~A967 & new_n1295;
  assign new_n1297 = ~new_n1293 & ~new_n1296;
  assign new_n1298 = ~A971 & ~A972;
  assign new_n1299 = A971 & A972;
  assign new_n1300 = ~new_n1298 & ~new_n1299;
  assign new_n1301 = ~A970 & new_n1300;
  assign new_n1302 = ~new_n1298 & ~new_n1301;
  assign new_n1303 = ~new_n1297 & ~new_n1302;
  assign new_n1304 = new_n1297 & new_n1302;
  assign new_n1305 = ~new_n1303 & ~new_n1304;
  assign new_n1306 = A967 & ~new_n1295;
  assign new_n1307 = ~new_n1296 & ~new_n1306;
  assign new_n1308 = A970 & ~new_n1300;
  assign new_n1309 = ~new_n1301 & ~new_n1308;
  assign new_n1310 = ~new_n1307 & ~new_n1309;
  assign new_n1311 = new_n1305 & ~new_n1310;
  assign new_n1312 = ~new_n1303 & ~new_n1311;
  assign new_n1313 = ~A977 & ~A978;
  assign new_n1314 = A973 & A974;
  assign new_n1315 = A975 & A976;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = ~A975 & ~A976;
  assign new_n1318 = ~A973 & ~A974;
  assign new_n1319 = ~new_n1317 & ~new_n1318;
  assign new_n1320 = ~new_n1313 & ~new_n1316;
  assign new_n1321 = new_n1319 & new_n1320;
  assign new_n1322 = new_n1316 & ~new_n1319;
  assign new_n1323 = new_n1314 & new_n1315;
  assign new_n1324 = ~new_n1322 & ~new_n1323;
  assign new_n1325 = ~new_n1313 & ~new_n1324;
  assign new_n1326 = A977 & A978;
  assign new_n1327 = ~new_n1323 & ~new_n1326;
  assign new_n1328 = ~new_n1325 & ~new_n1327;
  assign new_n1329 = ~new_n1321 & ~new_n1328;
  assign new_n1330 = ~new_n1312 & new_n1329;
  assign new_n1331 = new_n1307 & new_n1309;
  assign new_n1332 = ~new_n1310 & ~new_n1331;
  assign new_n1333 = ~new_n1315 & ~new_n1317;
  assign new_n1334 = ~new_n1313 & ~new_n1326;
  assign new_n1335 = new_n1333 & ~new_n1334;
  assign new_n1336 = ~new_n1333 & new_n1334;
  assign new_n1337 = ~new_n1335 & ~new_n1336;
  assign new_n1338 = ~new_n1314 & ~new_n1318;
  assign new_n1339 = ~new_n1337 & new_n1338;
  assign new_n1340 = new_n1337 & ~new_n1338;
  assign new_n1341 = ~new_n1339 & ~new_n1340;
  assign new_n1342 = new_n1332 & ~new_n1341;
  assign new_n1343 = ~new_n1331 & ~new_n1342;
  assign new_n1344 = ~new_n1305 & new_n1343;
  assign new_n1345 = new_n1305 & ~new_n1343;
  assign new_n1346 = ~new_n1344 & ~new_n1345;
  assign new_n1347 = new_n1317 & new_n1318;
  assign new_n1348 = ~new_n1321 & ~new_n1347;
  assign new_n1349 = ~new_n1326 & ~new_n1348;
  assign new_n1350 = new_n1313 & ~new_n1324;
  assign new_n1351 = ~new_n1328 & ~new_n1350;
  assign new_n1352 = ~new_n1349 & new_n1351;
  assign new_n1353 = ~new_n1346 & ~new_n1352;
  assign new_n1354 = ~new_n1311 & ~new_n1344;
  assign new_n1355 = ~new_n1353 & ~new_n1354;
  assign new_n1356 = new_n1312 & ~new_n1329;
  assign new_n1357 = ~new_n1330 & ~new_n1356;
  assign new_n1358 = ~new_n1355 & new_n1357;
  assign new_n1359 = ~new_n1330 & ~new_n1358;
  assign new_n1360 = new_n1292 & ~new_n1359;
  assign new_n1361 = new_n1288 & ~new_n1290;
  assign new_n1362 = ~new_n1291 & ~new_n1361;
  assign new_n1363 = ~new_n1282 & ~new_n1284;
  assign new_n1364 = ~new_n1285 & ~new_n1363;
  assign new_n1365 = ~new_n1332 & new_n1341;
  assign new_n1366 = ~new_n1342 & ~new_n1365;
  assign new_n1367 = new_n1364 & ~new_n1366;
  assign new_n1368 = ~new_n1263 & ~new_n1285;
  assign new_n1369 = new_n1265 & new_n1279;
  assign new_n1370 = ~new_n1286 & ~new_n1369;
  assign new_n1371 = new_n1368 & ~new_n1370;
  assign new_n1372 = ~new_n1368 & new_n1370;
  assign new_n1373 = ~new_n1371 & ~new_n1372;
  assign new_n1374 = new_n1367 & new_n1373;
  assign new_n1375 = new_n1346 & new_n1352;
  assign new_n1376 = ~new_n1353 & ~new_n1375;
  assign new_n1377 = ~new_n1367 & ~new_n1373;
  assign new_n1378 = ~new_n1374 & ~new_n1377;
  assign new_n1379 = ~new_n1376 & new_n1378;
  assign new_n1380 = ~new_n1374 & ~new_n1379;
  assign new_n1381 = new_n1362 & ~new_n1380;
  assign new_n1382 = new_n1355 & ~new_n1357;
  assign new_n1383 = ~new_n1358 & ~new_n1382;
  assign new_n1384 = ~new_n1362 & new_n1380;
  assign new_n1385 = ~new_n1381 & ~new_n1384;
  assign new_n1386 = ~new_n1383 & new_n1385;
  assign new_n1387 = ~new_n1381 & ~new_n1386;
  assign new_n1388 = ~new_n1292 & new_n1359;
  assign new_n1389 = ~new_n1360 & ~new_n1388;
  assign new_n1390 = new_n1387 & new_n1389;
  assign new_n1391 = ~new_n1360 & ~new_n1390;
  assign new_n1392 = new_n1218 & ~new_n1391;
  assign new_n1393 = ~new_n1218 & new_n1391;
  assign new_n1394 = ~new_n1392 & ~new_n1393;
  assign new_n1395 = ~new_n1193 & new_n1216;
  assign new_n1396 = ~new_n1217 & ~new_n1395;
  assign new_n1397 = ~new_n1387 & ~new_n1389;
  assign new_n1398 = ~new_n1390 & ~new_n1397;
  assign new_n1399 = new_n1396 & ~new_n1398;
  assign new_n1400 = ~new_n1396 & new_n1398;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = new_n1212 & ~new_n1214;
  assign new_n1403 = ~new_n1215 & ~new_n1402;
  assign new_n1404 = new_n1376 & ~new_n1378;
  assign new_n1405 = ~new_n1379 & ~new_n1404;
  assign new_n1406 = new_n1205 & ~new_n1207;
  assign new_n1407 = ~new_n1208 & ~new_n1406;
  assign new_n1408 = ~new_n1405 & new_n1407;
  assign new_n1409 = ~new_n1202 & ~new_n1204;
  assign new_n1410 = ~new_n1205 & ~new_n1409;
  assign new_n1411 = ~new_n1364 & new_n1366;
  assign new_n1412 = ~new_n1367 & ~new_n1411;
  assign new_n1413 = new_n1410 & new_n1412;
  assign new_n1414 = new_n1405 & ~new_n1407;
  assign new_n1415 = ~new_n1408 & ~new_n1414;
  assign new_n1416 = ~new_n1413 & new_n1415;
  assign new_n1417 = ~new_n1408 & ~new_n1416;
  assign new_n1418 = ~new_n1403 & ~new_n1417;
  assign new_n1419 = new_n1383 & ~new_n1385;
  assign new_n1420 = ~new_n1386 & ~new_n1419;
  assign new_n1421 = new_n1403 & new_n1417;
  assign new_n1422 = ~new_n1418 & ~new_n1421;
  assign new_n1423 = ~new_n1420 & new_n1422;
  assign new_n1424 = ~new_n1418 & ~new_n1423;
  assign new_n1425 = new_n1401 & new_n1424;
  assign new_n1426 = ~new_n1399 & ~new_n1425;
  assign new_n1427 = new_n1394 & new_n1426;
  assign new_n1428 = ~new_n1394 & ~new_n1426;
  assign new_n1429 = ~new_n1427 & ~new_n1428;
  assign new_n1430 = A5 & A6;
  assign new_n1431 = ~A5 & ~A6;
  assign new_n1432 = ~new_n1430 & ~new_n1431;
  assign new_n1433 = ~A3 & ~A4;
  assign new_n1434 = A3 & A4;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = A1 & A2;
  assign new_n1437 = ~A1 & ~A2;
  assign new_n1438 = ~new_n1436 & ~new_n1437;
  assign new_n1439 = A0 & ~new_n1438;
  assign new_n1440 = ~A0 & new_n1438;
  assign new_n1441 = ~new_n1439 & ~new_n1440;
  assign new_n1442 = new_n1435 & ~new_n1441;
  assign new_n1443 = ~new_n1435 & new_n1441;
  assign new_n1444 = ~new_n1442 & ~new_n1443;
  assign new_n1445 = new_n1432 & new_n1444;
  assign new_n1446 = ~new_n1432 & ~new_n1444;
  assign new_n1447 = ~new_n1445 & ~new_n1446;
  assign new_n1448 = A999 & new_n1447;
  assign new_n1449 = ~A999 & ~new_n1447;
  assign new_n1450 = ~new_n1448 & ~new_n1449;
  assign new_n1451 = A997 & A998;
  assign new_n1452 = ~A997 & ~A998;
  assign new_n1453 = ~new_n1451 & ~new_n1452;
  assign new_n1454 = ~new_n1450 & new_n1453;
  assign new_n1455 = new_n1450 & ~new_n1453;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = A995 & A996;
  assign new_n1458 = ~A995 & ~A996;
  assign new_n1459 = ~A992 & ~A993;
  assign new_n1460 = A992 & A993;
  assign new_n1461 = ~new_n1459 & ~new_n1460;
  assign new_n1462 = ~A991 & new_n1461;
  assign new_n1463 = ~new_n1459 & ~new_n1462;
  assign new_n1464 = ~new_n1458 & new_n1463;
  assign new_n1465 = ~new_n1457 & new_n1464;
  assign new_n1466 = ~A994 & new_n1465;
  assign new_n1467 = A991 & ~new_n1461;
  assign new_n1468 = ~new_n1462 & ~new_n1467;
  assign new_n1469 = ~A994 & new_n1468;
  assign new_n1470 = ~new_n1457 & ~new_n1463;
  assign new_n1471 = ~new_n1469 & ~new_n1470;
  assign new_n1472 = A994 & ~new_n1468;
  assign new_n1473 = ~new_n1458 & new_n1472;
  assign new_n1474 = ~new_n1471 & ~new_n1473;
  assign new_n1475 = ~new_n1464 & ~new_n1474;
  assign new_n1476 = ~new_n1466 & ~new_n1475;
  assign new_n1477 = ~new_n1456 & ~new_n1476;
  assign new_n1478 = ~new_n1469 & ~new_n1472;
  assign new_n1479 = new_n1465 & new_n1478;
  assign new_n1480 = ~new_n1456 & new_n1478;
  assign new_n1481 = new_n1458 & ~new_n1463;
  assign new_n1482 = ~new_n1472 & new_n1481;
  assign new_n1483 = ~new_n1480 & new_n1482;
  assign new_n1484 = new_n1464 & ~new_n1469;
  assign new_n1485 = new_n1457 & new_n1463;
  assign new_n1486 = ~new_n1472 & ~new_n1485;
  assign new_n1487 = ~new_n1470 & ~new_n1486;
  assign new_n1488 = ~new_n1484 & new_n1487;
  assign new_n1489 = new_n1469 & new_n1470;
  assign new_n1490 = ~new_n1467 & new_n1485;
  assign new_n1491 = A994 & new_n1457;
  assign new_n1492 = ~new_n1468 & ~new_n1491;
  assign new_n1493 = new_n1464 & new_n1492;
  assign new_n1494 = ~new_n1489 & ~new_n1490;
  assign new_n1495 = ~new_n1493 & new_n1494;
  assign new_n1496 = new_n1456 & ~new_n1495;
  assign new_n1497 = ~new_n1479 & ~new_n1488;
  assign new_n1498 = ~new_n1496 & new_n1497;
  assign new_n1499 = ~new_n1483 & new_n1498;
  assign new_n1500 = ~new_n1477 & new_n1499;
  assign new_n1501 = ~new_n1437 & ~new_n1440;
  assign new_n1502 = ~new_n1431 & ~new_n1433;
  assign new_n1503 = ~new_n1430 & new_n1441;
  assign new_n1504 = new_n1431 & new_n1433;
  assign new_n1505 = ~new_n1503 & ~new_n1504;
  assign new_n1506 = ~new_n1434 & ~new_n1502;
  assign new_n1507 = ~new_n1505 & new_n1506;
  assign new_n1508 = new_n1430 & ~new_n1441;
  assign new_n1509 = ~new_n1434 & ~new_n1508;
  assign new_n1510 = new_n1502 & ~new_n1503;
  assign new_n1511 = ~new_n1509 & new_n1510;
  assign new_n1512 = ~new_n1507 & ~new_n1511;
  assign new_n1513 = ~new_n1501 & new_n1512;
  assign new_n1514 = new_n1501 & ~new_n1512;
  assign new_n1515 = ~new_n1513 & ~new_n1514;
  assign new_n1516 = new_n1448 & new_n1451;
  assign new_n1517 = ~new_n1452 & ~new_n1454;
  assign new_n1518 = ~new_n1448 & ~new_n1517;
  assign new_n1519 = ~new_n1516 & ~new_n1518;
  assign new_n1520 = new_n1515 & ~new_n1519;
  assign new_n1521 = ~new_n1515 & new_n1519;
  assign new_n1522 = ~new_n1520 & ~new_n1521;
  assign new_n1523 = new_n1500 & ~new_n1522;
  assign new_n1524 = ~new_n1500 & new_n1522;
  assign new_n1525 = ~new_n1523 & ~new_n1524;
  assign new_n1526 = ~A25 & ~A26;
  assign new_n1527 = A25 & A26;
  assign new_n1528 = ~A27 & ~new_n1527;
  assign new_n1529 = ~new_n1526 & ~new_n1528;
  assign new_n1530 = A27 & new_n1527;
  assign new_n1531 = ~A28 & ~new_n1530;
  assign new_n1532 = new_n1529 & ~new_n1531;
  assign new_n1533 = A29 & new_n1532;
  assign new_n1534 = A27 & A28;
  assign new_n1535 = new_n1527 & new_n1534;
  assign new_n1536 = ~new_n1533 & ~new_n1535;
  assign new_n1537 = ~A30 & ~new_n1536;
  assign new_n1538 = A29 & A30;
  assign new_n1539 = new_n1529 & new_n1538;
  assign new_n1540 = ~A29 & ~A30;
  assign new_n1541 = ~new_n1526 & ~new_n1540;
  assign new_n1542 = new_n1528 & ~new_n1538;
  assign new_n1543 = ~new_n1541 & new_n1542;
  assign new_n1544 = ~new_n1539 & ~new_n1543;
  assign new_n1545 = ~A28 & ~new_n1544;
  assign new_n1546 = ~A29 & A30;
  assign new_n1547 = new_n1532 & new_n1546;
  assign new_n1548 = new_n1526 & ~new_n1534;
  assign new_n1549 = A28 & new_n1538;
  assign new_n1550 = ~new_n1530 & new_n1549;
  assign new_n1551 = ~new_n1548 & new_n1550;
  assign new_n1552 = ~new_n1547 & ~new_n1551;
  assign new_n1553 = ~new_n1545 & new_n1552;
  assign new_n1554 = ~new_n1537 & new_n1553;
  assign new_n1555 = new_n1540 & new_n1548;
  assign new_n1556 = new_n1554 & ~new_n1555;
  assign new_n1557 = A22 & A23;
  assign new_n1558 = ~A22 & ~A23;
  assign new_n1559 = ~new_n1557 & ~new_n1558;
  assign new_n1560 = A19 & A20;
  assign new_n1561 = ~A19 & ~A20;
  assign new_n1562 = ~new_n1560 & ~new_n1561;
  assign new_n1563 = ~A21 & A24;
  assign new_n1564 = A21 & ~A24;
  assign new_n1565 = ~new_n1563 & ~new_n1564;
  assign new_n1566 = new_n1562 & ~new_n1565;
  assign new_n1567 = ~new_n1562 & new_n1565;
  assign new_n1568 = ~new_n1566 & ~new_n1567;
  assign new_n1569 = new_n1559 & new_n1568;
  assign new_n1570 = ~new_n1559 & ~new_n1568;
  assign new_n1571 = ~new_n1569 & ~new_n1570;
  assign new_n1572 = A27 & ~A30;
  assign new_n1573 = ~A27 & A30;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = ~new_n1526 & ~new_n1527;
  assign new_n1576 = ~A28 & ~A29;
  assign new_n1577 = A28 & A29;
  assign new_n1578 = ~new_n1576 & ~new_n1577;
  assign new_n1579 = new_n1575 & ~new_n1578;
  assign new_n1580 = ~new_n1575 & new_n1578;
  assign new_n1581 = ~new_n1579 & ~new_n1580;
  assign new_n1582 = new_n1574 & new_n1581;
  assign new_n1583 = ~new_n1574 & ~new_n1581;
  assign new_n1584 = ~new_n1582 & ~new_n1583;
  assign new_n1585 = new_n1571 & new_n1584;
  assign new_n1586 = new_n1557 & new_n1563;
  assign new_n1587 = A24 & ~new_n1559;
  assign new_n1588 = ~A21 & ~new_n1560;
  assign new_n1589 = ~A24 & ~new_n1557;
  assign new_n1590 = ~new_n1588 & ~new_n1589;
  assign new_n1591 = ~new_n1587 & new_n1590;
  assign new_n1592 = ~new_n1586 & ~new_n1591;
  assign new_n1593 = ~new_n1561 & ~new_n1592;
  assign new_n1594 = A21 & A24;
  assign new_n1595 = ~new_n1557 & ~new_n1560;
  assign new_n1596 = new_n1594 & ~new_n1595;
  assign new_n1597 = A23 & new_n1560;
  assign new_n1598 = new_n1596 & ~new_n1597;
  assign new_n1599 = new_n1558 & new_n1561;
  assign new_n1600 = ~new_n1594 & new_n1599;
  assign new_n1601 = ~new_n1558 & new_n1560;
  assign new_n1602 = new_n1564 & new_n1601;
  assign new_n1603 = ~new_n1600 & ~new_n1602;
  assign new_n1604 = ~new_n1598 & new_n1603;
  assign new_n1605 = ~new_n1593 & new_n1604;
  assign new_n1606 = new_n1588 & new_n1589;
  assign new_n1607 = ~new_n1569 & new_n1606;
  assign new_n1608 = new_n1605 & ~new_n1607;
  assign new_n1609 = ~new_n1585 & ~new_n1608;
  assign new_n1610 = new_n1585 & new_n1608;
  assign new_n1611 = ~new_n1609 & ~new_n1610;
  assign new_n1612 = ~new_n1556 & new_n1611;
  assign new_n1613 = new_n1556 & ~new_n1611;
  assign new_n1614 = ~new_n1612 & ~new_n1613;
  assign new_n1615 = A10 & A11;
  assign new_n1616 = ~A10 & ~A11;
  assign new_n1617 = ~new_n1615 & ~new_n1616;
  assign new_n1618 = A7 & A8;
  assign new_n1619 = ~A7 & ~A8;
  assign new_n1620 = ~new_n1618 & ~new_n1619;
  assign new_n1621 = ~A9 & A12;
  assign new_n1622 = A9 & ~A12;
  assign new_n1623 = ~new_n1621 & ~new_n1622;
  assign new_n1624 = new_n1620 & ~new_n1623;
  assign new_n1625 = ~new_n1620 & new_n1623;
  assign new_n1626 = ~new_n1624 & ~new_n1625;
  assign new_n1627 = new_n1617 & new_n1626;
  assign new_n1628 = ~new_n1617 & ~new_n1626;
  assign new_n1629 = ~new_n1627 & ~new_n1628;
  assign new_n1630 = A14 & A15;
  assign new_n1631 = ~A14 & ~A15;
  assign new_n1632 = ~new_n1630 & ~new_n1631;
  assign new_n1633 = A13 & ~new_n1632;
  assign new_n1634 = ~A13 & new_n1632;
  assign new_n1635 = ~new_n1633 & ~new_n1634;
  assign new_n1636 = A18 & ~new_n1635;
  assign new_n1637 = ~A18 & new_n1635;
  assign new_n1638 = ~new_n1636 & ~new_n1637;
  assign new_n1639 = A16 & A17;
  assign new_n1640 = ~A16 & ~A17;
  assign new_n1641 = ~new_n1639 & ~new_n1640;
  assign new_n1642 = new_n1638 & ~new_n1641;
  assign new_n1643 = ~new_n1638 & new_n1641;
  assign new_n1644 = ~new_n1642 & ~new_n1643;
  assign new_n1645 = new_n1629 & ~new_n1644;
  assign new_n1646 = new_n1615 & new_n1621;
  assign new_n1647 = A12 & ~new_n1617;
  assign new_n1648 = ~A9 & ~new_n1618;
  assign new_n1649 = ~A12 & ~new_n1615;
  assign new_n1650 = ~new_n1648 & ~new_n1649;
  assign new_n1651 = ~new_n1647 & new_n1650;
  assign new_n1652 = ~new_n1646 & ~new_n1651;
  assign new_n1653 = ~new_n1619 & ~new_n1652;
  assign new_n1654 = A9 & A12;
  assign new_n1655 = ~new_n1615 & ~new_n1618;
  assign new_n1656 = new_n1654 & ~new_n1655;
  assign new_n1657 = A11 & new_n1618;
  assign new_n1658 = new_n1656 & ~new_n1657;
  assign new_n1659 = new_n1616 & new_n1619;
  assign new_n1660 = ~new_n1654 & new_n1659;
  assign new_n1661 = ~new_n1616 & new_n1618;
  assign new_n1662 = new_n1622 & new_n1661;
  assign new_n1663 = ~new_n1660 & ~new_n1662;
  assign new_n1664 = ~new_n1658 & new_n1663;
  assign new_n1665 = ~new_n1653 & new_n1664;
  assign new_n1666 = new_n1648 & new_n1649;
  assign new_n1667 = ~new_n1627 & new_n1666;
  assign new_n1668 = new_n1665 & ~new_n1667;
  assign new_n1669 = ~new_n1631 & ~new_n1634;
  assign new_n1670 = new_n1640 & ~new_n1669;
  assign new_n1671 = ~new_n1636 & new_n1670;
  assign new_n1672 = ~new_n1640 & new_n1669;
  assign new_n1673 = ~A18 & ~new_n1639;
  assign new_n1674 = new_n1672 & ~new_n1673;
  assign new_n1675 = ~new_n1669 & new_n1673;
  assign new_n1676 = ~new_n1674 & ~new_n1675;
  assign new_n1677 = new_n1635 & ~new_n1676;
  assign new_n1678 = ~A18 & ~new_n1672;
  assign new_n1679 = ~new_n1639 & ~new_n1669;
  assign new_n1680 = new_n1639 & new_n1669;
  assign new_n1681 = ~new_n1679 & ~new_n1680;
  assign new_n1682 = A18 & ~new_n1681;
  assign new_n1683 = ~new_n1635 & ~new_n1678;
  assign new_n1684 = ~new_n1682 & new_n1683;
  assign new_n1685 = ~new_n1671 & ~new_n1677;
  assign new_n1686 = ~new_n1684 & new_n1685;
  assign new_n1687 = ~new_n1668 & ~new_n1686;
  assign new_n1688 = new_n1668 & new_n1686;
  assign new_n1689 = ~new_n1687 & ~new_n1688;
  assign new_n1690 = ~new_n1645 & new_n1689;
  assign new_n1691 = new_n1645 & ~new_n1689;
  assign new_n1692 = ~new_n1690 & ~new_n1691;
  assign new_n1693 = new_n1614 & new_n1692;
  assign new_n1694 = ~new_n1614 & ~new_n1692;
  assign new_n1695 = ~new_n1693 & ~new_n1694;
  assign new_n1696 = ~new_n1629 & new_n1644;
  assign new_n1697 = ~new_n1645 & ~new_n1696;
  assign new_n1698 = ~new_n1571 & ~new_n1584;
  assign new_n1699 = ~new_n1585 & ~new_n1698;
  assign new_n1700 = new_n1697 & new_n1699;
  assign new_n1701 = ~new_n1697 & ~new_n1699;
  assign new_n1702 = ~new_n1700 & ~new_n1701;
  assign new_n1703 = ~new_n1457 & ~new_n1458;
  assign new_n1704 = new_n1456 & ~new_n1478;
  assign new_n1705 = ~new_n1480 & ~new_n1704;
  assign new_n1706 = new_n1703 & ~new_n1705;
  assign new_n1707 = ~new_n1703 & new_n1705;
  assign new_n1708 = ~new_n1706 & ~new_n1707;
  assign new_n1709 = new_n1702 & ~new_n1708;
  assign new_n1710 = ~new_n1700 & ~new_n1709;
  assign new_n1711 = new_n1695 & ~new_n1710;
  assign new_n1712 = ~new_n1695 & new_n1710;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = ~new_n1525 & new_n1713;
  assign new_n1715 = new_n1695 & new_n1709;
  assign new_n1716 = ~new_n1714 & ~new_n1715;
  assign new_n1717 = ~new_n1609 & ~new_n1612;
  assign new_n1718 = ~new_n1531 & ~new_n1554;
  assign new_n1719 = ~new_n1539 & ~new_n1718;
  assign new_n1720 = ~new_n1561 & ~new_n1605;
  assign new_n1721 = ~new_n1596 & ~new_n1720;
  assign new_n1722 = new_n1719 & new_n1721;
  assign new_n1723 = ~new_n1719 & ~new_n1721;
  assign new_n1724 = ~new_n1722 & ~new_n1723;
  assign new_n1725 = new_n1717 & ~new_n1724;
  assign new_n1726 = ~new_n1717 & new_n1724;
  assign new_n1727 = ~new_n1725 & ~new_n1726;
  assign new_n1728 = ~new_n1687 & ~new_n1690;
  assign new_n1729 = ~new_n1619 & ~new_n1665;
  assign new_n1730 = ~new_n1656 & ~new_n1729;
  assign new_n1731 = ~new_n1674 & ~new_n1684;
  assign new_n1732 = new_n1730 & new_n1731;
  assign new_n1733 = ~new_n1730 & ~new_n1731;
  assign new_n1734 = ~new_n1732 & ~new_n1733;
  assign new_n1735 = new_n1728 & ~new_n1734;
  assign new_n1736 = ~new_n1728 & new_n1734;
  assign new_n1737 = ~new_n1735 & ~new_n1736;
  assign new_n1738 = ~new_n1694 & ~new_n1700;
  assign new_n1739 = ~new_n1693 & ~new_n1738;
  assign new_n1740 = ~new_n1737 & new_n1739;
  assign new_n1741 = new_n1737 & ~new_n1739;
  assign new_n1742 = ~new_n1740 & ~new_n1741;
  assign new_n1743 = ~new_n1727 & new_n1742;
  assign new_n1744 = new_n1727 & ~new_n1742;
  assign new_n1745 = ~new_n1743 & ~new_n1744;
  assign new_n1746 = ~new_n1716 & new_n1745;
  assign new_n1747 = ~new_n1507 & ~new_n1513;
  assign new_n1748 = ~new_n1484 & ~new_n1487;
  assign new_n1749 = new_n1747 & ~new_n1748;
  assign new_n1750 = ~new_n1747 & new_n1748;
  assign new_n1751 = ~new_n1749 & ~new_n1750;
  assign new_n1752 = new_n1499 & ~new_n1523;
  assign new_n1753 = ~A999 & ~new_n1451;
  assign new_n1754 = ~new_n1452 & ~new_n1753;
  assign new_n1755 = ~new_n1515 & new_n1754;
  assign new_n1756 = new_n1752 & new_n1755;
  assign new_n1757 = ~new_n1516 & ~new_n1521;
  assign new_n1758 = ~new_n1752 & new_n1757;
  assign new_n1759 = ~new_n1756 & ~new_n1758;
  assign new_n1760 = new_n1751 & ~new_n1759;
  assign new_n1761 = ~new_n1751 & new_n1759;
  assign new_n1762 = ~new_n1760 & ~new_n1761;
  assign new_n1763 = new_n1716 & ~new_n1745;
  assign new_n1764 = ~new_n1746 & ~new_n1763;
  assign new_n1765 = ~new_n1762 & new_n1764;
  assign new_n1766 = ~new_n1746 & ~new_n1765;
  assign new_n1767 = ~new_n1732 & ~new_n1736;
  assign new_n1768 = ~new_n1722 & ~new_n1726;
  assign new_n1769 = ~new_n1767 & ~new_n1768;
  assign new_n1770 = new_n1767 & new_n1768;
  assign new_n1771 = ~new_n1769 & ~new_n1770;
  assign new_n1772 = ~new_n1740 & ~new_n1743;
  assign new_n1773 = new_n1771 & ~new_n1772;
  assign new_n1774 = ~new_n1771 & new_n1772;
  assign new_n1775 = ~new_n1773 & ~new_n1774;
  assign new_n1776 = new_n1749 & new_n1756;
  assign new_n1777 = ~new_n1750 & ~new_n1760;
  assign new_n1778 = ~new_n1756 & ~new_n1777;
  assign new_n1779 = ~new_n1776 & ~new_n1778;
  assign new_n1780 = ~new_n1775 & ~new_n1779;
  assign new_n1781 = new_n1775 & new_n1779;
  assign new_n1782 = ~new_n1780 & ~new_n1781;
  assign new_n1783 = ~new_n1766 & new_n1782;
  assign new_n1784 = new_n1766 & ~new_n1782;
  assign new_n1785 = ~new_n1783 & ~new_n1784;
  assign new_n1786 = A56 & A57;
  assign new_n1787 = ~A56 & ~A57;
  assign new_n1788 = ~new_n1786 & ~new_n1787;
  assign new_n1789 = A55 & ~new_n1788;
  assign new_n1790 = ~A55 & new_n1788;
  assign new_n1791 = ~new_n1789 & ~new_n1790;
  assign new_n1792 = A60 & ~new_n1791;
  assign new_n1793 = ~A58 & ~A59;
  assign new_n1794 = ~A60 & new_n1791;
  assign new_n1795 = ~new_n1792 & ~new_n1794;
  assign new_n1796 = A58 & A59;
  assign new_n1797 = ~new_n1793 & ~new_n1796;
  assign new_n1798 = ~new_n1795 & new_n1797;
  assign new_n1799 = ~new_n1793 & ~new_n1798;
  assign new_n1800 = ~new_n1792 & ~new_n1799;
  assign new_n1801 = new_n1792 & new_n1796;
  assign new_n1802 = ~new_n1800 & ~new_n1801;
  assign new_n1803 = ~new_n1787 & ~new_n1790;
  assign new_n1804 = new_n1802 & ~new_n1803;
  assign new_n1805 = ~new_n1802 & new_n1803;
  assign new_n1806 = ~new_n1804 & ~new_n1805;
  assign new_n1807 = new_n1795 & ~new_n1797;
  assign new_n1808 = ~new_n1798 & ~new_n1807;
  assign new_n1809 = A64 & A65;
  assign new_n1810 = ~A64 & ~A65;
  assign new_n1811 = ~new_n1809 & ~new_n1810;
  assign new_n1812 = A61 & A62;
  assign new_n1813 = ~A61 & ~A62;
  assign new_n1814 = ~new_n1812 & ~new_n1813;
  assign new_n1815 = ~A63 & A66;
  assign new_n1816 = A63 & ~A66;
  assign new_n1817 = ~new_n1815 & ~new_n1816;
  assign new_n1818 = new_n1814 & ~new_n1817;
  assign new_n1819 = ~new_n1814 & new_n1817;
  assign new_n1820 = ~new_n1818 & ~new_n1819;
  assign new_n1821 = new_n1811 & new_n1820;
  assign new_n1822 = ~new_n1811 & ~new_n1820;
  assign new_n1823 = ~new_n1821 & ~new_n1822;
  assign new_n1824 = ~new_n1808 & new_n1823;
  assign new_n1825 = new_n1809 & new_n1815;
  assign new_n1826 = A66 & ~new_n1811;
  assign new_n1827 = ~A63 & ~new_n1812;
  assign new_n1828 = ~A66 & ~new_n1809;
  assign new_n1829 = ~new_n1827 & ~new_n1828;
  assign new_n1830 = ~new_n1826 & new_n1829;
  assign new_n1831 = ~new_n1825 & ~new_n1830;
  assign new_n1832 = ~new_n1813 & ~new_n1831;
  assign new_n1833 = A63 & A66;
  assign new_n1834 = ~new_n1809 & ~new_n1812;
  assign new_n1835 = new_n1833 & ~new_n1834;
  assign new_n1836 = A65 & new_n1812;
  assign new_n1837 = new_n1835 & ~new_n1836;
  assign new_n1838 = new_n1810 & new_n1813;
  assign new_n1839 = ~new_n1833 & new_n1838;
  assign new_n1840 = ~new_n1810 & new_n1812;
  assign new_n1841 = new_n1816 & new_n1840;
  assign new_n1842 = ~new_n1839 & ~new_n1841;
  assign new_n1843 = ~new_n1837 & new_n1842;
  assign new_n1844 = ~new_n1832 & new_n1843;
  assign new_n1845 = new_n1827 & new_n1828;
  assign new_n1846 = ~new_n1821 & new_n1845;
  assign new_n1847 = new_n1844 & ~new_n1846;
  assign new_n1848 = new_n1824 & new_n1847;
  assign new_n1849 = ~new_n1824 & ~new_n1847;
  assign new_n1850 = ~new_n1848 & ~new_n1849;
  assign new_n1851 = ~new_n1806 & new_n1850;
  assign new_n1852 = new_n1806 & ~new_n1850;
  assign new_n1853 = ~new_n1851 & ~new_n1852;
  assign new_n1854 = new_n1808 & ~new_n1823;
  assign new_n1855 = ~new_n1824 & ~new_n1854;
  assign new_n1856 = A76 & A77;
  assign new_n1857 = ~A76 & ~A77;
  assign new_n1858 = ~new_n1856 & ~new_n1857;
  assign new_n1859 = A73 & A74;
  assign new_n1860 = ~A73 & ~A74;
  assign new_n1861 = ~new_n1859 & ~new_n1860;
  assign new_n1862 = ~A75 & A78;
  assign new_n1863 = A75 & ~A78;
  assign new_n1864 = ~new_n1862 & ~new_n1863;
  assign new_n1865 = new_n1861 & ~new_n1864;
  assign new_n1866 = ~new_n1861 & new_n1864;
  assign new_n1867 = ~new_n1865 & ~new_n1866;
  assign new_n1868 = new_n1858 & new_n1867;
  assign new_n1869 = ~new_n1858 & ~new_n1867;
  assign new_n1870 = ~new_n1868 & ~new_n1869;
  assign new_n1871 = A69 & ~A72;
  assign new_n1872 = ~A69 & A72;
  assign new_n1873 = ~new_n1871 & ~new_n1872;
  assign new_n1874 = ~A67 & ~A68;
  assign new_n1875 = A67 & A68;
  assign new_n1876 = ~new_n1874 & ~new_n1875;
  assign new_n1877 = ~A70 & ~A71;
  assign new_n1878 = A70 & A71;
  assign new_n1879 = ~new_n1877 & ~new_n1878;
  assign new_n1880 = new_n1876 & ~new_n1879;
  assign new_n1881 = ~new_n1876 & new_n1879;
  assign new_n1882 = ~new_n1880 & ~new_n1881;
  assign new_n1883 = new_n1873 & new_n1882;
  assign new_n1884 = ~new_n1873 & ~new_n1882;
  assign new_n1885 = ~new_n1883 & ~new_n1884;
  assign new_n1886 = new_n1870 & new_n1885;
  assign new_n1887 = ~new_n1870 & ~new_n1885;
  assign new_n1888 = ~new_n1886 & ~new_n1887;
  assign new_n1889 = new_n1855 & new_n1888;
  assign new_n1890 = ~A69 & ~new_n1875;
  assign new_n1891 = ~new_n1874 & ~new_n1890;
  assign new_n1892 = A69 & new_n1875;
  assign new_n1893 = ~A70 & ~new_n1892;
  assign new_n1894 = new_n1891 & ~new_n1893;
  assign new_n1895 = A71 & new_n1894;
  assign new_n1896 = A69 & A70;
  assign new_n1897 = new_n1875 & new_n1896;
  assign new_n1898 = ~new_n1895 & ~new_n1897;
  assign new_n1899 = ~A72 & ~new_n1898;
  assign new_n1900 = A71 & A72;
  assign new_n1901 = new_n1874 & ~new_n1896;
  assign new_n1902 = ~new_n1892 & new_n1900;
  assign new_n1903 = ~new_n1901 & new_n1902;
  assign new_n1904 = A70 & ~new_n1903;
  assign new_n1905 = new_n1891 & new_n1900;
  assign new_n1906 = ~A71 & ~A72;
  assign new_n1907 = ~new_n1874 & ~new_n1906;
  assign new_n1908 = new_n1890 & ~new_n1900;
  assign new_n1909 = ~new_n1907 & new_n1908;
  assign new_n1910 = ~A70 & ~new_n1905;
  assign new_n1911 = ~new_n1909 & new_n1910;
  assign new_n1912 = ~new_n1904 & ~new_n1911;
  assign new_n1913 = ~A71 & A72;
  assign new_n1914 = new_n1894 & new_n1913;
  assign new_n1915 = ~new_n1899 & ~new_n1914;
  assign new_n1916 = ~new_n1912 & new_n1915;
  assign new_n1917 = new_n1901 & new_n1906;
  assign new_n1918 = new_n1916 & ~new_n1917;
  assign new_n1919 = new_n1856 & new_n1862;
  assign new_n1920 = A78 & ~new_n1858;
  assign new_n1921 = ~A75 & ~new_n1859;
  assign new_n1922 = ~A78 & ~new_n1856;
  assign new_n1923 = ~new_n1921 & ~new_n1922;
  assign new_n1924 = ~new_n1920 & new_n1923;
  assign new_n1925 = ~new_n1919 & ~new_n1924;
  assign new_n1926 = ~new_n1860 & ~new_n1925;
  assign new_n1927 = A75 & A78;
  assign new_n1928 = ~new_n1856 & ~new_n1859;
  assign new_n1929 = new_n1927 & ~new_n1928;
  assign new_n1930 = A77 & new_n1859;
  assign new_n1931 = new_n1929 & ~new_n1930;
  assign new_n1932 = new_n1857 & new_n1860;
  assign new_n1933 = ~new_n1927 & new_n1932;
  assign new_n1934 = ~new_n1857 & new_n1859;
  assign new_n1935 = new_n1863 & new_n1934;
  assign new_n1936 = ~new_n1933 & ~new_n1935;
  assign new_n1937 = ~new_n1931 & new_n1936;
  assign new_n1938 = ~new_n1926 & new_n1937;
  assign new_n1939 = new_n1921 & new_n1922;
  assign new_n1940 = ~new_n1868 & new_n1939;
  assign new_n1941 = new_n1938 & ~new_n1940;
  assign new_n1942 = ~new_n1886 & ~new_n1941;
  assign new_n1943 = new_n1886 & new_n1941;
  assign new_n1944 = ~new_n1942 & ~new_n1943;
  assign new_n1945 = ~new_n1918 & new_n1944;
  assign new_n1946 = new_n1918 & ~new_n1944;
  assign new_n1947 = ~new_n1945 & ~new_n1946;
  assign new_n1948 = ~new_n1889 & new_n1947;
  assign new_n1949 = new_n1889 & ~new_n1947;
  assign new_n1950 = ~new_n1948 & ~new_n1949;
  assign new_n1951 = ~new_n1853 & new_n1950;
  assign new_n1952 = new_n1853 & ~new_n1950;
  assign new_n1953 = ~new_n1951 & ~new_n1952;
  assign new_n1954 = A34 & A35;
  assign new_n1955 = ~A34 & ~A35;
  assign new_n1956 = ~new_n1954 & ~new_n1955;
  assign new_n1957 = A31 & A32;
  assign new_n1958 = ~A31 & ~A32;
  assign new_n1959 = ~new_n1957 & ~new_n1958;
  assign new_n1960 = ~A33 & A36;
  assign new_n1961 = A33 & ~A36;
  assign new_n1962 = ~new_n1960 & ~new_n1961;
  assign new_n1963 = new_n1959 & ~new_n1962;
  assign new_n1964 = ~new_n1959 & new_n1962;
  assign new_n1965 = ~new_n1963 & ~new_n1964;
  assign new_n1966 = new_n1956 & new_n1965;
  assign new_n1967 = ~new_n1956 & ~new_n1965;
  assign new_n1968 = ~new_n1966 & ~new_n1967;
  assign new_n1969 = A38 & A39;
  assign new_n1970 = ~A38 & ~A39;
  assign new_n1971 = ~new_n1969 & ~new_n1970;
  assign new_n1972 = A37 & ~new_n1971;
  assign new_n1973 = ~A37 & new_n1971;
  assign new_n1974 = ~new_n1972 & ~new_n1973;
  assign new_n1975 = A42 & ~new_n1974;
  assign new_n1976 = ~A42 & new_n1974;
  assign new_n1977 = ~new_n1975 & ~new_n1976;
  assign new_n1978 = A40 & A41;
  assign new_n1979 = ~A40 & ~A41;
  assign new_n1980 = ~new_n1978 & ~new_n1979;
  assign new_n1981 = new_n1977 & ~new_n1980;
  assign new_n1982 = ~new_n1977 & new_n1980;
  assign new_n1983 = ~new_n1981 & ~new_n1982;
  assign new_n1984 = new_n1968 & ~new_n1983;
  assign new_n1985 = ~new_n1968 & new_n1983;
  assign new_n1986 = ~new_n1984 & ~new_n1985;
  assign new_n1987 = A46 & A47;
  assign new_n1988 = ~A46 & ~A47;
  assign new_n1989 = ~new_n1987 & ~new_n1988;
  assign new_n1990 = ~A43 & ~A44;
  assign new_n1991 = A43 & A44;
  assign new_n1992 = ~new_n1990 & ~new_n1991;
  assign new_n1993 = ~A45 & A48;
  assign new_n1994 = A45 & ~A48;
  assign new_n1995 = ~new_n1993 & ~new_n1994;
  assign new_n1996 = new_n1992 & ~new_n1995;
  assign new_n1997 = ~new_n1992 & new_n1995;
  assign new_n1998 = ~new_n1996 & ~new_n1997;
  assign new_n1999 = new_n1989 & new_n1998;
  assign new_n2000 = ~new_n1989 & ~new_n1998;
  assign new_n2001 = ~new_n1999 & ~new_n2000;
  assign new_n2002 = A50 & A51;
  assign new_n2003 = ~A50 & ~A51;
  assign new_n2004 = ~new_n2002 & ~new_n2003;
  assign new_n2005 = A49 & ~new_n2004;
  assign new_n2006 = ~A49 & new_n2004;
  assign new_n2007 = ~new_n2005 & ~new_n2006;
  assign new_n2008 = A52 & A54;
  assign new_n2009 = ~A52 & ~A54;
  assign new_n2010 = ~new_n2008 & ~new_n2009;
  assign new_n2011 = A53 & ~new_n2010;
  assign new_n2012 = ~A53 & new_n2010;
  assign new_n2013 = ~new_n2011 & ~new_n2012;
  assign new_n2014 = ~new_n2007 & ~new_n2013;
  assign new_n2015 = new_n2007 & new_n2013;
  assign new_n2016 = ~new_n2014 & ~new_n2015;
  assign new_n2017 = new_n2001 & new_n2016;
  assign new_n2018 = ~new_n2001 & ~new_n2016;
  assign new_n2019 = ~new_n2017 & ~new_n2018;
  assign new_n2020 = new_n1986 & new_n2019;
  assign new_n2021 = ~new_n1984 & ~new_n2020;
  assign new_n2022 = new_n1954 & new_n1960;
  assign new_n2023 = A36 & ~new_n1956;
  assign new_n2024 = ~A33 & ~new_n1957;
  assign new_n2025 = ~A36 & ~new_n1954;
  assign new_n2026 = ~new_n2024 & ~new_n2025;
  assign new_n2027 = ~new_n2023 & new_n2026;
  assign new_n2028 = ~new_n2022 & ~new_n2027;
  assign new_n2029 = ~new_n1958 & ~new_n2028;
  assign new_n2030 = A33 & A36;
  assign new_n2031 = ~new_n1954 & ~new_n1957;
  assign new_n2032 = new_n2030 & ~new_n2031;
  assign new_n2033 = A35 & new_n1957;
  assign new_n2034 = new_n2032 & ~new_n2033;
  assign new_n2035 = new_n1955 & new_n1958;
  assign new_n2036 = ~new_n2030 & new_n2035;
  assign new_n2037 = ~new_n1955 & new_n1957;
  assign new_n2038 = new_n1961 & new_n2037;
  assign new_n2039 = ~new_n2036 & ~new_n2038;
  assign new_n2040 = ~new_n2034 & new_n2039;
  assign new_n2041 = ~new_n2029 & new_n2040;
  assign new_n2042 = new_n2024 & new_n2025;
  assign new_n2043 = ~new_n1966 & new_n2042;
  assign new_n2044 = new_n2041 & ~new_n2043;
  assign new_n2045 = ~new_n1970 & ~new_n1973;
  assign new_n2046 = new_n1979 & ~new_n2045;
  assign new_n2047 = ~new_n1975 & new_n2046;
  assign new_n2048 = ~new_n1979 & new_n2045;
  assign new_n2049 = ~A42 & ~new_n1978;
  assign new_n2050 = new_n2048 & ~new_n2049;
  assign new_n2051 = ~new_n2045 & new_n2049;
  assign new_n2052 = ~new_n2050 & ~new_n2051;
  assign new_n2053 = new_n1974 & ~new_n2052;
  assign new_n2054 = ~A42 & ~new_n2048;
  assign new_n2055 = ~new_n1978 & ~new_n2045;
  assign new_n2056 = new_n1978 & new_n2045;
  assign new_n2057 = ~new_n2055 & ~new_n2056;
  assign new_n2058 = A42 & ~new_n2057;
  assign new_n2059 = ~new_n1974 & ~new_n2054;
  assign new_n2060 = ~new_n2058 & new_n2059;
  assign new_n2061 = ~new_n2047 & ~new_n2053;
  assign new_n2062 = ~new_n2060 & new_n2061;
  assign new_n2063 = ~new_n2044 & ~new_n2062;
  assign new_n2064 = new_n2044 & new_n2062;
  assign new_n2065 = ~new_n2063 & ~new_n2064;
  assign new_n2066 = ~new_n2014 & ~new_n2017;
  assign new_n2067 = ~new_n2009 & ~new_n2012;
  assign new_n2068 = ~new_n2003 & ~new_n2006;
  assign new_n2069 = new_n2067 & new_n2068;
  assign new_n2070 = ~new_n2067 & ~new_n2068;
  assign new_n2071 = ~new_n2069 & ~new_n2070;
  assign new_n2072 = new_n1987 & new_n1993;
  assign new_n2073 = A48 & ~new_n1989;
  assign new_n2074 = ~A45 & ~new_n1991;
  assign new_n2075 = ~A48 & ~new_n1987;
  assign new_n2076 = ~new_n2074 & ~new_n2075;
  assign new_n2077 = ~new_n2073 & new_n2076;
  assign new_n2078 = ~new_n2072 & ~new_n2077;
  assign new_n2079 = ~new_n1990 & ~new_n2078;
  assign new_n2080 = A45 & A48;
  assign new_n2081 = ~new_n1987 & ~new_n1991;
  assign new_n2082 = new_n2080 & ~new_n2081;
  assign new_n2083 = A47 & new_n1991;
  assign new_n2084 = new_n2082 & ~new_n2083;
  assign new_n2085 = new_n1988 & new_n1990;
  assign new_n2086 = ~new_n2080 & new_n2085;
  assign new_n2087 = ~new_n1988 & new_n1991;
  assign new_n2088 = new_n1994 & new_n2087;
  assign new_n2089 = ~new_n2086 & ~new_n2088;
  assign new_n2090 = ~new_n2084 & new_n2089;
  assign new_n2091 = ~new_n2079 & new_n2090;
  assign new_n2092 = new_n2074 & new_n2075;
  assign new_n2093 = ~new_n1999 & new_n2092;
  assign new_n2094 = new_n2091 & ~new_n2093;
  assign new_n2095 = ~new_n2071 & ~new_n2094;
  assign new_n2096 = new_n2071 & new_n2094;
  assign new_n2097 = ~new_n2095 & ~new_n2096;
  assign new_n2098 = new_n2066 & ~new_n2097;
  assign new_n2099 = ~new_n2066 & new_n2097;
  assign new_n2100 = ~new_n2098 & ~new_n2099;
  assign new_n2101 = ~new_n2065 & ~new_n2100;
  assign new_n2102 = new_n2065 & new_n2100;
  assign new_n2103 = ~new_n2101 & ~new_n2102;
  assign new_n2104 = new_n2021 & new_n2103;
  assign new_n2105 = ~new_n2021 & ~new_n2103;
  assign new_n2106 = ~new_n2104 & ~new_n2105;
  assign new_n2107 = new_n1953 & new_n2106;
  assign new_n2108 = ~new_n1986 & ~new_n2019;
  assign new_n2109 = ~new_n2020 & ~new_n2108;
  assign new_n2110 = ~new_n1855 & ~new_n1888;
  assign new_n2111 = ~new_n1889 & ~new_n2110;
  assign new_n2112 = new_n2109 & new_n2111;
  assign new_n2113 = ~new_n1953 & ~new_n2106;
  assign new_n2114 = ~new_n2107 & ~new_n2113;
  assign new_n2115 = ~new_n2112 & new_n2114;
  assign new_n2116 = ~new_n2107 & ~new_n2115;
  assign new_n2117 = ~new_n1958 & ~new_n2041;
  assign new_n2118 = ~new_n2032 & ~new_n2117;
  assign new_n2119 = ~new_n2050 & ~new_n2060;
  assign new_n2120 = new_n2118 & new_n2119;
  assign new_n2121 = ~new_n2118 & ~new_n2119;
  assign new_n2122 = ~new_n2120 & ~new_n2121;
  assign new_n2123 = ~new_n1984 & new_n2065;
  assign new_n2124 = ~new_n2063 & ~new_n2123;
  assign new_n2125 = ~new_n2122 & new_n2124;
  assign new_n2126 = new_n2122 & ~new_n2124;
  assign new_n2127 = ~new_n2125 & ~new_n2126;
  assign new_n2128 = new_n2014 & ~new_n2071;
  assign new_n2129 = ~new_n2014 & new_n2071;
  assign new_n2130 = ~new_n2128 & ~new_n2129;
  assign new_n2131 = new_n2094 & ~new_n2130;
  assign new_n2132 = new_n2017 & ~new_n2095;
  assign new_n2133 = ~new_n2131 & ~new_n2132;
  assign new_n2134 = ~new_n1990 & ~new_n2091;
  assign new_n2135 = ~new_n2082 & ~new_n2134;
  assign new_n2136 = ~new_n2070 & ~new_n2129;
  assign new_n2137 = new_n2135 & ~new_n2136;
  assign new_n2138 = ~new_n2135 & new_n2136;
  assign new_n2139 = ~new_n2137 & ~new_n2138;
  assign new_n2140 = new_n2133 & ~new_n2139;
  assign new_n2141 = ~new_n2133 & new_n2139;
  assign new_n2142 = ~new_n2140 & ~new_n2141;
  assign new_n2143 = new_n1984 & ~new_n2065;
  assign new_n2144 = ~new_n2123 & ~new_n2143;
  assign new_n2145 = new_n2100 & ~new_n2144;
  assign new_n2146 = new_n2020 & ~new_n2101;
  assign new_n2147 = ~new_n2145 & ~new_n2146;
  assign new_n2148 = ~new_n2142 & new_n2147;
  assign new_n2149 = new_n2142 & ~new_n2147;
  assign new_n2150 = ~new_n2148 & ~new_n2149;
  assign new_n2151 = new_n2127 & new_n2150;
  assign new_n2152 = ~new_n2127 & ~new_n2150;
  assign new_n2153 = ~new_n2151 & ~new_n2152;
  assign new_n2154 = ~new_n2116 & new_n2153;
  assign new_n2155 = ~new_n1942 & ~new_n1945;
  assign new_n2156 = ~new_n1893 & ~new_n1916;
  assign new_n2157 = ~new_n1905 & ~new_n2156;
  assign new_n2158 = ~new_n1860 & ~new_n1938;
  assign new_n2159 = ~new_n1929 & ~new_n2158;
  assign new_n2160 = new_n2157 & new_n2159;
  assign new_n2161 = ~new_n2157 & ~new_n2159;
  assign new_n2162 = ~new_n2160 & ~new_n2161;
  assign new_n2163 = new_n2155 & ~new_n2162;
  assign new_n2164 = ~new_n2155 & new_n2162;
  assign new_n2165 = ~new_n2163 & ~new_n2164;
  assign new_n2166 = ~new_n1813 & ~new_n1844;
  assign new_n2167 = ~new_n1835 & ~new_n2166;
  assign new_n2168 = ~new_n1800 & ~new_n1804;
  assign new_n2169 = new_n2167 & ~new_n2168;
  assign new_n2170 = ~new_n2167 & new_n2168;
  assign new_n2171 = ~new_n2169 & ~new_n2170;
  assign new_n2172 = ~new_n1848 & ~new_n1851;
  assign new_n2173 = new_n2171 & new_n2172;
  assign new_n2174 = ~new_n2171 & ~new_n2172;
  assign new_n2175 = ~new_n2173 & ~new_n2174;
  assign new_n2176 = ~new_n1948 & ~new_n1951;
  assign new_n2177 = ~new_n2175 & new_n2176;
  assign new_n2178 = new_n2175 & ~new_n2176;
  assign new_n2179 = ~new_n2177 & ~new_n2178;
  assign new_n2180 = ~new_n2165 & new_n2179;
  assign new_n2181 = new_n2165 & ~new_n2179;
  assign new_n2182 = ~new_n2180 & ~new_n2181;
  assign new_n2183 = new_n2116 & ~new_n2153;
  assign new_n2184 = ~new_n2154 & ~new_n2183;
  assign new_n2185 = ~new_n2182 & new_n2184;
  assign new_n2186 = ~new_n2154 & ~new_n2185;
  assign new_n2187 = ~new_n2169 & ~new_n2173;
  assign new_n2188 = ~new_n2160 & ~new_n2164;
  assign new_n2189 = ~new_n2187 & ~new_n2188;
  assign new_n2190 = new_n2187 & new_n2188;
  assign new_n2191 = ~new_n2189 & ~new_n2190;
  assign new_n2192 = ~new_n2177 & ~new_n2180;
  assign new_n2193 = new_n2191 & new_n2192;
  assign new_n2194 = ~new_n2191 & ~new_n2192;
  assign new_n2195 = ~new_n2193 & ~new_n2194;
  assign new_n2196 = ~new_n2138 & ~new_n2141;
  assign new_n2197 = ~new_n2120 & ~new_n2126;
  assign new_n2198 = new_n2196 & ~new_n2197;
  assign new_n2199 = ~new_n2196 & new_n2197;
  assign new_n2200 = ~new_n2198 & ~new_n2199;
  assign new_n2201 = ~new_n2148 & ~new_n2151;
  assign new_n2202 = new_n2200 & new_n2201;
  assign new_n2203 = ~new_n2200 & ~new_n2201;
  assign new_n2204 = ~new_n2202 & ~new_n2203;
  assign new_n2205 = ~new_n2195 & new_n2204;
  assign new_n2206 = new_n2195 & ~new_n2204;
  assign new_n2207 = ~new_n2205 & ~new_n2206;
  assign new_n2208 = new_n2186 & new_n2207;
  assign new_n2209 = ~new_n2186 & ~new_n2207;
  assign new_n2210 = ~new_n2208 & ~new_n2209;
  assign new_n2211 = new_n1785 & new_n2210;
  assign new_n2212 = ~new_n1785 & ~new_n2210;
  assign new_n2213 = ~new_n2211 & ~new_n2212;
  assign new_n2214 = new_n1762 & ~new_n1764;
  assign new_n2215 = ~new_n1765 & ~new_n2214;
  assign new_n2216 = new_n2182 & ~new_n2184;
  assign new_n2217 = ~new_n2185 & ~new_n2216;
  assign new_n2218 = ~new_n2215 & new_n2217;
  assign new_n2219 = new_n1525 & ~new_n1713;
  assign new_n2220 = ~new_n1714 & ~new_n2219;
  assign new_n2221 = ~new_n2109 & ~new_n2111;
  assign new_n2222 = ~new_n1702 & new_n1708;
  assign new_n2223 = ~new_n1709 & ~new_n2222;
  assign new_n2224 = ~new_n2112 & ~new_n2221;
  assign new_n2225 = ~new_n2223 & new_n2224;
  assign new_n2226 = ~new_n2221 & ~new_n2225;
  assign new_n2227 = ~new_n2220 & ~new_n2226;
  assign new_n2228 = new_n2220 & new_n2226;
  assign new_n2229 = ~new_n2227 & ~new_n2228;
  assign new_n2230 = ~new_n2114 & ~new_n2229;
  assign new_n2231 = ~new_n2115 & ~new_n2230;
  assign new_n2232 = ~new_n2227 & ~new_n2231;
  assign new_n2233 = new_n2215 & ~new_n2217;
  assign new_n2234 = ~new_n2218 & ~new_n2233;
  assign new_n2235 = ~new_n2232 & new_n2234;
  assign new_n2236 = ~new_n2218 & ~new_n2235;
  assign new_n2237 = new_n2213 & new_n2236;
  assign new_n2238 = ~new_n2213 & ~new_n2236;
  assign new_n2239 = ~new_n2237 & ~new_n2238;
  assign new_n2240 = ~new_n1401 & ~new_n1424;
  assign new_n2241 = ~new_n1425 & ~new_n2240;
  assign new_n2242 = new_n2239 & new_n2241;
  assign new_n2243 = new_n1420 & ~new_n1422;
  assign new_n2244 = ~new_n1423 & ~new_n2243;
  assign new_n2245 = new_n1413 & ~new_n1415;
  assign new_n2246 = new_n2223 & ~new_n2224;
  assign new_n2247 = ~new_n2225 & ~new_n2246;
  assign new_n2248 = ~new_n1410 & ~new_n1412;
  assign new_n2249 = ~new_n1413 & ~new_n2248;
  assign new_n2250 = ~new_n2247 & new_n2249;
  assign new_n2251 = ~new_n1416 & ~new_n2245;
  assign new_n2252 = ~new_n2250 & new_n2251;
  assign new_n2253 = new_n2114 & new_n2229;
  assign new_n2254 = ~new_n2230 & ~new_n2253;
  assign new_n2255 = new_n1415 & new_n2250;
  assign new_n2256 = ~new_n2252 & ~new_n2255;
  assign new_n2257 = ~new_n2254 & new_n2256;
  assign new_n2258 = ~new_n2252 & ~new_n2257;
  assign new_n2259 = new_n2244 & ~new_n2258;
  assign new_n2260 = new_n2232 & ~new_n2234;
  assign new_n2261 = ~new_n2235 & ~new_n2260;
  assign new_n2262 = ~new_n2244 & new_n2258;
  assign new_n2263 = ~new_n2259 & ~new_n2262;
  assign new_n2264 = new_n2261 & new_n2263;
  assign new_n2265 = ~new_n2259 & ~new_n2264;
  assign new_n2266 = ~new_n2239 & ~new_n2241;
  assign new_n2267 = ~new_n2242 & ~new_n2266;
  assign new_n2268 = new_n2265 & new_n2267;
  assign new_n2269 = ~new_n2242 & ~new_n2268;
  assign new_n2270 = new_n1429 & new_n2269;
  assign new_n2271 = ~new_n2211 & ~new_n2237;
  assign new_n2272 = ~new_n1770 & ~new_n1773;
  assign new_n2273 = new_n1776 & ~new_n2272;
  assign new_n2274 = ~new_n1776 & new_n2272;
  assign new_n2275 = ~new_n2273 & ~new_n2274;
  assign new_n2276 = ~new_n1781 & ~new_n1783;
  assign new_n2277 = new_n2275 & new_n2276;
  assign new_n2278 = ~new_n2275 & ~new_n2276;
  assign new_n2279 = ~new_n2277 & ~new_n2278;
  assign new_n2280 = ~new_n2189 & ~new_n2193;
  assign new_n2281 = ~new_n2199 & ~new_n2202;
  assign new_n2282 = ~new_n2280 & new_n2281;
  assign new_n2283 = new_n2280 & ~new_n2281;
  assign new_n2284 = ~new_n2282 & ~new_n2283;
  assign new_n2285 = ~new_n2205 & ~new_n2208;
  assign new_n2286 = new_n2284 & new_n2285;
  assign new_n2287 = ~new_n2284 & ~new_n2285;
  assign new_n2288 = ~new_n2286 & ~new_n2287;
  assign new_n2289 = new_n2279 & new_n2288;
  assign new_n2290 = ~new_n2279 & ~new_n2288;
  assign new_n2291 = ~new_n2289 & ~new_n2290;
  assign new_n2292 = new_n2271 & new_n2291;
  assign new_n2293 = ~new_n2271 & ~new_n2291;
  assign new_n2294 = ~new_n2292 & ~new_n2293;
  assign new_n2295 = ~new_n1429 & ~new_n2269;
  assign new_n2296 = ~new_n2270 & ~new_n2295;
  assign new_n2297 = new_n2294 & new_n2296;
  assign new_n2298 = ~new_n2270 & ~new_n2297;
  assign new_n2299 = ~new_n1392 & ~new_n1427;
  assign new_n2300 = ~new_n2282 & ~new_n2286;
  assign new_n2301 = ~new_n2274 & ~new_n2277;
  assign new_n2302 = ~new_n2300 & ~new_n2301;
  assign new_n2303 = ~new_n2289 & ~new_n2292;
  assign new_n2304 = new_n2302 & ~new_n2303;
  assign new_n2305 = new_n2300 & new_n2301;
  assign new_n2306 = ~new_n2303 & ~new_n2305;
  assign new_n2307 = ~new_n2302 & ~new_n2306;
  assign new_n2308 = ~new_n2304 & ~new_n2307;
  assign new_n2309 = new_n2299 & new_n2308;
  assign new_n2310 = ~new_n2299 & ~new_n2308;
  assign new_n2311 = ~new_n2309 & ~new_n2310;
  assign new_n2312 = ~new_n2298 & ~new_n2311;
  assign new_n2313 = new_n2298 & new_n2311;
  assign new_n2314 = ~new_n2312 & ~new_n2313;
  assign new_n2315 = ~new_n2265 & ~new_n2267;
  assign new_n2316 = ~new_n2268 & ~new_n2315;
  assign new_n2317 = A916 & A917;
  assign new_n2318 = A913 & A914;
  assign new_n2319 = ~new_n2317 & ~new_n2318;
  assign new_n2320 = A915 & A918;
  assign new_n2321 = ~new_n2319 & new_n2320;
  assign new_n2322 = ~A913 & ~A914;
  assign new_n2323 = ~A915 & A918;
  assign new_n2324 = new_n2317 & new_n2323;
  assign new_n2325 = ~A915 & ~new_n2318;
  assign new_n2326 = ~A916 & ~A917;
  assign new_n2327 = ~new_n2317 & ~new_n2326;
  assign new_n2328 = A918 & ~new_n2327;
  assign new_n2329 = ~A918 & ~new_n2317;
  assign new_n2330 = ~new_n2325 & ~new_n2329;
  assign new_n2331 = ~new_n2328 & new_n2330;
  assign new_n2332 = ~new_n2324 & ~new_n2331;
  assign new_n2333 = ~new_n2322 & ~new_n2332;
  assign new_n2334 = A917 & new_n2318;
  assign new_n2335 = new_n2321 & ~new_n2334;
  assign new_n2336 = ~new_n2320 & new_n2322;
  assign new_n2337 = new_n2326 & new_n2336;
  assign new_n2338 = A915 & ~A918;
  assign new_n2339 = new_n2318 & ~new_n2326;
  assign new_n2340 = new_n2338 & new_n2339;
  assign new_n2341 = ~new_n2337 & ~new_n2340;
  assign new_n2342 = ~new_n2335 & new_n2341;
  assign new_n2343 = ~new_n2333 & new_n2342;
  assign new_n2344 = ~new_n2322 & ~new_n2343;
  assign new_n2345 = ~new_n2321 & ~new_n2344;
  assign new_n2346 = ~A911 & ~A912;
  assign new_n2347 = A911 & A912;
  assign new_n2348 = ~new_n2346 & ~new_n2347;
  assign new_n2349 = ~A910 & new_n2348;
  assign new_n2350 = ~new_n2346 & ~new_n2349;
  assign new_n2351 = ~A908 & ~A909;
  assign new_n2352 = A908 & A909;
  assign new_n2353 = ~new_n2351 & ~new_n2352;
  assign new_n2354 = ~A907 & new_n2353;
  assign new_n2355 = ~new_n2351 & ~new_n2354;
  assign new_n2356 = new_n2350 & new_n2355;
  assign new_n2357 = ~new_n2350 & ~new_n2355;
  assign new_n2358 = ~new_n2356 & ~new_n2357;
  assign new_n2359 = A907 & ~new_n2353;
  assign new_n2360 = ~new_n2354 & ~new_n2359;
  assign new_n2361 = A910 & ~new_n2348;
  assign new_n2362 = ~new_n2349 & ~new_n2361;
  assign new_n2363 = ~new_n2360 & ~new_n2362;
  assign new_n2364 = new_n2358 & new_n2363;
  assign new_n2365 = ~new_n2356 & ~new_n2364;
  assign new_n2366 = ~new_n2345 & ~new_n2365;
  assign new_n2367 = new_n2345 & new_n2365;
  assign new_n2368 = ~new_n2366 & ~new_n2367;
  assign new_n2369 = new_n2360 & new_n2362;
  assign new_n2370 = ~new_n2318 & ~new_n2322;
  assign new_n2371 = ~new_n2323 & ~new_n2338;
  assign new_n2372 = new_n2370 & ~new_n2371;
  assign new_n2373 = ~new_n2370 & new_n2371;
  assign new_n2374 = ~new_n2372 & ~new_n2373;
  assign new_n2375 = new_n2327 & new_n2374;
  assign new_n2376 = ~new_n2327 & ~new_n2374;
  assign new_n2377 = ~new_n2375 & ~new_n2376;
  assign new_n2378 = ~new_n2363 & ~new_n2369;
  assign new_n2379 = ~new_n2377 & new_n2378;
  assign new_n2380 = ~new_n2369 & ~new_n2379;
  assign new_n2381 = new_n2325 & new_n2329;
  assign new_n2382 = ~new_n2375 & new_n2381;
  assign new_n2383 = new_n2343 & ~new_n2382;
  assign new_n2384 = ~new_n2380 & ~new_n2383;
  assign new_n2385 = new_n2380 & new_n2383;
  assign new_n2386 = ~new_n2384 & ~new_n2385;
  assign new_n2387 = ~new_n2358 & new_n2386;
  assign new_n2388 = ~new_n2364 & ~new_n2384;
  assign new_n2389 = ~new_n2387 & new_n2388;
  assign new_n2390 = new_n2368 & new_n2389;
  assign new_n2391 = ~new_n2368 & ~new_n2389;
  assign new_n2392 = ~new_n2390 & ~new_n2391;
  assign new_n2393 = ~A901 & ~A902;
  assign new_n2394 = A904 & A905;
  assign new_n2395 = ~A903 & A906;
  assign new_n2396 = new_n2394 & new_n2395;
  assign new_n2397 = A901 & A902;
  assign new_n2398 = ~A903 & ~new_n2397;
  assign new_n2399 = ~A904 & ~A905;
  assign new_n2400 = ~new_n2394 & ~new_n2399;
  assign new_n2401 = A906 & ~new_n2400;
  assign new_n2402 = ~A906 & ~new_n2394;
  assign new_n2403 = ~new_n2398 & ~new_n2402;
  assign new_n2404 = ~new_n2401 & new_n2403;
  assign new_n2405 = ~new_n2396 & ~new_n2404;
  assign new_n2406 = ~new_n2393 & ~new_n2405;
  assign new_n2407 = A903 & A906;
  assign new_n2408 = ~new_n2394 & ~new_n2397;
  assign new_n2409 = new_n2407 & ~new_n2408;
  assign new_n2410 = A905 & new_n2397;
  assign new_n2411 = new_n2409 & ~new_n2410;
  assign new_n2412 = new_n2393 & new_n2399;
  assign new_n2413 = ~new_n2407 & new_n2412;
  assign new_n2414 = A903 & ~A906;
  assign new_n2415 = new_n2397 & ~new_n2399;
  assign new_n2416 = new_n2414 & new_n2415;
  assign new_n2417 = ~new_n2413 & ~new_n2416;
  assign new_n2418 = ~new_n2411 & new_n2417;
  assign new_n2419 = ~new_n2406 & new_n2418;
  assign new_n2420 = ~new_n2393 & ~new_n2397;
  assign new_n2421 = ~new_n2395 & ~new_n2414;
  assign new_n2422 = new_n2420 & ~new_n2421;
  assign new_n2423 = ~new_n2420 & new_n2421;
  assign new_n2424 = ~new_n2422 & ~new_n2423;
  assign new_n2425 = new_n2400 & new_n2424;
  assign new_n2426 = new_n2398 & new_n2402;
  assign new_n2427 = ~new_n2425 & new_n2426;
  assign new_n2428 = new_n2419 & ~new_n2427;
  assign new_n2429 = ~A895 & ~A896;
  assign new_n2430 = A898 & A899;
  assign new_n2431 = ~A897 & A900;
  assign new_n2432 = new_n2430 & new_n2431;
  assign new_n2433 = A895 & A896;
  assign new_n2434 = ~A897 & ~new_n2433;
  assign new_n2435 = ~A898 & ~A899;
  assign new_n2436 = ~new_n2430 & ~new_n2435;
  assign new_n2437 = A900 & ~new_n2436;
  assign new_n2438 = ~A900 & ~new_n2430;
  assign new_n2439 = ~new_n2434 & ~new_n2438;
  assign new_n2440 = ~new_n2437 & new_n2439;
  assign new_n2441 = ~new_n2432 & ~new_n2440;
  assign new_n2442 = ~new_n2429 & ~new_n2441;
  assign new_n2443 = A897 & A900;
  assign new_n2444 = ~new_n2430 & ~new_n2433;
  assign new_n2445 = new_n2443 & ~new_n2444;
  assign new_n2446 = A899 & new_n2433;
  assign new_n2447 = new_n2445 & ~new_n2446;
  assign new_n2448 = new_n2429 & new_n2435;
  assign new_n2449 = ~new_n2443 & new_n2448;
  assign new_n2450 = A897 & ~A900;
  assign new_n2451 = new_n2433 & ~new_n2435;
  assign new_n2452 = new_n2450 & new_n2451;
  assign new_n2453 = ~new_n2449 & ~new_n2452;
  assign new_n2454 = ~new_n2447 & new_n2453;
  assign new_n2455 = ~new_n2442 & new_n2454;
  assign new_n2456 = ~new_n2429 & ~new_n2433;
  assign new_n2457 = ~new_n2431 & ~new_n2450;
  assign new_n2458 = new_n2456 & ~new_n2457;
  assign new_n2459 = ~new_n2456 & new_n2457;
  assign new_n2460 = ~new_n2458 & ~new_n2459;
  assign new_n2461 = new_n2436 & new_n2460;
  assign new_n2462 = new_n2434 & new_n2438;
  assign new_n2463 = ~new_n2461 & new_n2462;
  assign new_n2464 = new_n2455 & ~new_n2463;
  assign new_n2465 = ~new_n2428 & ~new_n2464;
  assign new_n2466 = ~new_n2436 & ~new_n2460;
  assign new_n2467 = ~new_n2461 & ~new_n2466;
  assign new_n2468 = ~new_n2400 & ~new_n2424;
  assign new_n2469 = ~new_n2425 & ~new_n2468;
  assign new_n2470 = new_n2467 & new_n2469;
  assign new_n2471 = new_n2428 & new_n2464;
  assign new_n2472 = ~new_n2465 & ~new_n2471;
  assign new_n2473 = ~new_n2470 & new_n2472;
  assign new_n2474 = ~new_n2465 & ~new_n2473;
  assign new_n2475 = ~new_n2429 & ~new_n2455;
  assign new_n2476 = ~new_n2445 & ~new_n2475;
  assign new_n2477 = ~new_n2393 & ~new_n2419;
  assign new_n2478 = ~new_n2409 & ~new_n2477;
  assign new_n2479 = new_n2476 & new_n2478;
  assign new_n2480 = ~new_n2476 & ~new_n2478;
  assign new_n2481 = ~new_n2479 & ~new_n2480;
  assign new_n2482 = ~new_n2474 & new_n2481;
  assign new_n2483 = new_n2474 & ~new_n2481;
  assign new_n2484 = ~new_n2482 & ~new_n2483;
  assign new_n2485 = new_n2358 & ~new_n2386;
  assign new_n2486 = ~new_n2387 & ~new_n2485;
  assign new_n2487 = new_n2470 & ~new_n2472;
  assign new_n2488 = ~new_n2473 & ~new_n2487;
  assign new_n2489 = ~new_n2486 & ~new_n2488;
  assign new_n2490 = ~new_n2467 & ~new_n2469;
  assign new_n2491 = ~new_n2470 & ~new_n2490;
  assign new_n2492 = new_n2377 & ~new_n2378;
  assign new_n2493 = ~new_n2379 & ~new_n2492;
  assign new_n2494 = new_n2491 & ~new_n2493;
  assign new_n2495 = new_n2486 & new_n2488;
  assign new_n2496 = ~new_n2489 & ~new_n2495;
  assign new_n2497 = new_n2494 & new_n2496;
  assign new_n2498 = ~new_n2489 & ~new_n2497;
  assign new_n2499 = new_n2484 & new_n2498;
  assign new_n2500 = ~new_n2484 & ~new_n2498;
  assign new_n2501 = ~new_n2499 & ~new_n2500;
  assign new_n2502 = ~new_n2392 & new_n2501;
  assign new_n2503 = new_n2392 & ~new_n2501;
  assign new_n2504 = ~new_n2502 & ~new_n2503;
  assign new_n2505 = ~A937 & ~A938;
  assign new_n2506 = A937 & A938;
  assign new_n2507 = ~A939 & ~new_n2506;
  assign new_n2508 = ~new_n2505 & ~new_n2507;
  assign new_n2509 = A939 & new_n2506;
  assign new_n2510 = ~A940 & ~new_n2509;
  assign new_n2511 = new_n2508 & ~new_n2510;
  assign new_n2512 = A941 & new_n2511;
  assign new_n2513 = A939 & A940;
  assign new_n2514 = new_n2506 & new_n2513;
  assign new_n2515 = ~new_n2512 & ~new_n2514;
  assign new_n2516 = ~A942 & ~new_n2515;
  assign new_n2517 = new_n2505 & ~new_n2513;
  assign new_n2518 = A941 & A942;
  assign new_n2519 = ~new_n2509 & new_n2518;
  assign new_n2520 = ~new_n2517 & new_n2519;
  assign new_n2521 = A940 & ~new_n2520;
  assign new_n2522 = new_n2508 & new_n2518;
  assign new_n2523 = ~A941 & ~A942;
  assign new_n2524 = ~new_n2505 & ~new_n2523;
  assign new_n2525 = new_n2507 & ~new_n2518;
  assign new_n2526 = ~new_n2524 & new_n2525;
  assign new_n2527 = ~A940 & ~new_n2522;
  assign new_n2528 = ~new_n2526 & new_n2527;
  assign new_n2529 = ~new_n2521 & ~new_n2528;
  assign new_n2530 = ~A941 & A942;
  assign new_n2531 = new_n2511 & new_n2530;
  assign new_n2532 = ~new_n2516 & ~new_n2531;
  assign new_n2533 = ~new_n2529 & new_n2532;
  assign new_n2534 = new_n2517 & new_n2523;
  assign new_n2535 = new_n2533 & ~new_n2534;
  assign new_n2536 = A934 & A935;
  assign new_n2537 = ~A934 & ~A935;
  assign new_n2538 = ~new_n2536 & ~new_n2537;
  assign new_n2539 = A931 & A932;
  assign new_n2540 = ~A931 & ~A932;
  assign new_n2541 = ~new_n2539 & ~new_n2540;
  assign new_n2542 = ~A933 & A936;
  assign new_n2543 = A933 & ~A936;
  assign new_n2544 = ~new_n2542 & ~new_n2543;
  assign new_n2545 = new_n2541 & ~new_n2544;
  assign new_n2546 = ~new_n2541 & new_n2544;
  assign new_n2547 = ~new_n2545 & ~new_n2546;
  assign new_n2548 = new_n2538 & new_n2547;
  assign new_n2549 = ~new_n2538 & ~new_n2547;
  assign new_n2550 = ~new_n2548 & ~new_n2549;
  assign new_n2551 = A939 & ~A942;
  assign new_n2552 = ~A939 & A942;
  assign new_n2553 = ~new_n2551 & ~new_n2552;
  assign new_n2554 = ~new_n2505 & ~new_n2506;
  assign new_n2555 = ~A940 & ~A941;
  assign new_n2556 = A940 & A941;
  assign new_n2557 = ~new_n2555 & ~new_n2556;
  assign new_n2558 = new_n2554 & ~new_n2557;
  assign new_n2559 = ~new_n2554 & new_n2557;
  assign new_n2560 = ~new_n2558 & ~new_n2559;
  assign new_n2561 = new_n2553 & new_n2560;
  assign new_n2562 = ~new_n2553 & ~new_n2560;
  assign new_n2563 = ~new_n2561 & ~new_n2562;
  assign new_n2564 = new_n2550 & new_n2563;
  assign new_n2565 = new_n2536 & new_n2542;
  assign new_n2566 = ~A933 & ~new_n2539;
  assign new_n2567 = A936 & ~new_n2538;
  assign new_n2568 = ~A936 & ~new_n2536;
  assign new_n2569 = ~new_n2566 & ~new_n2568;
  assign new_n2570 = ~new_n2567 & new_n2569;
  assign new_n2571 = ~new_n2565 & ~new_n2570;
  assign new_n2572 = ~new_n2540 & ~new_n2571;
  assign new_n2573 = A933 & A936;
  assign new_n2574 = ~new_n2536 & ~new_n2539;
  assign new_n2575 = new_n2573 & ~new_n2574;
  assign new_n2576 = A935 & new_n2539;
  assign new_n2577 = new_n2575 & ~new_n2576;
  assign new_n2578 = new_n2537 & new_n2540;
  assign new_n2579 = ~new_n2573 & new_n2578;
  assign new_n2580 = ~new_n2537 & new_n2539;
  assign new_n2581 = new_n2543 & new_n2580;
  assign new_n2582 = ~new_n2579 & ~new_n2581;
  assign new_n2583 = ~new_n2577 & new_n2582;
  assign new_n2584 = ~new_n2572 & new_n2583;
  assign new_n2585 = new_n2566 & new_n2568;
  assign new_n2586 = ~new_n2548 & new_n2585;
  assign new_n2587 = new_n2584 & ~new_n2586;
  assign new_n2588 = ~new_n2564 & ~new_n2587;
  assign new_n2589 = new_n2564 & new_n2587;
  assign new_n2590 = ~new_n2588 & ~new_n2589;
  assign new_n2591 = ~new_n2535 & new_n2590;
  assign new_n2592 = new_n2535 & ~new_n2590;
  assign new_n2593 = ~new_n2591 & ~new_n2592;
  assign new_n2594 = A922 & A923;
  assign new_n2595 = ~A922 & ~A923;
  assign new_n2596 = ~new_n2594 & ~new_n2595;
  assign new_n2597 = A919 & A920;
  assign new_n2598 = ~A919 & ~A920;
  assign new_n2599 = ~new_n2597 & ~new_n2598;
  assign new_n2600 = ~A921 & A924;
  assign new_n2601 = A921 & ~A924;
  assign new_n2602 = ~new_n2600 & ~new_n2601;
  assign new_n2603 = new_n2599 & ~new_n2602;
  assign new_n2604 = ~new_n2599 & new_n2602;
  assign new_n2605 = ~new_n2603 & ~new_n2604;
  assign new_n2606 = new_n2596 & new_n2605;
  assign new_n2607 = ~new_n2596 & ~new_n2605;
  assign new_n2608 = ~new_n2606 & ~new_n2607;
  assign new_n2609 = A928 & A929;
  assign new_n2610 = ~A928 & ~A929;
  assign new_n2611 = ~new_n2609 & ~new_n2610;
  assign new_n2612 = A925 & A926;
  assign new_n2613 = ~A925 & ~A926;
  assign new_n2614 = ~new_n2612 & ~new_n2613;
  assign new_n2615 = ~A927 & A930;
  assign new_n2616 = A927 & ~A930;
  assign new_n2617 = ~new_n2615 & ~new_n2616;
  assign new_n2618 = new_n2614 & ~new_n2617;
  assign new_n2619 = ~new_n2614 & new_n2617;
  assign new_n2620 = ~new_n2618 & ~new_n2619;
  assign new_n2621 = new_n2611 & new_n2620;
  assign new_n2622 = ~new_n2611 & ~new_n2620;
  assign new_n2623 = ~new_n2621 & ~new_n2622;
  assign new_n2624 = new_n2608 & new_n2623;
  assign new_n2625 = new_n2609 & new_n2615;
  assign new_n2626 = A930 & ~new_n2611;
  assign new_n2627 = ~A927 & ~new_n2612;
  assign new_n2628 = ~A930 & ~new_n2609;
  assign new_n2629 = ~new_n2627 & ~new_n2628;
  assign new_n2630 = ~new_n2626 & new_n2629;
  assign new_n2631 = ~new_n2625 & ~new_n2630;
  assign new_n2632 = ~new_n2613 & ~new_n2631;
  assign new_n2633 = A927 & A930;
  assign new_n2634 = ~new_n2609 & ~new_n2612;
  assign new_n2635 = new_n2633 & ~new_n2634;
  assign new_n2636 = A929 & new_n2612;
  assign new_n2637 = new_n2635 & ~new_n2636;
  assign new_n2638 = new_n2610 & new_n2613;
  assign new_n2639 = ~new_n2633 & new_n2638;
  assign new_n2640 = ~new_n2610 & new_n2612;
  assign new_n2641 = new_n2616 & new_n2640;
  assign new_n2642 = ~new_n2639 & ~new_n2641;
  assign new_n2643 = ~new_n2637 & new_n2642;
  assign new_n2644 = ~new_n2632 & new_n2643;
  assign new_n2645 = new_n2627 & new_n2628;
  assign new_n2646 = ~new_n2621 & new_n2645;
  assign new_n2647 = new_n2644 & ~new_n2646;
  assign new_n2648 = new_n2594 & new_n2600;
  assign new_n2649 = ~A921 & ~new_n2597;
  assign new_n2650 = A924 & ~new_n2596;
  assign new_n2651 = ~A924 & ~new_n2594;
  assign new_n2652 = ~new_n2649 & ~new_n2651;
  assign new_n2653 = ~new_n2650 & new_n2652;
  assign new_n2654 = ~new_n2648 & ~new_n2653;
  assign new_n2655 = ~new_n2598 & ~new_n2654;
  assign new_n2656 = A921 & A924;
  assign new_n2657 = ~new_n2594 & ~new_n2597;
  assign new_n2658 = new_n2656 & ~new_n2657;
  assign new_n2659 = A923 & new_n2597;
  assign new_n2660 = new_n2658 & ~new_n2659;
  assign new_n2661 = new_n2595 & new_n2598;
  assign new_n2662 = ~new_n2656 & new_n2661;
  assign new_n2663 = ~new_n2595 & new_n2597;
  assign new_n2664 = new_n2601 & new_n2663;
  assign new_n2665 = ~new_n2662 & ~new_n2664;
  assign new_n2666 = ~new_n2660 & new_n2665;
  assign new_n2667 = ~new_n2655 & new_n2666;
  assign new_n2668 = new_n2649 & new_n2651;
  assign new_n2669 = ~new_n2606 & new_n2668;
  assign new_n2670 = new_n2667 & ~new_n2669;
  assign new_n2671 = ~new_n2647 & ~new_n2670;
  assign new_n2672 = new_n2647 & new_n2670;
  assign new_n2673 = ~new_n2671 & ~new_n2672;
  assign new_n2674 = ~new_n2624 & new_n2673;
  assign new_n2675 = new_n2624 & ~new_n2673;
  assign new_n2676 = ~new_n2674 & ~new_n2675;
  assign new_n2677 = ~new_n2593 & ~new_n2676;
  assign new_n2678 = ~new_n2608 & ~new_n2623;
  assign new_n2679 = ~new_n2624 & ~new_n2678;
  assign new_n2680 = ~new_n2550 & ~new_n2563;
  assign new_n2681 = ~new_n2564 & ~new_n2680;
  assign new_n2682 = new_n2679 & new_n2681;
  assign new_n2683 = new_n2593 & ~new_n2673;
  assign new_n2684 = new_n2682 & ~new_n2683;
  assign new_n2685 = ~new_n2677 & ~new_n2684;
  assign new_n2686 = ~new_n2588 & ~new_n2591;
  assign new_n2687 = ~new_n2510 & ~new_n2533;
  assign new_n2688 = ~new_n2522 & ~new_n2687;
  assign new_n2689 = ~new_n2540 & ~new_n2584;
  assign new_n2690 = ~new_n2575 & ~new_n2689;
  assign new_n2691 = new_n2688 & new_n2690;
  assign new_n2692 = ~new_n2688 & ~new_n2690;
  assign new_n2693 = ~new_n2691 & ~new_n2692;
  assign new_n2694 = ~new_n2686 & new_n2693;
  assign new_n2695 = new_n2686 & ~new_n2693;
  assign new_n2696 = ~new_n2694 & ~new_n2695;
  assign new_n2697 = ~new_n2671 & ~new_n2674;
  assign new_n2698 = ~new_n2598 & ~new_n2667;
  assign new_n2699 = ~new_n2658 & ~new_n2698;
  assign new_n2700 = ~new_n2613 & ~new_n2644;
  assign new_n2701 = ~new_n2635 & ~new_n2700;
  assign new_n2702 = new_n2699 & new_n2701;
  assign new_n2703 = ~new_n2699 & ~new_n2701;
  assign new_n2704 = ~new_n2702 & ~new_n2703;
  assign new_n2705 = ~new_n2697 & new_n2704;
  assign new_n2706 = new_n2697 & ~new_n2704;
  assign new_n2707 = ~new_n2705 & ~new_n2706;
  assign new_n2708 = ~new_n2696 & ~new_n2707;
  assign new_n2709 = new_n2696 & new_n2707;
  assign new_n2710 = ~new_n2708 & ~new_n2709;
  assign new_n2711 = ~new_n2685 & new_n2710;
  assign new_n2712 = new_n2685 & ~new_n2710;
  assign new_n2713 = ~new_n2711 & ~new_n2712;
  assign new_n2714 = ~new_n2491 & new_n2493;
  assign new_n2715 = ~new_n2494 & ~new_n2714;
  assign new_n2716 = ~new_n2679 & ~new_n2681;
  assign new_n2717 = ~new_n2682 & ~new_n2716;
  assign new_n2718 = new_n2715 & new_n2717;
  assign new_n2719 = ~new_n2494 & ~new_n2718;
  assign new_n2720 = ~new_n2496 & new_n2719;
  assign new_n2721 = new_n2496 & ~new_n2719;
  assign new_n2722 = ~new_n2720 & ~new_n2721;
  assign new_n2723 = ~new_n2593 & new_n2673;
  assign new_n2724 = ~new_n2683 & ~new_n2723;
  assign new_n2725 = ~new_n2624 & ~new_n2682;
  assign new_n2726 = ~new_n2724 & new_n2725;
  assign new_n2727 = new_n2724 & ~new_n2725;
  assign new_n2728 = ~new_n2726 & ~new_n2727;
  assign new_n2729 = new_n2722 & ~new_n2728;
  assign new_n2730 = ~new_n2497 & ~new_n2720;
  assign new_n2731 = ~new_n2729 & new_n2730;
  assign new_n2732 = ~new_n2713 & ~new_n2731;
  assign new_n2733 = new_n2713 & new_n2731;
  assign new_n2734 = ~new_n2732 & ~new_n2733;
  assign new_n2735 = new_n2504 & new_n2734;
  assign new_n2736 = ~new_n2504 & ~new_n2734;
  assign new_n2737 = ~new_n2735 & ~new_n2736;
  assign new_n2738 = ~A865 & ~A866;
  assign new_n2739 = A865 & A866;
  assign new_n2740 = ~A867 & ~new_n2739;
  assign new_n2741 = ~new_n2738 & ~new_n2740;
  assign new_n2742 = A867 & new_n2739;
  assign new_n2743 = ~A868 & ~new_n2742;
  assign new_n2744 = new_n2741 & ~new_n2743;
  assign new_n2745 = A869 & new_n2744;
  assign new_n2746 = A867 & A868;
  assign new_n2747 = new_n2739 & new_n2746;
  assign new_n2748 = ~new_n2745 & ~new_n2747;
  assign new_n2749 = ~A870 & ~new_n2748;
  assign new_n2750 = A869 & A870;
  assign new_n2751 = new_n2741 & new_n2750;
  assign new_n2752 = ~A869 & ~A870;
  assign new_n2753 = ~new_n2738 & ~new_n2752;
  assign new_n2754 = new_n2740 & ~new_n2750;
  assign new_n2755 = ~new_n2753 & new_n2754;
  assign new_n2756 = ~new_n2751 & ~new_n2755;
  assign new_n2757 = ~A868 & ~new_n2756;
  assign new_n2758 = new_n2738 & ~new_n2746;
  assign new_n2759 = A868 & new_n2750;
  assign new_n2760 = ~new_n2742 & new_n2759;
  assign new_n2761 = ~new_n2758 & new_n2760;
  assign new_n2762 = ~A869 & A870;
  assign new_n2763 = new_n2744 & new_n2762;
  assign new_n2764 = ~new_n2761 & ~new_n2763;
  assign new_n2765 = ~new_n2757 & new_n2764;
  assign new_n2766 = ~new_n2749 & new_n2765;
  assign new_n2767 = new_n2752 & new_n2758;
  assign new_n2768 = new_n2766 & ~new_n2767;
  assign new_n2769 = A862 & A863;
  assign new_n2770 = ~A862 & ~A863;
  assign new_n2771 = ~new_n2769 & ~new_n2770;
  assign new_n2772 = A859 & A860;
  assign new_n2773 = ~A859 & ~A860;
  assign new_n2774 = ~new_n2772 & ~new_n2773;
  assign new_n2775 = ~A861 & A864;
  assign new_n2776 = A861 & ~A864;
  assign new_n2777 = ~new_n2775 & ~new_n2776;
  assign new_n2778 = new_n2774 & ~new_n2777;
  assign new_n2779 = ~new_n2774 & new_n2777;
  assign new_n2780 = ~new_n2778 & ~new_n2779;
  assign new_n2781 = new_n2771 & new_n2780;
  assign new_n2782 = ~new_n2771 & ~new_n2780;
  assign new_n2783 = ~new_n2781 & ~new_n2782;
  assign new_n2784 = A867 & ~A870;
  assign new_n2785 = ~A867 & A870;
  assign new_n2786 = ~new_n2784 & ~new_n2785;
  assign new_n2787 = ~new_n2738 & ~new_n2739;
  assign new_n2788 = ~A868 & ~A869;
  assign new_n2789 = A868 & A869;
  assign new_n2790 = ~new_n2788 & ~new_n2789;
  assign new_n2791 = new_n2787 & ~new_n2790;
  assign new_n2792 = ~new_n2787 & new_n2790;
  assign new_n2793 = ~new_n2791 & ~new_n2792;
  assign new_n2794 = new_n2786 & new_n2793;
  assign new_n2795 = ~new_n2786 & ~new_n2793;
  assign new_n2796 = ~new_n2794 & ~new_n2795;
  assign new_n2797 = new_n2783 & new_n2796;
  assign new_n2798 = new_n2769 & new_n2775;
  assign new_n2799 = ~A861 & ~new_n2772;
  assign new_n2800 = A864 & ~new_n2771;
  assign new_n2801 = ~A864 & ~new_n2769;
  assign new_n2802 = ~new_n2799 & ~new_n2801;
  assign new_n2803 = ~new_n2800 & new_n2802;
  assign new_n2804 = ~new_n2798 & ~new_n2803;
  assign new_n2805 = ~new_n2773 & ~new_n2804;
  assign new_n2806 = ~new_n2769 & ~new_n2772;
  assign new_n2807 = A861 & A864;
  assign new_n2808 = ~new_n2806 & new_n2807;
  assign new_n2809 = A863 & new_n2772;
  assign new_n2810 = new_n2808 & ~new_n2809;
  assign new_n2811 = new_n2770 & new_n2773;
  assign new_n2812 = ~new_n2807 & new_n2811;
  assign new_n2813 = ~new_n2770 & new_n2772;
  assign new_n2814 = new_n2776 & new_n2813;
  assign new_n2815 = ~new_n2812 & ~new_n2814;
  assign new_n2816 = ~new_n2810 & new_n2815;
  assign new_n2817 = ~new_n2805 & new_n2816;
  assign new_n2818 = new_n2799 & new_n2801;
  assign new_n2819 = ~new_n2781 & new_n2818;
  assign new_n2820 = new_n2817 & ~new_n2819;
  assign new_n2821 = ~new_n2797 & ~new_n2820;
  assign new_n2822 = new_n2797 & new_n2820;
  assign new_n2823 = ~new_n2821 & ~new_n2822;
  assign new_n2824 = ~new_n2768 & new_n2823;
  assign new_n2825 = new_n2768 & ~new_n2823;
  assign new_n2826 = ~new_n2824 & ~new_n2825;
  assign new_n2827 = ~A848 & ~A849;
  assign new_n2828 = A848 & A849;
  assign new_n2829 = ~new_n2827 & ~new_n2828;
  assign new_n2830 = A847 & ~new_n2829;
  assign new_n2831 = ~A847 & new_n2829;
  assign new_n2832 = ~new_n2830 & ~new_n2831;
  assign new_n2833 = A852 & ~new_n2832;
  assign new_n2834 = ~A850 & ~A851;
  assign new_n2835 = ~A852 & new_n2832;
  assign new_n2836 = ~new_n2833 & ~new_n2835;
  assign new_n2837 = A850 & A851;
  assign new_n2838 = ~new_n2834 & ~new_n2837;
  assign new_n2839 = ~new_n2836 & new_n2838;
  assign new_n2840 = ~new_n2834 & ~new_n2839;
  assign new_n2841 = ~new_n2833 & ~new_n2840;
  assign new_n2842 = new_n2833 & new_n2837;
  assign new_n2843 = ~new_n2841 & ~new_n2842;
  assign new_n2844 = ~new_n2827 & ~new_n2831;
  assign new_n2845 = new_n2843 & ~new_n2844;
  assign new_n2846 = ~new_n2843 & new_n2844;
  assign new_n2847 = ~new_n2845 & ~new_n2846;
  assign new_n2848 = new_n2836 & ~new_n2838;
  assign new_n2849 = ~new_n2839 & ~new_n2848;
  assign new_n2850 = A856 & A857;
  assign new_n2851 = ~A856 & ~A857;
  assign new_n2852 = ~new_n2850 & ~new_n2851;
  assign new_n2853 = A853 & A854;
  assign new_n2854 = ~A853 & ~A854;
  assign new_n2855 = ~new_n2853 & ~new_n2854;
  assign new_n2856 = ~A855 & A858;
  assign new_n2857 = A855 & ~A858;
  assign new_n2858 = ~new_n2856 & ~new_n2857;
  assign new_n2859 = new_n2855 & ~new_n2858;
  assign new_n2860 = ~new_n2855 & new_n2858;
  assign new_n2861 = ~new_n2859 & ~new_n2860;
  assign new_n2862 = new_n2852 & new_n2861;
  assign new_n2863 = ~new_n2852 & ~new_n2861;
  assign new_n2864 = ~new_n2862 & ~new_n2863;
  assign new_n2865 = ~new_n2849 & new_n2864;
  assign new_n2866 = new_n2850 & new_n2856;
  assign new_n2867 = ~A855 & ~new_n2853;
  assign new_n2868 = A858 & ~new_n2852;
  assign new_n2869 = ~A858 & ~new_n2850;
  assign new_n2870 = ~new_n2867 & ~new_n2869;
  assign new_n2871 = ~new_n2868 & new_n2870;
  assign new_n2872 = ~new_n2866 & ~new_n2871;
  assign new_n2873 = ~new_n2854 & ~new_n2872;
  assign new_n2874 = ~new_n2850 & ~new_n2853;
  assign new_n2875 = A855 & A858;
  assign new_n2876 = ~new_n2874 & new_n2875;
  assign new_n2877 = A857 & new_n2853;
  assign new_n2878 = new_n2876 & ~new_n2877;
  assign new_n2879 = new_n2851 & new_n2854;
  assign new_n2880 = ~new_n2875 & new_n2879;
  assign new_n2881 = ~new_n2851 & new_n2853;
  assign new_n2882 = new_n2857 & new_n2881;
  assign new_n2883 = ~new_n2880 & ~new_n2882;
  assign new_n2884 = ~new_n2878 & new_n2883;
  assign new_n2885 = ~new_n2873 & new_n2884;
  assign new_n2886 = new_n2867 & new_n2869;
  assign new_n2887 = ~new_n2862 & new_n2886;
  assign new_n2888 = new_n2885 & ~new_n2887;
  assign new_n2889 = new_n2865 & new_n2888;
  assign new_n2890 = ~new_n2865 & ~new_n2888;
  assign new_n2891 = ~new_n2889 & ~new_n2890;
  assign new_n2892 = ~new_n2847 & new_n2891;
  assign new_n2893 = new_n2847 & ~new_n2891;
  assign new_n2894 = ~new_n2892 & ~new_n2893;
  assign new_n2895 = new_n2826 & ~new_n2894;
  assign new_n2896 = ~new_n2826 & new_n2894;
  assign new_n2897 = ~new_n2895 & ~new_n2896;
  assign new_n2898 = ~A890 & ~A891;
  assign new_n2899 = A890 & A891;
  assign new_n2900 = ~new_n2898 & ~new_n2899;
  assign new_n2901 = ~A889 & new_n2900;
  assign new_n2902 = ~new_n2898 & ~new_n2901;
  assign new_n2903 = ~A892 & ~A894;
  assign new_n2904 = A892 & A894;
  assign new_n2905 = ~new_n2903 & ~new_n2904;
  assign new_n2906 = ~A893 & new_n2905;
  assign new_n2907 = ~new_n2903 & ~new_n2906;
  assign new_n2908 = ~new_n2902 & ~new_n2907;
  assign new_n2909 = new_n2902 & new_n2907;
  assign new_n2910 = ~new_n2908 & ~new_n2909;
  assign new_n2911 = ~A887 & ~A888;
  assign new_n2912 = A883 & A884;
  assign new_n2913 = A885 & A886;
  assign new_n2914 = ~new_n2912 & new_n2913;
  assign new_n2915 = ~A885 & ~A886;
  assign new_n2916 = ~new_n2913 & ~new_n2915;
  assign new_n2917 = ~A883 & ~A884;
  assign new_n2918 = ~new_n2912 & ~new_n2917;
  assign new_n2919 = ~new_n2916 & new_n2918;
  assign new_n2920 = ~new_n2913 & ~new_n2917;
  assign new_n2921 = ~new_n2919 & new_n2920;
  assign new_n2922 = ~new_n2914 & ~new_n2921;
  assign new_n2923 = new_n2911 & new_n2922;
  assign new_n2924 = A887 & A888;
  assign new_n2925 = ~new_n2912 & ~new_n2919;
  assign new_n2926 = ~new_n2911 & ~new_n2915;
  assign new_n2927 = ~new_n2925 & new_n2926;
  assign new_n2928 = ~new_n2924 & new_n2927;
  assign new_n2929 = new_n2912 & new_n2923;
  assign new_n2930 = ~new_n2922 & new_n2924;
  assign new_n2931 = ~new_n2929 & ~new_n2930;
  assign new_n2932 = new_n2915 & new_n2917;
  assign new_n2933 = ~new_n2924 & new_n2932;
  assign new_n2934 = ~new_n2923 & ~new_n2933;
  assign new_n2935 = ~new_n2928 & new_n2934;
  assign new_n2936 = new_n2931 & new_n2935;
  assign new_n2937 = ~new_n2910 & new_n2936;
  assign new_n2938 = new_n2910 & ~new_n2936;
  assign new_n2939 = ~new_n2937 & ~new_n2938;
  assign new_n2940 = A893 & ~new_n2905;
  assign new_n2941 = ~new_n2906 & ~new_n2940;
  assign new_n2942 = A889 & ~new_n2900;
  assign new_n2943 = ~new_n2901 & ~new_n2942;
  assign new_n2944 = new_n2941 & new_n2943;
  assign new_n2945 = ~new_n2941 & ~new_n2943;
  assign new_n2946 = ~new_n2944 & ~new_n2945;
  assign new_n2947 = ~new_n2911 & ~new_n2924;
  assign new_n2948 = new_n2916 & ~new_n2918;
  assign new_n2949 = ~new_n2919 & ~new_n2948;
  assign new_n2950 = new_n2947 & ~new_n2949;
  assign new_n2951 = ~new_n2947 & new_n2949;
  assign new_n2952 = ~new_n2950 & ~new_n2951;
  assign new_n2953 = new_n2946 & ~new_n2952;
  assign new_n2954 = ~new_n2944 & ~new_n2953;
  assign new_n2955 = ~new_n2939 & ~new_n2954;
  assign new_n2956 = new_n2939 & new_n2954;
  assign new_n2957 = ~new_n2955 & ~new_n2956;
  assign new_n2958 = A881 & A882;
  assign new_n2959 = ~A877 & ~A878;
  assign new_n2960 = ~A879 & ~A880;
  assign new_n2961 = new_n2959 & new_n2960;
  assign new_n2962 = A877 & A878;
  assign new_n2963 = A879 & A880;
  assign new_n2964 = ~new_n2962 & ~new_n2963;
  assign new_n2965 = ~A881 & ~A882;
  assign new_n2966 = ~new_n2959 & ~new_n2960;
  assign new_n2967 = ~new_n2964 & ~new_n2965;
  assign new_n2968 = new_n2966 & new_n2967;
  assign new_n2969 = ~new_n2961 & ~new_n2968;
  assign new_n2970 = ~new_n2958 & ~new_n2969;
  assign new_n2971 = new_n2964 & ~new_n2966;
  assign new_n2972 = new_n2962 & new_n2963;
  assign new_n2973 = ~new_n2971 & ~new_n2972;
  assign new_n2974 = new_n2965 & ~new_n2973;
  assign new_n2975 = ~new_n2965 & ~new_n2973;
  assign new_n2976 = ~new_n2958 & ~new_n2972;
  assign new_n2977 = ~new_n2975 & ~new_n2976;
  assign new_n2978 = ~new_n2970 & ~new_n2974;
  assign new_n2979 = ~new_n2977 & new_n2978;
  assign new_n2980 = ~A872 & ~A873;
  assign new_n2981 = A872 & A873;
  assign new_n2982 = ~new_n2980 & ~new_n2981;
  assign new_n2983 = A871 & ~new_n2982;
  assign new_n2984 = A874 & A875;
  assign new_n2985 = ~A871 & new_n2982;
  assign new_n2986 = ~new_n2980 & ~new_n2985;
  assign new_n2987 = new_n2984 & new_n2986;
  assign new_n2988 = ~new_n2983 & new_n2987;
  assign new_n2989 = ~new_n2983 & ~new_n2985;
  assign new_n2990 = A876 & ~new_n2989;
  assign new_n2991 = ~new_n2984 & ~new_n2986;
  assign new_n2992 = ~new_n2987 & new_n2990;
  assign new_n2993 = ~new_n2991 & new_n2992;
  assign new_n2994 = ~A876 & new_n2989;
  assign new_n2995 = ~new_n2990 & ~new_n2994;
  assign new_n2996 = ~A874 & ~A875;
  assign new_n2997 = new_n2986 & ~new_n2996;
  assign new_n2998 = new_n2995 & new_n2997;
  assign new_n2999 = ~new_n2993 & ~new_n2998;
  assign new_n3000 = ~new_n2984 & ~new_n2996;
  assign new_n3001 = new_n2995 & new_n3000;
  assign new_n3002 = ~new_n2990 & new_n2991;
  assign new_n3003 = ~new_n3001 & new_n3002;
  assign new_n3004 = ~new_n2988 & new_n2999;
  assign new_n3005 = ~new_n3003 & new_n3004;
  assign new_n3006 = ~new_n2979 & ~new_n3005;
  assign new_n3007 = new_n2979 & new_n3005;
  assign new_n3008 = ~new_n3006 & ~new_n3007;
  assign new_n3009 = ~new_n2995 & ~new_n3000;
  assign new_n3010 = ~new_n3001 & ~new_n3009;
  assign new_n3011 = ~new_n2958 & ~new_n2965;
  assign new_n3012 = ~new_n2960 & ~new_n2963;
  assign new_n3013 = ~new_n3011 & new_n3012;
  assign new_n3014 = new_n3011 & ~new_n3012;
  assign new_n3015 = ~new_n3013 & ~new_n3014;
  assign new_n3016 = ~new_n2959 & ~new_n2962;
  assign new_n3017 = ~new_n3015 & new_n3016;
  assign new_n3018 = new_n3015 & ~new_n3016;
  assign new_n3019 = ~new_n3017 & ~new_n3018;
  assign new_n3020 = ~new_n3010 & ~new_n3019;
  assign new_n3021 = ~new_n2946 & new_n2952;
  assign new_n3022 = ~new_n2953 & ~new_n3021;
  assign new_n3023 = new_n3010 & new_n3019;
  assign new_n3024 = ~new_n3020 & ~new_n3023;
  assign new_n3025 = new_n3022 & new_n3024;
  assign new_n3026 = ~new_n3020 & ~new_n3025;
  assign new_n3027 = new_n3008 & new_n3026;
  assign new_n3028 = ~new_n3008 & ~new_n3026;
  assign new_n3029 = ~new_n3027 & ~new_n3028;
  assign new_n3030 = ~new_n2957 & new_n3029;
  assign new_n3031 = new_n2957 & ~new_n3029;
  assign new_n3032 = ~new_n3030 & ~new_n3031;
  assign new_n3033 = ~new_n2897 & new_n3032;
  assign new_n3034 = new_n2897 & ~new_n3032;
  assign new_n3035 = ~new_n3033 & ~new_n3034;
  assign new_n3036 = new_n2849 & ~new_n2864;
  assign new_n3037 = ~new_n2865 & ~new_n3036;
  assign new_n3038 = ~new_n2783 & ~new_n2796;
  assign new_n3039 = ~new_n2797 & ~new_n3038;
  assign new_n3040 = new_n3037 & new_n3039;
  assign new_n3041 = ~new_n3022 & ~new_n3024;
  assign new_n3042 = ~new_n3025 & ~new_n3041;
  assign new_n3043 = ~new_n3037 & ~new_n3039;
  assign new_n3044 = ~new_n3040 & ~new_n3043;
  assign new_n3045 = ~new_n3042 & new_n3044;
  assign new_n3046 = ~new_n3040 & ~new_n3045;
  assign new_n3047 = ~new_n3035 & new_n3046;
  assign new_n3048 = new_n3035 & ~new_n3046;
  assign new_n3049 = ~new_n3047 & ~new_n3048;
  assign new_n3050 = ~new_n2722 & new_n2728;
  assign new_n3051 = ~new_n2729 & ~new_n3050;
  assign new_n3052 = ~new_n3049 & ~new_n3051;
  assign new_n3053 = new_n3049 & new_n3051;
  assign new_n3054 = ~new_n3052 & ~new_n3053;
  assign new_n3055 = new_n3042 & ~new_n3044;
  assign new_n3056 = ~new_n3045 & ~new_n3055;
  assign new_n3057 = ~new_n2715 & ~new_n2717;
  assign new_n3058 = ~new_n2718 & ~new_n3057;
  assign new_n3059 = new_n3056 & new_n3058;
  assign new_n3060 = new_n3054 & new_n3059;
  assign new_n3061 = ~new_n3052 & ~new_n3060;
  assign new_n3062 = new_n2897 & ~new_n3040;
  assign new_n3063 = ~new_n3033 & ~new_n3062;
  assign new_n3064 = ~new_n3047 & ~new_n3063;
  assign new_n3065 = ~new_n3023 & new_n3027;
  assign new_n3066 = ~new_n3030 & ~new_n3065;
  assign new_n3067 = new_n2910 & ~new_n2945;
  assign new_n3068 = ~new_n2937 & ~new_n3067;
  assign new_n3069 = ~new_n2955 & ~new_n3068;
  assign new_n3070 = ~new_n2908 & ~new_n3067;
  assign new_n3071 = ~new_n2927 & new_n2931;
  assign new_n3072 = ~new_n3070 & new_n3071;
  assign new_n3073 = new_n3070 & ~new_n3071;
  assign new_n3074 = ~new_n3072 & ~new_n3073;
  assign new_n3075 = ~new_n3069 & new_n3074;
  assign new_n3076 = new_n3069 & ~new_n3074;
  assign new_n3077 = ~new_n3075 & ~new_n3076;
  assign new_n3078 = ~new_n3007 & ~new_n3023;
  assign new_n3079 = ~new_n3006 & ~new_n3078;
  assign new_n3080 = ~new_n2987 & new_n2999;
  assign new_n3081 = ~new_n2968 & ~new_n2977;
  assign new_n3082 = new_n3080 & new_n3081;
  assign new_n3083 = ~new_n3080 & ~new_n3081;
  assign new_n3084 = ~new_n3082 & ~new_n3083;
  assign new_n3085 = ~new_n3079 & new_n3084;
  assign new_n3086 = new_n3079 & ~new_n3084;
  assign new_n3087 = ~new_n3085 & ~new_n3086;
  assign new_n3088 = ~new_n3077 & ~new_n3087;
  assign new_n3089 = new_n3077 & new_n3087;
  assign new_n3090 = ~new_n3088 & ~new_n3089;
  assign new_n3091 = ~new_n3066 & new_n3090;
  assign new_n3092 = new_n3066 & ~new_n3090;
  assign new_n3093 = ~new_n3091 & ~new_n3092;
  assign new_n3094 = ~new_n2821 & ~new_n2824;
  assign new_n3095 = ~new_n2743 & ~new_n2766;
  assign new_n3096 = ~new_n2751 & ~new_n3095;
  assign new_n3097 = ~new_n2773 & ~new_n2817;
  assign new_n3098 = ~new_n2808 & ~new_n3097;
  assign new_n3099 = new_n3096 & new_n3098;
  assign new_n3100 = ~new_n3096 & ~new_n3098;
  assign new_n3101 = ~new_n3099 & ~new_n3100;
  assign new_n3102 = ~new_n3094 & new_n3101;
  assign new_n3103 = new_n3094 & ~new_n3101;
  assign new_n3104 = ~new_n3102 & ~new_n3103;
  assign new_n3105 = ~new_n2854 & ~new_n2885;
  assign new_n3106 = ~new_n2876 & ~new_n3105;
  assign new_n3107 = ~new_n2841 & ~new_n2845;
  assign new_n3108 = new_n3106 & ~new_n3107;
  assign new_n3109 = ~new_n3106 & new_n3107;
  assign new_n3110 = ~new_n3108 & ~new_n3109;
  assign new_n3111 = ~new_n2889 & ~new_n2892;
  assign new_n3112 = new_n3110 & new_n3111;
  assign new_n3113 = ~new_n3110 & ~new_n3111;
  assign new_n3114 = ~new_n3112 & ~new_n3113;
  assign new_n3115 = ~new_n2895 & ~new_n3062;
  assign new_n3116 = ~new_n3114 & new_n3115;
  assign new_n3117 = new_n3114 & ~new_n3115;
  assign new_n3118 = ~new_n3116 & ~new_n3117;
  assign new_n3119 = ~new_n3104 & new_n3118;
  assign new_n3120 = new_n3104 & ~new_n3118;
  assign new_n3121 = ~new_n3119 & ~new_n3120;
  assign new_n3122 = new_n3093 & new_n3121;
  assign new_n3123 = ~new_n3093 & ~new_n3121;
  assign new_n3124 = ~new_n3122 & ~new_n3123;
  assign new_n3125 = new_n3064 & new_n3124;
  assign new_n3126 = ~new_n3064 & ~new_n3124;
  assign new_n3127 = ~new_n3125 & ~new_n3126;
  assign new_n3128 = ~new_n3061 & new_n3127;
  assign new_n3129 = new_n3061 & ~new_n3127;
  assign new_n3130 = ~new_n3128 & ~new_n3129;
  assign new_n3131 = ~new_n2737 & new_n3130;
  assign new_n3132 = new_n2737 & ~new_n3130;
  assign new_n3133 = ~new_n3131 & ~new_n3132;
  assign new_n3134 = ~new_n3056 & ~new_n3058;
  assign new_n3135 = new_n2247 & ~new_n2249;
  assign new_n3136 = ~new_n2250 & ~new_n3135;
  assign new_n3137 = ~new_n3059 & ~new_n3134;
  assign new_n3138 = ~new_n3136 & new_n3137;
  assign new_n3139 = ~new_n3134 & ~new_n3138;
  assign new_n3140 = ~new_n3054 & ~new_n3139;
  assign new_n3141 = new_n2254 & ~new_n2256;
  assign new_n3142 = ~new_n2257 & ~new_n3141;
  assign new_n3143 = new_n3054 & new_n3139;
  assign new_n3144 = ~new_n3140 & ~new_n3143;
  assign new_n3145 = new_n3142 & new_n3144;
  assign new_n3146 = ~new_n3060 & ~new_n3140;
  assign new_n3147 = ~new_n3145 & new_n3146;
  assign new_n3148 = new_n3133 & new_n3147;
  assign new_n3149 = ~new_n2261 & ~new_n2263;
  assign new_n3150 = ~new_n2264 & ~new_n3149;
  assign new_n3151 = ~new_n3133 & ~new_n3147;
  assign new_n3152 = ~new_n3148 & ~new_n3151;
  assign new_n3153 = ~new_n3150 & new_n3152;
  assign new_n3154 = ~new_n3148 & ~new_n3153;
  assign new_n3155 = ~new_n2316 & new_n3154;
  assign new_n3156 = ~new_n2708 & ~new_n2711;
  assign new_n3157 = ~new_n2691 & ~new_n2694;
  assign new_n3158 = ~new_n2702 & ~new_n2705;
  assign new_n3159 = new_n3157 & new_n3158;
  assign new_n3160 = ~new_n3157 & ~new_n3158;
  assign new_n3161 = ~new_n3159 & ~new_n3160;
  assign new_n3162 = ~new_n3156 & new_n3161;
  assign new_n3163 = new_n3156 & ~new_n3161;
  assign new_n3164 = ~new_n3162 & ~new_n3163;
  assign new_n3165 = ~new_n2366 & ~new_n2390;
  assign new_n3166 = ~new_n2479 & ~new_n2482;
  assign new_n3167 = new_n3165 & ~new_n3166;
  assign new_n3168 = ~new_n3165 & new_n3166;
  assign new_n3169 = ~new_n3167 & ~new_n3168;
  assign new_n3170 = ~new_n2499 & ~new_n2502;
  assign new_n3171 = new_n3169 & ~new_n3170;
  assign new_n3172 = ~new_n3169 & new_n3170;
  assign new_n3173 = ~new_n3171 & ~new_n3172;
  assign new_n3174 = new_n3164 & ~new_n3173;
  assign new_n3175 = ~new_n3164 & new_n3173;
  assign new_n3176 = ~new_n3174 & ~new_n3175;
  assign new_n3177 = ~new_n2732 & ~new_n2735;
  assign new_n3178 = new_n3176 & new_n3177;
  assign new_n3179 = ~new_n3176 & ~new_n3177;
  assign new_n3180 = ~new_n3178 & ~new_n3179;
  assign new_n3181 = ~new_n3116 & ~new_n3119;
  assign new_n3182 = ~new_n3108 & ~new_n3112;
  assign new_n3183 = ~new_n3099 & ~new_n3102;
  assign new_n3184 = new_n3182 & new_n3183;
  assign new_n3185 = ~new_n3182 & ~new_n3183;
  assign new_n3186 = ~new_n3184 & ~new_n3185;
  assign new_n3187 = ~new_n3181 & new_n3186;
  assign new_n3188 = new_n3181 & ~new_n3186;
  assign new_n3189 = ~new_n3187 & ~new_n3188;
  assign new_n3190 = ~new_n3082 & ~new_n3085;
  assign new_n3191 = ~new_n3072 & ~new_n3075;
  assign new_n3192 = ~new_n3190 & ~new_n3191;
  assign new_n3193 = new_n3190 & new_n3191;
  assign new_n3194 = ~new_n3192 & ~new_n3193;
  assign new_n3195 = ~new_n3088 & ~new_n3091;
  assign new_n3196 = new_n3194 & new_n3195;
  assign new_n3197 = ~new_n3194 & ~new_n3195;
  assign new_n3198 = ~new_n3196 & ~new_n3197;
  assign new_n3199 = new_n3189 & ~new_n3198;
  assign new_n3200 = ~new_n3189 & new_n3198;
  assign new_n3201 = ~new_n3199 & ~new_n3200;
  assign new_n3202 = ~new_n3122 & ~new_n3125;
  assign new_n3203 = new_n3201 & ~new_n3202;
  assign new_n3204 = ~new_n3201 & new_n3202;
  assign new_n3205 = ~new_n3203 & ~new_n3204;
  assign new_n3206 = ~new_n3180 & ~new_n3205;
  assign new_n3207 = new_n3180 & new_n3205;
  assign new_n3208 = ~new_n3206 & ~new_n3207;
  assign new_n3209 = ~new_n3128 & ~new_n3131;
  assign new_n3210 = new_n3208 & new_n3209;
  assign new_n3211 = ~new_n3208 & ~new_n3209;
  assign new_n3212 = ~new_n3210 & ~new_n3211;
  assign new_n3213 = new_n2316 & ~new_n3154;
  assign new_n3214 = ~new_n3155 & ~new_n3213;
  assign new_n3215 = new_n3212 & new_n3214;
  assign new_n3216 = ~new_n3155 & ~new_n3215;
  assign new_n3217 = ~new_n2294 & ~new_n2296;
  assign new_n3218 = ~new_n2297 & ~new_n3217;
  assign new_n3219 = ~new_n3216 & new_n3218;
  assign new_n3220 = ~new_n3167 & ~new_n3171;
  assign new_n3221 = ~new_n3159 & ~new_n3162;
  assign new_n3222 = ~new_n3220 & new_n3221;
  assign new_n3223 = new_n3220 & ~new_n3221;
  assign new_n3224 = ~new_n3222 & ~new_n3223;
  assign new_n3225 = ~new_n3174 & ~new_n3178;
  assign new_n3226 = new_n3224 & new_n3225;
  assign new_n3227 = ~new_n3224 & ~new_n3225;
  assign new_n3228 = ~new_n3226 & ~new_n3227;
  assign new_n3229 = ~new_n3192 & ~new_n3196;
  assign new_n3230 = ~new_n3184 & ~new_n3187;
  assign new_n3231 = ~new_n3229 & new_n3230;
  assign new_n3232 = new_n3229 & ~new_n3230;
  assign new_n3233 = ~new_n3231 & ~new_n3232;
  assign new_n3234 = ~new_n3199 & ~new_n3203;
  assign new_n3235 = new_n3233 & new_n3234;
  assign new_n3236 = ~new_n3233 & ~new_n3234;
  assign new_n3237 = ~new_n3235 & ~new_n3236;
  assign new_n3238 = new_n3228 & new_n3237;
  assign new_n3239 = ~new_n3228 & ~new_n3237;
  assign new_n3240 = ~new_n3238 & ~new_n3239;
  assign new_n3241 = ~new_n3206 & ~new_n3210;
  assign new_n3242 = new_n3240 & ~new_n3241;
  assign new_n3243 = ~new_n3240 & new_n3241;
  assign new_n3244 = ~new_n3242 & ~new_n3243;
  assign new_n3245 = new_n3216 & ~new_n3218;
  assign new_n3246 = ~new_n3219 & ~new_n3245;
  assign new_n3247 = new_n3244 & new_n3246;
  assign new_n3248 = ~new_n3219 & ~new_n3247;
  assign new_n3249 = ~new_n2314 & ~new_n3248;
  assign new_n3250 = ~new_n3222 & ~new_n3226;
  assign new_n3251 = ~new_n3231 & ~new_n3235;
  assign new_n3252 = ~new_n3250 & ~new_n3251;
  assign new_n3253 = new_n3250 & new_n3251;
  assign new_n3254 = ~new_n3252 & ~new_n3253;
  assign new_n3255 = ~new_n3238 & ~new_n3242;
  assign new_n3256 = new_n3254 & new_n3255;
  assign new_n3257 = ~new_n3254 & ~new_n3255;
  assign new_n3258 = ~new_n3256 & ~new_n3257;
  assign new_n3259 = new_n2314 & new_n3248;
  assign new_n3260 = ~new_n3249 & ~new_n3259;
  assign new_n3261 = ~new_n3258 & new_n3260;
  assign new_n3262 = ~new_n3249 & ~new_n3261;
  assign new_n3263 = ~new_n2309 & ~new_n2313;
  assign new_n3264 = new_n3262 & ~new_n3263;
  assign new_n3265 = ~new_n3253 & ~new_n3256;
  assign new_n3266 = ~new_n2307 & new_n3265;
  assign new_n3267 = ~new_n3262 & new_n3263;
  assign new_n3268 = ~new_n3264 & ~new_n3267;
  assign new_n3269 = new_n2307 & ~new_n3265;
  assign new_n3270 = ~new_n3266 & ~new_n3269;
  assign new_n3271 = ~new_n3268 & new_n3270;
  assign new_n3272 = ~new_n3266 & ~new_n3271;
  assign new_n3273 = ~new_n3264 & ~new_n3272;
  assign new_n3274 = ~A199 & ~A200;
  assign new_n3275 = A202 & A203;
  assign new_n3276 = ~A201 & A204;
  assign new_n3277 = new_n3275 & new_n3276;
  assign new_n3278 = A199 & A200;
  assign new_n3279 = ~A201 & ~new_n3278;
  assign new_n3280 = ~A202 & ~A203;
  assign new_n3281 = ~new_n3275 & ~new_n3280;
  assign new_n3282 = A204 & ~new_n3281;
  assign new_n3283 = ~A204 & ~new_n3275;
  assign new_n3284 = ~new_n3279 & ~new_n3283;
  assign new_n3285 = ~new_n3282 & new_n3284;
  assign new_n3286 = ~new_n3277 & ~new_n3285;
  assign new_n3287 = ~new_n3274 & ~new_n3286;
  assign new_n3288 = ~new_n3275 & ~new_n3278;
  assign new_n3289 = A201 & A204;
  assign new_n3290 = ~new_n3288 & new_n3289;
  assign new_n3291 = A203 & new_n3278;
  assign new_n3292 = new_n3290 & ~new_n3291;
  assign new_n3293 = new_n3274 & new_n3280;
  assign new_n3294 = ~new_n3289 & new_n3293;
  assign new_n3295 = A201 & ~A204;
  assign new_n3296 = new_n3278 & ~new_n3280;
  assign new_n3297 = new_n3295 & new_n3296;
  assign new_n3298 = ~new_n3294 & ~new_n3297;
  assign new_n3299 = ~new_n3292 & new_n3298;
  assign new_n3300 = ~new_n3287 & new_n3299;
  assign new_n3301 = ~new_n3274 & ~new_n3278;
  assign new_n3302 = ~new_n3276 & ~new_n3295;
  assign new_n3303 = new_n3301 & ~new_n3302;
  assign new_n3304 = ~new_n3301 & new_n3302;
  assign new_n3305 = ~new_n3303 & ~new_n3304;
  assign new_n3306 = new_n3281 & new_n3305;
  assign new_n3307 = new_n3279 & new_n3283;
  assign new_n3308 = ~new_n3306 & new_n3307;
  assign new_n3309 = new_n3300 & ~new_n3308;
  assign new_n3310 = ~A208 & ~A209;
  assign new_n3311 = ~A206 & ~A207;
  assign new_n3312 = A206 & A207;
  assign new_n3313 = ~new_n3311 & ~new_n3312;
  assign new_n3314 = ~A205 & new_n3313;
  assign new_n3315 = ~new_n3311 & ~new_n3314;
  assign new_n3316 = A205 & ~new_n3313;
  assign new_n3317 = ~new_n3314 & ~new_n3316;
  assign new_n3318 = A210 & ~new_n3317;
  assign new_n3319 = new_n3310 & ~new_n3315;
  assign new_n3320 = ~new_n3318 & new_n3319;
  assign new_n3321 = ~new_n3310 & new_n3315;
  assign new_n3322 = A208 & A209;
  assign new_n3323 = ~A210 & ~new_n3322;
  assign new_n3324 = new_n3321 & ~new_n3323;
  assign new_n3325 = ~new_n3315 & new_n3323;
  assign new_n3326 = ~new_n3324 & ~new_n3325;
  assign new_n3327 = new_n3317 & ~new_n3326;
  assign new_n3328 = ~A210 & ~new_n3321;
  assign new_n3329 = ~new_n3315 & ~new_n3322;
  assign new_n3330 = new_n3315 & new_n3322;
  assign new_n3331 = ~new_n3329 & ~new_n3330;
  assign new_n3332 = A210 & ~new_n3331;
  assign new_n3333 = ~new_n3317 & ~new_n3328;
  assign new_n3334 = ~new_n3332 & new_n3333;
  assign new_n3335 = ~new_n3320 & ~new_n3327;
  assign new_n3336 = ~new_n3334 & new_n3335;
  assign new_n3337 = ~new_n3309 & ~new_n3336;
  assign new_n3338 = ~new_n3281 & ~new_n3305;
  assign new_n3339 = ~new_n3306 & ~new_n3338;
  assign new_n3340 = ~A210 & new_n3317;
  assign new_n3341 = ~new_n3318 & ~new_n3340;
  assign new_n3342 = ~new_n3310 & ~new_n3322;
  assign new_n3343 = ~new_n3341 & new_n3342;
  assign new_n3344 = new_n3341 & ~new_n3342;
  assign new_n3345 = ~new_n3343 & ~new_n3344;
  assign new_n3346 = new_n3339 & ~new_n3345;
  assign new_n3347 = new_n3309 & new_n3336;
  assign new_n3348 = ~new_n3337 & ~new_n3347;
  assign new_n3349 = ~new_n3346 & new_n3348;
  assign new_n3350 = ~new_n3337 & ~new_n3349;
  assign new_n3351 = ~new_n3274 & ~new_n3300;
  assign new_n3352 = ~new_n3290 & ~new_n3351;
  assign new_n3353 = ~new_n3324 & ~new_n3334;
  assign new_n3354 = new_n3352 & new_n3353;
  assign new_n3355 = ~new_n3352 & ~new_n3353;
  assign new_n3356 = ~new_n3354 & ~new_n3355;
  assign new_n3357 = ~new_n3350 & new_n3356;
  assign new_n3358 = new_n3350 & ~new_n3356;
  assign new_n3359 = ~new_n3357 & ~new_n3358;
  assign new_n3360 = A214 & A215;
  assign new_n3361 = ~A214 & ~A215;
  assign new_n3362 = ~new_n3360 & ~new_n3361;
  assign new_n3363 = A211 & A212;
  assign new_n3364 = ~A211 & ~A212;
  assign new_n3365 = ~new_n3363 & ~new_n3364;
  assign new_n3366 = ~A213 & A216;
  assign new_n3367 = A213 & ~A216;
  assign new_n3368 = ~new_n3366 & ~new_n3367;
  assign new_n3369 = new_n3365 & ~new_n3368;
  assign new_n3370 = ~new_n3365 & new_n3368;
  assign new_n3371 = ~new_n3369 & ~new_n3370;
  assign new_n3372 = new_n3362 & new_n3371;
  assign new_n3373 = ~new_n3362 & ~new_n3371;
  assign new_n3374 = ~new_n3372 & ~new_n3373;
  assign new_n3375 = ~A218 & ~A219;
  assign new_n3376 = A218 & A219;
  assign new_n3377 = ~new_n3375 & ~new_n3376;
  assign new_n3378 = ~A217 & new_n3377;
  assign new_n3379 = A217 & ~new_n3377;
  assign new_n3380 = ~new_n3378 & ~new_n3379;
  assign new_n3381 = A222 & ~new_n3380;
  assign new_n3382 = ~A222 & new_n3380;
  assign new_n3383 = ~new_n3381 & ~new_n3382;
  assign new_n3384 = ~A220 & ~A221;
  assign new_n3385 = A220 & A221;
  assign new_n3386 = ~new_n3384 & ~new_n3385;
  assign new_n3387 = ~new_n3383 & new_n3386;
  assign new_n3388 = new_n3383 & ~new_n3386;
  assign new_n3389 = ~new_n3387 & ~new_n3388;
  assign new_n3390 = new_n3374 & ~new_n3389;
  assign new_n3391 = ~new_n3374 & new_n3389;
  assign new_n3392 = ~new_n3390 & ~new_n3391;
  assign new_n3393 = ~new_n3339 & new_n3345;
  assign new_n3394 = ~new_n3346 & ~new_n3393;
  assign new_n3395 = new_n3392 & new_n3394;
  assign new_n3396 = new_n3348 & new_n3395;
  assign new_n3397 = new_n3360 & new_n3366;
  assign new_n3398 = ~A213 & ~new_n3363;
  assign new_n3399 = A216 & ~new_n3362;
  assign new_n3400 = ~A216 & ~new_n3360;
  assign new_n3401 = ~new_n3398 & ~new_n3400;
  assign new_n3402 = ~new_n3399 & new_n3401;
  assign new_n3403 = ~new_n3397 & ~new_n3402;
  assign new_n3404 = ~new_n3364 & ~new_n3403;
  assign new_n3405 = A213 & A216;
  assign new_n3406 = ~new_n3360 & ~new_n3363;
  assign new_n3407 = new_n3405 & ~new_n3406;
  assign new_n3408 = A215 & new_n3363;
  assign new_n3409 = new_n3407 & ~new_n3408;
  assign new_n3410 = new_n3361 & new_n3364;
  assign new_n3411 = ~new_n3405 & new_n3410;
  assign new_n3412 = ~new_n3361 & new_n3363;
  assign new_n3413 = new_n3367 & new_n3412;
  assign new_n3414 = ~new_n3411 & ~new_n3413;
  assign new_n3415 = ~new_n3409 & new_n3414;
  assign new_n3416 = ~new_n3404 & new_n3415;
  assign new_n3417 = new_n3398 & new_n3400;
  assign new_n3418 = ~new_n3372 & new_n3417;
  assign new_n3419 = new_n3416 & ~new_n3418;
  assign new_n3420 = ~new_n3375 & ~new_n3378;
  assign new_n3421 = new_n3384 & ~new_n3420;
  assign new_n3422 = ~new_n3381 & new_n3421;
  assign new_n3423 = ~new_n3384 & new_n3420;
  assign new_n3424 = ~A222 & ~new_n3385;
  assign new_n3425 = new_n3423 & ~new_n3424;
  assign new_n3426 = ~new_n3420 & new_n3424;
  assign new_n3427 = ~new_n3425 & ~new_n3426;
  assign new_n3428 = new_n3380 & ~new_n3427;
  assign new_n3429 = ~A222 & ~new_n3423;
  assign new_n3430 = ~new_n3385 & ~new_n3420;
  assign new_n3431 = new_n3385 & new_n3420;
  assign new_n3432 = ~new_n3430 & ~new_n3431;
  assign new_n3433 = A222 & ~new_n3432;
  assign new_n3434 = ~new_n3380 & ~new_n3429;
  assign new_n3435 = ~new_n3433 & new_n3434;
  assign new_n3436 = ~new_n3422 & ~new_n3428;
  assign new_n3437 = ~new_n3435 & new_n3436;
  assign new_n3438 = ~new_n3419 & ~new_n3437;
  assign new_n3439 = new_n3419 & new_n3437;
  assign new_n3440 = ~new_n3438 & ~new_n3439;
  assign new_n3441 = ~new_n3390 & new_n3440;
  assign new_n3442 = new_n3390 & ~new_n3440;
  assign new_n3443 = ~new_n3441 & ~new_n3442;
  assign new_n3444 = ~new_n3346 & ~new_n3395;
  assign new_n3445 = new_n3348 & ~new_n3444;
  assign new_n3446 = ~new_n3348 & new_n3444;
  assign new_n3447 = ~new_n3445 & ~new_n3446;
  assign new_n3448 = ~new_n3443 & new_n3447;
  assign new_n3449 = ~new_n3396 & ~new_n3448;
  assign new_n3450 = ~new_n3359 & ~new_n3449;
  assign new_n3451 = ~new_n3438 & ~new_n3441;
  assign new_n3452 = ~new_n3364 & ~new_n3416;
  assign new_n3453 = ~new_n3407 & ~new_n3452;
  assign new_n3454 = ~new_n3425 & ~new_n3435;
  assign new_n3455 = new_n3453 & new_n3454;
  assign new_n3456 = ~new_n3453 & ~new_n3454;
  assign new_n3457 = ~new_n3455 & ~new_n3456;
  assign new_n3458 = ~new_n3451 & new_n3457;
  assign new_n3459 = new_n3451 & ~new_n3457;
  assign new_n3460 = ~new_n3458 & ~new_n3459;
  assign new_n3461 = new_n3359 & new_n3449;
  assign new_n3462 = ~new_n3450 & ~new_n3461;
  assign new_n3463 = ~new_n3460 & new_n3462;
  assign new_n3464 = ~new_n3450 & ~new_n3463;
  assign new_n3465 = ~new_n3455 & ~new_n3458;
  assign new_n3466 = ~new_n3354 & ~new_n3357;
  assign new_n3467 = new_n3465 & new_n3466;
  assign new_n3468 = ~new_n3465 & ~new_n3466;
  assign new_n3469 = ~new_n3467 & ~new_n3468;
  assign new_n3470 = ~new_n3464 & new_n3469;
  assign new_n3471 = new_n3464 & ~new_n3469;
  assign new_n3472 = ~new_n3470 & ~new_n3471;
  assign new_n3473 = new_n3460 & ~new_n3462;
  assign new_n3474 = ~new_n3463 & ~new_n3473;
  assign new_n3475 = new_n3443 & ~new_n3447;
  assign new_n3476 = ~new_n3448 & ~new_n3475;
  assign new_n3477 = A184 & A185;
  assign new_n3478 = ~A184 & ~A185;
  assign new_n3479 = ~new_n3477 & ~new_n3478;
  assign new_n3480 = A181 & A182;
  assign new_n3481 = ~A181 & ~A182;
  assign new_n3482 = ~new_n3480 & ~new_n3481;
  assign new_n3483 = ~A183 & A186;
  assign new_n3484 = A183 & ~A186;
  assign new_n3485 = ~new_n3483 & ~new_n3484;
  assign new_n3486 = new_n3482 & ~new_n3485;
  assign new_n3487 = ~new_n3482 & new_n3485;
  assign new_n3488 = ~new_n3486 & ~new_n3487;
  assign new_n3489 = new_n3479 & new_n3488;
  assign new_n3490 = ~new_n3479 & ~new_n3488;
  assign new_n3491 = ~new_n3489 & ~new_n3490;
  assign new_n3492 = ~A179 & ~A180;
  assign new_n3493 = A179 & A180;
  assign new_n3494 = ~new_n3492 & ~new_n3493;
  assign new_n3495 = ~A178 & new_n3494;
  assign new_n3496 = A178 & ~new_n3494;
  assign new_n3497 = ~new_n3495 & ~new_n3496;
  assign new_n3498 = ~A176 & ~A177;
  assign new_n3499 = A176 & A177;
  assign new_n3500 = ~new_n3498 & ~new_n3499;
  assign new_n3501 = ~A175 & new_n3500;
  assign new_n3502 = A175 & ~new_n3500;
  assign new_n3503 = ~new_n3501 & ~new_n3502;
  assign new_n3504 = ~new_n3497 & ~new_n3503;
  assign new_n3505 = new_n3497 & new_n3503;
  assign new_n3506 = ~new_n3504 & ~new_n3505;
  assign new_n3507 = ~new_n3491 & new_n3506;
  assign new_n3508 = new_n3491 & ~new_n3506;
  assign new_n3509 = ~new_n3507 & ~new_n3508;
  assign new_n3510 = ~A194 & ~A195;
  assign new_n3511 = A194 & A195;
  assign new_n3512 = ~new_n3510 & ~new_n3511;
  assign new_n3513 = A193 & new_n3512;
  assign new_n3514 = ~A193 & ~new_n3512;
  assign new_n3515 = ~new_n3513 & ~new_n3514;
  assign new_n3516 = A197 & A198;
  assign new_n3517 = ~A197 & ~A198;
  assign new_n3518 = ~new_n3516 & ~new_n3517;
  assign new_n3519 = A196 & ~new_n3518;
  assign new_n3520 = ~A196 & new_n3518;
  assign new_n3521 = ~new_n3519 & ~new_n3520;
  assign new_n3522 = ~new_n3515 & ~new_n3521;
  assign new_n3523 = new_n3515 & new_n3521;
  assign new_n3524 = ~new_n3522 & ~new_n3523;
  assign new_n3525 = ~A188 & ~A189;
  assign new_n3526 = A188 & A189;
  assign new_n3527 = ~new_n3525 & ~new_n3526;
  assign new_n3528 = ~A187 & new_n3527;
  assign new_n3529 = A187 & ~new_n3527;
  assign new_n3530 = ~new_n3528 & ~new_n3529;
  assign new_n3531 = ~A191 & ~A192;
  assign new_n3532 = A191 & A192;
  assign new_n3533 = ~new_n3531 & ~new_n3532;
  assign new_n3534 = ~A190 & new_n3533;
  assign new_n3535 = A190 & ~new_n3533;
  assign new_n3536 = ~new_n3534 & ~new_n3535;
  assign new_n3537 = ~new_n3530 & ~new_n3536;
  assign new_n3538 = new_n3530 & new_n3536;
  assign new_n3539 = ~new_n3537 & ~new_n3538;
  assign new_n3540 = ~new_n3524 & new_n3539;
  assign new_n3541 = new_n3524 & ~new_n3539;
  assign new_n3542 = ~new_n3540 & ~new_n3541;
  assign new_n3543 = ~new_n3509 & new_n3542;
  assign new_n3544 = ~new_n3498 & ~new_n3501;
  assign new_n3545 = ~new_n3492 & ~new_n3495;
  assign new_n3546 = new_n3544 & new_n3545;
  assign new_n3547 = ~new_n3544 & ~new_n3545;
  assign new_n3548 = ~new_n3546 & ~new_n3547;
  assign new_n3549 = ~new_n3505 & ~new_n3507;
  assign new_n3550 = new_n3477 & new_n3483;
  assign new_n3551 = ~A183 & ~new_n3480;
  assign new_n3552 = A186 & ~new_n3479;
  assign new_n3553 = ~A186 & ~new_n3477;
  assign new_n3554 = ~new_n3551 & ~new_n3553;
  assign new_n3555 = ~new_n3552 & new_n3554;
  assign new_n3556 = ~new_n3550 & ~new_n3555;
  assign new_n3557 = ~new_n3481 & ~new_n3556;
  assign new_n3558 = A183 & A186;
  assign new_n3559 = ~new_n3477 & ~new_n3480;
  assign new_n3560 = new_n3558 & ~new_n3559;
  assign new_n3561 = A185 & new_n3480;
  assign new_n3562 = new_n3560 & ~new_n3561;
  assign new_n3563 = new_n3478 & new_n3481;
  assign new_n3564 = ~new_n3558 & new_n3563;
  assign new_n3565 = ~new_n3478 & new_n3480;
  assign new_n3566 = new_n3484 & new_n3565;
  assign new_n3567 = ~new_n3564 & ~new_n3566;
  assign new_n3568 = ~new_n3562 & new_n3567;
  assign new_n3569 = ~new_n3557 & new_n3568;
  assign new_n3570 = new_n3551 & new_n3553;
  assign new_n3571 = ~new_n3489 & new_n3570;
  assign new_n3572 = new_n3569 & ~new_n3571;
  assign new_n3573 = ~new_n3549 & ~new_n3572;
  assign new_n3574 = new_n3549 & new_n3572;
  assign new_n3575 = ~new_n3573 & ~new_n3574;
  assign new_n3576 = ~new_n3548 & new_n3575;
  assign new_n3577 = new_n3548 & ~new_n3575;
  assign new_n3578 = ~new_n3576 & ~new_n3577;
  assign new_n3579 = ~new_n3537 & ~new_n3540;
  assign new_n3580 = ~new_n3525 & ~new_n3528;
  assign new_n3581 = ~new_n3531 & ~new_n3534;
  assign new_n3582 = new_n3580 & new_n3581;
  assign new_n3583 = ~new_n3580 & ~new_n3581;
  assign new_n3584 = ~new_n3582 & ~new_n3583;
  assign new_n3585 = ~new_n3511 & ~new_n3513;
  assign new_n3586 = new_n3516 & ~new_n3585;
  assign new_n3587 = A193 & A194;
  assign new_n3588 = ~new_n3516 & ~new_n3587;
  assign new_n3589 = ~A193 & ~A194;
  assign new_n3590 = ~new_n3517 & ~new_n3589;
  assign new_n3591 = ~A195 & new_n3588;
  assign new_n3592 = ~new_n3590 & new_n3591;
  assign new_n3593 = ~new_n3586 & ~new_n3592;
  assign new_n3594 = ~A196 & ~new_n3593;
  assign new_n3595 = A195 & A196;
  assign new_n3596 = ~new_n3588 & new_n3595;
  assign new_n3597 = A198 & new_n3587;
  assign new_n3598 = new_n3596 & ~new_n3597;
  assign new_n3599 = new_n3517 & new_n3589;
  assign new_n3600 = ~new_n3595 & new_n3599;
  assign new_n3601 = ~A195 & new_n3590;
  assign new_n3602 = new_n3519 & new_n3601;
  assign new_n3603 = new_n3518 & ~new_n3585;
  assign new_n3604 = ~new_n3522 & new_n3603;
  assign new_n3605 = ~new_n3598 & ~new_n3600;
  assign new_n3606 = ~new_n3602 & new_n3605;
  assign new_n3607 = ~new_n3604 & new_n3606;
  assign new_n3608 = ~new_n3594 & new_n3607;
  assign new_n3609 = ~new_n3584 & ~new_n3608;
  assign new_n3610 = new_n3584 & new_n3608;
  assign new_n3611 = ~new_n3609 & ~new_n3610;
  assign new_n3612 = new_n3579 & new_n3611;
  assign new_n3613 = ~new_n3579 & ~new_n3611;
  assign new_n3614 = ~new_n3612 & ~new_n3613;
  assign new_n3615 = new_n3578 & new_n3614;
  assign new_n3616 = ~new_n3578 & ~new_n3614;
  assign new_n3617 = ~new_n3615 & ~new_n3616;
  assign new_n3618 = ~new_n3543 & new_n3617;
  assign new_n3619 = new_n3543 & ~new_n3617;
  assign new_n3620 = ~new_n3618 & ~new_n3619;
  assign new_n3621 = new_n3476 & ~new_n3620;
  assign new_n3622 = ~new_n3392 & ~new_n3394;
  assign new_n3623 = ~new_n3395 & ~new_n3622;
  assign new_n3624 = new_n3509 & ~new_n3542;
  assign new_n3625 = ~new_n3543 & ~new_n3624;
  assign new_n3626 = new_n3623 & new_n3625;
  assign new_n3627 = ~new_n3476 & new_n3620;
  assign new_n3628 = new_n3626 & ~new_n3627;
  assign new_n3629 = ~new_n3621 & ~new_n3628;
  assign new_n3630 = new_n3474 & ~new_n3629;
  assign new_n3631 = ~new_n3481 & ~new_n3569;
  assign new_n3632 = ~new_n3560 & ~new_n3631;
  assign new_n3633 = new_n3504 & new_n3548;
  assign new_n3634 = ~new_n3546 & ~new_n3633;
  assign new_n3635 = ~new_n3632 & ~new_n3634;
  assign new_n3636 = new_n3632 & new_n3634;
  assign new_n3637 = ~new_n3635 & ~new_n3636;
  assign new_n3638 = ~new_n3573 & ~new_n3633;
  assign new_n3639 = ~new_n3576 & new_n3638;
  assign new_n3640 = new_n3637 & new_n3639;
  assign new_n3641 = ~new_n3637 & ~new_n3639;
  assign new_n3642 = ~new_n3640 & ~new_n3641;
  assign new_n3643 = new_n3590 & ~new_n3608;
  assign new_n3644 = ~new_n3596 & ~new_n3643;
  assign new_n3645 = new_n3537 & new_n3584;
  assign new_n3646 = ~new_n3582 & ~new_n3645;
  assign new_n3647 = ~new_n3644 & ~new_n3646;
  assign new_n3648 = new_n3644 & new_n3646;
  assign new_n3649 = ~new_n3647 & ~new_n3648;
  assign new_n3650 = ~new_n3609 & ~new_n3645;
  assign new_n3651 = ~new_n3612 & new_n3650;
  assign new_n3652 = new_n3649 & new_n3651;
  assign new_n3653 = ~new_n3649 & ~new_n3651;
  assign new_n3654 = ~new_n3652 & ~new_n3653;
  assign new_n3655 = ~new_n3615 & ~new_n3618;
  assign new_n3656 = ~new_n3654 & ~new_n3655;
  assign new_n3657 = new_n3654 & new_n3655;
  assign new_n3658 = ~new_n3656 & ~new_n3657;
  assign new_n3659 = ~new_n3642 & new_n3658;
  assign new_n3660 = new_n3642 & ~new_n3658;
  assign new_n3661 = ~new_n3659 & ~new_n3660;
  assign new_n3662 = ~new_n3474 & new_n3629;
  assign new_n3663 = ~new_n3630 & ~new_n3662;
  assign new_n3664 = ~new_n3661 & new_n3663;
  assign new_n3665 = ~new_n3630 & ~new_n3664;
  assign new_n3666 = new_n3472 & ~new_n3665;
  assign new_n3667 = ~new_n3656 & ~new_n3659;
  assign new_n3668 = ~new_n3635 & ~new_n3640;
  assign new_n3669 = ~new_n3647 & ~new_n3652;
  assign new_n3670 = new_n3668 & new_n3669;
  assign new_n3671 = ~new_n3668 & ~new_n3669;
  assign new_n3672 = ~new_n3670 & ~new_n3671;
  assign new_n3673 = ~new_n3667 & new_n3672;
  assign new_n3674 = new_n3667 & ~new_n3672;
  assign new_n3675 = ~new_n3673 & ~new_n3674;
  assign new_n3676 = ~new_n3472 & new_n3665;
  assign new_n3677 = ~new_n3666 & ~new_n3676;
  assign new_n3678 = ~new_n3675 & new_n3677;
  assign new_n3679 = ~new_n3666 & ~new_n3678;
  assign new_n3680 = ~new_n3670 & ~new_n3673;
  assign new_n3681 = ~new_n3467 & ~new_n3470;
  assign new_n3682 = ~new_n3680 & new_n3681;
  assign new_n3683 = new_n3680 & ~new_n3681;
  assign new_n3684 = ~new_n3682 & ~new_n3683;
  assign new_n3685 = new_n3679 & new_n3684;
  assign new_n3686 = ~new_n3679 & ~new_n3684;
  assign new_n3687 = ~new_n3685 & ~new_n3686;
  assign new_n3688 = ~A235 & ~A236;
  assign new_n3689 = A238 & A239;
  assign new_n3690 = ~A237 & A240;
  assign new_n3691 = new_n3689 & new_n3690;
  assign new_n3692 = A235 & A236;
  assign new_n3693 = ~A237 & ~new_n3692;
  assign new_n3694 = ~A238 & ~A239;
  assign new_n3695 = ~new_n3689 & ~new_n3694;
  assign new_n3696 = A240 & ~new_n3695;
  assign new_n3697 = ~A240 & ~new_n3689;
  assign new_n3698 = ~new_n3693 & ~new_n3697;
  assign new_n3699 = ~new_n3696 & new_n3698;
  assign new_n3700 = ~new_n3691 & ~new_n3699;
  assign new_n3701 = ~new_n3688 & ~new_n3700;
  assign new_n3702 = ~new_n3689 & ~new_n3692;
  assign new_n3703 = A237 & A240;
  assign new_n3704 = ~new_n3702 & new_n3703;
  assign new_n3705 = A239 & new_n3692;
  assign new_n3706 = new_n3704 & ~new_n3705;
  assign new_n3707 = A237 & ~A240;
  assign new_n3708 = new_n3692 & ~new_n3694;
  assign new_n3709 = new_n3707 & new_n3708;
  assign new_n3710 = new_n3688 & new_n3694;
  assign new_n3711 = ~new_n3703 & new_n3710;
  assign new_n3712 = ~new_n3709 & ~new_n3711;
  assign new_n3713 = ~new_n3706 & new_n3712;
  assign new_n3714 = ~new_n3701 & new_n3713;
  assign new_n3715 = ~new_n3688 & ~new_n3692;
  assign new_n3716 = ~new_n3690 & ~new_n3707;
  assign new_n3717 = new_n3715 & ~new_n3716;
  assign new_n3718 = ~new_n3715 & new_n3716;
  assign new_n3719 = ~new_n3717 & ~new_n3718;
  assign new_n3720 = new_n3695 & new_n3719;
  assign new_n3721 = new_n3693 & new_n3697;
  assign new_n3722 = ~new_n3720 & new_n3721;
  assign new_n3723 = new_n3714 & ~new_n3722;
  assign new_n3724 = ~A244 & ~A245;
  assign new_n3725 = ~A242 & ~A243;
  assign new_n3726 = A242 & A243;
  assign new_n3727 = ~new_n3725 & ~new_n3726;
  assign new_n3728 = ~A241 & new_n3727;
  assign new_n3729 = ~new_n3725 & ~new_n3728;
  assign new_n3730 = A241 & ~new_n3727;
  assign new_n3731 = ~new_n3728 & ~new_n3730;
  assign new_n3732 = A246 & ~new_n3731;
  assign new_n3733 = new_n3724 & ~new_n3729;
  assign new_n3734 = ~new_n3732 & new_n3733;
  assign new_n3735 = ~new_n3724 & new_n3729;
  assign new_n3736 = A244 & A245;
  assign new_n3737 = ~A246 & ~new_n3736;
  assign new_n3738 = new_n3735 & ~new_n3737;
  assign new_n3739 = ~new_n3729 & new_n3737;
  assign new_n3740 = ~new_n3738 & ~new_n3739;
  assign new_n3741 = new_n3731 & ~new_n3740;
  assign new_n3742 = ~A246 & ~new_n3735;
  assign new_n3743 = ~new_n3729 & ~new_n3736;
  assign new_n3744 = new_n3729 & new_n3736;
  assign new_n3745 = ~new_n3743 & ~new_n3744;
  assign new_n3746 = A246 & ~new_n3745;
  assign new_n3747 = ~new_n3731 & ~new_n3742;
  assign new_n3748 = ~new_n3746 & new_n3747;
  assign new_n3749 = ~new_n3734 & ~new_n3741;
  assign new_n3750 = ~new_n3748 & new_n3749;
  assign new_n3751 = ~new_n3723 & ~new_n3750;
  assign new_n3752 = ~new_n3695 & ~new_n3719;
  assign new_n3753 = ~new_n3720 & ~new_n3752;
  assign new_n3754 = ~A246 & new_n3731;
  assign new_n3755 = ~new_n3732 & ~new_n3754;
  assign new_n3756 = ~new_n3724 & ~new_n3736;
  assign new_n3757 = ~new_n3755 & new_n3756;
  assign new_n3758 = new_n3755 & ~new_n3756;
  assign new_n3759 = ~new_n3757 & ~new_n3758;
  assign new_n3760 = new_n3753 & ~new_n3759;
  assign new_n3761 = new_n3723 & new_n3750;
  assign new_n3762 = ~new_n3751 & ~new_n3761;
  assign new_n3763 = ~new_n3760 & new_n3762;
  assign new_n3764 = ~new_n3751 & ~new_n3763;
  assign new_n3765 = ~new_n3688 & ~new_n3714;
  assign new_n3766 = ~new_n3704 & ~new_n3765;
  assign new_n3767 = ~new_n3738 & ~new_n3748;
  assign new_n3768 = new_n3766 & new_n3767;
  assign new_n3769 = ~new_n3766 & ~new_n3767;
  assign new_n3770 = ~new_n3768 & ~new_n3769;
  assign new_n3771 = ~new_n3764 & new_n3770;
  assign new_n3772 = new_n3764 & ~new_n3770;
  assign new_n3773 = ~new_n3771 & ~new_n3772;
  assign new_n3774 = ~new_n3753 & new_n3759;
  assign new_n3775 = ~new_n3760 & ~new_n3774;
  assign new_n3776 = A232 & A233;
  assign new_n3777 = ~A232 & ~A233;
  assign new_n3778 = ~new_n3776 & ~new_n3777;
  assign new_n3779 = A229 & A230;
  assign new_n3780 = ~A229 & ~A230;
  assign new_n3781 = ~new_n3779 & ~new_n3780;
  assign new_n3782 = ~A231 & A234;
  assign new_n3783 = A231 & ~A234;
  assign new_n3784 = ~new_n3782 & ~new_n3783;
  assign new_n3785 = new_n3781 & ~new_n3784;
  assign new_n3786 = ~new_n3781 & new_n3784;
  assign new_n3787 = ~new_n3785 & ~new_n3786;
  assign new_n3788 = new_n3778 & new_n3787;
  assign new_n3789 = ~new_n3778 & ~new_n3787;
  assign new_n3790 = ~new_n3788 & ~new_n3789;
  assign new_n3791 = ~A224 & ~A225;
  assign new_n3792 = A224 & A225;
  assign new_n3793 = ~new_n3791 & ~new_n3792;
  assign new_n3794 = ~A223 & new_n3793;
  assign new_n3795 = A223 & ~new_n3793;
  assign new_n3796 = ~new_n3794 & ~new_n3795;
  assign new_n3797 = ~A227 & ~A228;
  assign new_n3798 = A227 & A228;
  assign new_n3799 = ~new_n3797 & ~new_n3798;
  assign new_n3800 = ~A226 & new_n3799;
  assign new_n3801 = A226 & ~new_n3799;
  assign new_n3802 = ~new_n3800 & ~new_n3801;
  assign new_n3803 = ~new_n3796 & ~new_n3802;
  assign new_n3804 = new_n3796 & new_n3802;
  assign new_n3805 = ~new_n3803 & ~new_n3804;
  assign new_n3806 = ~new_n3790 & new_n3805;
  assign new_n3807 = new_n3790 & ~new_n3805;
  assign new_n3808 = ~new_n3806 & ~new_n3807;
  assign new_n3809 = new_n3775 & ~new_n3808;
  assign new_n3810 = new_n3762 & new_n3809;
  assign new_n3811 = ~new_n3791 & ~new_n3794;
  assign new_n3812 = ~new_n3797 & ~new_n3800;
  assign new_n3813 = new_n3811 & new_n3812;
  assign new_n3814 = ~new_n3811 & ~new_n3812;
  assign new_n3815 = ~new_n3813 & ~new_n3814;
  assign new_n3816 = ~new_n3804 & ~new_n3806;
  assign new_n3817 = new_n3776 & new_n3782;
  assign new_n3818 = ~A231 & ~new_n3779;
  assign new_n3819 = A234 & ~new_n3778;
  assign new_n3820 = ~A234 & ~new_n3776;
  assign new_n3821 = ~new_n3818 & ~new_n3820;
  assign new_n3822 = ~new_n3819 & new_n3821;
  assign new_n3823 = ~new_n3817 & ~new_n3822;
  assign new_n3824 = ~new_n3780 & ~new_n3823;
  assign new_n3825 = A231 & A234;
  assign new_n3826 = ~new_n3776 & ~new_n3779;
  assign new_n3827 = new_n3825 & ~new_n3826;
  assign new_n3828 = A233 & new_n3779;
  assign new_n3829 = new_n3827 & ~new_n3828;
  assign new_n3830 = new_n3777 & new_n3780;
  assign new_n3831 = ~new_n3825 & new_n3830;
  assign new_n3832 = ~new_n3777 & new_n3779;
  assign new_n3833 = new_n3783 & new_n3832;
  assign new_n3834 = ~new_n3831 & ~new_n3833;
  assign new_n3835 = ~new_n3829 & new_n3834;
  assign new_n3836 = ~new_n3824 & new_n3835;
  assign new_n3837 = new_n3818 & new_n3820;
  assign new_n3838 = ~new_n3788 & new_n3837;
  assign new_n3839 = new_n3836 & ~new_n3838;
  assign new_n3840 = ~new_n3816 & ~new_n3839;
  assign new_n3841 = new_n3816 & new_n3839;
  assign new_n3842 = ~new_n3840 & ~new_n3841;
  assign new_n3843 = ~new_n3815 & new_n3842;
  assign new_n3844 = new_n3815 & ~new_n3842;
  assign new_n3845 = ~new_n3843 & ~new_n3844;
  assign new_n3846 = ~new_n3760 & ~new_n3809;
  assign new_n3847 = new_n3762 & ~new_n3846;
  assign new_n3848 = ~new_n3762 & new_n3846;
  assign new_n3849 = ~new_n3847 & ~new_n3848;
  assign new_n3850 = ~new_n3845 & new_n3849;
  assign new_n3851 = ~new_n3810 & ~new_n3850;
  assign new_n3852 = new_n3773 & new_n3851;
  assign new_n3853 = ~new_n3780 & ~new_n3836;
  assign new_n3854 = ~new_n3827 & ~new_n3853;
  assign new_n3855 = new_n3803 & new_n3815;
  assign new_n3856 = ~new_n3813 & ~new_n3855;
  assign new_n3857 = ~new_n3854 & ~new_n3856;
  assign new_n3858 = new_n3854 & new_n3856;
  assign new_n3859 = ~new_n3857 & ~new_n3858;
  assign new_n3860 = ~new_n3840 & ~new_n3855;
  assign new_n3861 = ~new_n3843 & new_n3860;
  assign new_n3862 = new_n3859 & new_n3861;
  assign new_n3863 = ~new_n3859 & ~new_n3861;
  assign new_n3864 = ~new_n3862 & ~new_n3863;
  assign new_n3865 = ~new_n3773 & ~new_n3851;
  assign new_n3866 = ~new_n3852 & ~new_n3865;
  assign new_n3867 = ~new_n3864 & new_n3866;
  assign new_n3868 = ~new_n3852 & ~new_n3867;
  assign new_n3869 = ~new_n3857 & ~new_n3862;
  assign new_n3870 = ~new_n3768 & ~new_n3771;
  assign new_n3871 = ~new_n3869 & new_n3870;
  assign new_n3872 = new_n3869 & ~new_n3870;
  assign new_n3873 = ~new_n3871 & ~new_n3872;
  assign new_n3874 = new_n3868 & new_n3873;
  assign new_n3875 = ~new_n3868 & ~new_n3873;
  assign new_n3876 = ~new_n3874 & ~new_n3875;
  assign new_n3877 = A267 & A268;
  assign new_n3878 = ~A267 & ~A268;
  assign new_n3879 = ~new_n3877 & ~new_n3878;
  assign new_n3880 = ~A269 & ~A270;
  assign new_n3881 = A269 & A270;
  assign new_n3882 = ~new_n3880 & ~new_n3881;
  assign new_n3883 = new_n3879 & ~new_n3882;
  assign new_n3884 = ~new_n3879 & new_n3882;
  assign new_n3885 = ~new_n3883 & ~new_n3884;
  assign new_n3886 = A265 & A266;
  assign new_n3887 = ~A265 & ~A266;
  assign new_n3888 = ~new_n3886 & ~new_n3887;
  assign new_n3889 = ~new_n3885 & new_n3888;
  assign new_n3890 = new_n3885 & ~new_n3888;
  assign new_n3891 = ~new_n3889 & ~new_n3890;
  assign new_n3892 = ~A260 & ~A261;
  assign new_n3893 = A260 & A261;
  assign new_n3894 = ~new_n3892 & ~new_n3893;
  assign new_n3895 = ~A259 & new_n3894;
  assign new_n3896 = A259 & ~new_n3894;
  assign new_n3897 = ~new_n3895 & ~new_n3896;
  assign new_n3898 = ~A262 & new_n3897;
  assign new_n3899 = ~new_n3892 & ~new_n3895;
  assign new_n3900 = A263 & A264;
  assign new_n3901 = ~new_n3899 & ~new_n3900;
  assign new_n3902 = new_n3898 & new_n3901;
  assign new_n3903 = new_n3899 & new_n3900;
  assign new_n3904 = ~new_n3896 & new_n3903;
  assign new_n3905 = ~A263 & ~A264;
  assign new_n3906 = new_n3899 & ~new_n3905;
  assign new_n3907 = A262 & new_n3900;
  assign new_n3908 = ~new_n3897 & ~new_n3907;
  assign new_n3909 = new_n3906 & new_n3908;
  assign new_n3910 = ~new_n3902 & ~new_n3904;
  assign new_n3911 = ~new_n3909 & new_n3910;
  assign new_n3912 = ~new_n3891 & ~new_n3911;
  assign new_n3913 = A262 & ~new_n3897;
  assign new_n3914 = ~new_n3898 & ~new_n3913;
  assign new_n3915 = ~new_n3900 & new_n3906;
  assign new_n3916 = new_n3914 & new_n3915;
  assign new_n3917 = ~new_n3898 & new_n3906;
  assign new_n3918 = ~new_n3903 & ~new_n3913;
  assign new_n3919 = ~new_n3901 & ~new_n3918;
  assign new_n3920 = ~new_n3917 & new_n3919;
  assign new_n3921 = new_n3891 & ~new_n3898;
  assign new_n3922 = ~new_n3899 & new_n3905;
  assign new_n3923 = ~new_n3913 & new_n3922;
  assign new_n3924 = ~new_n3921 & new_n3923;
  assign new_n3925 = ~new_n3916 & ~new_n3920;
  assign new_n3926 = ~new_n3924 & new_n3925;
  assign new_n3927 = ~new_n3912 & new_n3926;
  assign new_n3928 = ~A262 & new_n3915;
  assign new_n3929 = ~new_n3900 & ~new_n3905;
  assign new_n3930 = ~new_n3914 & new_n3929;
  assign new_n3931 = new_n3901 & ~new_n3930;
  assign new_n3932 = ~new_n3898 & ~new_n3906;
  assign new_n3933 = ~new_n3931 & new_n3932;
  assign new_n3934 = ~new_n3928 & ~new_n3933;
  assign new_n3935 = new_n3891 & ~new_n3934;
  assign new_n3936 = new_n3927 & ~new_n3935;
  assign new_n3937 = ~new_n3877 & ~new_n3886;
  assign new_n3938 = A268 & new_n3886;
  assign new_n3939 = ~new_n3937 & ~new_n3938;
  assign new_n3940 = new_n3879 & ~new_n3887;
  assign new_n3941 = ~new_n3939 & ~new_n3940;
  assign new_n3942 = new_n3880 & new_n3941;
  assign new_n3943 = ~new_n3878 & ~new_n3880;
  assign new_n3944 = ~new_n3887 & new_n3943;
  assign new_n3945 = ~new_n3937 & new_n3944;
  assign new_n3946 = ~new_n3881 & new_n3945;
  assign new_n3947 = new_n3886 & new_n3942;
  assign new_n3948 = new_n3881 & ~new_n3941;
  assign new_n3949 = ~new_n3947 & ~new_n3948;
  assign new_n3950 = new_n3878 & ~new_n3881;
  assign new_n3951 = new_n3887 & new_n3950;
  assign new_n3952 = ~new_n3942 & ~new_n3951;
  assign new_n3953 = ~new_n3946 & new_n3952;
  assign new_n3954 = new_n3949 & new_n3953;
  assign new_n3955 = new_n3936 & ~new_n3954;
  assign new_n3956 = new_n3927 & ~new_n3955;
  assign new_n3957 = ~new_n3917 & ~new_n3919;
  assign new_n3958 = ~new_n3945 & new_n3949;
  assign new_n3959 = new_n3957 & new_n3958;
  assign new_n3960 = ~new_n3957 & ~new_n3958;
  assign new_n3961 = ~new_n3959 & ~new_n3960;
  assign new_n3962 = ~new_n3956 & new_n3961;
  assign new_n3963 = new_n3956 & ~new_n3961;
  assign new_n3964 = ~new_n3962 & ~new_n3963;
  assign new_n3965 = ~A254 & ~A255;
  assign new_n3966 = A254 & A255;
  assign new_n3967 = ~new_n3965 & ~new_n3966;
  assign new_n3968 = ~A253 & new_n3967;
  assign new_n3969 = A253 & ~new_n3967;
  assign new_n3970 = ~new_n3968 & ~new_n3969;
  assign new_n3971 = A258 & ~new_n3970;
  assign new_n3972 = ~A258 & new_n3970;
  assign new_n3973 = ~new_n3971 & ~new_n3972;
  assign new_n3974 = A256 & A257;
  assign new_n3975 = ~A256 & ~A257;
  assign new_n3976 = ~new_n3974 & ~new_n3975;
  assign new_n3977 = new_n3973 & new_n3976;
  assign new_n3978 = ~new_n3973 & ~new_n3976;
  assign new_n3979 = ~new_n3977 & ~new_n3978;
  assign new_n3980 = A250 & A251;
  assign new_n3981 = ~A250 & ~A251;
  assign new_n3982 = ~new_n3980 & ~new_n3981;
  assign new_n3983 = A247 & A248;
  assign new_n3984 = ~A247 & ~A248;
  assign new_n3985 = ~new_n3983 & ~new_n3984;
  assign new_n3986 = ~A249 & A252;
  assign new_n3987 = A249 & ~A252;
  assign new_n3988 = ~new_n3986 & ~new_n3987;
  assign new_n3989 = new_n3985 & ~new_n3988;
  assign new_n3990 = ~new_n3985 & new_n3988;
  assign new_n3991 = ~new_n3989 & ~new_n3990;
  assign new_n3992 = new_n3982 & new_n3991;
  assign new_n3993 = ~new_n3982 & ~new_n3991;
  assign new_n3994 = ~new_n3992 & ~new_n3993;
  assign new_n3995 = new_n3979 & new_n3994;
  assign new_n3996 = ~new_n3965 & ~new_n3968;
  assign new_n3997 = new_n3974 & new_n3996;
  assign new_n3998 = ~new_n3969 & new_n3997;
  assign new_n3999 = ~new_n3974 & ~new_n3996;
  assign new_n4000 = new_n3971 & ~new_n3997;
  assign new_n4001 = ~new_n3999 & new_n4000;
  assign new_n4002 = ~new_n3975 & new_n3996;
  assign new_n4003 = new_n3973 & new_n4002;
  assign new_n4004 = ~new_n4001 & ~new_n4003;
  assign new_n4005 = ~new_n3971 & new_n3999;
  assign new_n4006 = ~new_n3977 & new_n4005;
  assign new_n4007 = ~new_n3998 & new_n4004;
  assign new_n4008 = ~new_n4006 & new_n4007;
  assign new_n4009 = ~new_n3995 & ~new_n4008;
  assign new_n4010 = new_n3995 & new_n4008;
  assign new_n4011 = ~new_n4009 & ~new_n4010;
  assign new_n4012 = new_n3980 & new_n3986;
  assign new_n4013 = ~A249 & ~new_n3983;
  assign new_n4014 = A252 & ~new_n3982;
  assign new_n4015 = ~A252 & ~new_n3980;
  assign new_n4016 = ~new_n4013 & ~new_n4015;
  assign new_n4017 = ~new_n4014 & new_n4016;
  assign new_n4018 = ~new_n4012 & ~new_n4017;
  assign new_n4019 = ~new_n3984 & ~new_n4018;
  assign new_n4020 = A249 & A252;
  assign new_n4021 = ~new_n3980 & ~new_n3983;
  assign new_n4022 = new_n4020 & ~new_n4021;
  assign new_n4023 = A251 & new_n3983;
  assign new_n4024 = new_n4022 & ~new_n4023;
  assign new_n4025 = new_n3981 & new_n3984;
  assign new_n4026 = ~new_n4020 & new_n4025;
  assign new_n4027 = ~new_n3981 & new_n3983;
  assign new_n4028 = new_n3987 & new_n4027;
  assign new_n4029 = ~new_n4026 & ~new_n4028;
  assign new_n4030 = ~new_n4024 & new_n4029;
  assign new_n4031 = ~new_n4019 & new_n4030;
  assign new_n4032 = new_n4013 & new_n4015;
  assign new_n4033 = ~new_n3992 & new_n4032;
  assign new_n4034 = new_n4031 & ~new_n4033;
  assign new_n4035 = new_n4011 & ~new_n4034;
  assign new_n4036 = ~new_n4011 & new_n4034;
  assign new_n4037 = ~new_n4035 & ~new_n4036;
  assign new_n4038 = ~new_n3936 & new_n3954;
  assign new_n4039 = ~new_n3955 & ~new_n4038;
  assign new_n4040 = ~new_n4037 & ~new_n4039;
  assign new_n4041 = ~new_n3979 & ~new_n3994;
  assign new_n4042 = ~new_n3995 & ~new_n4041;
  assign new_n4043 = new_n3914 & ~new_n3929;
  assign new_n4044 = ~new_n3930 & ~new_n4043;
  assign new_n4045 = new_n3891 & new_n4044;
  assign new_n4046 = ~new_n3891 & ~new_n4044;
  assign new_n4047 = ~new_n4045 & ~new_n4046;
  assign new_n4048 = new_n4042 & ~new_n4047;
  assign new_n4049 = new_n4037 & new_n4039;
  assign new_n4050 = ~new_n4040 & ~new_n4049;
  assign new_n4051 = new_n4048 & new_n4050;
  assign new_n4052 = ~new_n4040 & ~new_n4051;
  assign new_n4053 = ~new_n3964 & ~new_n4052;
  assign new_n4054 = ~new_n4009 & ~new_n4035;
  assign new_n4055 = ~new_n3984 & ~new_n4031;
  assign new_n4056 = ~new_n4022 & ~new_n4055;
  assign new_n4057 = ~new_n3997 & new_n4004;
  assign new_n4058 = new_n4056 & new_n4057;
  assign new_n4059 = ~new_n4056 & ~new_n4057;
  assign new_n4060 = ~new_n4058 & ~new_n4059;
  assign new_n4061 = ~new_n4054 & new_n4060;
  assign new_n4062 = new_n4054 & ~new_n4060;
  assign new_n4063 = ~new_n4061 & ~new_n4062;
  assign new_n4064 = new_n3964 & new_n4052;
  assign new_n4065 = ~new_n4053 & ~new_n4064;
  assign new_n4066 = ~new_n4063 & new_n4065;
  assign new_n4067 = ~new_n4053 & ~new_n4066;
  assign new_n4068 = ~new_n4058 & ~new_n4061;
  assign new_n4069 = ~new_n3959 & ~new_n3962;
  assign new_n4070 = new_n4068 & new_n4069;
  assign new_n4071 = ~new_n4068 & ~new_n4069;
  assign new_n4072 = ~new_n4070 & ~new_n4071;
  assign new_n4073 = ~new_n4067 & new_n4072;
  assign new_n4074 = new_n4067 & ~new_n4072;
  assign new_n4075 = ~new_n4073 & ~new_n4074;
  assign new_n4076 = new_n4063 & ~new_n4065;
  assign new_n4077 = ~new_n4066 & ~new_n4076;
  assign new_n4078 = ~new_n3775 & new_n3808;
  assign new_n4079 = ~new_n3809 & ~new_n4078;
  assign new_n4080 = ~new_n4042 & new_n4047;
  assign new_n4081 = ~new_n4048 & ~new_n4080;
  assign new_n4082 = new_n4079 & new_n4081;
  assign new_n4083 = ~new_n4048 & ~new_n4082;
  assign new_n4084 = ~new_n4050 & new_n4083;
  assign new_n4085 = new_n3845 & ~new_n3849;
  assign new_n4086 = ~new_n3850 & ~new_n4085;
  assign new_n4087 = new_n4050 & ~new_n4083;
  assign new_n4088 = ~new_n4084 & ~new_n4087;
  assign new_n4089 = ~new_n4086 & new_n4088;
  assign new_n4090 = ~new_n4051 & ~new_n4084;
  assign new_n4091 = ~new_n4089 & new_n4090;
  assign new_n4092 = ~new_n4077 & ~new_n4091;
  assign new_n4093 = new_n3864 & ~new_n3866;
  assign new_n4094 = ~new_n3867 & ~new_n4093;
  assign new_n4095 = new_n4077 & new_n4091;
  assign new_n4096 = ~new_n4092 & ~new_n4095;
  assign new_n4097 = new_n4094 & new_n4096;
  assign new_n4098 = ~new_n4092 & ~new_n4097;
  assign new_n4099 = ~new_n4075 & ~new_n4098;
  assign new_n4100 = new_n4075 & new_n4098;
  assign new_n4101 = ~new_n4099 & ~new_n4100;
  assign new_n4102 = ~new_n3876 & new_n4101;
  assign new_n4103 = new_n3876 & ~new_n4101;
  assign new_n4104 = ~new_n4102 & ~new_n4103;
  assign new_n4105 = new_n3675 & ~new_n3677;
  assign new_n4106 = ~new_n3678 & ~new_n4105;
  assign new_n4107 = ~new_n4104 & new_n4106;
  assign new_n4108 = new_n4104 & ~new_n4106;
  assign new_n4109 = ~new_n4107 & ~new_n4108;
  assign new_n4110 = new_n3661 & ~new_n3663;
  assign new_n4111 = ~new_n3664 & ~new_n4110;
  assign new_n4112 = new_n4086 & ~new_n4088;
  assign new_n4113 = ~new_n4089 & ~new_n4112;
  assign new_n4114 = ~new_n3621 & ~new_n3627;
  assign new_n4115 = ~new_n4079 & ~new_n4081;
  assign new_n4116 = ~new_n4082 & ~new_n4115;
  assign new_n4117 = ~new_n3623 & ~new_n3625;
  assign new_n4118 = ~new_n3626 & ~new_n4117;
  assign new_n4119 = new_n4116 & new_n4118;
  assign new_n4120 = ~new_n3626 & ~new_n4119;
  assign new_n4121 = new_n4114 & new_n4120;
  assign new_n4122 = ~new_n4114 & ~new_n4120;
  assign new_n4123 = ~new_n4121 & ~new_n4122;
  assign new_n4124 = ~new_n4113 & ~new_n4123;
  assign new_n4125 = new_n4114 & new_n4119;
  assign new_n4126 = ~new_n4124 & ~new_n4125;
  assign new_n4127 = new_n4111 & ~new_n4126;
  assign new_n4128 = ~new_n4094 & ~new_n4096;
  assign new_n4129 = ~new_n4097 & ~new_n4128;
  assign new_n4130 = ~new_n4111 & new_n4126;
  assign new_n4131 = ~new_n4127 & ~new_n4130;
  assign new_n4132 = ~new_n4129 & new_n4131;
  assign new_n4133 = ~new_n4127 & ~new_n4132;
  assign new_n4134 = new_n4109 & ~new_n4133;
  assign new_n4135 = ~new_n4107 & ~new_n4134;
  assign new_n4136 = new_n3687 & new_n4135;
  assign new_n4137 = ~new_n3871 & ~new_n3874;
  assign new_n4138 = ~new_n4070 & ~new_n4073;
  assign new_n4139 = ~new_n4137 & ~new_n4138;
  assign new_n4140 = new_n4137 & new_n4138;
  assign new_n4141 = ~new_n4139 & ~new_n4140;
  assign new_n4142 = ~new_n4099 & ~new_n4102;
  assign new_n4143 = new_n4141 & new_n4142;
  assign new_n4144 = ~new_n4141 & ~new_n4142;
  assign new_n4145 = ~new_n4143 & ~new_n4144;
  assign new_n4146 = ~new_n3687 & ~new_n4135;
  assign new_n4147 = ~new_n4136 & ~new_n4146;
  assign new_n4148 = ~new_n4145 & new_n4147;
  assign new_n4149 = ~new_n4136 & ~new_n4148;
  assign new_n4150 = ~new_n4139 & ~new_n4143;
  assign new_n4151 = ~new_n3682 & ~new_n3685;
  assign new_n4152 = ~new_n4150 & new_n4151;
  assign new_n4153 = new_n4150 & ~new_n4151;
  assign new_n4154 = ~new_n4152 & ~new_n4153;
  assign new_n4155 = new_n4149 & new_n4154;
  assign new_n4156 = ~new_n4149 & ~new_n4154;
  assign new_n4157 = ~new_n4155 & ~new_n4156;
  assign new_n4158 = new_n4145 & ~new_n4147;
  assign new_n4159 = ~new_n4148 & ~new_n4158;
  assign new_n4160 = A97 & A98;
  assign new_n4161 = A100 & A101;
  assign new_n4162 = ~new_n4160 & ~new_n4161;
  assign new_n4163 = A99 & A102;
  assign new_n4164 = ~new_n4162 & new_n4163;
  assign new_n4165 = ~A97 & ~A98;
  assign new_n4166 = ~A99 & A102;
  assign new_n4167 = new_n4161 & new_n4166;
  assign new_n4168 = ~A99 & ~new_n4160;
  assign new_n4169 = ~A100 & ~A101;
  assign new_n4170 = ~new_n4161 & ~new_n4169;
  assign new_n4171 = A102 & ~new_n4170;
  assign new_n4172 = ~A102 & ~new_n4161;
  assign new_n4173 = ~new_n4168 & ~new_n4172;
  assign new_n4174 = ~new_n4171 & new_n4173;
  assign new_n4175 = ~new_n4167 & ~new_n4174;
  assign new_n4176 = ~new_n4165 & ~new_n4175;
  assign new_n4177 = A101 & new_n4160;
  assign new_n4178 = new_n4164 & ~new_n4177;
  assign new_n4179 = ~new_n4163 & new_n4165;
  assign new_n4180 = new_n4169 & new_n4179;
  assign new_n4181 = A99 & ~A102;
  assign new_n4182 = new_n4160 & ~new_n4169;
  assign new_n4183 = new_n4181 & new_n4182;
  assign new_n4184 = ~new_n4180 & ~new_n4183;
  assign new_n4185 = ~new_n4178 & new_n4184;
  assign new_n4186 = ~new_n4176 & new_n4185;
  assign new_n4187 = ~new_n4165 & ~new_n4186;
  assign new_n4188 = ~new_n4164 & ~new_n4187;
  assign new_n4189 = ~A95 & ~A96;
  assign new_n4190 = A95 & A96;
  assign new_n4191 = ~new_n4189 & ~new_n4190;
  assign new_n4192 = ~A94 & new_n4191;
  assign new_n4193 = ~new_n4189 & ~new_n4192;
  assign new_n4194 = ~A92 & ~A93;
  assign new_n4195 = A92 & A93;
  assign new_n4196 = ~new_n4194 & ~new_n4195;
  assign new_n4197 = ~A91 & new_n4196;
  assign new_n4198 = ~new_n4194 & ~new_n4197;
  assign new_n4199 = new_n4193 & new_n4198;
  assign new_n4200 = A91 & ~new_n4196;
  assign new_n4201 = ~new_n4197 & ~new_n4200;
  assign new_n4202 = A94 & ~new_n4191;
  assign new_n4203 = ~new_n4192 & ~new_n4202;
  assign new_n4204 = ~new_n4201 & ~new_n4203;
  assign new_n4205 = ~new_n4193 & ~new_n4198;
  assign new_n4206 = ~new_n4199 & ~new_n4205;
  assign new_n4207 = new_n4204 & new_n4206;
  assign new_n4208 = ~new_n4199 & ~new_n4207;
  assign new_n4209 = ~new_n4188 & ~new_n4208;
  assign new_n4210 = new_n4188 & new_n4208;
  assign new_n4211 = ~new_n4209 & ~new_n4210;
  assign new_n4212 = new_n4201 & new_n4203;
  assign new_n4213 = ~new_n4160 & ~new_n4165;
  assign new_n4214 = ~new_n4166 & ~new_n4181;
  assign new_n4215 = new_n4213 & ~new_n4214;
  assign new_n4216 = ~new_n4213 & new_n4214;
  assign new_n4217 = ~new_n4215 & ~new_n4216;
  assign new_n4218 = new_n4170 & new_n4217;
  assign new_n4219 = ~new_n4170 & ~new_n4217;
  assign new_n4220 = ~new_n4218 & ~new_n4219;
  assign new_n4221 = ~new_n4204 & ~new_n4212;
  assign new_n4222 = ~new_n4220 & new_n4221;
  assign new_n4223 = ~new_n4212 & ~new_n4222;
  assign new_n4224 = new_n4168 & new_n4172;
  assign new_n4225 = ~new_n4218 & new_n4224;
  assign new_n4226 = new_n4186 & ~new_n4225;
  assign new_n4227 = ~new_n4223 & ~new_n4226;
  assign new_n4228 = new_n4223 & new_n4226;
  assign new_n4229 = ~new_n4227 & ~new_n4228;
  assign new_n4230 = ~new_n4206 & new_n4229;
  assign new_n4231 = ~new_n4207 & ~new_n4227;
  assign new_n4232 = ~new_n4230 & new_n4231;
  assign new_n4233 = new_n4211 & new_n4232;
  assign new_n4234 = ~new_n4209 & ~new_n4233;
  assign new_n4235 = A89 & A90;
  assign new_n4236 = A86 & A87;
  assign new_n4237 = ~A86 & ~A87;
  assign new_n4238 = ~new_n4236 & ~new_n4237;
  assign new_n4239 = A85 & new_n4238;
  assign new_n4240 = ~new_n4236 & ~new_n4239;
  assign new_n4241 = new_n4235 & ~new_n4240;
  assign new_n4242 = ~A89 & ~A90;
  assign new_n4243 = ~A85 & ~A86;
  assign new_n4244 = ~new_n4242 & ~new_n4243;
  assign new_n4245 = ~new_n4235 & ~new_n4242;
  assign new_n4246 = A88 & ~new_n4245;
  assign new_n4247 = ~A87 & new_n4244;
  assign new_n4248 = new_n4246 & new_n4247;
  assign new_n4249 = A85 & A86;
  assign new_n4250 = A90 & new_n4249;
  assign new_n4251 = ~new_n4235 & ~new_n4249;
  assign new_n4252 = A87 & A88;
  assign new_n4253 = ~new_n4250 & new_n4252;
  assign new_n4254 = ~new_n4251 & new_n4253;
  assign new_n4255 = ~A85 & ~new_n4238;
  assign new_n4256 = ~new_n4239 & ~new_n4255;
  assign new_n4257 = ~A88 & new_n4245;
  assign new_n4258 = ~new_n4246 & ~new_n4257;
  assign new_n4259 = ~new_n4256 & ~new_n4258;
  assign new_n4260 = ~new_n4240 & new_n4245;
  assign new_n4261 = ~new_n4259 & new_n4260;
  assign new_n4262 = ~new_n4248 & ~new_n4254;
  assign new_n4263 = ~new_n4261 & new_n4262;
  assign new_n4264 = ~new_n4241 & new_n4263;
  assign new_n4265 = ~A83 & ~A84;
  assign new_n4266 = A83 & A84;
  assign new_n4267 = ~new_n4265 & ~new_n4266;
  assign new_n4268 = ~A82 & new_n4267;
  assign new_n4269 = ~new_n4265 & ~new_n4268;
  assign new_n4270 = ~A80 & ~A81;
  assign new_n4271 = A80 & A81;
  assign new_n4272 = ~new_n4270 & ~new_n4271;
  assign new_n4273 = ~A79 & new_n4272;
  assign new_n4274 = ~new_n4270 & ~new_n4273;
  assign new_n4275 = new_n4269 & new_n4274;
  assign new_n4276 = A79 & ~new_n4272;
  assign new_n4277 = ~new_n4273 & ~new_n4276;
  assign new_n4278 = A82 & ~new_n4267;
  assign new_n4279 = ~new_n4268 & ~new_n4278;
  assign new_n4280 = ~new_n4277 & ~new_n4279;
  assign new_n4281 = ~new_n4269 & ~new_n4274;
  assign new_n4282 = ~new_n4275 & ~new_n4281;
  assign new_n4283 = new_n4280 & new_n4282;
  assign new_n4284 = ~new_n4275 & ~new_n4283;
  assign new_n4285 = new_n4264 & new_n4284;
  assign new_n4286 = ~new_n4264 & ~new_n4284;
  assign new_n4287 = ~new_n4285 & ~new_n4286;
  assign new_n4288 = new_n4242 & new_n4243;
  assign new_n4289 = ~new_n4252 & new_n4288;
  assign new_n4290 = ~A87 & ~new_n4244;
  assign new_n4291 = new_n4251 & new_n4290;
  assign new_n4292 = ~new_n4241 & ~new_n4291;
  assign new_n4293 = ~A88 & ~new_n4292;
  assign new_n4294 = new_n4263 & ~new_n4289;
  assign new_n4295 = ~new_n4293 & new_n4294;
  assign new_n4296 = ~new_n4282 & ~new_n4295;
  assign new_n4297 = new_n4256 & new_n4258;
  assign new_n4298 = ~new_n4259 & ~new_n4297;
  assign new_n4299 = new_n4277 & new_n4279;
  assign new_n4300 = ~new_n4280 & ~new_n4299;
  assign new_n4301 = ~new_n4298 & new_n4300;
  assign new_n4302 = ~new_n4280 & ~new_n4301;
  assign new_n4303 = new_n4282 & new_n4295;
  assign new_n4304 = ~new_n4296 & ~new_n4303;
  assign new_n4305 = new_n4302 & new_n4304;
  assign new_n4306 = ~new_n4283 & ~new_n4296;
  assign new_n4307 = ~new_n4305 & new_n4306;
  assign new_n4308 = new_n4287 & ~new_n4307;
  assign new_n4309 = ~new_n4285 & ~new_n4308;
  assign new_n4310 = ~new_n4234 & new_n4309;
  assign new_n4311 = new_n4234 & ~new_n4309;
  assign new_n4312 = ~new_n4310 & ~new_n4311;
  assign new_n4313 = ~new_n4287 & new_n4307;
  assign new_n4314 = ~new_n4308 & ~new_n4313;
  assign new_n4315 = new_n4206 & ~new_n4229;
  assign new_n4316 = ~new_n4230 & ~new_n4315;
  assign new_n4317 = ~new_n4302 & ~new_n4304;
  assign new_n4318 = ~new_n4305 & ~new_n4317;
  assign new_n4319 = ~new_n4316 & ~new_n4318;
  assign new_n4320 = new_n4316 & new_n4318;
  assign new_n4321 = new_n4220 & ~new_n4221;
  assign new_n4322 = ~new_n4222 & ~new_n4321;
  assign new_n4323 = new_n4298 & ~new_n4300;
  assign new_n4324 = ~new_n4301 & ~new_n4323;
  assign new_n4325 = ~new_n4322 & new_n4324;
  assign new_n4326 = ~new_n4320 & new_n4325;
  assign new_n4327 = ~new_n4319 & ~new_n4326;
  assign new_n4328 = new_n4314 & new_n4327;
  assign new_n4329 = ~new_n4211 & ~new_n4232;
  assign new_n4330 = ~new_n4233 & ~new_n4329;
  assign new_n4331 = ~new_n4314 & ~new_n4327;
  assign new_n4332 = ~new_n4328 & ~new_n4331;
  assign new_n4333 = ~new_n4330 & new_n4332;
  assign new_n4334 = ~new_n4328 & ~new_n4333;
  assign new_n4335 = new_n4312 & new_n4334;
  assign new_n4336 = ~new_n4310 & ~new_n4335;
  assign new_n4337 = ~A119 & ~A120;
  assign new_n4338 = A119 & A120;
  assign new_n4339 = ~new_n4337 & ~new_n4338;
  assign new_n4340 = ~A118 & new_n4339;
  assign new_n4341 = ~new_n4337 & ~new_n4340;
  assign new_n4342 = ~A115 & ~A117;
  assign new_n4343 = A115 & A117;
  assign new_n4344 = ~new_n4342 & ~new_n4343;
  assign new_n4345 = ~A116 & new_n4344;
  assign new_n4346 = ~new_n4342 & ~new_n4345;
  assign new_n4347 = new_n4341 & new_n4346;
  assign new_n4348 = A116 & ~new_n4344;
  assign new_n4349 = ~new_n4345 & ~new_n4348;
  assign new_n4350 = A118 & ~new_n4339;
  assign new_n4351 = ~new_n4340 & ~new_n4350;
  assign new_n4352 = ~new_n4349 & ~new_n4351;
  assign new_n4353 = ~new_n4341 & ~new_n4346;
  assign new_n4354 = ~new_n4347 & ~new_n4353;
  assign new_n4355 = new_n4352 & new_n4354;
  assign new_n4356 = ~new_n4347 & ~new_n4355;
  assign new_n4357 = ~A125 & ~A126;
  assign new_n4358 = A121 & A122;
  assign new_n4359 = A123 & A124;
  assign new_n4360 = ~new_n4358 & ~new_n4359;
  assign new_n4361 = ~A121 & ~A122;
  assign new_n4362 = ~A123 & ~A124;
  assign new_n4363 = ~new_n4361 & ~new_n4362;
  assign new_n4364 = ~new_n4357 & ~new_n4360;
  assign new_n4365 = new_n4363 & new_n4364;
  assign new_n4366 = new_n4360 & ~new_n4363;
  assign new_n4367 = new_n4358 & new_n4359;
  assign new_n4368 = ~new_n4366 & ~new_n4367;
  assign new_n4369 = ~new_n4357 & ~new_n4368;
  assign new_n4370 = A125 & A126;
  assign new_n4371 = ~new_n4367 & ~new_n4370;
  assign new_n4372 = ~new_n4369 & ~new_n4371;
  assign new_n4373 = ~new_n4365 & ~new_n4372;
  assign new_n4374 = ~new_n4356 & ~new_n4373;
  assign new_n4375 = new_n4356 & new_n4373;
  assign new_n4376 = ~new_n4374 & ~new_n4375;
  assign new_n4377 = new_n4361 & new_n4362;
  assign new_n4378 = ~new_n4365 & ~new_n4377;
  assign new_n4379 = ~new_n4370 & ~new_n4378;
  assign new_n4380 = new_n4357 & ~new_n4368;
  assign new_n4381 = ~new_n4372 & ~new_n4380;
  assign new_n4382 = ~new_n4379 & new_n4381;
  assign new_n4383 = ~new_n4354 & ~new_n4382;
  assign new_n4384 = new_n4349 & new_n4351;
  assign new_n4385 = ~new_n4352 & ~new_n4384;
  assign new_n4386 = ~new_n4357 & ~new_n4370;
  assign new_n4387 = ~new_n4359 & ~new_n4362;
  assign new_n4388 = ~new_n4386 & new_n4387;
  assign new_n4389 = new_n4386 & ~new_n4387;
  assign new_n4390 = ~new_n4388 & ~new_n4389;
  assign new_n4391 = ~new_n4358 & ~new_n4361;
  assign new_n4392 = ~new_n4390 & new_n4391;
  assign new_n4393 = new_n4390 & ~new_n4391;
  assign new_n4394 = ~new_n4392 & ~new_n4393;
  assign new_n4395 = new_n4385 & ~new_n4394;
  assign new_n4396 = ~new_n4384 & ~new_n4395;
  assign new_n4397 = new_n4354 & new_n4382;
  assign new_n4398 = ~new_n4383 & ~new_n4397;
  assign new_n4399 = ~new_n4396 & new_n4398;
  assign new_n4400 = ~new_n4355 & ~new_n4383;
  assign new_n4401 = ~new_n4399 & new_n4400;
  assign new_n4402 = new_n4376 & new_n4401;
  assign new_n4403 = ~new_n4374 & ~new_n4402;
  assign new_n4404 = A113 & A114;
  assign new_n4405 = A110 & A111;
  assign new_n4406 = ~A110 & ~A111;
  assign new_n4407 = ~new_n4405 & ~new_n4406;
  assign new_n4408 = A109 & new_n4407;
  assign new_n4409 = ~new_n4405 & ~new_n4408;
  assign new_n4410 = new_n4404 & ~new_n4409;
  assign new_n4411 = ~A113 & ~A114;
  assign new_n4412 = ~A109 & ~A110;
  assign new_n4413 = ~new_n4411 & ~new_n4412;
  assign new_n4414 = ~new_n4404 & ~new_n4411;
  assign new_n4415 = A112 & ~new_n4414;
  assign new_n4416 = ~A111 & new_n4413;
  assign new_n4417 = new_n4415 & new_n4416;
  assign new_n4418 = A109 & A110;
  assign new_n4419 = A114 & new_n4418;
  assign new_n4420 = ~new_n4404 & ~new_n4418;
  assign new_n4421 = A111 & A112;
  assign new_n4422 = ~new_n4419 & new_n4421;
  assign new_n4423 = ~new_n4420 & new_n4422;
  assign new_n4424 = ~A109 & ~new_n4407;
  assign new_n4425 = ~new_n4408 & ~new_n4424;
  assign new_n4426 = ~A112 & new_n4414;
  assign new_n4427 = ~new_n4415 & ~new_n4426;
  assign new_n4428 = ~new_n4425 & ~new_n4427;
  assign new_n4429 = ~new_n4409 & new_n4414;
  assign new_n4430 = ~new_n4428 & new_n4429;
  assign new_n4431 = ~new_n4417 & ~new_n4423;
  assign new_n4432 = ~new_n4430 & new_n4431;
  assign new_n4433 = ~new_n4410 & new_n4432;
  assign new_n4434 = ~A104 & ~A105;
  assign new_n4435 = A104 & A105;
  assign new_n4436 = ~new_n4434 & ~new_n4435;
  assign new_n4437 = ~A103 & new_n4436;
  assign new_n4438 = ~new_n4434 & ~new_n4437;
  assign new_n4439 = ~A107 & ~A108;
  assign new_n4440 = A107 & A108;
  assign new_n4441 = ~new_n4439 & ~new_n4440;
  assign new_n4442 = ~A106 & new_n4441;
  assign new_n4443 = ~new_n4439 & ~new_n4442;
  assign new_n4444 = new_n4438 & new_n4443;
  assign new_n4445 = A103 & ~new_n4436;
  assign new_n4446 = ~new_n4437 & ~new_n4445;
  assign new_n4447 = A106 & ~new_n4441;
  assign new_n4448 = ~new_n4442 & ~new_n4447;
  assign new_n4449 = ~new_n4446 & ~new_n4448;
  assign new_n4450 = ~new_n4438 & ~new_n4443;
  assign new_n4451 = ~new_n4444 & ~new_n4450;
  assign new_n4452 = new_n4449 & new_n4451;
  assign new_n4453 = ~new_n4444 & ~new_n4452;
  assign new_n4454 = new_n4433 & new_n4453;
  assign new_n4455 = ~new_n4433 & ~new_n4453;
  assign new_n4456 = ~new_n4454 & ~new_n4455;
  assign new_n4457 = new_n4411 & new_n4412;
  assign new_n4458 = ~new_n4421 & new_n4457;
  assign new_n4459 = ~A111 & ~new_n4413;
  assign new_n4460 = new_n4420 & new_n4459;
  assign new_n4461 = ~new_n4410 & ~new_n4460;
  assign new_n4462 = ~A112 & ~new_n4461;
  assign new_n4463 = new_n4432 & ~new_n4458;
  assign new_n4464 = ~new_n4462 & new_n4463;
  assign new_n4465 = ~new_n4451 & ~new_n4464;
  assign new_n4466 = new_n4425 & new_n4427;
  assign new_n4467 = ~new_n4428 & ~new_n4466;
  assign new_n4468 = new_n4446 & new_n4448;
  assign new_n4469 = ~new_n4449 & ~new_n4468;
  assign new_n4470 = ~new_n4467 & new_n4469;
  assign new_n4471 = ~new_n4449 & ~new_n4470;
  assign new_n4472 = new_n4451 & new_n4464;
  assign new_n4473 = ~new_n4465 & ~new_n4472;
  assign new_n4474 = new_n4471 & new_n4473;
  assign new_n4475 = ~new_n4452 & ~new_n4465;
  assign new_n4476 = ~new_n4474 & new_n4475;
  assign new_n4477 = new_n4456 & ~new_n4476;
  assign new_n4478 = ~new_n4454 & ~new_n4477;
  assign new_n4479 = ~new_n4403 & new_n4478;
  assign new_n4480 = new_n4403 & ~new_n4478;
  assign new_n4481 = ~new_n4479 & ~new_n4480;
  assign new_n4482 = ~new_n4385 & new_n4394;
  assign new_n4483 = ~new_n4395 & ~new_n4482;
  assign new_n4484 = new_n4467 & ~new_n4469;
  assign new_n4485 = ~new_n4470 & ~new_n4484;
  assign new_n4486 = ~new_n4483 & new_n4485;
  assign new_n4487 = ~new_n4471 & ~new_n4473;
  assign new_n4488 = ~new_n4474 & ~new_n4487;
  assign new_n4489 = new_n4486 & ~new_n4488;
  assign new_n4490 = new_n4396 & ~new_n4398;
  assign new_n4491 = ~new_n4399 & ~new_n4490;
  assign new_n4492 = ~new_n4486 & new_n4488;
  assign new_n4493 = ~new_n4489 & ~new_n4492;
  assign new_n4494 = ~new_n4491 & new_n4493;
  assign new_n4495 = ~new_n4489 & ~new_n4494;
  assign new_n4496 = ~new_n4456 & new_n4476;
  assign new_n4497 = ~new_n4477 & ~new_n4496;
  assign new_n4498 = ~new_n4495 & ~new_n4497;
  assign new_n4499 = ~new_n4376 & ~new_n4401;
  assign new_n4500 = ~new_n4402 & ~new_n4499;
  assign new_n4501 = new_n4495 & new_n4497;
  assign new_n4502 = ~new_n4498 & ~new_n4501;
  assign new_n4503 = new_n4500 & new_n4502;
  assign new_n4504 = ~new_n4498 & ~new_n4503;
  assign new_n4505 = new_n4481 & ~new_n4504;
  assign new_n4506 = ~new_n4479 & ~new_n4505;
  assign new_n4507 = new_n4336 & new_n4506;
  assign new_n4508 = ~new_n4336 & ~new_n4506;
  assign new_n4509 = ~new_n4507 & ~new_n4508;
  assign new_n4510 = ~new_n4481 & new_n4504;
  assign new_n4511 = ~new_n4505 & ~new_n4510;
  assign new_n4512 = new_n4491 & ~new_n4493;
  assign new_n4513 = ~new_n4494 & ~new_n4512;
  assign new_n4514 = ~new_n4319 & ~new_n4320;
  assign new_n4515 = new_n4483 & ~new_n4485;
  assign new_n4516 = ~new_n4486 & ~new_n4515;
  assign new_n4517 = new_n4322 & ~new_n4324;
  assign new_n4518 = ~new_n4325 & ~new_n4517;
  assign new_n4519 = new_n4516 & new_n4518;
  assign new_n4520 = ~new_n4325 & ~new_n4519;
  assign new_n4521 = new_n4514 & ~new_n4520;
  assign new_n4522 = ~new_n4514 & new_n4520;
  assign new_n4523 = ~new_n4521 & ~new_n4522;
  assign new_n4524 = new_n4513 & new_n4523;
  assign new_n4525 = new_n4514 & new_n4519;
  assign new_n4526 = ~new_n4524 & ~new_n4525;
  assign new_n4527 = ~new_n4500 & ~new_n4502;
  assign new_n4528 = ~new_n4503 & ~new_n4527;
  assign new_n4529 = ~new_n4526 & new_n4528;
  assign new_n4530 = new_n4330 & ~new_n4332;
  assign new_n4531 = ~new_n4333 & ~new_n4530;
  assign new_n4532 = new_n4526 & ~new_n4528;
  assign new_n4533 = ~new_n4529 & ~new_n4532;
  assign new_n4534 = ~new_n4531 & new_n4533;
  assign new_n4535 = ~new_n4529 & ~new_n4534;
  assign new_n4536 = new_n4511 & ~new_n4535;
  assign new_n4537 = ~new_n4312 & ~new_n4334;
  assign new_n4538 = ~new_n4335 & ~new_n4537;
  assign new_n4539 = ~new_n4511 & new_n4535;
  assign new_n4540 = ~new_n4536 & ~new_n4539;
  assign new_n4541 = new_n4538 & new_n4540;
  assign new_n4542 = ~new_n4536 & ~new_n4541;
  assign new_n4543 = new_n4509 & new_n4542;
  assign new_n4544 = ~new_n4509 & ~new_n4542;
  assign new_n4545 = ~new_n4543 & ~new_n4544;
  assign new_n4546 = A157 & A158;
  assign new_n4547 = A160 & A161;
  assign new_n4548 = ~new_n4546 & ~new_n4547;
  assign new_n4549 = A159 & A162;
  assign new_n4550 = ~new_n4548 & new_n4549;
  assign new_n4551 = ~A157 & ~A158;
  assign new_n4552 = ~A159 & A162;
  assign new_n4553 = new_n4547 & new_n4552;
  assign new_n4554 = ~A159 & ~new_n4546;
  assign new_n4555 = ~A160 & ~A161;
  assign new_n4556 = ~new_n4547 & ~new_n4555;
  assign new_n4557 = A162 & ~new_n4556;
  assign new_n4558 = ~A162 & ~new_n4547;
  assign new_n4559 = ~new_n4554 & ~new_n4558;
  assign new_n4560 = ~new_n4557 & new_n4559;
  assign new_n4561 = ~new_n4553 & ~new_n4560;
  assign new_n4562 = ~new_n4551 & ~new_n4561;
  assign new_n4563 = A161 & new_n4546;
  assign new_n4564 = new_n4550 & ~new_n4563;
  assign new_n4565 = ~new_n4549 & new_n4551;
  assign new_n4566 = new_n4555 & new_n4565;
  assign new_n4567 = A159 & ~A162;
  assign new_n4568 = new_n4546 & ~new_n4555;
  assign new_n4569 = new_n4567 & new_n4568;
  assign new_n4570 = ~new_n4566 & ~new_n4569;
  assign new_n4571 = ~new_n4564 & new_n4570;
  assign new_n4572 = ~new_n4562 & new_n4571;
  assign new_n4573 = ~new_n4551 & ~new_n4572;
  assign new_n4574 = ~new_n4550 & ~new_n4573;
  assign new_n4575 = ~A155 & ~A156;
  assign new_n4576 = A155 & A156;
  assign new_n4577 = ~new_n4575 & ~new_n4576;
  assign new_n4578 = ~A154 & new_n4577;
  assign new_n4579 = ~new_n4575 & ~new_n4578;
  assign new_n4580 = ~A152 & ~A153;
  assign new_n4581 = A152 & A153;
  assign new_n4582 = ~new_n4580 & ~new_n4581;
  assign new_n4583 = ~A151 & new_n4582;
  assign new_n4584 = ~new_n4580 & ~new_n4583;
  assign new_n4585 = new_n4579 & new_n4584;
  assign new_n4586 = A151 & ~new_n4582;
  assign new_n4587 = ~new_n4583 & ~new_n4586;
  assign new_n4588 = A154 & ~new_n4577;
  assign new_n4589 = ~new_n4578 & ~new_n4588;
  assign new_n4590 = ~new_n4587 & ~new_n4589;
  assign new_n4591 = ~new_n4579 & ~new_n4584;
  assign new_n4592 = ~new_n4585 & ~new_n4591;
  assign new_n4593 = new_n4590 & new_n4592;
  assign new_n4594 = ~new_n4585 & ~new_n4593;
  assign new_n4595 = ~new_n4574 & ~new_n4594;
  assign new_n4596 = new_n4574 & new_n4594;
  assign new_n4597 = ~new_n4595 & ~new_n4596;
  assign new_n4598 = new_n4587 & new_n4589;
  assign new_n4599 = ~new_n4546 & ~new_n4551;
  assign new_n4600 = ~new_n4552 & ~new_n4567;
  assign new_n4601 = new_n4599 & ~new_n4600;
  assign new_n4602 = ~new_n4599 & new_n4600;
  assign new_n4603 = ~new_n4601 & ~new_n4602;
  assign new_n4604 = new_n4556 & new_n4603;
  assign new_n4605 = ~new_n4556 & ~new_n4603;
  assign new_n4606 = ~new_n4604 & ~new_n4605;
  assign new_n4607 = ~new_n4590 & ~new_n4598;
  assign new_n4608 = ~new_n4606 & new_n4607;
  assign new_n4609 = ~new_n4598 & ~new_n4608;
  assign new_n4610 = new_n4554 & new_n4558;
  assign new_n4611 = ~new_n4604 & new_n4610;
  assign new_n4612 = new_n4572 & ~new_n4611;
  assign new_n4613 = ~new_n4609 & ~new_n4612;
  assign new_n4614 = new_n4609 & new_n4612;
  assign new_n4615 = ~new_n4613 & ~new_n4614;
  assign new_n4616 = ~new_n4592 & new_n4615;
  assign new_n4617 = ~new_n4593 & ~new_n4613;
  assign new_n4618 = ~new_n4616 & new_n4617;
  assign new_n4619 = new_n4597 & new_n4618;
  assign new_n4620 = ~new_n4595 & ~new_n4619;
  assign new_n4621 = A173 & A174;
  assign new_n4622 = A170 & A171;
  assign new_n4623 = ~A170 & ~A171;
  assign new_n4624 = ~new_n4622 & ~new_n4623;
  assign new_n4625 = A169 & new_n4624;
  assign new_n4626 = ~new_n4622 & ~new_n4625;
  assign new_n4627 = new_n4621 & ~new_n4626;
  assign new_n4628 = ~A173 & ~A174;
  assign new_n4629 = ~A169 & ~A170;
  assign new_n4630 = ~new_n4628 & ~new_n4629;
  assign new_n4631 = ~new_n4621 & ~new_n4628;
  assign new_n4632 = A172 & ~new_n4631;
  assign new_n4633 = ~A171 & new_n4630;
  assign new_n4634 = new_n4632 & new_n4633;
  assign new_n4635 = A169 & A170;
  assign new_n4636 = A174 & new_n4635;
  assign new_n4637 = ~new_n4621 & ~new_n4635;
  assign new_n4638 = A171 & A172;
  assign new_n4639 = ~new_n4636 & new_n4638;
  assign new_n4640 = ~new_n4637 & new_n4639;
  assign new_n4641 = ~A169 & ~new_n4624;
  assign new_n4642 = ~new_n4625 & ~new_n4641;
  assign new_n4643 = ~A172 & new_n4631;
  assign new_n4644 = ~new_n4632 & ~new_n4643;
  assign new_n4645 = ~new_n4642 & ~new_n4644;
  assign new_n4646 = ~new_n4626 & new_n4631;
  assign new_n4647 = ~new_n4645 & new_n4646;
  assign new_n4648 = ~new_n4634 & ~new_n4640;
  assign new_n4649 = ~new_n4647 & new_n4648;
  assign new_n4650 = ~new_n4627 & new_n4649;
  assign new_n4651 = ~A167 & ~A168;
  assign new_n4652 = A167 & A168;
  assign new_n4653 = ~new_n4651 & ~new_n4652;
  assign new_n4654 = ~A166 & new_n4653;
  assign new_n4655 = ~new_n4651 & ~new_n4654;
  assign new_n4656 = ~A164 & ~A165;
  assign new_n4657 = A164 & A165;
  assign new_n4658 = ~new_n4656 & ~new_n4657;
  assign new_n4659 = ~A163 & new_n4658;
  assign new_n4660 = ~new_n4656 & ~new_n4659;
  assign new_n4661 = new_n4655 & new_n4660;
  assign new_n4662 = A163 & ~new_n4658;
  assign new_n4663 = ~new_n4659 & ~new_n4662;
  assign new_n4664 = A166 & ~new_n4653;
  assign new_n4665 = ~new_n4654 & ~new_n4664;
  assign new_n4666 = ~new_n4663 & ~new_n4665;
  assign new_n4667 = ~new_n4655 & ~new_n4660;
  assign new_n4668 = ~new_n4661 & ~new_n4667;
  assign new_n4669 = new_n4666 & new_n4668;
  assign new_n4670 = ~new_n4661 & ~new_n4669;
  assign new_n4671 = new_n4650 & new_n4670;
  assign new_n4672 = ~new_n4650 & ~new_n4670;
  assign new_n4673 = ~new_n4671 & ~new_n4672;
  assign new_n4674 = new_n4628 & new_n4629;
  assign new_n4675 = ~new_n4638 & new_n4674;
  assign new_n4676 = ~A171 & ~new_n4630;
  assign new_n4677 = new_n4637 & new_n4676;
  assign new_n4678 = ~new_n4627 & ~new_n4677;
  assign new_n4679 = ~A172 & ~new_n4678;
  assign new_n4680 = new_n4649 & ~new_n4675;
  assign new_n4681 = ~new_n4679 & new_n4680;
  assign new_n4682 = ~new_n4668 & ~new_n4681;
  assign new_n4683 = new_n4642 & new_n4644;
  assign new_n4684 = ~new_n4645 & ~new_n4683;
  assign new_n4685 = new_n4663 & new_n4665;
  assign new_n4686 = ~new_n4666 & ~new_n4685;
  assign new_n4687 = ~new_n4684 & new_n4686;
  assign new_n4688 = ~new_n4666 & ~new_n4687;
  assign new_n4689 = new_n4668 & new_n4681;
  assign new_n4690 = ~new_n4682 & ~new_n4689;
  assign new_n4691 = new_n4688 & new_n4690;
  assign new_n4692 = ~new_n4669 & ~new_n4682;
  assign new_n4693 = ~new_n4691 & new_n4692;
  assign new_n4694 = new_n4673 & ~new_n4693;
  assign new_n4695 = ~new_n4671 & ~new_n4694;
  assign new_n4696 = ~new_n4620 & new_n4695;
  assign new_n4697 = new_n4620 & ~new_n4695;
  assign new_n4698 = ~new_n4696 & ~new_n4697;
  assign new_n4699 = ~new_n4688 & ~new_n4690;
  assign new_n4700 = ~new_n4691 & ~new_n4699;
  assign new_n4701 = new_n4606 & ~new_n4607;
  assign new_n4702 = ~new_n4608 & ~new_n4701;
  assign new_n4703 = new_n4684 & ~new_n4686;
  assign new_n4704 = ~new_n4687 & ~new_n4703;
  assign new_n4705 = ~new_n4702 & new_n4704;
  assign new_n4706 = ~new_n4700 & new_n4705;
  assign new_n4707 = new_n4592 & ~new_n4615;
  assign new_n4708 = ~new_n4616 & ~new_n4707;
  assign new_n4709 = new_n4700 & ~new_n4705;
  assign new_n4710 = ~new_n4706 & ~new_n4709;
  assign new_n4711 = ~new_n4708 & new_n4710;
  assign new_n4712 = ~new_n4706 & ~new_n4711;
  assign new_n4713 = ~new_n4673 & new_n4693;
  assign new_n4714 = ~new_n4694 & ~new_n4713;
  assign new_n4715 = new_n4712 & new_n4714;
  assign new_n4716 = ~new_n4597 & ~new_n4618;
  assign new_n4717 = ~new_n4619 & ~new_n4716;
  assign new_n4718 = ~new_n4712 & ~new_n4714;
  assign new_n4719 = ~new_n4715 & ~new_n4718;
  assign new_n4720 = ~new_n4717 & new_n4719;
  assign new_n4721 = ~new_n4715 & ~new_n4720;
  assign new_n4722 = new_n4698 & new_n4721;
  assign new_n4723 = ~new_n4696 & ~new_n4722;
  assign new_n4724 = ~A131 & ~A132;
  assign new_n4725 = A131 & A132;
  assign new_n4726 = ~new_n4724 & ~new_n4725;
  assign new_n4727 = A129 & A130;
  assign new_n4728 = A127 & A128;
  assign new_n4729 = new_n4727 & ~new_n4728;
  assign new_n4730 = ~A129 & ~A130;
  assign new_n4731 = ~new_n4727 & ~new_n4730;
  assign new_n4732 = ~A127 & ~A128;
  assign new_n4733 = ~new_n4728 & ~new_n4732;
  assign new_n4734 = ~new_n4731 & new_n4733;
  assign new_n4735 = ~new_n4727 & ~new_n4732;
  assign new_n4736 = ~new_n4734 & new_n4735;
  assign new_n4737 = ~new_n4729 & ~new_n4736;
  assign new_n4738 = new_n4724 & new_n4737;
  assign new_n4739 = ~new_n4726 & ~new_n4738;
  assign new_n4740 = new_n4731 & ~new_n4733;
  assign new_n4741 = ~new_n4727 & ~new_n4740;
  assign new_n4742 = ~new_n4732 & ~new_n4741;
  assign new_n4743 = ~new_n4739 & new_n4742;
  assign new_n4744 = new_n4725 & ~new_n4737;
  assign new_n4745 = ~new_n4743 & ~new_n4744;
  assign new_n4746 = ~new_n4724 & new_n4742;
  assign new_n4747 = new_n4745 & ~new_n4746;
  assign new_n4748 = ~A137 & ~A138;
  assign new_n4749 = A137 & A138;
  assign new_n4750 = ~new_n4748 & ~new_n4749;
  assign new_n4751 = ~A136 & new_n4750;
  assign new_n4752 = ~new_n4748 & ~new_n4751;
  assign new_n4753 = ~A134 & ~A135;
  assign new_n4754 = A134 & A135;
  assign new_n4755 = ~new_n4753 & ~new_n4754;
  assign new_n4756 = ~A133 & new_n4755;
  assign new_n4757 = ~new_n4753 & ~new_n4756;
  assign new_n4758 = ~new_n4752 & ~new_n4757;
  assign new_n4759 = A136 & ~new_n4750;
  assign new_n4760 = ~new_n4751 & ~new_n4759;
  assign new_n4761 = A133 & ~new_n4755;
  assign new_n4762 = ~new_n4756 & ~new_n4761;
  assign new_n4763 = ~new_n4760 & ~new_n4762;
  assign new_n4764 = new_n4752 & new_n4757;
  assign new_n4765 = ~new_n4763 & ~new_n4764;
  assign new_n4766 = ~new_n4758 & ~new_n4765;
  assign new_n4767 = ~new_n4747 & new_n4766;
  assign new_n4768 = new_n4760 & new_n4762;
  assign new_n4769 = ~new_n4763 & ~new_n4768;
  assign new_n4770 = ~new_n4734 & ~new_n4740;
  assign new_n4771 = new_n4726 & ~new_n4770;
  assign new_n4772 = ~new_n4726 & new_n4770;
  assign new_n4773 = ~new_n4771 & ~new_n4772;
  assign new_n4774 = new_n4769 & new_n4773;
  assign new_n4775 = ~new_n4763 & ~new_n4774;
  assign new_n4776 = ~new_n4758 & ~new_n4764;
  assign new_n4777 = ~new_n4775 & new_n4776;
  assign new_n4778 = new_n4775 & ~new_n4776;
  assign new_n4779 = ~new_n4777 & ~new_n4778;
  assign new_n4780 = ~new_n4725 & new_n4730;
  assign new_n4781 = new_n4732 & new_n4780;
  assign new_n4782 = ~new_n4738 & ~new_n4781;
  assign new_n4783 = new_n4745 & new_n4782;
  assign new_n4784 = new_n4779 & new_n4783;
  assign new_n4785 = new_n4774 & new_n4776;
  assign new_n4786 = ~new_n4784 & ~new_n4785;
  assign new_n4787 = new_n4747 & ~new_n4766;
  assign new_n4788 = ~new_n4767 & ~new_n4787;
  assign new_n4789 = ~new_n4786 & new_n4788;
  assign new_n4790 = ~new_n4767 & ~new_n4789;
  assign new_n4791 = ~A145 & ~A147;
  assign new_n4792 = A145 & A147;
  assign new_n4793 = ~new_n4791 & ~new_n4792;
  assign new_n4794 = ~A146 & new_n4793;
  assign new_n4795 = ~new_n4791 & ~new_n4794;
  assign new_n4796 = ~A148 & ~A149;
  assign new_n4797 = A146 & ~new_n4793;
  assign new_n4798 = ~new_n4794 & ~new_n4797;
  assign new_n4799 = A150 & ~new_n4798;
  assign new_n4800 = ~A150 & new_n4798;
  assign new_n4801 = ~new_n4799 & ~new_n4800;
  assign new_n4802 = A148 & A149;
  assign new_n4803 = ~new_n4796 & ~new_n4802;
  assign new_n4804 = ~new_n4801 & new_n4803;
  assign new_n4805 = ~new_n4796 & ~new_n4799;
  assign new_n4806 = ~new_n4804 & new_n4805;
  assign new_n4807 = new_n4795 & new_n4806;
  assign new_n4808 = ~new_n4795 & ~new_n4802;
  assign new_n4809 = new_n4799 & ~new_n4808;
  assign new_n4810 = ~new_n4807 & ~new_n4809;
  assign new_n4811 = ~A143 & ~A144;
  assign new_n4812 = A143 & A144;
  assign new_n4813 = ~new_n4811 & ~new_n4812;
  assign new_n4814 = ~A142 & new_n4813;
  assign new_n4815 = ~new_n4811 & ~new_n4814;
  assign new_n4816 = ~A140 & ~A141;
  assign new_n4817 = A140 & A141;
  assign new_n4818 = ~new_n4816 & ~new_n4817;
  assign new_n4819 = ~A139 & new_n4818;
  assign new_n4820 = ~new_n4816 & ~new_n4819;
  assign new_n4821 = new_n4815 & new_n4820;
  assign new_n4822 = A139 & ~new_n4818;
  assign new_n4823 = ~new_n4819 & ~new_n4822;
  assign new_n4824 = A142 & ~new_n4813;
  assign new_n4825 = ~new_n4814 & ~new_n4824;
  assign new_n4826 = ~new_n4823 & ~new_n4825;
  assign new_n4827 = ~new_n4815 & ~new_n4820;
  assign new_n4828 = ~new_n4821 & ~new_n4827;
  assign new_n4829 = new_n4826 & new_n4828;
  assign new_n4830 = ~new_n4821 & ~new_n4829;
  assign new_n4831 = ~new_n4810 & ~new_n4830;
  assign new_n4832 = new_n4810 & new_n4830;
  assign new_n4833 = ~new_n4831 & ~new_n4832;
  assign new_n4834 = new_n4801 & ~new_n4803;
  assign new_n4835 = ~new_n4804 & ~new_n4834;
  assign new_n4836 = new_n4823 & new_n4825;
  assign new_n4837 = ~new_n4826 & ~new_n4836;
  assign new_n4838 = ~new_n4835 & new_n4837;
  assign new_n4839 = ~new_n4826 & ~new_n4838;
  assign new_n4840 = new_n4795 & new_n4802;
  assign new_n4841 = ~new_n4807 & new_n4840;
  assign new_n4842 = ~new_n4810 & ~new_n4841;
  assign new_n4843 = ~new_n4795 & ~new_n4799;
  assign new_n4844 = ~new_n4806 & new_n4843;
  assign new_n4845 = ~new_n4842 & ~new_n4844;
  assign new_n4846 = new_n4839 & ~new_n4845;
  assign new_n4847 = ~new_n4839 & new_n4845;
  assign new_n4848 = ~new_n4846 & ~new_n4847;
  assign new_n4849 = ~new_n4828 & new_n4848;
  assign new_n4850 = ~new_n4829 & ~new_n4846;
  assign new_n4851 = ~new_n4849 & new_n4850;
  assign new_n4852 = new_n4833 & new_n4851;
  assign new_n4853 = ~new_n4831 & ~new_n4852;
  assign new_n4854 = new_n4790 & new_n4853;
  assign new_n4855 = ~new_n4790 & ~new_n4853;
  assign new_n4856 = ~new_n4854 & ~new_n4855;
  assign new_n4857 = new_n4786 & ~new_n4788;
  assign new_n4858 = ~new_n4789 & ~new_n4857;
  assign new_n4859 = ~new_n4779 & ~new_n4783;
  assign new_n4860 = ~new_n4784 & ~new_n4859;
  assign new_n4861 = new_n4835 & ~new_n4837;
  assign new_n4862 = ~new_n4838 & ~new_n4861;
  assign new_n4863 = ~new_n4769 & ~new_n4773;
  assign new_n4864 = ~new_n4774 & ~new_n4863;
  assign new_n4865 = new_n4862 & new_n4864;
  assign new_n4866 = ~new_n4860 & ~new_n4865;
  assign new_n4867 = new_n4828 & ~new_n4848;
  assign new_n4868 = ~new_n4849 & ~new_n4867;
  assign new_n4869 = new_n4860 & new_n4865;
  assign new_n4870 = ~new_n4866 & ~new_n4869;
  assign new_n4871 = new_n4868 & new_n4870;
  assign new_n4872 = ~new_n4866 & ~new_n4871;
  assign new_n4873 = ~new_n4858 & ~new_n4872;
  assign new_n4874 = ~new_n4833 & ~new_n4851;
  assign new_n4875 = ~new_n4852 & ~new_n4874;
  assign new_n4876 = new_n4858 & new_n4872;
  assign new_n4877 = ~new_n4873 & ~new_n4876;
  assign new_n4878 = ~new_n4875 & new_n4877;
  assign new_n4879 = ~new_n4873 & ~new_n4878;
  assign new_n4880 = new_n4856 & ~new_n4879;
  assign new_n4881 = ~new_n4854 & ~new_n4880;
  assign new_n4882 = new_n4723 & ~new_n4881;
  assign new_n4883 = ~new_n4723 & new_n4881;
  assign new_n4884 = ~new_n4882 & ~new_n4883;
  assign new_n4885 = ~new_n4698 & ~new_n4721;
  assign new_n4886 = ~new_n4722 & ~new_n4885;
  assign new_n4887 = new_n4717 & ~new_n4719;
  assign new_n4888 = ~new_n4720 & ~new_n4887;
  assign new_n4889 = ~new_n4868 & ~new_n4870;
  assign new_n4890 = ~new_n4871 & ~new_n4889;
  assign new_n4891 = new_n4708 & ~new_n4710;
  assign new_n4892 = ~new_n4711 & ~new_n4891;
  assign new_n4893 = new_n4890 & ~new_n4892;
  assign new_n4894 = ~new_n4890 & new_n4892;
  assign new_n4895 = ~new_n4862 & ~new_n4864;
  assign new_n4896 = ~new_n4865 & ~new_n4895;
  assign new_n4897 = new_n4702 & ~new_n4704;
  assign new_n4898 = ~new_n4705 & ~new_n4897;
  assign new_n4899 = new_n4896 & new_n4898;
  assign new_n4900 = ~new_n4894 & ~new_n4899;
  assign new_n4901 = ~new_n4893 & ~new_n4900;
  assign new_n4902 = new_n4888 & ~new_n4901;
  assign new_n4903 = new_n4875 & ~new_n4877;
  assign new_n4904 = ~new_n4878 & ~new_n4903;
  assign new_n4905 = ~new_n4888 & new_n4901;
  assign new_n4906 = ~new_n4902 & ~new_n4905;
  assign new_n4907 = new_n4904 & new_n4906;
  assign new_n4908 = ~new_n4902 & ~new_n4907;
  assign new_n4909 = new_n4886 & new_n4908;
  assign new_n4910 = ~new_n4856 & new_n4879;
  assign new_n4911 = ~new_n4880 & ~new_n4910;
  assign new_n4912 = ~new_n4886 & ~new_n4908;
  assign new_n4913 = ~new_n4909 & ~new_n4912;
  assign new_n4914 = ~new_n4911 & new_n4913;
  assign new_n4915 = ~new_n4909 & ~new_n4914;
  assign new_n4916 = new_n4884 & new_n4915;
  assign new_n4917 = ~new_n4884 & ~new_n4915;
  assign new_n4918 = ~new_n4916 & ~new_n4917;
  assign new_n4919 = ~new_n4538 & ~new_n4540;
  assign new_n4920 = ~new_n4541 & ~new_n4919;
  assign new_n4921 = new_n4911 & ~new_n4913;
  assign new_n4922 = ~new_n4914 & ~new_n4921;
  assign new_n4923 = ~new_n4920 & ~new_n4922;
  assign new_n4924 = ~new_n4904 & ~new_n4906;
  assign new_n4925 = ~new_n4907 & ~new_n4924;
  assign new_n4926 = new_n4531 & ~new_n4533;
  assign new_n4927 = ~new_n4534 & ~new_n4926;
  assign new_n4928 = ~new_n4925 & new_n4927;
  assign new_n4929 = new_n4925 & ~new_n4927;
  assign new_n4930 = ~new_n4928 & ~new_n4929;
  assign new_n4931 = ~new_n4513 & ~new_n4523;
  assign new_n4932 = ~new_n4524 & ~new_n4931;
  assign new_n4933 = ~new_n4893 & ~new_n4894;
  assign new_n4934 = ~new_n4896 & ~new_n4898;
  assign new_n4935 = ~new_n4899 & ~new_n4934;
  assign new_n4936 = ~new_n4516 & ~new_n4518;
  assign new_n4937 = ~new_n4519 & ~new_n4936;
  assign new_n4938 = new_n4935 & new_n4937;
  assign new_n4939 = ~new_n4899 & ~new_n4938;
  assign new_n4940 = new_n4933 & ~new_n4939;
  assign new_n4941 = ~new_n4933 & new_n4939;
  assign new_n4942 = ~new_n4940 & ~new_n4941;
  assign new_n4943 = ~new_n4932 & new_n4942;
  assign new_n4944 = ~new_n4938 & ~new_n4942;
  assign new_n4945 = ~new_n4943 & ~new_n4944;
  assign new_n4946 = new_n4930 & new_n4945;
  assign new_n4947 = ~new_n4928 & ~new_n4946;
  assign new_n4948 = new_n4920 & new_n4922;
  assign new_n4949 = ~new_n4923 & ~new_n4948;
  assign new_n4950 = new_n4947 & new_n4949;
  assign new_n4951 = ~new_n4923 & ~new_n4950;
  assign new_n4952 = ~new_n4918 & new_n4951;
  assign new_n4953 = new_n4918 & ~new_n4951;
  assign new_n4954 = ~new_n4952 & ~new_n4953;
  assign new_n4955 = ~new_n4545 & new_n4954;
  assign new_n4956 = new_n4545 & ~new_n4954;
  assign new_n4957 = ~new_n4955 & ~new_n4956;
  assign new_n4958 = new_n4159 & ~new_n4957;
  assign new_n4959 = ~new_n4159 & new_n4957;
  assign new_n4960 = ~new_n4958 & ~new_n4959;
  assign new_n4961 = ~new_n4109 & new_n4133;
  assign new_n4962 = ~new_n4134 & ~new_n4961;
  assign new_n4963 = ~new_n4947 & ~new_n4949;
  assign new_n4964 = ~new_n4950 & ~new_n4963;
  assign new_n4965 = new_n4962 & ~new_n4964;
  assign new_n4966 = new_n4129 & ~new_n4131;
  assign new_n4967 = ~new_n4132 & ~new_n4966;
  assign new_n4968 = new_n4932 & ~new_n4942;
  assign new_n4969 = ~new_n4943 & ~new_n4968;
  assign new_n4970 = ~new_n4116 & ~new_n4118;
  assign new_n4971 = ~new_n4119 & ~new_n4970;
  assign new_n4972 = ~new_n4935 & ~new_n4937;
  assign new_n4973 = ~new_n4938 & ~new_n4972;
  assign new_n4974 = new_n4971 & new_n4973;
  assign new_n4975 = new_n4969 & ~new_n4974;
  assign new_n4976 = new_n4113 & new_n4123;
  assign new_n4977 = ~new_n4124 & ~new_n4976;
  assign new_n4978 = ~new_n4969 & new_n4974;
  assign new_n4979 = ~new_n4975 & ~new_n4978;
  assign new_n4980 = ~new_n4977 & new_n4979;
  assign new_n4981 = ~new_n4975 & ~new_n4980;
  assign new_n4982 = ~new_n4967 & ~new_n4981;
  assign new_n4983 = ~new_n4930 & ~new_n4945;
  assign new_n4984 = ~new_n4946 & ~new_n4983;
  assign new_n4985 = new_n4967 & new_n4981;
  assign new_n4986 = ~new_n4982 & ~new_n4985;
  assign new_n4987 = ~new_n4984 & new_n4986;
  assign new_n4988 = ~new_n4982 & ~new_n4987;
  assign new_n4989 = ~new_n4962 & new_n4964;
  assign new_n4990 = ~new_n4965 & ~new_n4989;
  assign new_n4991 = new_n4988 & new_n4990;
  assign new_n4992 = ~new_n4965 & ~new_n4991;
  assign new_n4993 = new_n4960 & new_n4992;
  assign new_n4994 = ~new_n4958 & ~new_n4993;
  assign new_n4995 = ~new_n4157 & ~new_n4994;
  assign new_n4996 = ~new_n4507 & ~new_n4543;
  assign new_n4997 = ~new_n4882 & ~new_n4916;
  assign new_n4998 = ~new_n4996 & ~new_n4997;
  assign new_n4999 = new_n4996 & new_n4997;
  assign new_n5000 = ~new_n4998 & ~new_n4999;
  assign new_n5001 = ~new_n4952 & ~new_n4955;
  assign new_n5002 = new_n5000 & new_n5001;
  assign new_n5003 = ~new_n5000 & ~new_n5001;
  assign new_n5004 = ~new_n5002 & ~new_n5003;
  assign new_n5005 = new_n4157 & new_n4994;
  assign new_n5006 = ~new_n4995 & ~new_n5005;
  assign new_n5007 = new_n5004 & new_n5006;
  assign new_n5008 = ~new_n4995 & ~new_n5007;
  assign new_n5009 = ~new_n4998 & ~new_n5002;
  assign new_n5010 = ~new_n4152 & ~new_n4155;
  assign new_n5011 = new_n5009 & ~new_n5010;
  assign new_n5012 = ~new_n5009 & new_n5010;
  assign new_n5013 = ~new_n5011 & ~new_n5012;
  assign new_n5014 = new_n5008 & new_n5013;
  assign new_n5015 = ~new_n5008 & ~new_n5013;
  assign new_n5016 = ~new_n5014 & ~new_n5015;
  assign new_n5017 = A277 & A278;
  assign new_n5018 = A280 & A281;
  assign new_n5019 = ~new_n5017 & ~new_n5018;
  assign new_n5020 = A279 & A282;
  assign new_n5021 = ~new_n5019 & new_n5020;
  assign new_n5022 = ~A277 & ~A278;
  assign new_n5023 = ~A279 & A282;
  assign new_n5024 = new_n5018 & new_n5023;
  assign new_n5025 = ~A279 & ~new_n5017;
  assign new_n5026 = ~A280 & ~A281;
  assign new_n5027 = ~new_n5018 & ~new_n5026;
  assign new_n5028 = A282 & ~new_n5027;
  assign new_n5029 = ~A282 & ~new_n5018;
  assign new_n5030 = ~new_n5025 & ~new_n5029;
  assign new_n5031 = ~new_n5028 & new_n5030;
  assign new_n5032 = ~new_n5024 & ~new_n5031;
  assign new_n5033 = ~new_n5022 & ~new_n5032;
  assign new_n5034 = A281 & new_n5017;
  assign new_n5035 = new_n5021 & ~new_n5034;
  assign new_n5036 = ~new_n5020 & new_n5022;
  assign new_n5037 = new_n5026 & new_n5036;
  assign new_n5038 = A279 & ~A282;
  assign new_n5039 = new_n5017 & ~new_n5026;
  assign new_n5040 = new_n5038 & new_n5039;
  assign new_n5041 = ~new_n5037 & ~new_n5040;
  assign new_n5042 = ~new_n5035 & new_n5041;
  assign new_n5043 = ~new_n5033 & new_n5042;
  assign new_n5044 = ~new_n5022 & ~new_n5043;
  assign new_n5045 = ~new_n5021 & ~new_n5044;
  assign new_n5046 = ~A271 & ~A273;
  assign new_n5047 = A271 & A273;
  assign new_n5048 = ~new_n5046 & ~new_n5047;
  assign new_n5049 = ~A272 & new_n5048;
  assign new_n5050 = ~new_n5046 & ~new_n5049;
  assign new_n5051 = ~A275 & ~A276;
  assign new_n5052 = A275 & A276;
  assign new_n5053 = ~new_n5051 & ~new_n5052;
  assign new_n5054 = ~A274 & new_n5053;
  assign new_n5055 = ~new_n5051 & ~new_n5054;
  assign new_n5056 = new_n5050 & new_n5055;
  assign new_n5057 = A272 & ~new_n5048;
  assign new_n5058 = ~new_n5049 & ~new_n5057;
  assign new_n5059 = A274 & ~new_n5053;
  assign new_n5060 = ~new_n5054 & ~new_n5059;
  assign new_n5061 = ~new_n5058 & ~new_n5060;
  assign new_n5062 = ~new_n5050 & ~new_n5055;
  assign new_n5063 = ~new_n5056 & ~new_n5062;
  assign new_n5064 = new_n5061 & new_n5063;
  assign new_n5065 = ~new_n5056 & ~new_n5064;
  assign new_n5066 = ~new_n5045 & ~new_n5065;
  assign new_n5067 = new_n5045 & new_n5065;
  assign new_n5068 = ~new_n5066 & ~new_n5067;
  assign new_n5069 = new_n5058 & new_n5060;
  assign new_n5070 = ~new_n5017 & ~new_n5022;
  assign new_n5071 = ~new_n5023 & ~new_n5038;
  assign new_n5072 = new_n5070 & ~new_n5071;
  assign new_n5073 = ~new_n5070 & new_n5071;
  assign new_n5074 = ~new_n5072 & ~new_n5073;
  assign new_n5075 = new_n5027 & new_n5074;
  assign new_n5076 = ~new_n5027 & ~new_n5074;
  assign new_n5077 = ~new_n5075 & ~new_n5076;
  assign new_n5078 = ~new_n5061 & ~new_n5069;
  assign new_n5079 = ~new_n5077 & new_n5078;
  assign new_n5080 = ~new_n5069 & ~new_n5079;
  assign new_n5081 = new_n5025 & new_n5029;
  assign new_n5082 = ~new_n5075 & new_n5081;
  assign new_n5083 = new_n5043 & ~new_n5082;
  assign new_n5084 = ~new_n5080 & ~new_n5083;
  assign new_n5085 = new_n5080 & new_n5083;
  assign new_n5086 = ~new_n5084 & ~new_n5085;
  assign new_n5087 = ~new_n5063 & new_n5086;
  assign new_n5088 = ~new_n5064 & ~new_n5084;
  assign new_n5089 = ~new_n5087 & new_n5088;
  assign new_n5090 = new_n5068 & new_n5089;
  assign new_n5091 = ~new_n5066 & ~new_n5090;
  assign new_n5092 = A289 & A290;
  assign new_n5093 = A292 & A293;
  assign new_n5094 = ~new_n5092 & ~new_n5093;
  assign new_n5095 = A291 & A294;
  assign new_n5096 = ~new_n5094 & new_n5095;
  assign new_n5097 = ~A289 & ~A290;
  assign new_n5098 = ~A291 & A294;
  assign new_n5099 = new_n5093 & new_n5098;
  assign new_n5100 = ~A291 & ~new_n5092;
  assign new_n5101 = ~A292 & ~A293;
  assign new_n5102 = ~new_n5093 & ~new_n5101;
  assign new_n5103 = A294 & ~new_n5102;
  assign new_n5104 = ~A294 & ~new_n5093;
  assign new_n5105 = ~new_n5100 & ~new_n5104;
  assign new_n5106 = ~new_n5103 & new_n5105;
  assign new_n5107 = ~new_n5099 & ~new_n5106;
  assign new_n5108 = ~new_n5097 & ~new_n5107;
  assign new_n5109 = A293 & new_n5092;
  assign new_n5110 = new_n5096 & ~new_n5109;
  assign new_n5111 = ~new_n5095 & new_n5097;
  assign new_n5112 = new_n5101 & new_n5111;
  assign new_n5113 = A291 & ~A294;
  assign new_n5114 = new_n5092 & ~new_n5101;
  assign new_n5115 = new_n5113 & new_n5114;
  assign new_n5116 = ~new_n5112 & ~new_n5115;
  assign new_n5117 = ~new_n5110 & new_n5116;
  assign new_n5118 = ~new_n5108 & new_n5117;
  assign new_n5119 = ~new_n5097 & ~new_n5118;
  assign new_n5120 = ~new_n5096 & ~new_n5119;
  assign new_n5121 = ~A287 & ~A288;
  assign new_n5122 = A287 & A288;
  assign new_n5123 = ~new_n5121 & ~new_n5122;
  assign new_n5124 = ~A286 & new_n5123;
  assign new_n5125 = ~new_n5121 & ~new_n5124;
  assign new_n5126 = ~A283 & ~A285;
  assign new_n5127 = A283 & A285;
  assign new_n5128 = ~new_n5126 & ~new_n5127;
  assign new_n5129 = ~A284 & new_n5128;
  assign new_n5130 = ~new_n5126 & ~new_n5129;
  assign new_n5131 = new_n5125 & new_n5130;
  assign new_n5132 = A284 & ~new_n5128;
  assign new_n5133 = ~new_n5129 & ~new_n5132;
  assign new_n5134 = A286 & ~new_n5123;
  assign new_n5135 = ~new_n5124 & ~new_n5134;
  assign new_n5136 = ~new_n5133 & ~new_n5135;
  assign new_n5137 = ~new_n5125 & ~new_n5130;
  assign new_n5138 = ~new_n5131 & ~new_n5137;
  assign new_n5139 = new_n5136 & new_n5138;
  assign new_n5140 = ~new_n5131 & ~new_n5139;
  assign new_n5141 = ~new_n5120 & ~new_n5140;
  assign new_n5142 = new_n5120 & new_n5140;
  assign new_n5143 = ~new_n5141 & ~new_n5142;
  assign new_n5144 = new_n5133 & new_n5135;
  assign new_n5145 = ~new_n5092 & ~new_n5097;
  assign new_n5146 = ~new_n5098 & ~new_n5113;
  assign new_n5147 = new_n5145 & ~new_n5146;
  assign new_n5148 = ~new_n5145 & new_n5146;
  assign new_n5149 = ~new_n5147 & ~new_n5148;
  assign new_n5150 = new_n5102 & new_n5149;
  assign new_n5151 = ~new_n5102 & ~new_n5149;
  assign new_n5152 = ~new_n5150 & ~new_n5151;
  assign new_n5153 = ~new_n5136 & ~new_n5144;
  assign new_n5154 = ~new_n5152 & new_n5153;
  assign new_n5155 = ~new_n5144 & ~new_n5154;
  assign new_n5156 = new_n5100 & new_n5104;
  assign new_n5157 = ~new_n5150 & new_n5156;
  assign new_n5158 = new_n5118 & ~new_n5157;
  assign new_n5159 = ~new_n5155 & ~new_n5158;
  assign new_n5160 = new_n5155 & new_n5158;
  assign new_n5161 = ~new_n5159 & ~new_n5160;
  assign new_n5162 = ~new_n5138 & new_n5161;
  assign new_n5163 = ~new_n5139 & ~new_n5159;
  assign new_n5164 = ~new_n5162 & new_n5163;
  assign new_n5165 = new_n5143 & new_n5164;
  assign new_n5166 = ~new_n5141 & ~new_n5165;
  assign new_n5167 = ~new_n5091 & ~new_n5166;
  assign new_n5168 = new_n5091 & new_n5166;
  assign new_n5169 = ~new_n5167 & ~new_n5168;
  assign new_n5170 = ~new_n5068 & ~new_n5089;
  assign new_n5171 = ~new_n5090 & ~new_n5170;
  assign new_n5172 = new_n5138 & ~new_n5161;
  assign new_n5173 = ~new_n5162 & ~new_n5172;
  assign new_n5174 = new_n5063 & ~new_n5086;
  assign new_n5175 = ~new_n5087 & ~new_n5174;
  assign new_n5176 = new_n5173 & new_n5175;
  assign new_n5177 = new_n5077 & ~new_n5078;
  assign new_n5178 = ~new_n5079 & ~new_n5177;
  assign new_n5179 = new_n5152 & ~new_n5153;
  assign new_n5180 = ~new_n5154 & ~new_n5179;
  assign new_n5181 = ~new_n5178 & ~new_n5180;
  assign new_n5182 = ~new_n5173 & ~new_n5175;
  assign new_n5183 = ~new_n5176 & ~new_n5182;
  assign new_n5184 = ~new_n5181 & new_n5183;
  assign new_n5185 = ~new_n5176 & ~new_n5184;
  assign new_n5186 = new_n5171 & new_n5185;
  assign new_n5187 = ~new_n5143 & ~new_n5164;
  assign new_n5188 = ~new_n5165 & ~new_n5187;
  assign new_n5189 = ~new_n5171 & ~new_n5185;
  assign new_n5190 = ~new_n5186 & ~new_n5189;
  assign new_n5191 = new_n5188 & new_n5190;
  assign new_n5192 = ~new_n5186 & ~new_n5191;
  assign new_n5193 = new_n5169 & ~new_n5192;
  assign new_n5194 = ~new_n5167 & ~new_n5193;
  assign new_n5195 = ~A299 & ~A300;
  assign new_n5196 = A299 & A300;
  assign new_n5197 = ~new_n5195 & ~new_n5196;
  assign new_n5198 = ~A298 & new_n5197;
  assign new_n5199 = ~new_n5195 & ~new_n5198;
  assign new_n5200 = ~A296 & ~A297;
  assign new_n5201 = A296 & A297;
  assign new_n5202 = ~new_n5200 & ~new_n5201;
  assign new_n5203 = ~A295 & new_n5202;
  assign new_n5204 = ~new_n5200 & ~new_n5203;
  assign new_n5205 = new_n5199 & new_n5204;
  assign new_n5206 = A295 & ~new_n5202;
  assign new_n5207 = ~new_n5203 & ~new_n5206;
  assign new_n5208 = A298 & ~new_n5197;
  assign new_n5209 = ~new_n5198 & ~new_n5208;
  assign new_n5210 = ~new_n5207 & ~new_n5209;
  assign new_n5211 = ~new_n5199 & ~new_n5204;
  assign new_n5212 = ~new_n5205 & ~new_n5211;
  assign new_n5213 = new_n5210 & new_n5212;
  assign new_n5214 = ~new_n5205 & ~new_n5213;
  assign new_n5215 = ~A305 & ~A306;
  assign new_n5216 = A301 & A302;
  assign new_n5217 = A303 & A304;
  assign new_n5218 = ~new_n5216 & ~new_n5217;
  assign new_n5219 = ~A301 & ~A302;
  assign new_n5220 = ~A303 & ~A304;
  assign new_n5221 = ~new_n5219 & ~new_n5220;
  assign new_n5222 = ~new_n5215 & ~new_n5218;
  assign new_n5223 = new_n5221 & new_n5222;
  assign new_n5224 = new_n5218 & ~new_n5221;
  assign new_n5225 = new_n5216 & new_n5217;
  assign new_n5226 = ~new_n5224 & ~new_n5225;
  assign new_n5227 = ~new_n5215 & ~new_n5226;
  assign new_n5228 = A305 & A306;
  assign new_n5229 = ~new_n5225 & ~new_n5228;
  assign new_n5230 = ~new_n5227 & ~new_n5229;
  assign new_n5231 = ~new_n5223 & ~new_n5230;
  assign new_n5232 = ~new_n5214 & ~new_n5231;
  assign new_n5233 = new_n5214 & new_n5231;
  assign new_n5234 = ~new_n5232 & ~new_n5233;
  assign new_n5235 = new_n5207 & new_n5209;
  assign new_n5236 = ~new_n5210 & ~new_n5235;
  assign new_n5237 = ~new_n5217 & ~new_n5220;
  assign new_n5238 = ~new_n5215 & ~new_n5228;
  assign new_n5239 = new_n5237 & ~new_n5238;
  assign new_n5240 = ~new_n5237 & new_n5238;
  assign new_n5241 = ~new_n5239 & ~new_n5240;
  assign new_n5242 = ~new_n5216 & ~new_n5219;
  assign new_n5243 = ~new_n5241 & new_n5242;
  assign new_n5244 = new_n5241 & ~new_n5242;
  assign new_n5245 = ~new_n5243 & ~new_n5244;
  assign new_n5246 = new_n5236 & ~new_n5245;
  assign new_n5247 = ~new_n5235 & ~new_n5246;
  assign new_n5248 = new_n5219 & new_n5220;
  assign new_n5249 = ~new_n5223 & ~new_n5248;
  assign new_n5250 = ~new_n5228 & ~new_n5249;
  assign new_n5251 = new_n5215 & ~new_n5226;
  assign new_n5252 = ~new_n5230 & ~new_n5251;
  assign new_n5253 = ~new_n5250 & new_n5252;
  assign new_n5254 = ~new_n5247 & ~new_n5253;
  assign new_n5255 = new_n5247 & new_n5253;
  assign new_n5256 = ~new_n5254 & ~new_n5255;
  assign new_n5257 = ~new_n5212 & new_n5256;
  assign new_n5258 = ~new_n5213 & ~new_n5254;
  assign new_n5259 = ~new_n5257 & new_n5258;
  assign new_n5260 = new_n5234 & new_n5259;
  assign new_n5261 = ~new_n5232 & ~new_n5260;
  assign new_n5262 = A313 & A314;
  assign new_n5263 = A316 & A317;
  assign new_n5264 = ~new_n5262 & ~new_n5263;
  assign new_n5265 = A315 & A318;
  assign new_n5266 = ~new_n5264 & new_n5265;
  assign new_n5267 = ~A313 & ~A314;
  assign new_n5268 = ~A315 & A318;
  assign new_n5269 = new_n5263 & new_n5268;
  assign new_n5270 = ~A315 & ~new_n5262;
  assign new_n5271 = ~A316 & ~A317;
  assign new_n5272 = ~new_n5263 & ~new_n5271;
  assign new_n5273 = A318 & ~new_n5272;
  assign new_n5274 = ~A318 & ~new_n5263;
  assign new_n5275 = ~new_n5270 & ~new_n5274;
  assign new_n5276 = ~new_n5273 & new_n5275;
  assign new_n5277 = ~new_n5269 & ~new_n5276;
  assign new_n5278 = ~new_n5267 & ~new_n5277;
  assign new_n5279 = A317 & new_n5262;
  assign new_n5280 = new_n5266 & ~new_n5279;
  assign new_n5281 = ~new_n5265 & new_n5267;
  assign new_n5282 = new_n5271 & new_n5281;
  assign new_n5283 = A315 & ~A318;
  assign new_n5284 = new_n5262 & ~new_n5271;
  assign new_n5285 = new_n5283 & new_n5284;
  assign new_n5286 = ~new_n5282 & ~new_n5285;
  assign new_n5287 = ~new_n5280 & new_n5286;
  assign new_n5288 = ~new_n5278 & new_n5287;
  assign new_n5289 = ~new_n5267 & ~new_n5288;
  assign new_n5290 = ~new_n5266 & ~new_n5289;
  assign new_n5291 = ~A308 & ~A309;
  assign new_n5292 = A308 & A309;
  assign new_n5293 = ~new_n5291 & ~new_n5292;
  assign new_n5294 = ~A307 & new_n5293;
  assign new_n5295 = ~new_n5291 & ~new_n5294;
  assign new_n5296 = ~A310 & ~A311;
  assign new_n5297 = new_n5295 & ~new_n5296;
  assign new_n5298 = A310 & A311;
  assign new_n5299 = ~A312 & ~new_n5298;
  assign new_n5300 = new_n5297 & ~new_n5299;
  assign new_n5301 = ~A312 & ~new_n5297;
  assign new_n5302 = A307 & ~new_n5293;
  assign new_n5303 = ~new_n5294 & ~new_n5302;
  assign new_n5304 = ~new_n5295 & ~new_n5298;
  assign new_n5305 = new_n5295 & new_n5298;
  assign new_n5306 = ~new_n5304 & ~new_n5305;
  assign new_n5307 = A312 & ~new_n5306;
  assign new_n5308 = ~new_n5301 & ~new_n5303;
  assign new_n5309 = ~new_n5307 & new_n5308;
  assign new_n5310 = ~new_n5300 & ~new_n5309;
  assign new_n5311 = new_n5290 & new_n5310;
  assign new_n5312 = ~new_n5262 & ~new_n5267;
  assign new_n5313 = ~new_n5268 & ~new_n5283;
  assign new_n5314 = new_n5312 & ~new_n5313;
  assign new_n5315 = ~new_n5312 & new_n5313;
  assign new_n5316 = ~new_n5314 & ~new_n5315;
  assign new_n5317 = new_n5272 & new_n5316;
  assign new_n5318 = new_n5270 & new_n5274;
  assign new_n5319 = ~new_n5317 & new_n5318;
  assign new_n5320 = new_n5288 & ~new_n5319;
  assign new_n5321 = A312 & ~new_n5303;
  assign new_n5322 = ~new_n5295 & new_n5296;
  assign new_n5323 = ~new_n5321 & new_n5322;
  assign new_n5324 = ~new_n5295 & new_n5299;
  assign new_n5325 = ~new_n5300 & ~new_n5324;
  assign new_n5326 = new_n5303 & ~new_n5325;
  assign new_n5327 = ~new_n5309 & ~new_n5323;
  assign new_n5328 = ~new_n5326 & new_n5327;
  assign new_n5329 = ~new_n5320 & ~new_n5328;
  assign new_n5330 = ~new_n5272 & ~new_n5316;
  assign new_n5331 = ~new_n5317 & ~new_n5330;
  assign new_n5332 = ~A312 & new_n5303;
  assign new_n5333 = ~new_n5321 & ~new_n5332;
  assign new_n5334 = ~new_n5296 & ~new_n5298;
  assign new_n5335 = ~new_n5333 & new_n5334;
  assign new_n5336 = new_n5333 & ~new_n5334;
  assign new_n5337 = ~new_n5335 & ~new_n5336;
  assign new_n5338 = new_n5331 & ~new_n5337;
  assign new_n5339 = new_n5320 & new_n5328;
  assign new_n5340 = ~new_n5329 & ~new_n5339;
  assign new_n5341 = ~new_n5338 & new_n5340;
  assign new_n5342 = ~new_n5329 & ~new_n5341;
  assign new_n5343 = ~new_n5290 & ~new_n5310;
  assign new_n5344 = ~new_n5311 & ~new_n5343;
  assign new_n5345 = ~new_n5342 & new_n5344;
  assign new_n5346 = ~new_n5311 & ~new_n5345;
  assign new_n5347 = ~new_n5261 & new_n5346;
  assign new_n5348 = new_n5261 & ~new_n5346;
  assign new_n5349 = ~new_n5347 & ~new_n5348;
  assign new_n5350 = new_n5342 & ~new_n5344;
  assign new_n5351 = ~new_n5345 & ~new_n5350;
  assign new_n5352 = ~new_n5331 & new_n5337;
  assign new_n5353 = ~new_n5338 & ~new_n5352;
  assign new_n5354 = ~new_n5236 & new_n5245;
  assign new_n5355 = ~new_n5246 & ~new_n5354;
  assign new_n5356 = new_n5353 & ~new_n5355;
  assign new_n5357 = new_n5340 & new_n5356;
  assign new_n5358 = new_n5212 & ~new_n5256;
  assign new_n5359 = ~new_n5257 & ~new_n5358;
  assign new_n5360 = ~new_n5338 & ~new_n5356;
  assign new_n5361 = new_n5340 & ~new_n5360;
  assign new_n5362 = ~new_n5340 & new_n5360;
  assign new_n5363 = ~new_n5361 & ~new_n5362;
  assign new_n5364 = ~new_n5359 & new_n5363;
  assign new_n5365 = ~new_n5357 & ~new_n5364;
  assign new_n5366 = new_n5351 & new_n5365;
  assign new_n5367 = ~new_n5234 & ~new_n5259;
  assign new_n5368 = ~new_n5260 & ~new_n5367;
  assign new_n5369 = ~new_n5351 & ~new_n5365;
  assign new_n5370 = ~new_n5366 & ~new_n5369;
  assign new_n5371 = ~new_n5368 & new_n5370;
  assign new_n5372 = ~new_n5366 & ~new_n5371;
  assign new_n5373 = new_n5349 & new_n5372;
  assign new_n5374 = ~new_n5347 & ~new_n5373;
  assign new_n5375 = ~new_n5194 & ~new_n5374;
  assign new_n5376 = new_n5194 & new_n5374;
  assign new_n5377 = ~new_n5375 & ~new_n5376;
  assign new_n5378 = ~new_n5169 & new_n5192;
  assign new_n5379 = ~new_n5193 & ~new_n5378;
  assign new_n5380 = ~new_n5188 & ~new_n5190;
  assign new_n5381 = ~new_n5191 & ~new_n5380;
  assign new_n5382 = new_n5359 & ~new_n5363;
  assign new_n5383 = ~new_n5364 & ~new_n5382;
  assign new_n5384 = new_n5181 & ~new_n5183;
  assign new_n5385 = ~new_n5184 & ~new_n5384;
  assign new_n5386 = new_n5383 & ~new_n5385;
  assign new_n5387 = ~new_n5353 & new_n5355;
  assign new_n5388 = ~new_n5356 & ~new_n5387;
  assign new_n5389 = new_n5178 & new_n5180;
  assign new_n5390 = ~new_n5181 & ~new_n5389;
  assign new_n5391 = new_n5388 & new_n5390;
  assign new_n5392 = ~new_n5383 & new_n5385;
  assign new_n5393 = ~new_n5386 & ~new_n5392;
  assign new_n5394 = new_n5391 & new_n5393;
  assign new_n5395 = ~new_n5386 & ~new_n5394;
  assign new_n5396 = new_n5381 & ~new_n5395;
  assign new_n5397 = new_n5368 & ~new_n5370;
  assign new_n5398 = ~new_n5371 & ~new_n5397;
  assign new_n5399 = ~new_n5381 & new_n5395;
  assign new_n5400 = ~new_n5396 & ~new_n5399;
  assign new_n5401 = ~new_n5398 & new_n5400;
  assign new_n5402 = ~new_n5396 & ~new_n5401;
  assign new_n5403 = new_n5379 & ~new_n5402;
  assign new_n5404 = ~new_n5349 & ~new_n5372;
  assign new_n5405 = ~new_n5373 & ~new_n5404;
  assign new_n5406 = ~new_n5379 & new_n5402;
  assign new_n5407 = ~new_n5403 & ~new_n5406;
  assign new_n5408 = new_n5405 & new_n5407;
  assign new_n5409 = ~new_n5403 & ~new_n5408;
  assign new_n5410 = new_n5377 & ~new_n5409;
  assign new_n5411 = ~new_n5377 & new_n5409;
  assign new_n5412 = ~new_n5410 & ~new_n5411;
  assign new_n5413 = ~new_n5405 & ~new_n5407;
  assign new_n5414 = ~new_n5408 & ~new_n5413;
  assign new_n5415 = ~A320 & ~A321;
  assign new_n5416 = A320 & A321;
  assign new_n5417 = ~new_n5415 & ~new_n5416;
  assign new_n5418 = ~A319 & new_n5417;
  assign new_n5419 = ~new_n5415 & ~new_n5418;
  assign new_n5420 = ~A323 & ~A324;
  assign new_n5421 = A323 & A324;
  assign new_n5422 = ~new_n5420 & ~new_n5421;
  assign new_n5423 = ~A322 & new_n5422;
  assign new_n5424 = ~new_n5420 & ~new_n5423;
  assign new_n5425 = new_n5419 & new_n5424;
  assign new_n5426 = A322 & ~new_n5422;
  assign new_n5427 = ~new_n5423 & ~new_n5426;
  assign new_n5428 = A319 & ~new_n5417;
  assign new_n5429 = ~new_n5418 & ~new_n5428;
  assign new_n5430 = ~new_n5427 & ~new_n5429;
  assign new_n5431 = ~new_n5419 & ~new_n5424;
  assign new_n5432 = ~new_n5425 & ~new_n5431;
  assign new_n5433 = new_n5430 & new_n5432;
  assign new_n5434 = ~new_n5425 & ~new_n5433;
  assign new_n5435 = ~A329 & ~A330;
  assign new_n5436 = A325 & A326;
  assign new_n5437 = A327 & A328;
  assign new_n5438 = ~new_n5436 & ~new_n5437;
  assign new_n5439 = ~A325 & ~A326;
  assign new_n5440 = ~A327 & ~A328;
  assign new_n5441 = ~new_n5439 & ~new_n5440;
  assign new_n5442 = ~new_n5435 & ~new_n5438;
  assign new_n5443 = new_n5441 & new_n5442;
  assign new_n5444 = new_n5438 & ~new_n5441;
  assign new_n5445 = new_n5436 & new_n5437;
  assign new_n5446 = ~new_n5444 & ~new_n5445;
  assign new_n5447 = ~new_n5435 & ~new_n5446;
  assign new_n5448 = A329 & A330;
  assign new_n5449 = ~new_n5445 & ~new_n5448;
  assign new_n5450 = ~new_n5447 & ~new_n5449;
  assign new_n5451 = ~new_n5443 & ~new_n5450;
  assign new_n5452 = ~new_n5434 & ~new_n5451;
  assign new_n5453 = new_n5434 & new_n5451;
  assign new_n5454 = ~new_n5452 & ~new_n5453;
  assign new_n5455 = new_n5439 & new_n5440;
  assign new_n5456 = ~new_n5443 & ~new_n5455;
  assign new_n5457 = ~new_n5448 & ~new_n5456;
  assign new_n5458 = new_n5435 & ~new_n5446;
  assign new_n5459 = ~new_n5450 & ~new_n5458;
  assign new_n5460 = ~new_n5457 & new_n5459;
  assign new_n5461 = ~new_n5432 & ~new_n5460;
  assign new_n5462 = new_n5427 & new_n5429;
  assign new_n5463 = ~new_n5430 & ~new_n5462;
  assign new_n5464 = ~new_n5435 & ~new_n5448;
  assign new_n5465 = ~new_n5437 & ~new_n5440;
  assign new_n5466 = ~new_n5464 & new_n5465;
  assign new_n5467 = new_n5464 & ~new_n5465;
  assign new_n5468 = ~new_n5466 & ~new_n5467;
  assign new_n5469 = ~new_n5436 & ~new_n5439;
  assign new_n5470 = ~new_n5468 & new_n5469;
  assign new_n5471 = new_n5468 & ~new_n5469;
  assign new_n5472 = ~new_n5470 & ~new_n5471;
  assign new_n5473 = new_n5463 & ~new_n5472;
  assign new_n5474 = ~new_n5462 & ~new_n5473;
  assign new_n5475 = new_n5432 & new_n5460;
  assign new_n5476 = ~new_n5461 & ~new_n5475;
  assign new_n5477 = ~new_n5474 & new_n5476;
  assign new_n5478 = ~new_n5433 & ~new_n5461;
  assign new_n5479 = ~new_n5477 & new_n5478;
  assign new_n5480 = new_n5454 & new_n5479;
  assign new_n5481 = ~new_n5454 & ~new_n5479;
  assign new_n5482 = ~new_n5480 & ~new_n5481;
  assign new_n5483 = ~A331 & ~A332;
  assign new_n5484 = A334 & A335;
  assign new_n5485 = ~A333 & A336;
  assign new_n5486 = new_n5484 & new_n5485;
  assign new_n5487 = A331 & A332;
  assign new_n5488 = ~A333 & ~new_n5487;
  assign new_n5489 = ~A334 & ~A335;
  assign new_n5490 = ~new_n5484 & ~new_n5489;
  assign new_n5491 = A336 & ~new_n5490;
  assign new_n5492 = ~A336 & ~new_n5484;
  assign new_n5493 = ~new_n5488 & ~new_n5492;
  assign new_n5494 = ~new_n5491 & new_n5493;
  assign new_n5495 = ~new_n5486 & ~new_n5494;
  assign new_n5496 = ~new_n5483 & ~new_n5495;
  assign new_n5497 = ~new_n5484 & ~new_n5487;
  assign new_n5498 = A333 & A336;
  assign new_n5499 = ~new_n5497 & new_n5498;
  assign new_n5500 = A335 & new_n5487;
  assign new_n5501 = new_n5499 & ~new_n5500;
  assign new_n5502 = new_n5483 & new_n5489;
  assign new_n5503 = ~new_n5498 & new_n5502;
  assign new_n5504 = A333 & ~A336;
  assign new_n5505 = new_n5487 & ~new_n5489;
  assign new_n5506 = new_n5504 & new_n5505;
  assign new_n5507 = ~new_n5503 & ~new_n5506;
  assign new_n5508 = ~new_n5501 & new_n5507;
  assign new_n5509 = ~new_n5496 & new_n5508;
  assign new_n5510 = ~new_n5483 & ~new_n5487;
  assign new_n5511 = ~new_n5485 & ~new_n5504;
  assign new_n5512 = new_n5510 & ~new_n5511;
  assign new_n5513 = ~new_n5510 & new_n5511;
  assign new_n5514 = ~new_n5512 & ~new_n5513;
  assign new_n5515 = new_n5490 & new_n5514;
  assign new_n5516 = new_n5488 & new_n5492;
  assign new_n5517 = ~new_n5515 & new_n5516;
  assign new_n5518 = new_n5509 & ~new_n5517;
  assign new_n5519 = ~A340 & ~A341;
  assign new_n5520 = ~A337 & ~A338;
  assign new_n5521 = A337 & A338;
  assign new_n5522 = ~new_n5520 & ~new_n5521;
  assign new_n5523 = ~A339 & new_n5522;
  assign new_n5524 = ~new_n5520 & ~new_n5523;
  assign new_n5525 = A339 & ~new_n5522;
  assign new_n5526 = ~new_n5523 & ~new_n5525;
  assign new_n5527 = A342 & ~new_n5526;
  assign new_n5528 = new_n5519 & ~new_n5524;
  assign new_n5529 = ~new_n5527 & new_n5528;
  assign new_n5530 = ~new_n5519 & new_n5524;
  assign new_n5531 = A340 & A341;
  assign new_n5532 = ~A342 & ~new_n5531;
  assign new_n5533 = new_n5530 & ~new_n5532;
  assign new_n5534 = ~new_n5524 & new_n5532;
  assign new_n5535 = ~new_n5533 & ~new_n5534;
  assign new_n5536 = new_n5526 & ~new_n5535;
  assign new_n5537 = ~A342 & ~new_n5530;
  assign new_n5538 = ~new_n5524 & ~new_n5531;
  assign new_n5539 = new_n5524 & new_n5531;
  assign new_n5540 = ~new_n5538 & ~new_n5539;
  assign new_n5541 = A342 & ~new_n5540;
  assign new_n5542 = ~new_n5526 & ~new_n5537;
  assign new_n5543 = ~new_n5541 & new_n5542;
  assign new_n5544 = ~new_n5529 & ~new_n5536;
  assign new_n5545 = ~new_n5543 & new_n5544;
  assign new_n5546 = ~new_n5518 & ~new_n5545;
  assign new_n5547 = ~new_n5490 & ~new_n5514;
  assign new_n5548 = ~new_n5515 & ~new_n5547;
  assign new_n5549 = ~A342 & new_n5526;
  assign new_n5550 = ~new_n5527 & ~new_n5549;
  assign new_n5551 = ~new_n5519 & ~new_n5531;
  assign new_n5552 = ~new_n5550 & new_n5551;
  assign new_n5553 = new_n5550 & ~new_n5551;
  assign new_n5554 = ~new_n5552 & ~new_n5553;
  assign new_n5555 = new_n5548 & ~new_n5554;
  assign new_n5556 = new_n5518 & new_n5545;
  assign new_n5557 = ~new_n5546 & ~new_n5556;
  assign new_n5558 = ~new_n5555 & new_n5557;
  assign new_n5559 = ~new_n5546 & ~new_n5558;
  assign new_n5560 = ~new_n5483 & ~new_n5509;
  assign new_n5561 = ~new_n5499 & ~new_n5560;
  assign new_n5562 = ~new_n5533 & ~new_n5543;
  assign new_n5563 = new_n5561 & new_n5562;
  assign new_n5564 = ~new_n5561 & ~new_n5562;
  assign new_n5565 = ~new_n5563 & ~new_n5564;
  assign new_n5566 = ~new_n5559 & new_n5565;
  assign new_n5567 = new_n5559 & ~new_n5565;
  assign new_n5568 = ~new_n5566 & ~new_n5567;
  assign new_n5569 = new_n5474 & ~new_n5476;
  assign new_n5570 = ~new_n5477 & ~new_n5569;
  assign new_n5571 = new_n5555 & ~new_n5557;
  assign new_n5572 = ~new_n5558 & ~new_n5571;
  assign new_n5573 = ~new_n5570 & ~new_n5572;
  assign new_n5574 = new_n5570 & new_n5572;
  assign new_n5575 = ~new_n5548 & new_n5554;
  assign new_n5576 = ~new_n5555 & ~new_n5575;
  assign new_n5577 = ~new_n5463 & new_n5472;
  assign new_n5578 = ~new_n5473 & ~new_n5577;
  assign new_n5579 = new_n5576 & ~new_n5578;
  assign new_n5580 = ~new_n5574 & new_n5579;
  assign new_n5581 = ~new_n5573 & ~new_n5580;
  assign new_n5582 = new_n5568 & new_n5581;
  assign new_n5583 = ~new_n5568 & ~new_n5581;
  assign new_n5584 = ~new_n5582 & ~new_n5583;
  assign new_n5585 = ~new_n5482 & new_n5584;
  assign new_n5586 = new_n5482 & ~new_n5584;
  assign new_n5587 = ~new_n5585 & ~new_n5586;
  assign new_n5588 = ~A343 & ~A344;
  assign new_n5589 = A343 & A344;
  assign new_n5590 = ~A345 & ~new_n5589;
  assign new_n5591 = ~new_n5588 & ~new_n5590;
  assign new_n5592 = A345 & new_n5589;
  assign new_n5593 = ~A346 & ~new_n5592;
  assign new_n5594 = new_n5591 & ~new_n5593;
  assign new_n5595 = A347 & new_n5594;
  assign new_n5596 = A345 & A346;
  assign new_n5597 = new_n5589 & new_n5596;
  assign new_n5598 = ~new_n5595 & ~new_n5597;
  assign new_n5599 = ~A348 & ~new_n5598;
  assign new_n5600 = A347 & A348;
  assign new_n5601 = new_n5591 & new_n5600;
  assign new_n5602 = ~A347 & ~A348;
  assign new_n5603 = ~new_n5588 & ~new_n5602;
  assign new_n5604 = new_n5590 & ~new_n5600;
  assign new_n5605 = ~new_n5603 & new_n5604;
  assign new_n5606 = ~new_n5601 & ~new_n5605;
  assign new_n5607 = ~A346 & ~new_n5606;
  assign new_n5608 = ~A347 & A348;
  assign new_n5609 = new_n5594 & new_n5608;
  assign new_n5610 = new_n5588 & ~new_n5596;
  assign new_n5611 = A346 & new_n5600;
  assign new_n5612 = ~new_n5592 & new_n5611;
  assign new_n5613 = ~new_n5610 & new_n5612;
  assign new_n5614 = ~new_n5609 & ~new_n5613;
  assign new_n5615 = ~new_n5607 & new_n5614;
  assign new_n5616 = ~new_n5599 & new_n5615;
  assign new_n5617 = new_n5602 & new_n5610;
  assign new_n5618 = new_n5616 & ~new_n5617;
  assign new_n5619 = A346 & ~A348;
  assign new_n5620 = ~A346 & A348;
  assign new_n5621 = ~new_n5619 & ~new_n5620;
  assign new_n5622 = ~new_n5588 & ~new_n5589;
  assign new_n5623 = ~A345 & ~A347;
  assign new_n5624 = A345 & A347;
  assign new_n5625 = ~new_n5623 & ~new_n5624;
  assign new_n5626 = new_n5622 & ~new_n5625;
  assign new_n5627 = ~new_n5622 & new_n5625;
  assign new_n5628 = ~new_n5626 & ~new_n5627;
  assign new_n5629 = new_n5621 & new_n5628;
  assign new_n5630 = ~new_n5621 & ~new_n5628;
  assign new_n5631 = ~new_n5629 & ~new_n5630;
  assign new_n5632 = ~A349 & ~A351;
  assign new_n5633 = A349 & A351;
  assign new_n5634 = ~new_n5632 & ~new_n5633;
  assign new_n5635 = ~A350 & new_n5634;
  assign new_n5636 = A350 & ~new_n5634;
  assign new_n5637 = ~new_n5635 & ~new_n5636;
  assign new_n5638 = A354 & ~new_n5637;
  assign new_n5639 = ~A354 & new_n5637;
  assign new_n5640 = ~new_n5638 & ~new_n5639;
  assign new_n5641 = ~A352 & ~A353;
  assign new_n5642 = A352 & A353;
  assign new_n5643 = ~new_n5641 & ~new_n5642;
  assign new_n5644 = ~new_n5640 & new_n5643;
  assign new_n5645 = new_n5640 & ~new_n5643;
  assign new_n5646 = ~new_n5644 & ~new_n5645;
  assign new_n5647 = new_n5631 & ~new_n5646;
  assign new_n5648 = ~new_n5632 & ~new_n5635;
  assign new_n5649 = new_n5641 & ~new_n5648;
  assign new_n5650 = ~new_n5638 & new_n5649;
  assign new_n5651 = ~new_n5641 & new_n5648;
  assign new_n5652 = ~A354 & ~new_n5642;
  assign new_n5653 = new_n5651 & ~new_n5652;
  assign new_n5654 = ~new_n5642 & ~new_n5648;
  assign new_n5655 = ~A354 & new_n5654;
  assign new_n5656 = ~new_n5653 & ~new_n5655;
  assign new_n5657 = new_n5637 & ~new_n5656;
  assign new_n5658 = new_n5642 & new_n5648;
  assign new_n5659 = ~new_n5654 & ~new_n5658;
  assign new_n5660 = A354 & ~new_n5659;
  assign new_n5661 = ~A354 & ~new_n5651;
  assign new_n5662 = ~new_n5637 & ~new_n5661;
  assign new_n5663 = ~new_n5660 & new_n5662;
  assign new_n5664 = ~new_n5650 & ~new_n5657;
  assign new_n5665 = ~new_n5663 & new_n5664;
  assign new_n5666 = ~new_n5647 & ~new_n5665;
  assign new_n5667 = new_n5647 & new_n5665;
  assign new_n5668 = ~new_n5666 & ~new_n5667;
  assign new_n5669 = ~new_n5618 & new_n5668;
  assign new_n5670 = new_n5618 & ~new_n5668;
  assign new_n5671 = ~new_n5669 & ~new_n5670;
  assign new_n5672 = ~A361 & ~A362;
  assign new_n5673 = A364 & A365;
  assign new_n5674 = ~A363 & A366;
  assign new_n5675 = new_n5673 & new_n5674;
  assign new_n5676 = A361 & A362;
  assign new_n5677 = ~A363 & ~new_n5676;
  assign new_n5678 = ~A364 & ~A365;
  assign new_n5679 = ~new_n5673 & ~new_n5678;
  assign new_n5680 = A366 & ~new_n5679;
  assign new_n5681 = ~A366 & ~new_n5673;
  assign new_n5682 = ~new_n5677 & ~new_n5681;
  assign new_n5683 = ~new_n5680 & new_n5682;
  assign new_n5684 = ~new_n5675 & ~new_n5683;
  assign new_n5685 = ~new_n5672 & ~new_n5684;
  assign new_n5686 = ~new_n5673 & ~new_n5676;
  assign new_n5687 = A363 & A366;
  assign new_n5688 = ~new_n5686 & new_n5687;
  assign new_n5689 = A365 & new_n5676;
  assign new_n5690 = new_n5688 & ~new_n5689;
  assign new_n5691 = new_n5672 & new_n5678;
  assign new_n5692 = ~new_n5687 & new_n5691;
  assign new_n5693 = A363 & ~A366;
  assign new_n5694 = new_n5676 & ~new_n5678;
  assign new_n5695 = new_n5693 & new_n5694;
  assign new_n5696 = ~new_n5692 & ~new_n5695;
  assign new_n5697 = ~new_n5690 & new_n5696;
  assign new_n5698 = ~new_n5685 & new_n5697;
  assign new_n5699 = ~new_n5672 & ~new_n5676;
  assign new_n5700 = ~new_n5674 & ~new_n5693;
  assign new_n5701 = new_n5699 & ~new_n5700;
  assign new_n5702 = ~new_n5699 & new_n5700;
  assign new_n5703 = ~new_n5701 & ~new_n5702;
  assign new_n5704 = new_n5679 & new_n5703;
  assign new_n5705 = new_n5677 & new_n5681;
  assign new_n5706 = ~new_n5704 & new_n5705;
  assign new_n5707 = new_n5698 & ~new_n5706;
  assign new_n5708 = ~A358 & ~A359;
  assign new_n5709 = ~A356 & ~A357;
  assign new_n5710 = A356 & A357;
  assign new_n5711 = ~new_n5709 & ~new_n5710;
  assign new_n5712 = ~A355 & new_n5711;
  assign new_n5713 = ~new_n5709 & ~new_n5712;
  assign new_n5714 = A355 & ~new_n5711;
  assign new_n5715 = ~new_n5712 & ~new_n5714;
  assign new_n5716 = A360 & ~new_n5715;
  assign new_n5717 = new_n5708 & ~new_n5713;
  assign new_n5718 = ~new_n5716 & new_n5717;
  assign new_n5719 = ~new_n5708 & new_n5713;
  assign new_n5720 = A358 & A359;
  assign new_n5721 = ~A360 & ~new_n5720;
  assign new_n5722 = new_n5719 & ~new_n5721;
  assign new_n5723 = ~new_n5713 & new_n5721;
  assign new_n5724 = ~new_n5722 & ~new_n5723;
  assign new_n5725 = new_n5715 & ~new_n5724;
  assign new_n5726 = ~A360 & ~new_n5719;
  assign new_n5727 = ~new_n5713 & ~new_n5720;
  assign new_n5728 = new_n5713 & new_n5720;
  assign new_n5729 = ~new_n5727 & ~new_n5728;
  assign new_n5730 = A360 & ~new_n5729;
  assign new_n5731 = ~new_n5715 & ~new_n5726;
  assign new_n5732 = ~new_n5730 & new_n5731;
  assign new_n5733 = ~new_n5718 & ~new_n5725;
  assign new_n5734 = ~new_n5732 & new_n5733;
  assign new_n5735 = ~new_n5707 & ~new_n5734;
  assign new_n5736 = new_n5707 & new_n5734;
  assign new_n5737 = ~new_n5735 & ~new_n5736;
  assign new_n5738 = ~new_n5679 & ~new_n5703;
  assign new_n5739 = ~new_n5704 & ~new_n5738;
  assign new_n5740 = ~A360 & new_n5715;
  assign new_n5741 = ~new_n5716 & ~new_n5740;
  assign new_n5742 = ~new_n5708 & ~new_n5720;
  assign new_n5743 = ~new_n5741 & new_n5742;
  assign new_n5744 = new_n5741 & ~new_n5742;
  assign new_n5745 = ~new_n5743 & ~new_n5744;
  assign new_n5746 = new_n5739 & ~new_n5745;
  assign new_n5747 = ~new_n5739 & new_n5745;
  assign new_n5748 = ~new_n5746 & ~new_n5747;
  assign new_n5749 = ~new_n5631 & new_n5646;
  assign new_n5750 = ~new_n5647 & ~new_n5749;
  assign new_n5751 = new_n5748 & new_n5750;
  assign new_n5752 = ~new_n5746 & ~new_n5751;
  assign new_n5753 = new_n5737 & ~new_n5752;
  assign new_n5754 = ~new_n5737 & new_n5752;
  assign new_n5755 = ~new_n5753 & ~new_n5754;
  assign new_n5756 = ~new_n5671 & new_n5755;
  assign new_n5757 = new_n5671 & ~new_n5755;
  assign new_n5758 = ~new_n5756 & ~new_n5757;
  assign new_n5759 = ~new_n5573 & ~new_n5574;
  assign new_n5760 = ~new_n5576 & new_n5578;
  assign new_n5761 = ~new_n5579 & ~new_n5760;
  assign new_n5762 = ~new_n5748 & ~new_n5750;
  assign new_n5763 = ~new_n5751 & ~new_n5762;
  assign new_n5764 = new_n5761 & new_n5763;
  assign new_n5765 = ~new_n5579 & ~new_n5764;
  assign new_n5766 = new_n5759 & ~new_n5765;
  assign new_n5767 = ~new_n5759 & new_n5765;
  assign new_n5768 = ~new_n5766 & ~new_n5767;
  assign new_n5769 = new_n5758 & new_n5768;
  assign new_n5770 = new_n5759 & new_n5764;
  assign new_n5771 = ~new_n5769 & ~new_n5770;
  assign new_n5772 = ~new_n5666 & ~new_n5669;
  assign new_n5773 = ~new_n5593 & ~new_n5616;
  assign new_n5774 = ~new_n5601 & ~new_n5773;
  assign new_n5775 = ~new_n5653 & ~new_n5663;
  assign new_n5776 = new_n5774 & new_n5775;
  assign new_n5777 = ~new_n5774 & ~new_n5775;
  assign new_n5778 = ~new_n5776 & ~new_n5777;
  assign new_n5779 = ~new_n5772 & new_n5778;
  assign new_n5780 = new_n5772 & ~new_n5778;
  assign new_n5781 = ~new_n5779 & ~new_n5780;
  assign new_n5782 = new_n5737 & ~new_n5746;
  assign new_n5783 = ~new_n5735 & ~new_n5782;
  assign new_n5784 = ~new_n5672 & ~new_n5698;
  assign new_n5785 = ~new_n5688 & ~new_n5784;
  assign new_n5786 = ~new_n5722 & ~new_n5732;
  assign new_n5787 = new_n5785 & new_n5786;
  assign new_n5788 = ~new_n5785 & ~new_n5786;
  assign new_n5789 = ~new_n5787 & ~new_n5788;
  assign new_n5790 = ~new_n5783 & new_n5789;
  assign new_n5791 = new_n5783 & ~new_n5789;
  assign new_n5792 = ~new_n5790 & ~new_n5791;
  assign new_n5793 = new_n5737 & new_n5751;
  assign new_n5794 = ~new_n5756 & ~new_n5793;
  assign new_n5795 = ~new_n5792 & ~new_n5794;
  assign new_n5796 = new_n5792 & new_n5794;
  assign new_n5797 = ~new_n5795 & ~new_n5796;
  assign new_n5798 = ~new_n5781 & new_n5797;
  assign new_n5799 = new_n5781 & ~new_n5797;
  assign new_n5800 = ~new_n5798 & ~new_n5799;
  assign new_n5801 = ~new_n5771 & new_n5800;
  assign new_n5802 = new_n5771 & ~new_n5800;
  assign new_n5803 = ~new_n5801 & ~new_n5802;
  assign new_n5804 = ~new_n5587 & new_n5803;
  assign new_n5805 = new_n5587 & ~new_n5803;
  assign new_n5806 = ~new_n5804 & ~new_n5805;
  assign new_n5807 = ~new_n5758 & ~new_n5768;
  assign new_n5808 = ~new_n5769 & ~new_n5807;
  assign new_n5809 = ~new_n5761 & ~new_n5763;
  assign new_n5810 = ~new_n5764 & ~new_n5809;
  assign new_n5811 = ~new_n5388 & ~new_n5390;
  assign new_n5812 = ~new_n5391 & ~new_n5811;
  assign new_n5813 = new_n5810 & new_n5812;
  assign new_n5814 = ~new_n5808 & ~new_n5813;
  assign new_n5815 = ~new_n5391 & ~new_n5393;
  assign new_n5816 = ~new_n5394 & ~new_n5815;
  assign new_n5817 = new_n5808 & new_n5813;
  assign new_n5818 = ~new_n5814 & ~new_n5817;
  assign new_n5819 = ~new_n5816 & new_n5818;
  assign new_n5820 = ~new_n5814 & ~new_n5819;
  assign new_n5821 = new_n5806 & new_n5820;
  assign new_n5822 = new_n5398 & ~new_n5400;
  assign new_n5823 = ~new_n5401 & ~new_n5822;
  assign new_n5824 = ~new_n5806 & ~new_n5820;
  assign new_n5825 = ~new_n5821 & ~new_n5824;
  assign new_n5826 = new_n5823 & new_n5825;
  assign new_n5827 = ~new_n5821 & ~new_n5826;
  assign new_n5828 = new_n5414 & ~new_n5827;
  assign new_n5829 = ~new_n5795 & ~new_n5798;
  assign new_n5830 = ~new_n5776 & ~new_n5779;
  assign new_n5831 = ~new_n5787 & ~new_n5790;
  assign new_n5832 = new_n5830 & new_n5831;
  assign new_n5833 = ~new_n5830 & ~new_n5831;
  assign new_n5834 = ~new_n5832 & ~new_n5833;
  assign new_n5835 = ~new_n5829 & new_n5834;
  assign new_n5836 = new_n5829 & ~new_n5834;
  assign new_n5837 = ~new_n5835 & ~new_n5836;
  assign new_n5838 = ~new_n5582 & ~new_n5585;
  assign new_n5839 = ~new_n5452 & ~new_n5480;
  assign new_n5840 = ~new_n5563 & ~new_n5566;
  assign new_n5841 = new_n5839 & ~new_n5840;
  assign new_n5842 = ~new_n5839 & new_n5840;
  assign new_n5843 = ~new_n5841 & ~new_n5842;
  assign new_n5844 = ~new_n5838 & new_n5843;
  assign new_n5845 = new_n5838 & ~new_n5843;
  assign new_n5846 = ~new_n5844 & ~new_n5845;
  assign new_n5847 = ~new_n5801 & ~new_n5804;
  assign new_n5848 = new_n5846 & new_n5847;
  assign new_n5849 = ~new_n5846 & ~new_n5847;
  assign new_n5850 = ~new_n5848 & ~new_n5849;
  assign new_n5851 = ~new_n5837 & new_n5850;
  assign new_n5852 = new_n5837 & ~new_n5850;
  assign new_n5853 = ~new_n5851 & ~new_n5852;
  assign new_n5854 = ~new_n5414 & new_n5827;
  assign new_n5855 = ~new_n5828 & ~new_n5854;
  assign new_n5856 = ~new_n5853 & new_n5855;
  assign new_n5857 = ~new_n5828 & ~new_n5856;
  assign new_n5858 = ~new_n5412 & new_n5857;
  assign new_n5859 = ~new_n5841 & ~new_n5844;
  assign new_n5860 = ~new_n5832 & ~new_n5835;
  assign new_n5861 = new_n5859 & ~new_n5860;
  assign new_n5862 = ~new_n5859 & new_n5860;
  assign new_n5863 = ~new_n5861 & ~new_n5862;
  assign new_n5864 = ~new_n5848 & ~new_n5851;
  assign new_n5865 = new_n5863 & new_n5864;
  assign new_n5866 = ~new_n5863 & ~new_n5864;
  assign new_n5867 = ~new_n5865 & ~new_n5866;
  assign new_n5868 = new_n5412 & ~new_n5857;
  assign new_n5869 = ~new_n5858 & ~new_n5868;
  assign new_n5870 = ~new_n5867 & new_n5869;
  assign new_n5871 = ~new_n5858 & ~new_n5870;
  assign new_n5872 = ~new_n5861 & ~new_n5865;
  assign new_n5873 = ~new_n5375 & ~new_n5410;
  assign new_n5874 = new_n5872 & new_n5873;
  assign new_n5875 = ~new_n5872 & ~new_n5873;
  assign new_n5876 = ~new_n5874 & ~new_n5875;
  assign new_n5877 = ~new_n5871 & new_n5876;
  assign new_n5878 = new_n5871 & ~new_n5876;
  assign new_n5879 = ~new_n5877 & ~new_n5878;
  assign new_n5880 = A451 & A452;
  assign new_n5881 = A454 & A455;
  assign new_n5882 = ~new_n5880 & ~new_n5881;
  assign new_n5883 = A453 & A456;
  assign new_n5884 = ~new_n5882 & new_n5883;
  assign new_n5885 = ~A451 & ~A452;
  assign new_n5886 = ~A453 & A456;
  assign new_n5887 = new_n5881 & new_n5886;
  assign new_n5888 = ~A453 & ~new_n5880;
  assign new_n5889 = ~A454 & ~A455;
  assign new_n5890 = ~new_n5881 & ~new_n5889;
  assign new_n5891 = A456 & ~new_n5890;
  assign new_n5892 = ~A456 & ~new_n5881;
  assign new_n5893 = ~new_n5888 & ~new_n5892;
  assign new_n5894 = ~new_n5891 & new_n5893;
  assign new_n5895 = ~new_n5887 & ~new_n5894;
  assign new_n5896 = ~new_n5885 & ~new_n5895;
  assign new_n5897 = A455 & new_n5880;
  assign new_n5898 = new_n5884 & ~new_n5897;
  assign new_n5899 = ~new_n5883 & new_n5885;
  assign new_n5900 = new_n5889 & new_n5899;
  assign new_n5901 = A453 & ~A456;
  assign new_n5902 = new_n5880 & ~new_n5889;
  assign new_n5903 = new_n5901 & new_n5902;
  assign new_n5904 = ~new_n5900 & ~new_n5903;
  assign new_n5905 = ~new_n5898 & new_n5904;
  assign new_n5906 = ~new_n5896 & new_n5905;
  assign new_n5907 = ~new_n5885 & ~new_n5906;
  assign new_n5908 = ~new_n5884 & ~new_n5907;
  assign new_n5909 = ~A458 & ~A459;
  assign new_n5910 = A458 & A459;
  assign new_n5911 = ~new_n5909 & ~new_n5910;
  assign new_n5912 = ~A457 & new_n5911;
  assign new_n5913 = ~new_n5909 & ~new_n5912;
  assign new_n5914 = ~A460 & ~A461;
  assign new_n5915 = new_n5913 & ~new_n5914;
  assign new_n5916 = A460 & A461;
  assign new_n5917 = ~A462 & ~new_n5916;
  assign new_n5918 = new_n5915 & ~new_n5917;
  assign new_n5919 = ~A462 & ~new_n5915;
  assign new_n5920 = A457 & ~new_n5911;
  assign new_n5921 = ~new_n5912 & ~new_n5920;
  assign new_n5922 = ~new_n5913 & ~new_n5916;
  assign new_n5923 = new_n5913 & new_n5916;
  assign new_n5924 = ~new_n5922 & ~new_n5923;
  assign new_n5925 = A462 & ~new_n5924;
  assign new_n5926 = ~new_n5919 & ~new_n5921;
  assign new_n5927 = ~new_n5925 & new_n5926;
  assign new_n5928 = ~new_n5918 & ~new_n5927;
  assign new_n5929 = new_n5908 & new_n5928;
  assign new_n5930 = ~new_n5880 & ~new_n5885;
  assign new_n5931 = ~new_n5886 & ~new_n5901;
  assign new_n5932 = new_n5930 & ~new_n5931;
  assign new_n5933 = ~new_n5930 & new_n5931;
  assign new_n5934 = ~new_n5932 & ~new_n5933;
  assign new_n5935 = new_n5890 & new_n5934;
  assign new_n5936 = new_n5888 & new_n5892;
  assign new_n5937 = ~new_n5935 & new_n5936;
  assign new_n5938 = new_n5906 & ~new_n5937;
  assign new_n5939 = A462 & ~new_n5921;
  assign new_n5940 = ~new_n5913 & new_n5914;
  assign new_n5941 = ~new_n5939 & new_n5940;
  assign new_n5942 = ~new_n5913 & new_n5917;
  assign new_n5943 = ~new_n5918 & ~new_n5942;
  assign new_n5944 = new_n5921 & ~new_n5943;
  assign new_n5945 = ~new_n5927 & ~new_n5941;
  assign new_n5946 = ~new_n5944 & new_n5945;
  assign new_n5947 = ~new_n5938 & ~new_n5946;
  assign new_n5948 = ~new_n5890 & ~new_n5934;
  assign new_n5949 = ~new_n5935 & ~new_n5948;
  assign new_n5950 = ~A462 & new_n5921;
  assign new_n5951 = ~new_n5939 & ~new_n5950;
  assign new_n5952 = ~new_n5914 & ~new_n5916;
  assign new_n5953 = ~new_n5951 & new_n5952;
  assign new_n5954 = new_n5951 & ~new_n5952;
  assign new_n5955 = ~new_n5953 & ~new_n5954;
  assign new_n5956 = new_n5949 & ~new_n5955;
  assign new_n5957 = new_n5938 & new_n5946;
  assign new_n5958 = ~new_n5947 & ~new_n5957;
  assign new_n5959 = ~new_n5956 & new_n5958;
  assign new_n5960 = ~new_n5947 & ~new_n5959;
  assign new_n5961 = ~new_n5908 & ~new_n5928;
  assign new_n5962 = ~new_n5929 & ~new_n5961;
  assign new_n5963 = ~new_n5960 & new_n5962;
  assign new_n5964 = ~new_n5929 & ~new_n5963;
  assign new_n5965 = A445 & A446;
  assign new_n5966 = A448 & A449;
  assign new_n5967 = ~new_n5965 & ~new_n5966;
  assign new_n5968 = A447 & A450;
  assign new_n5969 = ~new_n5967 & new_n5968;
  assign new_n5970 = ~A445 & ~A446;
  assign new_n5971 = ~A447 & A450;
  assign new_n5972 = new_n5966 & new_n5971;
  assign new_n5973 = ~A447 & ~new_n5965;
  assign new_n5974 = ~A448 & ~A449;
  assign new_n5975 = ~new_n5966 & ~new_n5974;
  assign new_n5976 = A450 & ~new_n5975;
  assign new_n5977 = ~A450 & ~new_n5966;
  assign new_n5978 = ~new_n5973 & ~new_n5977;
  assign new_n5979 = ~new_n5976 & new_n5978;
  assign new_n5980 = ~new_n5972 & ~new_n5979;
  assign new_n5981 = ~new_n5970 & ~new_n5980;
  assign new_n5982 = A449 & new_n5965;
  assign new_n5983 = new_n5969 & ~new_n5982;
  assign new_n5984 = ~new_n5968 & new_n5970;
  assign new_n5985 = new_n5974 & new_n5984;
  assign new_n5986 = A447 & ~A450;
  assign new_n5987 = new_n5965 & ~new_n5974;
  assign new_n5988 = new_n5986 & new_n5987;
  assign new_n5989 = ~new_n5985 & ~new_n5988;
  assign new_n5990 = ~new_n5983 & new_n5989;
  assign new_n5991 = ~new_n5981 & new_n5990;
  assign new_n5992 = ~new_n5970 & ~new_n5991;
  assign new_n5993 = ~new_n5969 & ~new_n5992;
  assign new_n5994 = A439 & A440;
  assign new_n5995 = A442 & A443;
  assign new_n5996 = ~new_n5994 & ~new_n5995;
  assign new_n5997 = A441 & A444;
  assign new_n5998 = ~new_n5996 & new_n5997;
  assign new_n5999 = ~A439 & ~A440;
  assign new_n6000 = ~A441 & A444;
  assign new_n6001 = new_n5995 & new_n6000;
  assign new_n6002 = ~A441 & ~new_n5994;
  assign new_n6003 = ~A442 & ~A443;
  assign new_n6004 = ~new_n5995 & ~new_n6003;
  assign new_n6005 = A444 & ~new_n6004;
  assign new_n6006 = ~A444 & ~new_n5995;
  assign new_n6007 = ~new_n6002 & ~new_n6006;
  assign new_n6008 = ~new_n6005 & new_n6007;
  assign new_n6009 = ~new_n6001 & ~new_n6008;
  assign new_n6010 = ~new_n5999 & ~new_n6009;
  assign new_n6011 = A443 & new_n5994;
  assign new_n6012 = new_n5998 & ~new_n6011;
  assign new_n6013 = ~new_n5997 & new_n5999;
  assign new_n6014 = new_n6003 & new_n6013;
  assign new_n6015 = A441 & ~A444;
  assign new_n6016 = new_n5994 & ~new_n6003;
  assign new_n6017 = new_n6015 & new_n6016;
  assign new_n6018 = ~new_n6014 & ~new_n6017;
  assign new_n6019 = ~new_n6012 & new_n6018;
  assign new_n6020 = ~new_n6010 & new_n6019;
  assign new_n6021 = ~new_n5999 & ~new_n6020;
  assign new_n6022 = ~new_n5998 & ~new_n6021;
  assign new_n6023 = new_n5993 & new_n6022;
  assign new_n6024 = ~new_n5965 & ~new_n5970;
  assign new_n6025 = ~new_n5971 & ~new_n5986;
  assign new_n6026 = new_n6024 & ~new_n6025;
  assign new_n6027 = ~new_n6024 & new_n6025;
  assign new_n6028 = ~new_n6026 & ~new_n6027;
  assign new_n6029 = new_n5975 & new_n6028;
  assign new_n6030 = ~new_n5975 & ~new_n6028;
  assign new_n6031 = ~new_n6029 & ~new_n6030;
  assign new_n6032 = ~new_n5994 & ~new_n5999;
  assign new_n6033 = ~new_n6000 & ~new_n6015;
  assign new_n6034 = new_n6032 & ~new_n6033;
  assign new_n6035 = ~new_n6032 & new_n6033;
  assign new_n6036 = ~new_n6034 & ~new_n6035;
  assign new_n6037 = new_n6004 & new_n6036;
  assign new_n6038 = ~new_n6004 & ~new_n6036;
  assign new_n6039 = ~new_n6037 & ~new_n6038;
  assign new_n6040 = new_n6031 & new_n6039;
  assign new_n6041 = new_n5973 & new_n5977;
  assign new_n6042 = ~new_n6029 & new_n6041;
  assign new_n6043 = new_n5991 & ~new_n6042;
  assign new_n6044 = ~new_n6040 & ~new_n6043;
  assign new_n6045 = new_n6040 & new_n6043;
  assign new_n6046 = ~new_n6044 & ~new_n6045;
  assign new_n6047 = new_n6002 & new_n6006;
  assign new_n6048 = ~new_n6037 & new_n6047;
  assign new_n6049 = new_n6020 & ~new_n6048;
  assign new_n6050 = new_n6046 & ~new_n6049;
  assign new_n6051 = ~new_n6044 & ~new_n6050;
  assign new_n6052 = ~new_n5993 & ~new_n6022;
  assign new_n6053 = ~new_n6023 & ~new_n6052;
  assign new_n6054 = ~new_n6051 & new_n6053;
  assign new_n6055 = ~new_n6023 & ~new_n6054;
  assign new_n6056 = ~new_n5964 & ~new_n6055;
  assign new_n6057 = new_n5964 & new_n6055;
  assign new_n6058 = ~new_n6056 & ~new_n6057;
  assign new_n6059 = new_n5960 & ~new_n5962;
  assign new_n6060 = ~new_n5963 & ~new_n6059;
  assign new_n6061 = ~new_n6046 & new_n6049;
  assign new_n6062 = ~new_n6050 & ~new_n6061;
  assign new_n6063 = ~new_n6031 & ~new_n6039;
  assign new_n6064 = ~new_n6040 & ~new_n6063;
  assign new_n6065 = ~new_n5949 & new_n5955;
  assign new_n6066 = ~new_n5956 & ~new_n6065;
  assign new_n6067 = new_n6064 & new_n6066;
  assign new_n6068 = ~new_n6062 & new_n6067;
  assign new_n6069 = new_n5956 & ~new_n5958;
  assign new_n6070 = ~new_n5959 & ~new_n6069;
  assign new_n6071 = new_n6062 & ~new_n6067;
  assign new_n6072 = ~new_n6068 & ~new_n6071;
  assign new_n6073 = ~new_n6070 & new_n6072;
  assign new_n6074 = ~new_n6068 & ~new_n6073;
  assign new_n6075 = ~new_n6060 & ~new_n6074;
  assign new_n6076 = new_n6051 & ~new_n6053;
  assign new_n6077 = ~new_n6054 & ~new_n6076;
  assign new_n6078 = new_n6060 & new_n6074;
  assign new_n6079 = ~new_n6075 & ~new_n6078;
  assign new_n6080 = ~new_n6077 & new_n6079;
  assign new_n6081 = ~new_n6075 & ~new_n6080;
  assign new_n6082 = new_n6058 & new_n6081;
  assign new_n6083 = ~new_n6058 & ~new_n6081;
  assign new_n6084 = ~new_n6082 & ~new_n6083;
  assign new_n6085 = new_n6077 & ~new_n6079;
  assign new_n6086 = ~new_n6080 & ~new_n6085;
  assign new_n6087 = new_n6070 & ~new_n6072;
  assign new_n6088 = ~new_n6073 & ~new_n6087;
  assign new_n6089 = A424 & A425;
  assign new_n6090 = ~A424 & ~A425;
  assign new_n6091 = ~new_n6089 & ~new_n6090;
  assign new_n6092 = A421 & A422;
  assign new_n6093 = ~A421 & ~A422;
  assign new_n6094 = ~new_n6092 & ~new_n6093;
  assign new_n6095 = ~A423 & A426;
  assign new_n6096 = A423 & ~A426;
  assign new_n6097 = ~new_n6095 & ~new_n6096;
  assign new_n6098 = new_n6094 & ~new_n6097;
  assign new_n6099 = ~new_n6094 & new_n6097;
  assign new_n6100 = ~new_n6098 & ~new_n6099;
  assign new_n6101 = new_n6091 & new_n6100;
  assign new_n6102 = ~new_n6091 & ~new_n6100;
  assign new_n6103 = ~new_n6101 & ~new_n6102;
  assign new_n6104 = ~A415 & ~A417;
  assign new_n6105 = A415 & A417;
  assign new_n6106 = ~new_n6104 & ~new_n6105;
  assign new_n6107 = ~A416 & new_n6106;
  assign new_n6108 = A416 & ~new_n6106;
  assign new_n6109 = ~new_n6107 & ~new_n6108;
  assign new_n6110 = ~A419 & ~A420;
  assign new_n6111 = A419 & A420;
  assign new_n6112 = ~new_n6110 & ~new_n6111;
  assign new_n6113 = ~A418 & new_n6112;
  assign new_n6114 = A418 & ~new_n6112;
  assign new_n6115 = ~new_n6113 & ~new_n6114;
  assign new_n6116 = ~new_n6109 & ~new_n6115;
  assign new_n6117 = new_n6109 & new_n6115;
  assign new_n6118 = ~new_n6116 & ~new_n6117;
  assign new_n6119 = ~new_n6103 & new_n6118;
  assign new_n6120 = new_n6103 & ~new_n6118;
  assign new_n6121 = ~new_n6119 & ~new_n6120;
  assign new_n6122 = A436 & A437;
  assign new_n6123 = ~A436 & ~A437;
  assign new_n6124 = ~new_n6122 & ~new_n6123;
  assign new_n6125 = A433 & A434;
  assign new_n6126 = ~A433 & ~A434;
  assign new_n6127 = ~new_n6125 & ~new_n6126;
  assign new_n6128 = ~A435 & A438;
  assign new_n6129 = A435 & ~A438;
  assign new_n6130 = ~new_n6128 & ~new_n6129;
  assign new_n6131 = new_n6127 & ~new_n6130;
  assign new_n6132 = ~new_n6127 & new_n6130;
  assign new_n6133 = ~new_n6131 & ~new_n6132;
  assign new_n6134 = new_n6124 & new_n6133;
  assign new_n6135 = ~new_n6124 & ~new_n6133;
  assign new_n6136 = ~new_n6134 & ~new_n6135;
  assign new_n6137 = ~A428 & ~A429;
  assign new_n6138 = A428 & A429;
  assign new_n6139 = ~new_n6137 & ~new_n6138;
  assign new_n6140 = ~A427 & new_n6139;
  assign new_n6141 = A427 & ~new_n6139;
  assign new_n6142 = ~new_n6140 & ~new_n6141;
  assign new_n6143 = ~A431 & ~A432;
  assign new_n6144 = A431 & A432;
  assign new_n6145 = ~new_n6143 & ~new_n6144;
  assign new_n6146 = ~A430 & new_n6145;
  assign new_n6147 = A430 & ~new_n6145;
  assign new_n6148 = ~new_n6146 & ~new_n6147;
  assign new_n6149 = ~new_n6142 & ~new_n6148;
  assign new_n6150 = new_n6142 & new_n6148;
  assign new_n6151 = ~new_n6149 & ~new_n6150;
  assign new_n6152 = ~new_n6136 & new_n6151;
  assign new_n6153 = new_n6136 & ~new_n6151;
  assign new_n6154 = ~new_n6152 & ~new_n6153;
  assign new_n6155 = ~new_n6121 & ~new_n6154;
  assign new_n6156 = new_n6121 & new_n6154;
  assign new_n6157 = ~new_n6155 & ~new_n6156;
  assign new_n6158 = ~new_n6064 & ~new_n6066;
  assign new_n6159 = ~new_n6067 & ~new_n6158;
  assign new_n6160 = new_n6157 & new_n6159;
  assign new_n6161 = ~new_n6088 & ~new_n6160;
  assign new_n6162 = ~new_n6110 & ~new_n6113;
  assign new_n6163 = ~new_n6104 & ~new_n6107;
  assign new_n6164 = new_n6162 & new_n6163;
  assign new_n6165 = ~new_n6162 & ~new_n6163;
  assign new_n6166 = ~new_n6164 & ~new_n6165;
  assign new_n6167 = ~new_n6117 & ~new_n6119;
  assign new_n6168 = new_n6089 & new_n6095;
  assign new_n6169 = ~A423 & ~new_n6092;
  assign new_n6170 = A426 & ~new_n6091;
  assign new_n6171 = ~A426 & ~new_n6089;
  assign new_n6172 = ~new_n6169 & ~new_n6171;
  assign new_n6173 = ~new_n6170 & new_n6172;
  assign new_n6174 = ~new_n6168 & ~new_n6173;
  assign new_n6175 = ~new_n6093 & ~new_n6174;
  assign new_n6176 = A423 & A426;
  assign new_n6177 = ~new_n6089 & ~new_n6092;
  assign new_n6178 = new_n6176 & ~new_n6177;
  assign new_n6179 = A425 & new_n6092;
  assign new_n6180 = new_n6178 & ~new_n6179;
  assign new_n6181 = new_n6090 & new_n6093;
  assign new_n6182 = ~new_n6176 & new_n6181;
  assign new_n6183 = ~new_n6090 & new_n6092;
  assign new_n6184 = new_n6096 & new_n6183;
  assign new_n6185 = ~new_n6182 & ~new_n6184;
  assign new_n6186 = ~new_n6180 & new_n6185;
  assign new_n6187 = ~new_n6175 & new_n6186;
  assign new_n6188 = new_n6169 & new_n6171;
  assign new_n6189 = ~new_n6101 & new_n6188;
  assign new_n6190 = new_n6187 & ~new_n6189;
  assign new_n6191 = ~new_n6167 & ~new_n6190;
  assign new_n6192 = new_n6167 & new_n6190;
  assign new_n6193 = ~new_n6191 & ~new_n6192;
  assign new_n6194 = ~new_n6166 & new_n6193;
  assign new_n6195 = new_n6166 & ~new_n6193;
  assign new_n6196 = ~new_n6194 & ~new_n6195;
  assign new_n6197 = ~new_n6137 & ~new_n6140;
  assign new_n6198 = ~new_n6143 & ~new_n6146;
  assign new_n6199 = new_n6197 & new_n6198;
  assign new_n6200 = ~new_n6197 & ~new_n6198;
  assign new_n6201 = ~new_n6199 & ~new_n6200;
  assign new_n6202 = ~new_n6150 & ~new_n6152;
  assign new_n6203 = new_n6122 & new_n6128;
  assign new_n6204 = ~A435 & ~new_n6125;
  assign new_n6205 = A438 & ~new_n6124;
  assign new_n6206 = ~A438 & ~new_n6122;
  assign new_n6207 = ~new_n6204 & ~new_n6206;
  assign new_n6208 = ~new_n6205 & new_n6207;
  assign new_n6209 = ~new_n6203 & ~new_n6208;
  assign new_n6210 = ~new_n6126 & ~new_n6209;
  assign new_n6211 = A435 & A438;
  assign new_n6212 = ~new_n6122 & ~new_n6125;
  assign new_n6213 = new_n6211 & ~new_n6212;
  assign new_n6214 = A437 & new_n6125;
  assign new_n6215 = new_n6213 & ~new_n6214;
  assign new_n6216 = new_n6123 & new_n6126;
  assign new_n6217 = ~new_n6211 & new_n6216;
  assign new_n6218 = ~new_n6123 & new_n6125;
  assign new_n6219 = new_n6129 & new_n6218;
  assign new_n6220 = ~new_n6217 & ~new_n6219;
  assign new_n6221 = ~new_n6215 & new_n6220;
  assign new_n6222 = ~new_n6210 & new_n6221;
  assign new_n6223 = new_n6204 & new_n6206;
  assign new_n6224 = ~new_n6134 & new_n6223;
  assign new_n6225 = new_n6222 & ~new_n6224;
  assign new_n6226 = ~new_n6202 & ~new_n6225;
  assign new_n6227 = new_n6202 & new_n6225;
  assign new_n6228 = ~new_n6226 & ~new_n6227;
  assign new_n6229 = ~new_n6201 & new_n6228;
  assign new_n6230 = new_n6201 & ~new_n6228;
  assign new_n6231 = ~new_n6229 & ~new_n6230;
  assign new_n6232 = new_n6155 & ~new_n6231;
  assign new_n6233 = ~new_n6155 & new_n6231;
  assign new_n6234 = ~new_n6232 & ~new_n6233;
  assign new_n6235 = ~new_n6196 & new_n6234;
  assign new_n6236 = new_n6196 & ~new_n6234;
  assign new_n6237 = ~new_n6235 & ~new_n6236;
  assign new_n6238 = new_n6088 & new_n6160;
  assign new_n6239 = ~new_n6161 & ~new_n6238;
  assign new_n6240 = ~new_n6237 & new_n6239;
  assign new_n6241 = ~new_n6161 & ~new_n6240;
  assign new_n6242 = new_n6086 & new_n6241;
  assign new_n6243 = ~new_n6126 & ~new_n6222;
  assign new_n6244 = ~new_n6213 & ~new_n6243;
  assign new_n6245 = new_n6149 & new_n6201;
  assign new_n6246 = ~new_n6199 & ~new_n6245;
  assign new_n6247 = ~new_n6244 & ~new_n6246;
  assign new_n6248 = new_n6244 & new_n6246;
  assign new_n6249 = ~new_n6247 & ~new_n6248;
  assign new_n6250 = ~new_n6226 & ~new_n6245;
  assign new_n6251 = ~new_n6229 & new_n6250;
  assign new_n6252 = new_n6249 & new_n6251;
  assign new_n6253 = ~new_n6249 & ~new_n6251;
  assign new_n6254 = ~new_n6252 & ~new_n6253;
  assign new_n6255 = ~new_n6093 & ~new_n6187;
  assign new_n6256 = ~new_n6178 & ~new_n6255;
  assign new_n6257 = new_n6116 & new_n6166;
  assign new_n6258 = ~new_n6164 & ~new_n6257;
  assign new_n6259 = ~new_n6256 & ~new_n6258;
  assign new_n6260 = new_n6256 & new_n6258;
  assign new_n6261 = ~new_n6259 & ~new_n6260;
  assign new_n6262 = ~new_n6191 & ~new_n6257;
  assign new_n6263 = ~new_n6194 & new_n6262;
  assign new_n6264 = new_n6261 & new_n6263;
  assign new_n6265 = ~new_n6261 & ~new_n6263;
  assign new_n6266 = ~new_n6264 & ~new_n6265;
  assign new_n6267 = ~new_n6232 & ~new_n6235;
  assign new_n6268 = new_n6266 & ~new_n6267;
  assign new_n6269 = ~new_n6266 & new_n6267;
  assign new_n6270 = ~new_n6268 & ~new_n6269;
  assign new_n6271 = new_n6254 & new_n6270;
  assign new_n6272 = ~new_n6254 & ~new_n6270;
  assign new_n6273 = ~new_n6271 & ~new_n6272;
  assign new_n6274 = ~new_n6086 & ~new_n6241;
  assign new_n6275 = ~new_n6242 & ~new_n6274;
  assign new_n6276 = new_n6273 & new_n6275;
  assign new_n6277 = ~new_n6242 & ~new_n6276;
  assign new_n6278 = new_n6084 & new_n6277;
  assign new_n6279 = ~new_n6268 & ~new_n6271;
  assign new_n6280 = ~new_n6247 & ~new_n6252;
  assign new_n6281 = ~new_n6259 & ~new_n6264;
  assign new_n6282 = ~new_n6280 & ~new_n6281;
  assign new_n6283 = new_n6280 & new_n6281;
  assign new_n6284 = ~new_n6282 & ~new_n6283;
  assign new_n6285 = ~new_n6279 & new_n6284;
  assign new_n6286 = new_n6279 & ~new_n6284;
  assign new_n6287 = ~new_n6285 & ~new_n6286;
  assign new_n6288 = ~new_n6084 & ~new_n6277;
  assign new_n6289 = ~new_n6278 & ~new_n6288;
  assign new_n6290 = ~new_n6287 & new_n6289;
  assign new_n6291 = ~new_n6278 & ~new_n6290;
  assign new_n6292 = ~new_n6056 & ~new_n6082;
  assign new_n6293 = ~new_n6282 & ~new_n6285;
  assign new_n6294 = new_n6292 & ~new_n6293;
  assign new_n6295 = ~new_n6292 & new_n6293;
  assign new_n6296 = ~new_n6294 & ~new_n6295;
  assign new_n6297 = new_n6291 & new_n6296;
  assign new_n6298 = ~new_n6291 & ~new_n6296;
  assign new_n6299 = ~new_n6297 & ~new_n6298;
  assign new_n6300 = A385 & A386;
  assign new_n6301 = A388 & A389;
  assign new_n6302 = ~new_n6300 & ~new_n6301;
  assign new_n6303 = A387 & A390;
  assign new_n6304 = ~new_n6302 & new_n6303;
  assign new_n6305 = ~A385 & ~A386;
  assign new_n6306 = ~A387 & A390;
  assign new_n6307 = new_n6301 & new_n6306;
  assign new_n6308 = ~A387 & ~new_n6300;
  assign new_n6309 = ~A388 & ~A389;
  assign new_n6310 = ~new_n6301 & ~new_n6309;
  assign new_n6311 = A390 & ~new_n6310;
  assign new_n6312 = ~A390 & ~new_n6301;
  assign new_n6313 = ~new_n6308 & ~new_n6312;
  assign new_n6314 = ~new_n6311 & new_n6313;
  assign new_n6315 = ~new_n6307 & ~new_n6314;
  assign new_n6316 = ~new_n6305 & ~new_n6315;
  assign new_n6317 = A389 & new_n6300;
  assign new_n6318 = new_n6304 & ~new_n6317;
  assign new_n6319 = ~new_n6303 & new_n6305;
  assign new_n6320 = new_n6309 & new_n6319;
  assign new_n6321 = A387 & ~A390;
  assign new_n6322 = new_n6300 & ~new_n6309;
  assign new_n6323 = new_n6321 & new_n6322;
  assign new_n6324 = ~new_n6320 & ~new_n6323;
  assign new_n6325 = ~new_n6318 & new_n6324;
  assign new_n6326 = ~new_n6316 & new_n6325;
  assign new_n6327 = ~new_n6305 & ~new_n6326;
  assign new_n6328 = ~new_n6304 & ~new_n6327;
  assign new_n6329 = ~A380 & ~A381;
  assign new_n6330 = A380 & A381;
  assign new_n6331 = ~new_n6329 & ~new_n6330;
  assign new_n6332 = ~A379 & new_n6331;
  assign new_n6333 = ~new_n6329 & ~new_n6332;
  assign new_n6334 = ~A383 & ~A384;
  assign new_n6335 = A383 & A384;
  assign new_n6336 = ~new_n6334 & ~new_n6335;
  assign new_n6337 = ~A382 & new_n6336;
  assign new_n6338 = ~new_n6334 & ~new_n6337;
  assign new_n6339 = new_n6333 & new_n6338;
  assign new_n6340 = A379 & ~new_n6331;
  assign new_n6341 = ~new_n6332 & ~new_n6340;
  assign new_n6342 = A382 & ~new_n6336;
  assign new_n6343 = ~new_n6337 & ~new_n6342;
  assign new_n6344 = ~new_n6341 & ~new_n6343;
  assign new_n6345 = ~new_n6333 & ~new_n6338;
  assign new_n6346 = ~new_n6339 & ~new_n6345;
  assign new_n6347 = new_n6344 & new_n6346;
  assign new_n6348 = ~new_n6339 & ~new_n6347;
  assign new_n6349 = ~new_n6328 & ~new_n6348;
  assign new_n6350 = new_n6328 & new_n6348;
  assign new_n6351 = ~new_n6349 & ~new_n6350;
  assign new_n6352 = new_n6341 & new_n6343;
  assign new_n6353 = ~new_n6300 & ~new_n6305;
  assign new_n6354 = ~new_n6306 & ~new_n6321;
  assign new_n6355 = new_n6353 & ~new_n6354;
  assign new_n6356 = ~new_n6353 & new_n6354;
  assign new_n6357 = ~new_n6355 & ~new_n6356;
  assign new_n6358 = new_n6310 & new_n6357;
  assign new_n6359 = ~new_n6310 & ~new_n6357;
  assign new_n6360 = ~new_n6358 & ~new_n6359;
  assign new_n6361 = ~new_n6344 & ~new_n6352;
  assign new_n6362 = ~new_n6360 & new_n6361;
  assign new_n6363 = ~new_n6352 & ~new_n6362;
  assign new_n6364 = new_n6308 & new_n6312;
  assign new_n6365 = ~new_n6358 & new_n6364;
  assign new_n6366 = new_n6326 & ~new_n6365;
  assign new_n6367 = ~new_n6363 & ~new_n6366;
  assign new_n6368 = new_n6363 & new_n6366;
  assign new_n6369 = ~new_n6367 & ~new_n6368;
  assign new_n6370 = ~new_n6346 & new_n6369;
  assign new_n6371 = ~new_n6347 & ~new_n6367;
  assign new_n6372 = ~new_n6370 & new_n6371;
  assign new_n6373 = new_n6351 & new_n6372;
  assign new_n6374 = ~new_n6349 & ~new_n6373;
  assign new_n6375 = A373 & A374;
  assign new_n6376 = A376 & A377;
  assign new_n6377 = ~new_n6375 & ~new_n6376;
  assign new_n6378 = A375 & A378;
  assign new_n6379 = ~new_n6377 & new_n6378;
  assign new_n6380 = ~A373 & ~A374;
  assign new_n6381 = ~A375 & A378;
  assign new_n6382 = new_n6376 & new_n6381;
  assign new_n6383 = ~A375 & ~new_n6375;
  assign new_n6384 = ~A376 & ~A377;
  assign new_n6385 = ~new_n6376 & ~new_n6384;
  assign new_n6386 = A378 & ~new_n6385;
  assign new_n6387 = ~A378 & ~new_n6376;
  assign new_n6388 = ~new_n6383 & ~new_n6387;
  assign new_n6389 = ~new_n6386 & new_n6388;
  assign new_n6390 = ~new_n6382 & ~new_n6389;
  assign new_n6391 = ~new_n6380 & ~new_n6390;
  assign new_n6392 = A377 & new_n6375;
  assign new_n6393 = new_n6379 & ~new_n6392;
  assign new_n6394 = ~new_n6378 & new_n6380;
  assign new_n6395 = new_n6384 & new_n6394;
  assign new_n6396 = A375 & ~A378;
  assign new_n6397 = new_n6375 & ~new_n6384;
  assign new_n6398 = new_n6396 & new_n6397;
  assign new_n6399 = ~new_n6395 & ~new_n6398;
  assign new_n6400 = ~new_n6393 & new_n6399;
  assign new_n6401 = ~new_n6391 & new_n6400;
  assign new_n6402 = ~new_n6380 & ~new_n6401;
  assign new_n6403 = ~new_n6379 & ~new_n6402;
  assign new_n6404 = ~A368 & ~A369;
  assign new_n6405 = A368 & A369;
  assign new_n6406 = ~new_n6404 & ~new_n6405;
  assign new_n6407 = ~A367 & new_n6406;
  assign new_n6408 = ~new_n6404 & ~new_n6407;
  assign new_n6409 = ~A371 & ~A372;
  assign new_n6410 = A371 & A372;
  assign new_n6411 = ~new_n6409 & ~new_n6410;
  assign new_n6412 = ~A370 & new_n6411;
  assign new_n6413 = ~new_n6409 & ~new_n6412;
  assign new_n6414 = new_n6408 & new_n6413;
  assign new_n6415 = A367 & ~new_n6406;
  assign new_n6416 = ~new_n6407 & ~new_n6415;
  assign new_n6417 = A370 & ~new_n6411;
  assign new_n6418 = ~new_n6412 & ~new_n6417;
  assign new_n6419 = ~new_n6416 & ~new_n6418;
  assign new_n6420 = ~new_n6408 & ~new_n6413;
  assign new_n6421 = ~new_n6414 & ~new_n6420;
  assign new_n6422 = new_n6419 & new_n6421;
  assign new_n6423 = ~new_n6414 & ~new_n6422;
  assign new_n6424 = ~new_n6403 & ~new_n6423;
  assign new_n6425 = new_n6403 & new_n6423;
  assign new_n6426 = ~new_n6424 & ~new_n6425;
  assign new_n6427 = new_n6416 & new_n6418;
  assign new_n6428 = ~new_n6375 & ~new_n6380;
  assign new_n6429 = ~new_n6381 & ~new_n6396;
  assign new_n6430 = new_n6428 & ~new_n6429;
  assign new_n6431 = ~new_n6428 & new_n6429;
  assign new_n6432 = ~new_n6430 & ~new_n6431;
  assign new_n6433 = new_n6385 & new_n6432;
  assign new_n6434 = ~new_n6385 & ~new_n6432;
  assign new_n6435 = ~new_n6433 & ~new_n6434;
  assign new_n6436 = ~new_n6419 & ~new_n6427;
  assign new_n6437 = ~new_n6435 & new_n6436;
  assign new_n6438 = ~new_n6427 & ~new_n6437;
  assign new_n6439 = new_n6383 & new_n6387;
  assign new_n6440 = ~new_n6433 & new_n6439;
  assign new_n6441 = new_n6401 & ~new_n6440;
  assign new_n6442 = ~new_n6438 & ~new_n6441;
  assign new_n6443 = new_n6438 & new_n6441;
  assign new_n6444 = ~new_n6442 & ~new_n6443;
  assign new_n6445 = ~new_n6421 & new_n6444;
  assign new_n6446 = ~new_n6422 & ~new_n6442;
  assign new_n6447 = ~new_n6445 & new_n6446;
  assign new_n6448 = new_n6426 & new_n6447;
  assign new_n6449 = ~new_n6424 & ~new_n6448;
  assign new_n6450 = new_n6374 & new_n6449;
  assign new_n6451 = ~new_n6374 & ~new_n6449;
  assign new_n6452 = ~new_n6450 & ~new_n6451;
  assign new_n6453 = ~new_n6426 & ~new_n6447;
  assign new_n6454 = ~new_n6448 & ~new_n6453;
  assign new_n6455 = new_n6346 & ~new_n6369;
  assign new_n6456 = ~new_n6370 & ~new_n6455;
  assign new_n6457 = new_n6421 & ~new_n6444;
  assign new_n6458 = ~new_n6445 & ~new_n6457;
  assign new_n6459 = new_n6456 & new_n6458;
  assign new_n6460 = ~new_n6456 & ~new_n6458;
  assign new_n6461 = new_n6360 & ~new_n6361;
  assign new_n6462 = ~new_n6362 & ~new_n6461;
  assign new_n6463 = new_n6435 & ~new_n6436;
  assign new_n6464 = ~new_n6437 & ~new_n6463;
  assign new_n6465 = ~new_n6462 & ~new_n6464;
  assign new_n6466 = ~new_n6460 & ~new_n6465;
  assign new_n6467 = ~new_n6459 & ~new_n6466;
  assign new_n6468 = new_n6454 & new_n6467;
  assign new_n6469 = ~new_n6351 & ~new_n6372;
  assign new_n6470 = ~new_n6373 & ~new_n6469;
  assign new_n6471 = ~new_n6454 & ~new_n6467;
  assign new_n6472 = ~new_n6468 & ~new_n6471;
  assign new_n6473 = new_n6470 & new_n6472;
  assign new_n6474 = ~new_n6468 & ~new_n6473;
  assign new_n6475 = new_n6452 & new_n6474;
  assign new_n6476 = ~new_n6452 & ~new_n6474;
  assign new_n6477 = ~new_n6475 & ~new_n6476;
  assign new_n6478 = A411 & A414;
  assign new_n6479 = A409 & A410;
  assign new_n6480 = A412 & A413;
  assign new_n6481 = ~new_n6479 & ~new_n6480;
  assign new_n6482 = new_n6478 & ~new_n6481;
  assign new_n6483 = ~A409 & ~A410;
  assign new_n6484 = ~A411 & A414;
  assign new_n6485 = new_n6480 & new_n6484;
  assign new_n6486 = ~A411 & ~new_n6479;
  assign new_n6487 = ~A412 & ~A413;
  assign new_n6488 = ~new_n6480 & ~new_n6487;
  assign new_n6489 = A414 & ~new_n6488;
  assign new_n6490 = ~A414 & ~new_n6480;
  assign new_n6491 = ~new_n6486 & ~new_n6490;
  assign new_n6492 = ~new_n6489 & new_n6491;
  assign new_n6493 = ~new_n6485 & ~new_n6492;
  assign new_n6494 = ~new_n6483 & ~new_n6493;
  assign new_n6495 = A413 & new_n6479;
  assign new_n6496 = new_n6482 & ~new_n6495;
  assign new_n6497 = ~new_n6478 & new_n6483;
  assign new_n6498 = new_n6487 & new_n6497;
  assign new_n6499 = A411 & ~A414;
  assign new_n6500 = new_n6479 & ~new_n6487;
  assign new_n6501 = new_n6499 & new_n6500;
  assign new_n6502 = ~new_n6498 & ~new_n6501;
  assign new_n6503 = ~new_n6496 & new_n6502;
  assign new_n6504 = ~new_n6494 & new_n6503;
  assign new_n6505 = ~new_n6483 & ~new_n6504;
  assign new_n6506 = ~new_n6482 & ~new_n6505;
  assign new_n6507 = ~A404 & ~A405;
  assign new_n6508 = A404 & A405;
  assign new_n6509 = ~new_n6507 & ~new_n6508;
  assign new_n6510 = ~A403 & new_n6509;
  assign new_n6511 = ~new_n6507 & ~new_n6510;
  assign new_n6512 = ~A407 & ~A408;
  assign new_n6513 = A407 & A408;
  assign new_n6514 = ~new_n6512 & ~new_n6513;
  assign new_n6515 = ~A406 & new_n6514;
  assign new_n6516 = ~new_n6512 & ~new_n6515;
  assign new_n6517 = new_n6511 & new_n6516;
  assign new_n6518 = A403 & ~new_n6509;
  assign new_n6519 = ~new_n6510 & ~new_n6518;
  assign new_n6520 = A406 & ~new_n6514;
  assign new_n6521 = ~new_n6515 & ~new_n6520;
  assign new_n6522 = ~new_n6519 & ~new_n6521;
  assign new_n6523 = ~new_n6511 & ~new_n6516;
  assign new_n6524 = ~new_n6517 & ~new_n6523;
  assign new_n6525 = new_n6522 & new_n6524;
  assign new_n6526 = ~new_n6517 & ~new_n6525;
  assign new_n6527 = ~new_n6506 & ~new_n6526;
  assign new_n6528 = new_n6506 & new_n6526;
  assign new_n6529 = ~new_n6527 & ~new_n6528;
  assign new_n6530 = ~new_n6479 & ~new_n6483;
  assign new_n6531 = ~new_n6484 & ~new_n6499;
  assign new_n6532 = new_n6530 & ~new_n6531;
  assign new_n6533 = ~new_n6530 & new_n6531;
  assign new_n6534 = ~new_n6532 & ~new_n6533;
  assign new_n6535 = new_n6488 & new_n6534;
  assign new_n6536 = new_n6486 & new_n6490;
  assign new_n6537 = ~new_n6535 & new_n6536;
  assign new_n6538 = new_n6504 & ~new_n6537;
  assign new_n6539 = ~new_n6524 & ~new_n6538;
  assign new_n6540 = new_n6519 & new_n6521;
  assign new_n6541 = ~new_n6488 & ~new_n6534;
  assign new_n6542 = ~new_n6535 & ~new_n6541;
  assign new_n6543 = ~new_n6522 & ~new_n6540;
  assign new_n6544 = ~new_n6542 & new_n6543;
  assign new_n6545 = ~new_n6540 & ~new_n6544;
  assign new_n6546 = new_n6524 & new_n6538;
  assign new_n6547 = ~new_n6539 & ~new_n6546;
  assign new_n6548 = ~new_n6545 & new_n6547;
  assign new_n6549 = ~new_n6525 & ~new_n6539;
  assign new_n6550 = ~new_n6548 & new_n6549;
  assign new_n6551 = new_n6529 & new_n6550;
  assign new_n6552 = ~new_n6527 & ~new_n6551;
  assign new_n6553 = A393 & A396;
  assign new_n6554 = A391 & A392;
  assign new_n6555 = A394 & A395;
  assign new_n6556 = ~new_n6554 & ~new_n6555;
  assign new_n6557 = new_n6553 & ~new_n6556;
  assign new_n6558 = ~A391 & ~A392;
  assign new_n6559 = ~A393 & A396;
  assign new_n6560 = new_n6555 & new_n6559;
  assign new_n6561 = ~A393 & ~new_n6554;
  assign new_n6562 = ~A394 & ~A395;
  assign new_n6563 = ~new_n6555 & ~new_n6562;
  assign new_n6564 = A396 & ~new_n6563;
  assign new_n6565 = ~A396 & ~new_n6555;
  assign new_n6566 = ~new_n6561 & ~new_n6565;
  assign new_n6567 = ~new_n6564 & new_n6566;
  assign new_n6568 = ~new_n6560 & ~new_n6567;
  assign new_n6569 = ~new_n6558 & ~new_n6568;
  assign new_n6570 = A395 & new_n6554;
  assign new_n6571 = new_n6557 & ~new_n6570;
  assign new_n6572 = ~new_n6553 & new_n6558;
  assign new_n6573 = new_n6562 & new_n6572;
  assign new_n6574 = A393 & ~A396;
  assign new_n6575 = new_n6554 & ~new_n6562;
  assign new_n6576 = new_n6574 & new_n6575;
  assign new_n6577 = ~new_n6573 & ~new_n6576;
  assign new_n6578 = ~new_n6571 & new_n6577;
  assign new_n6579 = ~new_n6569 & new_n6578;
  assign new_n6580 = ~new_n6558 & ~new_n6579;
  assign new_n6581 = ~new_n6557 & ~new_n6580;
  assign new_n6582 = ~A397 & ~A399;
  assign new_n6583 = A397 & A399;
  assign new_n6584 = ~new_n6582 & ~new_n6583;
  assign new_n6585 = ~A398 & new_n6584;
  assign new_n6586 = ~new_n6582 & ~new_n6585;
  assign new_n6587 = ~A400 & ~A401;
  assign new_n6588 = new_n6586 & ~new_n6587;
  assign new_n6589 = A400 & A401;
  assign new_n6590 = ~A402 & ~new_n6589;
  assign new_n6591 = new_n6588 & ~new_n6590;
  assign new_n6592 = ~A402 & ~new_n6588;
  assign new_n6593 = A398 & ~new_n6584;
  assign new_n6594 = ~new_n6585 & ~new_n6593;
  assign new_n6595 = ~new_n6586 & ~new_n6589;
  assign new_n6596 = new_n6586 & new_n6589;
  assign new_n6597 = ~new_n6595 & ~new_n6596;
  assign new_n6598 = A402 & ~new_n6597;
  assign new_n6599 = ~new_n6592 & ~new_n6594;
  assign new_n6600 = ~new_n6598 & new_n6599;
  assign new_n6601 = ~new_n6591 & ~new_n6600;
  assign new_n6602 = new_n6581 & new_n6601;
  assign new_n6603 = ~new_n6554 & ~new_n6558;
  assign new_n6604 = ~new_n6559 & ~new_n6574;
  assign new_n6605 = new_n6603 & ~new_n6604;
  assign new_n6606 = ~new_n6603 & new_n6604;
  assign new_n6607 = ~new_n6605 & ~new_n6606;
  assign new_n6608 = new_n6563 & new_n6607;
  assign new_n6609 = new_n6561 & new_n6565;
  assign new_n6610 = ~new_n6608 & new_n6609;
  assign new_n6611 = new_n6579 & ~new_n6610;
  assign new_n6612 = A402 & ~new_n6594;
  assign new_n6613 = ~new_n6586 & new_n6587;
  assign new_n6614 = ~new_n6612 & new_n6613;
  assign new_n6615 = ~new_n6586 & new_n6590;
  assign new_n6616 = ~new_n6591 & ~new_n6615;
  assign new_n6617 = new_n6594 & ~new_n6616;
  assign new_n6618 = ~new_n6600 & ~new_n6614;
  assign new_n6619 = ~new_n6617 & new_n6618;
  assign new_n6620 = ~new_n6611 & ~new_n6619;
  assign new_n6621 = ~new_n6563 & ~new_n6607;
  assign new_n6622 = ~new_n6608 & ~new_n6621;
  assign new_n6623 = ~A402 & new_n6594;
  assign new_n6624 = ~new_n6612 & ~new_n6623;
  assign new_n6625 = ~new_n6587 & ~new_n6589;
  assign new_n6626 = ~new_n6624 & new_n6625;
  assign new_n6627 = new_n6624 & ~new_n6625;
  assign new_n6628 = ~new_n6626 & ~new_n6627;
  assign new_n6629 = new_n6622 & ~new_n6628;
  assign new_n6630 = new_n6611 & new_n6619;
  assign new_n6631 = ~new_n6620 & ~new_n6630;
  assign new_n6632 = ~new_n6629 & new_n6631;
  assign new_n6633 = ~new_n6620 & ~new_n6632;
  assign new_n6634 = ~new_n6581 & ~new_n6601;
  assign new_n6635 = ~new_n6602 & ~new_n6634;
  assign new_n6636 = ~new_n6633 & new_n6635;
  assign new_n6637 = ~new_n6602 & ~new_n6636;
  assign new_n6638 = ~new_n6552 & new_n6637;
  assign new_n6639 = new_n6552 & ~new_n6637;
  assign new_n6640 = ~new_n6638 & ~new_n6639;
  assign new_n6641 = new_n6633 & ~new_n6635;
  assign new_n6642 = ~new_n6636 & ~new_n6641;
  assign new_n6643 = ~new_n6622 & new_n6628;
  assign new_n6644 = ~new_n6629 & ~new_n6643;
  assign new_n6645 = new_n6542 & ~new_n6543;
  assign new_n6646 = ~new_n6544 & ~new_n6645;
  assign new_n6647 = new_n6644 & ~new_n6646;
  assign new_n6648 = new_n6631 & new_n6647;
  assign new_n6649 = new_n6545 & ~new_n6547;
  assign new_n6650 = ~new_n6548 & ~new_n6649;
  assign new_n6651 = ~new_n6629 & ~new_n6647;
  assign new_n6652 = new_n6631 & ~new_n6651;
  assign new_n6653 = ~new_n6631 & new_n6651;
  assign new_n6654 = ~new_n6652 & ~new_n6653;
  assign new_n6655 = ~new_n6650 & new_n6654;
  assign new_n6656 = ~new_n6648 & ~new_n6655;
  assign new_n6657 = ~new_n6642 & ~new_n6656;
  assign new_n6658 = ~new_n6529 & ~new_n6550;
  assign new_n6659 = ~new_n6551 & ~new_n6658;
  assign new_n6660 = new_n6642 & new_n6656;
  assign new_n6661 = ~new_n6657 & ~new_n6660;
  assign new_n6662 = new_n6659 & new_n6661;
  assign new_n6663 = ~new_n6657 & ~new_n6662;
  assign new_n6664 = new_n6640 & ~new_n6663;
  assign new_n6665 = ~new_n6640 & new_n6663;
  assign new_n6666 = ~new_n6664 & ~new_n6665;
  assign new_n6667 = new_n6650 & ~new_n6654;
  assign new_n6668 = ~new_n6655 & ~new_n6667;
  assign new_n6669 = ~new_n6459 & ~new_n6460;
  assign new_n6670 = ~new_n6644 & new_n6646;
  assign new_n6671 = ~new_n6647 & ~new_n6670;
  assign new_n6672 = new_n6462 & new_n6464;
  assign new_n6673 = ~new_n6465 & ~new_n6672;
  assign new_n6674 = new_n6671 & new_n6673;
  assign new_n6675 = ~new_n6465 & ~new_n6674;
  assign new_n6676 = new_n6669 & ~new_n6675;
  assign new_n6677 = ~new_n6669 & new_n6675;
  assign new_n6678 = ~new_n6676 & ~new_n6677;
  assign new_n6679 = ~new_n6668 & new_n6678;
  assign new_n6680 = ~new_n6674 & ~new_n6678;
  assign new_n6681 = ~new_n6679 & ~new_n6680;
  assign new_n6682 = ~new_n6659 & ~new_n6661;
  assign new_n6683 = ~new_n6662 & ~new_n6682;
  assign new_n6684 = ~new_n6681 & ~new_n6683;
  assign new_n6685 = ~new_n6470 & ~new_n6472;
  assign new_n6686 = ~new_n6473 & ~new_n6685;
  assign new_n6687 = new_n6681 & new_n6683;
  assign new_n6688 = ~new_n6684 & ~new_n6687;
  assign new_n6689 = ~new_n6686 & new_n6688;
  assign new_n6690 = ~new_n6684 & ~new_n6689;
  assign new_n6691 = ~new_n6666 & ~new_n6690;
  assign new_n6692 = new_n6666 & new_n6690;
  assign new_n6693 = ~new_n6691 & ~new_n6692;
  assign new_n6694 = new_n6477 & new_n6693;
  assign new_n6695 = ~new_n6477 & ~new_n6693;
  assign new_n6696 = ~new_n6694 & ~new_n6695;
  assign new_n6697 = new_n6287 & ~new_n6289;
  assign new_n6698 = ~new_n6290 & ~new_n6697;
  assign new_n6699 = ~new_n6696 & ~new_n6698;
  assign new_n6700 = new_n6696 & new_n6698;
  assign new_n6701 = ~new_n6699 & ~new_n6700;
  assign new_n6702 = ~new_n6273 & ~new_n6275;
  assign new_n6703 = ~new_n6276 & ~new_n6702;
  assign new_n6704 = new_n6668 & ~new_n6678;
  assign new_n6705 = ~new_n6679 & ~new_n6704;
  assign new_n6706 = new_n6237 & ~new_n6239;
  assign new_n6707 = ~new_n6240 & ~new_n6706;
  assign new_n6708 = ~new_n6705 & ~new_n6707;
  assign new_n6709 = new_n6705 & new_n6707;
  assign new_n6710 = ~new_n6671 & ~new_n6673;
  assign new_n6711 = ~new_n6674 & ~new_n6710;
  assign new_n6712 = ~new_n6157 & ~new_n6159;
  assign new_n6713 = ~new_n6160 & ~new_n6712;
  assign new_n6714 = new_n6711 & new_n6713;
  assign new_n6715 = ~new_n6709 & new_n6714;
  assign new_n6716 = ~new_n6708 & ~new_n6715;
  assign new_n6717 = new_n6703 & ~new_n6716;
  assign new_n6718 = new_n6686 & ~new_n6688;
  assign new_n6719 = ~new_n6689 & ~new_n6718;
  assign new_n6720 = ~new_n6703 & new_n6716;
  assign new_n6721 = ~new_n6717 & ~new_n6720;
  assign new_n6722 = ~new_n6719 & new_n6721;
  assign new_n6723 = ~new_n6717 & ~new_n6722;
  assign new_n6724 = new_n6701 & ~new_n6723;
  assign new_n6725 = ~new_n6699 & ~new_n6724;
  assign new_n6726 = new_n6299 & ~new_n6725;
  assign new_n6727 = ~new_n6691 & ~new_n6694;
  assign new_n6728 = ~new_n6450 & ~new_n6475;
  assign new_n6729 = ~new_n6638 & ~new_n6664;
  assign new_n6730 = new_n6728 & ~new_n6729;
  assign new_n6731 = ~new_n6728 & new_n6729;
  assign new_n6732 = ~new_n6730 & ~new_n6731;
  assign new_n6733 = new_n6727 & new_n6732;
  assign new_n6734 = ~new_n6727 & ~new_n6732;
  assign new_n6735 = ~new_n6733 & ~new_n6734;
  assign new_n6736 = ~new_n6299 & new_n6725;
  assign new_n6737 = ~new_n6726 & ~new_n6736;
  assign new_n6738 = new_n6735 & new_n6737;
  assign new_n6739 = ~new_n6726 & ~new_n6738;
  assign new_n6740 = ~new_n6294 & ~new_n6297;
  assign new_n6741 = ~new_n6730 & ~new_n6733;
  assign new_n6742 = ~new_n6740 & ~new_n6741;
  assign new_n6743 = new_n6740 & new_n6741;
  assign new_n6744 = ~new_n6742 & ~new_n6743;
  assign new_n6745 = ~new_n6739 & new_n6744;
  assign new_n6746 = new_n6739 & ~new_n6744;
  assign new_n6747 = ~new_n6745 & ~new_n6746;
  assign new_n6748 = ~new_n5879 & new_n6747;
  assign new_n6749 = new_n5879 & ~new_n6747;
  assign new_n6750 = ~new_n6748 & ~new_n6749;
  assign new_n6751 = ~new_n6735 & ~new_n6737;
  assign new_n6752 = ~new_n6738 & ~new_n6751;
  assign new_n6753 = new_n5867 & ~new_n5869;
  assign new_n6754 = ~new_n5870 & ~new_n6753;
  assign new_n6755 = ~new_n6752 & new_n6754;
  assign new_n6756 = new_n6752 & ~new_n6754;
  assign new_n6757 = ~new_n6755 & ~new_n6756;
  assign new_n6758 = ~new_n6701 & new_n6723;
  assign new_n6759 = ~new_n6724 & ~new_n6758;
  assign new_n6760 = new_n5853 & ~new_n5855;
  assign new_n6761 = ~new_n5856 & ~new_n6760;
  assign new_n6762 = new_n6759 & new_n6761;
  assign new_n6763 = ~new_n5823 & ~new_n5825;
  assign new_n6764 = ~new_n5826 & ~new_n6763;
  assign new_n6765 = new_n6719 & ~new_n6721;
  assign new_n6766 = ~new_n6722 & ~new_n6765;
  assign new_n6767 = ~new_n6764 & ~new_n6766;
  assign new_n6768 = new_n6764 & new_n6766;
  assign new_n6769 = ~new_n6767 & ~new_n6768;
  assign new_n6770 = new_n5816 & ~new_n5818;
  assign new_n6771 = ~new_n5819 & ~new_n6770;
  assign new_n6772 = ~new_n6708 & ~new_n6709;
  assign new_n6773 = ~new_n6711 & ~new_n6713;
  assign new_n6774 = ~new_n6714 & ~new_n6773;
  assign new_n6775 = ~new_n5810 & ~new_n5812;
  assign new_n6776 = ~new_n5813 & ~new_n6775;
  assign new_n6777 = new_n6774 & new_n6776;
  assign new_n6778 = ~new_n6714 & ~new_n6777;
  assign new_n6779 = new_n6772 & ~new_n6778;
  assign new_n6780 = ~new_n6772 & new_n6778;
  assign new_n6781 = ~new_n6779 & ~new_n6780;
  assign new_n6782 = ~new_n6771 & new_n6781;
  assign new_n6783 = new_n6772 & new_n6777;
  assign new_n6784 = ~new_n6782 & ~new_n6783;
  assign new_n6785 = new_n6769 & new_n6784;
  assign new_n6786 = ~new_n6767 & ~new_n6785;
  assign new_n6787 = ~new_n6759 & ~new_n6761;
  assign new_n6788 = ~new_n6762 & ~new_n6787;
  assign new_n6789 = new_n6786 & new_n6788;
  assign new_n6790 = ~new_n6762 & ~new_n6789;
  assign new_n6791 = new_n6757 & new_n6790;
  assign new_n6792 = ~new_n6755 & ~new_n6791;
  assign new_n6793 = new_n6750 & new_n6792;
  assign new_n6794 = ~new_n6750 & ~new_n6792;
  assign new_n6795 = ~new_n6793 & ~new_n6794;
  assign new_n6796 = ~new_n6757 & ~new_n6790;
  assign new_n6797 = ~new_n6791 & ~new_n6796;
  assign new_n6798 = ~new_n4988 & ~new_n4990;
  assign new_n6799 = ~new_n4991 & ~new_n6798;
  assign new_n6800 = ~new_n6786 & ~new_n6788;
  assign new_n6801 = ~new_n6789 & ~new_n6800;
  assign new_n6802 = new_n6799 & new_n6801;
  assign new_n6803 = ~new_n6799 & ~new_n6801;
  assign new_n6804 = ~new_n6802 & ~new_n6803;
  assign new_n6805 = new_n4984 & ~new_n4986;
  assign new_n6806 = ~new_n4987 & ~new_n6805;
  assign new_n6807 = new_n6771 & ~new_n6781;
  assign new_n6808 = ~new_n6782 & ~new_n6807;
  assign new_n6809 = new_n4977 & ~new_n4979;
  assign new_n6810 = ~new_n4980 & ~new_n6809;
  assign new_n6811 = ~new_n6808 & new_n6810;
  assign new_n6812 = new_n6808 & ~new_n6810;
  assign new_n6813 = ~new_n6774 & ~new_n6776;
  assign new_n6814 = ~new_n6777 & ~new_n6813;
  assign new_n6815 = ~new_n4971 & ~new_n4973;
  assign new_n6816 = ~new_n4974 & ~new_n6815;
  assign new_n6817 = new_n6814 & new_n6816;
  assign new_n6818 = ~new_n6812 & ~new_n6817;
  assign new_n6819 = ~new_n6811 & ~new_n6818;
  assign new_n6820 = new_n6806 & ~new_n6819;
  assign new_n6821 = ~new_n6769 & ~new_n6784;
  assign new_n6822 = ~new_n6785 & ~new_n6821;
  assign new_n6823 = ~new_n6806 & new_n6819;
  assign new_n6824 = ~new_n6820 & ~new_n6823;
  assign new_n6825 = new_n6822 & new_n6824;
  assign new_n6826 = ~new_n6820 & ~new_n6825;
  assign new_n6827 = new_n6804 & new_n6826;
  assign new_n6828 = ~new_n6802 & ~new_n6827;
  assign new_n6829 = new_n6797 & new_n6828;
  assign new_n6830 = ~new_n4960 & ~new_n4992;
  assign new_n6831 = ~new_n4993 & ~new_n6830;
  assign new_n6832 = ~new_n6797 & ~new_n6828;
  assign new_n6833 = ~new_n6829 & ~new_n6832;
  assign new_n6834 = new_n6831 & new_n6833;
  assign new_n6835 = ~new_n6829 & ~new_n6834;
  assign new_n6836 = new_n6795 & new_n6835;
  assign new_n6837 = ~new_n5004 & ~new_n5006;
  assign new_n6838 = ~new_n5007 & ~new_n6837;
  assign new_n6839 = ~new_n6795 & ~new_n6835;
  assign new_n6840 = ~new_n6836 & ~new_n6839;
  assign new_n6841 = ~new_n6838 & new_n6840;
  assign new_n6842 = ~new_n6836 & ~new_n6841;
  assign new_n6843 = new_n5016 & ~new_n6842;
  assign new_n6844 = ~new_n6748 & ~new_n6793;
  assign new_n6845 = ~new_n5874 & ~new_n5877;
  assign new_n6846 = ~new_n6742 & ~new_n6745;
  assign new_n6847 = new_n6845 & ~new_n6846;
  assign new_n6848 = ~new_n6845 & new_n6846;
  assign new_n6849 = ~new_n6847 & ~new_n6848;
  assign new_n6850 = ~new_n6844 & new_n6849;
  assign new_n6851 = new_n6844 & ~new_n6849;
  assign new_n6852 = ~new_n6850 & ~new_n6851;
  assign new_n6853 = ~new_n5016 & new_n6842;
  assign new_n6854 = ~new_n6843 & ~new_n6853;
  assign new_n6855 = new_n6852 & new_n6854;
  assign new_n6856 = ~new_n6843 & ~new_n6855;
  assign new_n6857 = ~new_n6847 & ~new_n6850;
  assign new_n6858 = ~new_n5011 & ~new_n5014;
  assign new_n6859 = new_n6857 & new_n6858;
  assign new_n6860 = ~new_n6857 & ~new_n6858;
  assign new_n6861 = ~new_n6859 & ~new_n6860;
  assign new_n6862 = new_n6856 & new_n6861;
  assign new_n6863 = ~new_n6856 & ~new_n6861;
  assign new_n6864 = ~new_n6862 & ~new_n6863;
  assign new_n6865 = new_n3273 & new_n6864;
  assign new_n6866 = ~new_n3273 & ~new_n6864;
  assign new_n6867 = ~new_n6865 & ~new_n6866;
  assign new_n6868 = ~new_n6852 & ~new_n6854;
  assign new_n6869 = ~new_n6855 & ~new_n6868;
  assign new_n6870 = new_n6838 & ~new_n6840;
  assign new_n6871 = ~new_n6841 & ~new_n6870;
  assign new_n6872 = ~new_n6831 & ~new_n6833;
  assign new_n6873 = ~new_n6834 & ~new_n6872;
  assign new_n6874 = ~new_n3244 & ~new_n3246;
  assign new_n6875 = ~new_n3247 & ~new_n6874;
  assign new_n6876 = ~new_n6873 & ~new_n6875;
  assign new_n6877 = new_n6873 & new_n6875;
  assign new_n6878 = ~new_n6876 & ~new_n6877;
  assign new_n6879 = ~new_n6804 & ~new_n6826;
  assign new_n6880 = ~new_n6827 & ~new_n6879;
  assign new_n6881 = ~new_n6822 & ~new_n6824;
  assign new_n6882 = ~new_n6825 & ~new_n6881;
  assign new_n6883 = new_n3150 & ~new_n3152;
  assign new_n6884 = ~new_n3153 & ~new_n6883;
  assign new_n6885 = new_n6882 & ~new_n6884;
  assign new_n6886 = ~new_n6882 & new_n6884;
  assign new_n6887 = ~new_n6885 & ~new_n6886;
  assign new_n6888 = ~new_n3142 & ~new_n3144;
  assign new_n6889 = ~new_n3145 & ~new_n6888;
  assign new_n6890 = ~new_n6811 & ~new_n6812;
  assign new_n6891 = ~new_n6814 & ~new_n6816;
  assign new_n6892 = ~new_n6817 & ~new_n6891;
  assign new_n6893 = new_n3136 & ~new_n3137;
  assign new_n6894 = ~new_n3138 & ~new_n6893;
  assign new_n6895 = new_n6892 & ~new_n6894;
  assign new_n6896 = ~new_n6817 & ~new_n6895;
  assign new_n6897 = new_n6890 & ~new_n6896;
  assign new_n6898 = ~new_n6890 & new_n6896;
  assign new_n6899 = ~new_n6897 & ~new_n6898;
  assign new_n6900 = ~new_n6889 & new_n6899;
  assign new_n6901 = new_n6890 & new_n6895;
  assign new_n6902 = ~new_n6900 & ~new_n6901;
  assign new_n6903 = new_n6887 & new_n6902;
  assign new_n6904 = ~new_n6885 & ~new_n6903;
  assign new_n6905 = new_n6880 & new_n6904;
  assign new_n6906 = ~new_n3212 & ~new_n3214;
  assign new_n6907 = ~new_n3215 & ~new_n6906;
  assign new_n6908 = ~new_n6880 & ~new_n6904;
  assign new_n6909 = ~new_n6905 & ~new_n6908;
  assign new_n6910 = ~new_n6907 & new_n6909;
  assign new_n6911 = ~new_n6905 & ~new_n6910;
  assign new_n6912 = new_n6878 & ~new_n6911;
  assign new_n6913 = ~new_n6876 & ~new_n6912;
  assign new_n6914 = new_n6871 & ~new_n6913;
  assign new_n6915 = new_n3258 & ~new_n3260;
  assign new_n6916 = ~new_n3261 & ~new_n6915;
  assign new_n6917 = ~new_n6871 & new_n6913;
  assign new_n6918 = ~new_n6914 & ~new_n6917;
  assign new_n6919 = ~new_n6916 & new_n6918;
  assign new_n6920 = ~new_n6914 & ~new_n6919;
  assign new_n6921 = new_n6869 & ~new_n6920;
  assign new_n6922 = new_n3268 & ~new_n3270;
  assign new_n6923 = ~new_n3271 & ~new_n6922;
  assign new_n6924 = ~new_n6869 & new_n6920;
  assign new_n6925 = ~new_n6921 & ~new_n6924;
  assign new_n6926 = ~new_n6923 & new_n6925;
  assign new_n6927 = ~new_n6921 & ~new_n6926;
  assign new_n6928 = new_n6867 & new_n6927;
  assign new_n6929 = ~new_n6865 & ~new_n6928;
  assign new_n6930 = ~new_n6867 & ~new_n6927;
  assign new_n6931 = ~new_n6928 & ~new_n6930;
  assign new_n6932 = ~A629 & ~A630;
  assign new_n6933 = A629 & A630;
  assign new_n6934 = ~new_n6932 & ~new_n6933;
  assign new_n6935 = ~A628 & new_n6934;
  assign new_n6936 = ~new_n6932 & ~new_n6935;
  assign new_n6937 = ~A626 & ~A627;
  assign new_n6938 = A626 & A627;
  assign new_n6939 = ~new_n6937 & ~new_n6938;
  assign new_n6940 = ~A625 & new_n6939;
  assign new_n6941 = ~new_n6937 & ~new_n6940;
  assign new_n6942 = ~new_n6936 & ~new_n6941;
  assign new_n6943 = A628 & ~new_n6934;
  assign new_n6944 = ~new_n6935 & ~new_n6943;
  assign new_n6945 = A625 & ~new_n6939;
  assign new_n6946 = ~new_n6940 & ~new_n6945;
  assign new_n6947 = ~new_n6944 & ~new_n6946;
  assign new_n6948 = new_n6936 & new_n6941;
  assign new_n6949 = ~new_n6942 & ~new_n6948;
  assign new_n6950 = ~new_n6947 & new_n6949;
  assign new_n6951 = ~new_n6942 & ~new_n6950;
  assign new_n6952 = A619 & A620;
  assign new_n6953 = ~A623 & ~A624;
  assign new_n6954 = A621 & A622;
  assign new_n6955 = ~new_n6952 & new_n6954;
  assign new_n6956 = ~A621 & ~A622;
  assign new_n6957 = ~new_n6954 & ~new_n6956;
  assign new_n6958 = ~A619 & ~A620;
  assign new_n6959 = ~new_n6952 & ~new_n6958;
  assign new_n6960 = ~new_n6957 & new_n6959;
  assign new_n6961 = ~new_n6954 & ~new_n6958;
  assign new_n6962 = ~new_n6960 & new_n6961;
  assign new_n6963 = ~new_n6955 & ~new_n6962;
  assign new_n6964 = new_n6953 & new_n6963;
  assign new_n6965 = new_n6952 & new_n6964;
  assign new_n6966 = A623 & A624;
  assign new_n6967 = ~new_n6963 & new_n6966;
  assign new_n6968 = ~new_n6965 & ~new_n6967;
  assign new_n6969 = ~new_n6952 & ~new_n6960;
  assign new_n6970 = ~new_n6953 & ~new_n6956;
  assign new_n6971 = ~new_n6969 & new_n6970;
  assign new_n6972 = new_n6968 & ~new_n6971;
  assign new_n6973 = ~new_n6951 & new_n6972;
  assign new_n6974 = ~new_n6966 & new_n6971;
  assign new_n6975 = new_n6956 & new_n6958;
  assign new_n6976 = ~new_n6966 & new_n6975;
  assign new_n6977 = ~new_n6964 & ~new_n6976;
  assign new_n6978 = ~new_n6974 & new_n6977;
  assign new_n6979 = new_n6968 & new_n6978;
  assign new_n6980 = ~new_n6949 & new_n6979;
  assign new_n6981 = new_n6949 & ~new_n6979;
  assign new_n6982 = ~new_n6980 & ~new_n6981;
  assign new_n6983 = new_n6944 & new_n6946;
  assign new_n6984 = ~new_n6947 & ~new_n6983;
  assign new_n6985 = ~new_n6953 & ~new_n6966;
  assign new_n6986 = new_n6957 & ~new_n6959;
  assign new_n6987 = ~new_n6960 & ~new_n6986;
  assign new_n6988 = new_n6985 & ~new_n6987;
  assign new_n6989 = ~new_n6985 & new_n6987;
  assign new_n6990 = ~new_n6988 & ~new_n6989;
  assign new_n6991 = new_n6984 & ~new_n6990;
  assign new_n6992 = ~new_n6983 & ~new_n6991;
  assign new_n6993 = ~new_n6982 & ~new_n6992;
  assign new_n6994 = ~new_n6950 & ~new_n6980;
  assign new_n6995 = ~new_n6993 & ~new_n6994;
  assign new_n6996 = new_n6951 & ~new_n6972;
  assign new_n6997 = ~new_n6973 & ~new_n6996;
  assign new_n6998 = ~new_n6995 & new_n6997;
  assign new_n6999 = ~new_n6973 & ~new_n6998;
  assign new_n7000 = A613 & A614;
  assign new_n7001 = A616 & A617;
  assign new_n7002 = ~new_n7000 & ~new_n7001;
  assign new_n7003 = A615 & A618;
  assign new_n7004 = ~new_n7002 & new_n7003;
  assign new_n7005 = ~A613 & ~A614;
  assign new_n7006 = ~A615 & A618;
  assign new_n7007 = new_n7001 & new_n7006;
  assign new_n7008 = ~A615 & ~new_n7000;
  assign new_n7009 = ~A616 & ~A617;
  assign new_n7010 = ~new_n7001 & ~new_n7009;
  assign new_n7011 = A618 & ~new_n7010;
  assign new_n7012 = ~A618 & ~new_n7001;
  assign new_n7013 = ~new_n7008 & ~new_n7012;
  assign new_n7014 = ~new_n7011 & new_n7013;
  assign new_n7015 = ~new_n7007 & ~new_n7014;
  assign new_n7016 = ~new_n7005 & ~new_n7015;
  assign new_n7017 = A617 & new_n7000;
  assign new_n7018 = new_n7004 & ~new_n7017;
  assign new_n7019 = ~new_n7003 & new_n7005;
  assign new_n7020 = new_n7009 & new_n7019;
  assign new_n7021 = A615 & ~A618;
  assign new_n7022 = new_n7000 & ~new_n7009;
  assign new_n7023 = new_n7021 & new_n7022;
  assign new_n7024 = ~new_n7020 & ~new_n7023;
  assign new_n7025 = ~new_n7018 & new_n7024;
  assign new_n7026 = ~new_n7016 & new_n7025;
  assign new_n7027 = ~new_n7005 & ~new_n7026;
  assign new_n7028 = ~new_n7004 & ~new_n7027;
  assign new_n7029 = ~A608 & ~A609;
  assign new_n7030 = A608 & A609;
  assign new_n7031 = ~new_n7029 & ~new_n7030;
  assign new_n7032 = ~A607 & new_n7031;
  assign new_n7033 = ~new_n7029 & ~new_n7032;
  assign new_n7034 = ~A610 & ~A611;
  assign new_n7035 = new_n7033 & ~new_n7034;
  assign new_n7036 = A610 & A611;
  assign new_n7037 = ~A612 & ~new_n7036;
  assign new_n7038 = new_n7035 & ~new_n7037;
  assign new_n7039 = ~A612 & ~new_n7035;
  assign new_n7040 = A607 & ~new_n7031;
  assign new_n7041 = ~new_n7032 & ~new_n7040;
  assign new_n7042 = ~new_n7033 & ~new_n7036;
  assign new_n7043 = new_n7033 & new_n7036;
  assign new_n7044 = ~new_n7042 & ~new_n7043;
  assign new_n7045 = A612 & ~new_n7044;
  assign new_n7046 = ~new_n7039 & ~new_n7041;
  assign new_n7047 = ~new_n7045 & new_n7046;
  assign new_n7048 = ~new_n7038 & ~new_n7047;
  assign new_n7049 = new_n7028 & new_n7048;
  assign new_n7050 = ~new_n7000 & ~new_n7005;
  assign new_n7051 = ~new_n7006 & ~new_n7021;
  assign new_n7052 = new_n7050 & ~new_n7051;
  assign new_n7053 = ~new_n7050 & new_n7051;
  assign new_n7054 = ~new_n7052 & ~new_n7053;
  assign new_n7055 = new_n7010 & new_n7054;
  assign new_n7056 = new_n7008 & new_n7012;
  assign new_n7057 = ~new_n7055 & new_n7056;
  assign new_n7058 = new_n7026 & ~new_n7057;
  assign new_n7059 = A612 & ~new_n7041;
  assign new_n7060 = ~new_n7033 & new_n7034;
  assign new_n7061 = ~new_n7059 & new_n7060;
  assign new_n7062 = ~new_n7033 & new_n7037;
  assign new_n7063 = ~new_n7038 & ~new_n7062;
  assign new_n7064 = new_n7041 & ~new_n7063;
  assign new_n7065 = ~new_n7047 & ~new_n7061;
  assign new_n7066 = ~new_n7064 & new_n7065;
  assign new_n7067 = ~new_n7058 & ~new_n7066;
  assign new_n7068 = ~new_n7010 & ~new_n7054;
  assign new_n7069 = ~new_n7055 & ~new_n7068;
  assign new_n7070 = ~A612 & new_n7041;
  assign new_n7071 = ~new_n7059 & ~new_n7070;
  assign new_n7072 = ~new_n7034 & ~new_n7036;
  assign new_n7073 = ~new_n7071 & new_n7072;
  assign new_n7074 = new_n7071 & ~new_n7072;
  assign new_n7075 = ~new_n7073 & ~new_n7074;
  assign new_n7076 = new_n7069 & ~new_n7075;
  assign new_n7077 = new_n7058 & new_n7066;
  assign new_n7078 = ~new_n7067 & ~new_n7077;
  assign new_n7079 = ~new_n7076 & new_n7078;
  assign new_n7080 = ~new_n7067 & ~new_n7079;
  assign new_n7081 = ~new_n7028 & ~new_n7048;
  assign new_n7082 = ~new_n7049 & ~new_n7081;
  assign new_n7083 = ~new_n7080 & new_n7082;
  assign new_n7084 = ~new_n7049 & ~new_n7083;
  assign new_n7085 = ~new_n6999 & ~new_n7084;
  assign new_n7086 = new_n6999 & new_n7084;
  assign new_n7087 = ~new_n7085 & ~new_n7086;
  assign new_n7088 = new_n7080 & ~new_n7082;
  assign new_n7089 = ~new_n7083 & ~new_n7088;
  assign new_n7090 = ~new_n7069 & new_n7075;
  assign new_n7091 = ~new_n7076 & ~new_n7090;
  assign new_n7092 = ~new_n6984 & new_n6990;
  assign new_n7093 = ~new_n6991 & ~new_n7092;
  assign new_n7094 = new_n7091 & ~new_n7093;
  assign new_n7095 = new_n7078 & new_n7094;
  assign new_n7096 = new_n6982 & new_n6992;
  assign new_n7097 = ~new_n6993 & ~new_n7096;
  assign new_n7098 = ~new_n7076 & ~new_n7094;
  assign new_n7099 = new_n7078 & ~new_n7098;
  assign new_n7100 = ~new_n7078 & new_n7098;
  assign new_n7101 = ~new_n7099 & ~new_n7100;
  assign new_n7102 = ~new_n7097 & new_n7101;
  assign new_n7103 = ~new_n7095 & ~new_n7102;
  assign new_n7104 = ~new_n7089 & ~new_n7103;
  assign new_n7105 = new_n6995 & ~new_n6997;
  assign new_n7106 = ~new_n6998 & ~new_n7105;
  assign new_n7107 = new_n7089 & new_n7103;
  assign new_n7108 = ~new_n7104 & ~new_n7107;
  assign new_n7109 = ~new_n7106 & new_n7108;
  assign new_n7110 = ~new_n7104 & ~new_n7109;
  assign new_n7111 = new_n7087 & new_n7110;
  assign new_n7112 = ~new_n7085 & ~new_n7111;
  assign new_n7113 = ~A635 & ~A636;
  assign new_n7114 = A635 & A636;
  assign new_n7115 = ~new_n7113 & ~new_n7114;
  assign new_n7116 = A633 & A634;
  assign new_n7117 = A631 & A632;
  assign new_n7118 = new_n7116 & ~new_n7117;
  assign new_n7119 = ~A633 & ~A634;
  assign new_n7120 = ~new_n7116 & ~new_n7119;
  assign new_n7121 = ~A631 & ~A632;
  assign new_n7122 = ~new_n7117 & ~new_n7121;
  assign new_n7123 = ~new_n7120 & new_n7122;
  assign new_n7124 = ~new_n7116 & ~new_n7121;
  assign new_n7125 = ~new_n7123 & new_n7124;
  assign new_n7126 = ~new_n7118 & ~new_n7125;
  assign new_n7127 = new_n7113 & new_n7126;
  assign new_n7128 = ~new_n7115 & ~new_n7127;
  assign new_n7129 = new_n7120 & ~new_n7122;
  assign new_n7130 = ~new_n7116 & ~new_n7129;
  assign new_n7131 = ~new_n7121 & ~new_n7130;
  assign new_n7132 = ~new_n7128 & new_n7131;
  assign new_n7133 = new_n7114 & ~new_n7126;
  assign new_n7134 = ~new_n7132 & ~new_n7133;
  assign new_n7135 = ~new_n7113 & new_n7131;
  assign new_n7136 = new_n7134 & ~new_n7135;
  assign new_n7137 = ~A640 & ~A641;
  assign new_n7138 = A640 & A641;
  assign new_n7139 = ~new_n7137 & ~new_n7138;
  assign new_n7140 = ~A642 & new_n7139;
  assign new_n7141 = ~new_n7137 & ~new_n7140;
  assign new_n7142 = ~A638 & ~A639;
  assign new_n7143 = A638 & A639;
  assign new_n7144 = ~new_n7142 & ~new_n7143;
  assign new_n7145 = ~A637 & new_n7144;
  assign new_n7146 = ~new_n7142 & ~new_n7145;
  assign new_n7147 = ~new_n7141 & ~new_n7146;
  assign new_n7148 = A642 & ~new_n7139;
  assign new_n7149 = ~new_n7140 & ~new_n7148;
  assign new_n7150 = A637 & ~new_n7144;
  assign new_n7151 = ~new_n7145 & ~new_n7150;
  assign new_n7152 = ~new_n7149 & ~new_n7151;
  assign new_n7153 = new_n7141 & new_n7146;
  assign new_n7154 = ~new_n7152 & ~new_n7153;
  assign new_n7155 = ~new_n7147 & ~new_n7154;
  assign new_n7156 = ~new_n7136 & new_n7155;
  assign new_n7157 = new_n7149 & new_n7151;
  assign new_n7158 = ~new_n7152 & ~new_n7157;
  assign new_n7159 = ~new_n7123 & ~new_n7129;
  assign new_n7160 = new_n7115 & ~new_n7159;
  assign new_n7161 = ~new_n7115 & new_n7159;
  assign new_n7162 = ~new_n7160 & ~new_n7161;
  assign new_n7163 = new_n7158 & new_n7162;
  assign new_n7164 = ~new_n7152 & ~new_n7163;
  assign new_n7165 = ~new_n7147 & ~new_n7153;
  assign new_n7166 = ~new_n7164 & new_n7165;
  assign new_n7167 = new_n7164 & ~new_n7165;
  assign new_n7168 = ~new_n7166 & ~new_n7167;
  assign new_n7169 = ~new_n7114 & new_n7119;
  assign new_n7170 = new_n7121 & new_n7169;
  assign new_n7171 = ~new_n7127 & ~new_n7170;
  assign new_n7172 = new_n7134 & new_n7171;
  assign new_n7173 = new_n7168 & new_n7172;
  assign new_n7174 = new_n7163 & new_n7165;
  assign new_n7175 = ~new_n7173 & ~new_n7174;
  assign new_n7176 = new_n7136 & ~new_n7155;
  assign new_n7177 = ~new_n7156 & ~new_n7176;
  assign new_n7178 = ~new_n7175 & new_n7177;
  assign new_n7179 = ~new_n7156 & ~new_n7178;
  assign new_n7180 = ~A653 & ~A654;
  assign new_n7181 = A653 & A654;
  assign new_n7182 = ~new_n7180 & ~new_n7181;
  assign new_n7183 = ~A652 & new_n7182;
  assign new_n7184 = ~new_n7180 & ~new_n7183;
  assign new_n7185 = ~A650 & ~A651;
  assign new_n7186 = A650 & A651;
  assign new_n7187 = ~new_n7185 & ~new_n7186;
  assign new_n7188 = ~A649 & new_n7187;
  assign new_n7189 = ~new_n7185 & ~new_n7188;
  assign new_n7190 = ~new_n7184 & ~new_n7189;
  assign new_n7191 = A649 & ~new_n7187;
  assign new_n7192 = ~new_n7188 & ~new_n7191;
  assign new_n7193 = A652 & ~new_n7182;
  assign new_n7194 = ~new_n7183 & ~new_n7193;
  assign new_n7195 = ~new_n7192 & ~new_n7194;
  assign new_n7196 = new_n7184 & new_n7189;
  assign new_n7197 = ~new_n7190 & ~new_n7196;
  assign new_n7198 = ~new_n7195 & new_n7197;
  assign new_n7199 = ~new_n7190 & ~new_n7198;
  assign new_n7200 = A643 & A644;
  assign new_n7201 = ~A647 & ~A648;
  assign new_n7202 = A645 & A646;
  assign new_n7203 = ~new_n7200 & new_n7202;
  assign new_n7204 = ~A645 & ~A646;
  assign new_n7205 = ~new_n7202 & ~new_n7204;
  assign new_n7206 = ~A643 & ~A644;
  assign new_n7207 = ~new_n7200 & ~new_n7206;
  assign new_n7208 = ~new_n7205 & new_n7207;
  assign new_n7209 = ~new_n7202 & ~new_n7206;
  assign new_n7210 = ~new_n7208 & new_n7209;
  assign new_n7211 = ~new_n7203 & ~new_n7210;
  assign new_n7212 = new_n7201 & new_n7211;
  assign new_n7213 = new_n7200 & new_n7212;
  assign new_n7214 = A647 & A648;
  assign new_n7215 = ~new_n7211 & new_n7214;
  assign new_n7216 = ~new_n7213 & ~new_n7215;
  assign new_n7217 = ~new_n7200 & ~new_n7208;
  assign new_n7218 = ~new_n7201 & ~new_n7204;
  assign new_n7219 = ~new_n7217 & new_n7218;
  assign new_n7220 = new_n7216 & ~new_n7219;
  assign new_n7221 = ~new_n7199 & new_n7220;
  assign new_n7222 = ~new_n7214 & new_n7219;
  assign new_n7223 = new_n7204 & new_n7206;
  assign new_n7224 = ~new_n7214 & new_n7223;
  assign new_n7225 = ~new_n7212 & ~new_n7224;
  assign new_n7226 = ~new_n7222 & new_n7225;
  assign new_n7227 = new_n7216 & new_n7226;
  assign new_n7228 = ~new_n7197 & new_n7227;
  assign new_n7229 = ~new_n7198 & ~new_n7228;
  assign new_n7230 = new_n7197 & ~new_n7227;
  assign new_n7231 = ~new_n7228 & ~new_n7230;
  assign new_n7232 = new_n7192 & new_n7194;
  assign new_n7233 = ~new_n7195 & ~new_n7232;
  assign new_n7234 = ~new_n7201 & ~new_n7214;
  assign new_n7235 = new_n7205 & ~new_n7207;
  assign new_n7236 = ~new_n7208 & ~new_n7235;
  assign new_n7237 = new_n7234 & ~new_n7236;
  assign new_n7238 = ~new_n7234 & new_n7236;
  assign new_n7239 = ~new_n7237 & ~new_n7238;
  assign new_n7240 = new_n7233 & new_n7239;
  assign new_n7241 = ~new_n7195 & ~new_n7240;
  assign new_n7242 = ~new_n7231 & new_n7241;
  assign new_n7243 = ~new_n7229 & ~new_n7242;
  assign new_n7244 = new_n7199 & ~new_n7220;
  assign new_n7245 = ~new_n7221 & ~new_n7244;
  assign new_n7246 = ~new_n7243 & new_n7245;
  assign new_n7247 = ~new_n7221 & ~new_n7246;
  assign new_n7248 = new_n7179 & ~new_n7247;
  assign new_n7249 = ~new_n7179 & new_n7247;
  assign new_n7250 = ~new_n7248 & ~new_n7249;
  assign new_n7251 = new_n7175 & ~new_n7177;
  assign new_n7252 = ~new_n7178 & ~new_n7251;
  assign new_n7253 = ~new_n7168 & ~new_n7172;
  assign new_n7254 = ~new_n7173 & ~new_n7253;
  assign new_n7255 = ~new_n7233 & ~new_n7239;
  assign new_n7256 = ~new_n7240 & ~new_n7255;
  assign new_n7257 = ~new_n7158 & ~new_n7162;
  assign new_n7258 = ~new_n7163 & ~new_n7257;
  assign new_n7259 = new_n7256 & new_n7258;
  assign new_n7260 = ~new_n7254 & ~new_n7259;
  assign new_n7261 = new_n7231 & ~new_n7241;
  assign new_n7262 = ~new_n7242 & ~new_n7261;
  assign new_n7263 = new_n7254 & new_n7259;
  assign new_n7264 = ~new_n7260 & ~new_n7263;
  assign new_n7265 = new_n7262 & new_n7264;
  assign new_n7266 = ~new_n7260 & ~new_n7265;
  assign new_n7267 = new_n7252 & new_n7266;
  assign new_n7268 = new_n7243 & ~new_n7245;
  assign new_n7269 = ~new_n7246 & ~new_n7268;
  assign new_n7270 = ~new_n7252 & ~new_n7266;
  assign new_n7271 = ~new_n7267 & ~new_n7270;
  assign new_n7272 = ~new_n7269 & new_n7271;
  assign new_n7273 = ~new_n7267 & ~new_n7272;
  assign new_n7274 = new_n7250 & new_n7273;
  assign new_n7275 = ~new_n7248 & ~new_n7274;
  assign new_n7276 = ~new_n7112 & ~new_n7275;
  assign new_n7277 = new_n7112 & new_n7275;
  assign new_n7278 = ~new_n7276 & ~new_n7277;
  assign new_n7279 = ~new_n7087 & ~new_n7110;
  assign new_n7280 = ~new_n7111 & ~new_n7279;
  assign new_n7281 = new_n7269 & ~new_n7271;
  assign new_n7282 = ~new_n7272 & ~new_n7281;
  assign new_n7283 = ~new_n7262 & ~new_n7264;
  assign new_n7284 = ~new_n7265 & ~new_n7283;
  assign new_n7285 = new_n7097 & ~new_n7101;
  assign new_n7286 = ~new_n7102 & ~new_n7285;
  assign new_n7287 = new_n7284 & ~new_n7286;
  assign new_n7288 = ~new_n7091 & new_n7093;
  assign new_n7289 = ~new_n7094 & ~new_n7288;
  assign new_n7290 = ~new_n7256 & ~new_n7258;
  assign new_n7291 = ~new_n7259 & ~new_n7290;
  assign new_n7292 = new_n7289 & new_n7291;
  assign new_n7293 = ~new_n7284 & new_n7286;
  assign new_n7294 = ~new_n7287 & ~new_n7293;
  assign new_n7295 = ~new_n7292 & new_n7294;
  assign new_n7296 = ~new_n7287 & ~new_n7295;
  assign new_n7297 = ~new_n7282 & ~new_n7296;
  assign new_n7298 = new_n7106 & ~new_n7108;
  assign new_n7299 = ~new_n7109 & ~new_n7298;
  assign new_n7300 = new_n7282 & new_n7296;
  assign new_n7301 = ~new_n7297 & ~new_n7300;
  assign new_n7302 = ~new_n7299 & new_n7301;
  assign new_n7303 = ~new_n7297 & ~new_n7302;
  assign new_n7304 = ~new_n7280 & new_n7303;
  assign new_n7305 = ~new_n7250 & ~new_n7273;
  assign new_n7306 = ~new_n7274 & ~new_n7305;
  assign new_n7307 = new_n7280 & ~new_n7303;
  assign new_n7308 = ~new_n7304 & ~new_n7307;
  assign new_n7309 = ~new_n7306 & new_n7308;
  assign new_n7310 = ~new_n7304 & ~new_n7309;
  assign new_n7311 = new_n7278 & new_n7310;
  assign new_n7312 = ~new_n7276 & ~new_n7311;
  assign new_n7313 = ~A575 & ~A576;
  assign new_n7314 = A575 & A576;
  assign new_n7315 = ~new_n7313 & ~new_n7314;
  assign new_n7316 = A573 & A574;
  assign new_n7317 = A571 & A572;
  assign new_n7318 = new_n7316 & ~new_n7317;
  assign new_n7319 = ~A573 & ~A574;
  assign new_n7320 = ~new_n7316 & ~new_n7319;
  assign new_n7321 = ~A571 & ~A572;
  assign new_n7322 = ~new_n7317 & ~new_n7321;
  assign new_n7323 = ~new_n7320 & new_n7322;
  assign new_n7324 = ~new_n7316 & ~new_n7321;
  assign new_n7325 = ~new_n7323 & new_n7324;
  assign new_n7326 = ~new_n7318 & ~new_n7325;
  assign new_n7327 = new_n7313 & new_n7326;
  assign new_n7328 = ~new_n7315 & ~new_n7327;
  assign new_n7329 = new_n7320 & ~new_n7322;
  assign new_n7330 = ~new_n7316 & ~new_n7329;
  assign new_n7331 = ~new_n7321 & ~new_n7330;
  assign new_n7332 = ~new_n7328 & new_n7331;
  assign new_n7333 = new_n7314 & ~new_n7326;
  assign new_n7334 = ~new_n7332 & ~new_n7333;
  assign new_n7335 = ~new_n7313 & new_n7331;
  assign new_n7336 = new_n7334 & ~new_n7335;
  assign new_n7337 = ~A581 & ~A582;
  assign new_n7338 = A581 & A582;
  assign new_n7339 = ~new_n7337 & ~new_n7338;
  assign new_n7340 = ~A580 & new_n7339;
  assign new_n7341 = ~new_n7337 & ~new_n7340;
  assign new_n7342 = ~A578 & ~A579;
  assign new_n7343 = A578 & A579;
  assign new_n7344 = ~new_n7342 & ~new_n7343;
  assign new_n7345 = ~A577 & new_n7344;
  assign new_n7346 = ~new_n7342 & ~new_n7345;
  assign new_n7347 = ~new_n7341 & ~new_n7346;
  assign new_n7348 = new_n7341 & new_n7346;
  assign new_n7349 = A580 & ~new_n7339;
  assign new_n7350 = ~new_n7340 & ~new_n7349;
  assign new_n7351 = A577 & ~new_n7344;
  assign new_n7352 = ~new_n7345 & ~new_n7351;
  assign new_n7353 = ~new_n7350 & ~new_n7352;
  assign new_n7354 = ~new_n7348 & ~new_n7353;
  assign new_n7355 = ~new_n7347 & ~new_n7354;
  assign new_n7356 = new_n7336 & ~new_n7355;
  assign new_n7357 = new_n7350 & new_n7352;
  assign new_n7358 = ~new_n7353 & ~new_n7357;
  assign new_n7359 = ~new_n7323 & ~new_n7329;
  assign new_n7360 = new_n7315 & ~new_n7359;
  assign new_n7361 = ~new_n7315 & new_n7359;
  assign new_n7362 = ~new_n7360 & ~new_n7361;
  assign new_n7363 = new_n7358 & new_n7362;
  assign new_n7364 = ~new_n7353 & ~new_n7363;
  assign new_n7365 = ~new_n7347 & ~new_n7348;
  assign new_n7366 = ~new_n7364 & new_n7365;
  assign new_n7367 = new_n7364 & ~new_n7365;
  assign new_n7368 = ~new_n7366 & ~new_n7367;
  assign new_n7369 = ~new_n7314 & new_n7319;
  assign new_n7370 = new_n7321 & new_n7369;
  assign new_n7371 = ~new_n7327 & ~new_n7370;
  assign new_n7372 = new_n7334 & new_n7371;
  assign new_n7373 = new_n7368 & new_n7372;
  assign new_n7374 = new_n7363 & new_n7365;
  assign new_n7375 = ~new_n7373 & ~new_n7374;
  assign new_n7376 = ~new_n7336 & new_n7355;
  assign new_n7377 = ~new_n7356 & ~new_n7376;
  assign new_n7378 = new_n7375 & new_n7377;
  assign new_n7379 = ~new_n7356 & ~new_n7378;
  assign new_n7380 = A559 & A560;
  assign new_n7381 = A562 & A563;
  assign new_n7382 = ~new_n7380 & ~new_n7381;
  assign new_n7383 = A561 & A564;
  assign new_n7384 = ~new_n7382 & new_n7383;
  assign new_n7385 = ~A559 & ~A560;
  assign new_n7386 = ~A561 & A564;
  assign new_n7387 = new_n7381 & new_n7386;
  assign new_n7388 = ~A561 & ~new_n7380;
  assign new_n7389 = ~A562 & ~A563;
  assign new_n7390 = ~new_n7381 & ~new_n7389;
  assign new_n7391 = A564 & ~new_n7390;
  assign new_n7392 = ~A564 & ~new_n7381;
  assign new_n7393 = ~new_n7388 & ~new_n7392;
  assign new_n7394 = ~new_n7391 & new_n7393;
  assign new_n7395 = ~new_n7387 & ~new_n7394;
  assign new_n7396 = ~new_n7385 & ~new_n7395;
  assign new_n7397 = A563 & new_n7380;
  assign new_n7398 = new_n7384 & ~new_n7397;
  assign new_n7399 = ~new_n7383 & new_n7385;
  assign new_n7400 = new_n7389 & new_n7399;
  assign new_n7401 = A561 & ~A564;
  assign new_n7402 = new_n7380 & ~new_n7389;
  assign new_n7403 = new_n7401 & new_n7402;
  assign new_n7404 = ~new_n7400 & ~new_n7403;
  assign new_n7405 = ~new_n7398 & new_n7404;
  assign new_n7406 = ~new_n7396 & new_n7405;
  assign new_n7407 = ~new_n7385 & ~new_n7406;
  assign new_n7408 = ~new_n7384 & ~new_n7407;
  assign new_n7409 = A565 & A566;
  assign new_n7410 = A568 & A569;
  assign new_n7411 = ~new_n7409 & ~new_n7410;
  assign new_n7412 = A567 & A570;
  assign new_n7413 = ~new_n7411 & new_n7412;
  assign new_n7414 = ~A565 & ~A566;
  assign new_n7415 = ~A567 & A570;
  assign new_n7416 = new_n7410 & new_n7415;
  assign new_n7417 = ~A567 & ~new_n7409;
  assign new_n7418 = ~A568 & ~A569;
  assign new_n7419 = ~new_n7410 & ~new_n7418;
  assign new_n7420 = A570 & ~new_n7419;
  assign new_n7421 = ~A570 & ~new_n7410;
  assign new_n7422 = ~new_n7417 & ~new_n7421;
  assign new_n7423 = ~new_n7420 & new_n7422;
  assign new_n7424 = ~new_n7416 & ~new_n7423;
  assign new_n7425 = ~new_n7414 & ~new_n7424;
  assign new_n7426 = A569 & new_n7409;
  assign new_n7427 = new_n7413 & ~new_n7426;
  assign new_n7428 = ~new_n7412 & new_n7414;
  assign new_n7429 = new_n7418 & new_n7428;
  assign new_n7430 = A567 & ~A570;
  assign new_n7431 = new_n7409 & ~new_n7418;
  assign new_n7432 = new_n7430 & new_n7431;
  assign new_n7433 = ~new_n7429 & ~new_n7432;
  assign new_n7434 = ~new_n7427 & new_n7433;
  assign new_n7435 = ~new_n7425 & new_n7434;
  assign new_n7436 = ~new_n7414 & ~new_n7435;
  assign new_n7437 = ~new_n7413 & ~new_n7436;
  assign new_n7438 = new_n7408 & new_n7437;
  assign new_n7439 = ~new_n7380 & ~new_n7385;
  assign new_n7440 = ~new_n7386 & ~new_n7401;
  assign new_n7441 = new_n7439 & ~new_n7440;
  assign new_n7442 = ~new_n7439 & new_n7440;
  assign new_n7443 = ~new_n7441 & ~new_n7442;
  assign new_n7444 = new_n7390 & new_n7443;
  assign new_n7445 = new_n7388 & new_n7392;
  assign new_n7446 = ~new_n7444 & new_n7445;
  assign new_n7447 = new_n7406 & ~new_n7446;
  assign new_n7448 = ~new_n7409 & ~new_n7414;
  assign new_n7449 = ~new_n7415 & ~new_n7430;
  assign new_n7450 = new_n7448 & ~new_n7449;
  assign new_n7451 = ~new_n7448 & new_n7449;
  assign new_n7452 = ~new_n7450 & ~new_n7451;
  assign new_n7453 = new_n7419 & new_n7452;
  assign new_n7454 = new_n7417 & new_n7421;
  assign new_n7455 = ~new_n7453 & new_n7454;
  assign new_n7456 = new_n7435 & ~new_n7455;
  assign new_n7457 = ~new_n7447 & ~new_n7456;
  assign new_n7458 = ~new_n7390 & ~new_n7443;
  assign new_n7459 = ~new_n7444 & ~new_n7458;
  assign new_n7460 = ~new_n7419 & ~new_n7452;
  assign new_n7461 = ~new_n7453 & ~new_n7460;
  assign new_n7462 = new_n7459 & new_n7461;
  assign new_n7463 = new_n7447 & new_n7456;
  assign new_n7464 = ~new_n7457 & ~new_n7463;
  assign new_n7465 = ~new_n7462 & new_n7464;
  assign new_n7466 = ~new_n7457 & ~new_n7465;
  assign new_n7467 = ~new_n7408 & ~new_n7437;
  assign new_n7468 = ~new_n7438 & ~new_n7467;
  assign new_n7469 = ~new_n7466 & new_n7468;
  assign new_n7470 = ~new_n7438 & ~new_n7469;
  assign new_n7471 = ~new_n7379 & ~new_n7470;
  assign new_n7472 = new_n7379 & new_n7470;
  assign new_n7473 = ~new_n7471 & ~new_n7472;
  assign new_n7474 = new_n7466 & ~new_n7468;
  assign new_n7475 = ~new_n7469 & ~new_n7474;
  assign new_n7476 = new_n7462 & ~new_n7464;
  assign new_n7477 = ~new_n7465 & ~new_n7476;
  assign new_n7478 = ~new_n7368 & ~new_n7372;
  assign new_n7479 = ~new_n7373 & ~new_n7478;
  assign new_n7480 = new_n7477 & ~new_n7479;
  assign new_n7481 = ~new_n7477 & new_n7479;
  assign new_n7482 = ~new_n7459 & ~new_n7461;
  assign new_n7483 = ~new_n7462 & ~new_n7482;
  assign new_n7484 = ~new_n7358 & ~new_n7362;
  assign new_n7485 = ~new_n7363 & ~new_n7484;
  assign new_n7486 = new_n7483 & new_n7485;
  assign new_n7487 = ~new_n7481 & ~new_n7486;
  assign new_n7488 = ~new_n7480 & ~new_n7487;
  assign new_n7489 = ~new_n7475 & new_n7488;
  assign new_n7490 = ~new_n7375 & ~new_n7377;
  assign new_n7491 = ~new_n7378 & ~new_n7490;
  assign new_n7492 = new_n7475 & ~new_n7488;
  assign new_n7493 = ~new_n7489 & ~new_n7492;
  assign new_n7494 = ~new_n7491 & new_n7493;
  assign new_n7495 = ~new_n7489 & ~new_n7494;
  assign new_n7496 = new_n7473 & new_n7495;
  assign new_n7497 = ~new_n7471 & ~new_n7496;
  assign new_n7498 = ~A599 & ~A600;
  assign new_n7499 = A599 & A600;
  assign new_n7500 = ~new_n7498 & ~new_n7499;
  assign new_n7501 = A597 & A598;
  assign new_n7502 = A595 & A596;
  assign new_n7503 = new_n7501 & ~new_n7502;
  assign new_n7504 = ~A597 & ~A598;
  assign new_n7505 = ~new_n7501 & ~new_n7504;
  assign new_n7506 = ~A595 & ~A596;
  assign new_n7507 = ~new_n7502 & ~new_n7506;
  assign new_n7508 = ~new_n7505 & new_n7507;
  assign new_n7509 = ~new_n7501 & ~new_n7506;
  assign new_n7510 = ~new_n7508 & new_n7509;
  assign new_n7511 = ~new_n7503 & ~new_n7510;
  assign new_n7512 = new_n7498 & new_n7511;
  assign new_n7513 = ~new_n7500 & ~new_n7512;
  assign new_n7514 = new_n7505 & ~new_n7507;
  assign new_n7515 = ~new_n7501 & ~new_n7514;
  assign new_n7516 = ~new_n7506 & ~new_n7515;
  assign new_n7517 = ~new_n7513 & new_n7516;
  assign new_n7518 = new_n7499 & ~new_n7511;
  assign new_n7519 = ~new_n7517 & ~new_n7518;
  assign new_n7520 = ~new_n7498 & new_n7516;
  assign new_n7521 = new_n7519 & ~new_n7520;
  assign new_n7522 = ~A605 & ~A606;
  assign new_n7523 = A605 & A606;
  assign new_n7524 = ~new_n7522 & ~new_n7523;
  assign new_n7525 = ~A604 & new_n7524;
  assign new_n7526 = ~new_n7522 & ~new_n7525;
  assign new_n7527 = ~A602 & ~A603;
  assign new_n7528 = A602 & A603;
  assign new_n7529 = ~new_n7527 & ~new_n7528;
  assign new_n7530 = ~A601 & new_n7529;
  assign new_n7531 = ~new_n7527 & ~new_n7530;
  assign new_n7532 = ~new_n7526 & ~new_n7531;
  assign new_n7533 = A604 & ~new_n7524;
  assign new_n7534 = ~new_n7525 & ~new_n7533;
  assign new_n7535 = A601 & ~new_n7529;
  assign new_n7536 = ~new_n7530 & ~new_n7535;
  assign new_n7537 = ~new_n7534 & ~new_n7536;
  assign new_n7538 = new_n7526 & new_n7531;
  assign new_n7539 = ~new_n7537 & ~new_n7538;
  assign new_n7540 = ~new_n7532 & ~new_n7539;
  assign new_n7541 = ~new_n7521 & new_n7540;
  assign new_n7542 = new_n7534 & new_n7536;
  assign new_n7543 = ~new_n7537 & ~new_n7542;
  assign new_n7544 = ~new_n7508 & ~new_n7514;
  assign new_n7545 = new_n7500 & ~new_n7544;
  assign new_n7546 = ~new_n7500 & new_n7544;
  assign new_n7547 = ~new_n7545 & ~new_n7546;
  assign new_n7548 = new_n7543 & new_n7547;
  assign new_n7549 = ~new_n7537 & ~new_n7548;
  assign new_n7550 = ~new_n7532 & ~new_n7538;
  assign new_n7551 = ~new_n7549 & new_n7550;
  assign new_n7552 = new_n7549 & ~new_n7550;
  assign new_n7553 = ~new_n7551 & ~new_n7552;
  assign new_n7554 = ~new_n7499 & new_n7504;
  assign new_n7555 = new_n7506 & new_n7554;
  assign new_n7556 = ~new_n7512 & ~new_n7555;
  assign new_n7557 = new_n7519 & new_n7556;
  assign new_n7558 = new_n7553 & new_n7557;
  assign new_n7559 = new_n7548 & new_n7550;
  assign new_n7560 = ~new_n7558 & ~new_n7559;
  assign new_n7561 = new_n7521 & ~new_n7540;
  assign new_n7562 = ~new_n7541 & ~new_n7561;
  assign new_n7563 = ~new_n7560 & new_n7562;
  assign new_n7564 = ~new_n7541 & ~new_n7563;
  assign new_n7565 = A583 & A584;
  assign new_n7566 = A586 & A587;
  assign new_n7567 = ~new_n7565 & ~new_n7566;
  assign new_n7568 = A585 & A588;
  assign new_n7569 = ~new_n7567 & new_n7568;
  assign new_n7570 = ~A583 & ~A584;
  assign new_n7571 = ~A585 & A588;
  assign new_n7572 = new_n7566 & new_n7571;
  assign new_n7573 = ~A585 & ~new_n7565;
  assign new_n7574 = ~A586 & ~A587;
  assign new_n7575 = ~new_n7566 & ~new_n7574;
  assign new_n7576 = A588 & ~new_n7575;
  assign new_n7577 = ~A588 & ~new_n7566;
  assign new_n7578 = ~new_n7573 & ~new_n7577;
  assign new_n7579 = ~new_n7576 & new_n7578;
  assign new_n7580 = ~new_n7572 & ~new_n7579;
  assign new_n7581 = ~new_n7570 & ~new_n7580;
  assign new_n7582 = A587 & new_n7565;
  assign new_n7583 = new_n7569 & ~new_n7582;
  assign new_n7584 = ~new_n7568 & new_n7570;
  assign new_n7585 = new_n7574 & new_n7584;
  assign new_n7586 = A585 & ~A588;
  assign new_n7587 = new_n7565 & ~new_n7574;
  assign new_n7588 = new_n7586 & new_n7587;
  assign new_n7589 = ~new_n7585 & ~new_n7588;
  assign new_n7590 = ~new_n7583 & new_n7589;
  assign new_n7591 = ~new_n7581 & new_n7590;
  assign new_n7592 = ~new_n7570 & ~new_n7591;
  assign new_n7593 = ~new_n7569 & ~new_n7592;
  assign new_n7594 = A589 & A590;
  assign new_n7595 = A592 & A593;
  assign new_n7596 = ~new_n7594 & ~new_n7595;
  assign new_n7597 = A591 & A594;
  assign new_n7598 = ~new_n7596 & new_n7597;
  assign new_n7599 = ~A589 & ~A590;
  assign new_n7600 = ~A591 & A594;
  assign new_n7601 = new_n7595 & new_n7600;
  assign new_n7602 = ~A591 & ~new_n7594;
  assign new_n7603 = ~A592 & ~A593;
  assign new_n7604 = ~new_n7595 & ~new_n7603;
  assign new_n7605 = A594 & ~new_n7604;
  assign new_n7606 = ~A594 & ~new_n7595;
  assign new_n7607 = ~new_n7602 & ~new_n7606;
  assign new_n7608 = ~new_n7605 & new_n7607;
  assign new_n7609 = ~new_n7601 & ~new_n7608;
  assign new_n7610 = ~new_n7599 & ~new_n7609;
  assign new_n7611 = A593 & new_n7594;
  assign new_n7612 = new_n7598 & ~new_n7611;
  assign new_n7613 = ~new_n7597 & new_n7599;
  assign new_n7614 = new_n7603 & new_n7613;
  assign new_n7615 = A591 & ~A594;
  assign new_n7616 = new_n7594 & ~new_n7603;
  assign new_n7617 = new_n7615 & new_n7616;
  assign new_n7618 = ~new_n7614 & ~new_n7617;
  assign new_n7619 = ~new_n7612 & new_n7618;
  assign new_n7620 = ~new_n7610 & new_n7619;
  assign new_n7621 = ~new_n7599 & ~new_n7620;
  assign new_n7622 = ~new_n7598 & ~new_n7621;
  assign new_n7623 = new_n7593 & new_n7622;
  assign new_n7624 = ~new_n7565 & ~new_n7570;
  assign new_n7625 = ~new_n7571 & ~new_n7586;
  assign new_n7626 = new_n7624 & ~new_n7625;
  assign new_n7627 = ~new_n7624 & new_n7625;
  assign new_n7628 = ~new_n7626 & ~new_n7627;
  assign new_n7629 = new_n7575 & new_n7628;
  assign new_n7630 = new_n7573 & new_n7577;
  assign new_n7631 = ~new_n7629 & new_n7630;
  assign new_n7632 = new_n7591 & ~new_n7631;
  assign new_n7633 = ~new_n7594 & ~new_n7599;
  assign new_n7634 = ~new_n7600 & ~new_n7615;
  assign new_n7635 = new_n7633 & ~new_n7634;
  assign new_n7636 = ~new_n7633 & new_n7634;
  assign new_n7637 = ~new_n7635 & ~new_n7636;
  assign new_n7638 = new_n7604 & new_n7637;
  assign new_n7639 = new_n7602 & new_n7606;
  assign new_n7640 = ~new_n7638 & new_n7639;
  assign new_n7641 = new_n7620 & ~new_n7640;
  assign new_n7642 = ~new_n7632 & ~new_n7641;
  assign new_n7643 = ~new_n7575 & ~new_n7628;
  assign new_n7644 = ~new_n7629 & ~new_n7643;
  assign new_n7645 = ~new_n7604 & ~new_n7637;
  assign new_n7646 = ~new_n7638 & ~new_n7645;
  assign new_n7647 = new_n7644 & new_n7646;
  assign new_n7648 = new_n7632 & new_n7641;
  assign new_n7649 = ~new_n7642 & ~new_n7648;
  assign new_n7650 = ~new_n7647 & new_n7649;
  assign new_n7651 = ~new_n7642 & ~new_n7650;
  assign new_n7652 = ~new_n7593 & ~new_n7622;
  assign new_n7653 = ~new_n7623 & ~new_n7652;
  assign new_n7654 = ~new_n7651 & new_n7653;
  assign new_n7655 = ~new_n7623 & ~new_n7654;
  assign new_n7656 = new_n7564 & ~new_n7655;
  assign new_n7657 = ~new_n7564 & new_n7655;
  assign new_n7658 = ~new_n7656 & ~new_n7657;
  assign new_n7659 = new_n7651 & ~new_n7653;
  assign new_n7660 = ~new_n7654 & ~new_n7659;
  assign new_n7661 = ~new_n7644 & ~new_n7646;
  assign new_n7662 = ~new_n7647 & ~new_n7661;
  assign new_n7663 = ~new_n7543 & ~new_n7547;
  assign new_n7664 = ~new_n7548 & ~new_n7663;
  assign new_n7665 = new_n7662 & new_n7664;
  assign new_n7666 = new_n7647 & ~new_n7649;
  assign new_n7667 = ~new_n7650 & ~new_n7665;
  assign new_n7668 = ~new_n7666 & new_n7667;
  assign new_n7669 = ~new_n7553 & ~new_n7557;
  assign new_n7670 = ~new_n7558 & ~new_n7669;
  assign new_n7671 = new_n7649 & new_n7665;
  assign new_n7672 = ~new_n7668 & ~new_n7671;
  assign new_n7673 = ~new_n7670 & new_n7672;
  assign new_n7674 = ~new_n7668 & ~new_n7673;
  assign new_n7675 = new_n7660 & ~new_n7674;
  assign new_n7676 = new_n7560 & ~new_n7562;
  assign new_n7677 = ~new_n7563 & ~new_n7676;
  assign new_n7678 = ~new_n7660 & new_n7674;
  assign new_n7679 = ~new_n7675 & ~new_n7678;
  assign new_n7680 = ~new_n7677 & new_n7679;
  assign new_n7681 = ~new_n7675 & ~new_n7680;
  assign new_n7682 = new_n7658 & ~new_n7681;
  assign new_n7683 = ~new_n7656 & ~new_n7682;
  assign new_n7684 = ~new_n7497 & ~new_n7683;
  assign new_n7685 = ~new_n7658 & new_n7681;
  assign new_n7686 = ~new_n7682 & ~new_n7685;
  assign new_n7687 = ~new_n7473 & ~new_n7495;
  assign new_n7688 = ~new_n7496 & ~new_n7687;
  assign new_n7689 = ~new_n7686 & ~new_n7688;
  assign new_n7690 = new_n7686 & new_n7688;
  assign new_n7691 = ~new_n7689 & ~new_n7690;
  assign new_n7692 = new_n7677 & ~new_n7679;
  assign new_n7693 = ~new_n7680 & ~new_n7692;
  assign new_n7694 = new_n7491 & ~new_n7493;
  assign new_n7695 = ~new_n7494 & ~new_n7694;
  assign new_n7696 = ~new_n7693 & new_n7695;
  assign new_n7697 = new_n7693 & ~new_n7695;
  assign new_n7698 = ~new_n7696 & ~new_n7697;
  assign new_n7699 = new_n7670 & ~new_n7672;
  assign new_n7700 = ~new_n7673 & ~new_n7699;
  assign new_n7701 = ~new_n7480 & ~new_n7481;
  assign new_n7702 = ~new_n7662 & ~new_n7664;
  assign new_n7703 = ~new_n7665 & ~new_n7702;
  assign new_n7704 = ~new_n7483 & ~new_n7485;
  assign new_n7705 = ~new_n7486 & ~new_n7704;
  assign new_n7706 = new_n7703 & new_n7705;
  assign new_n7707 = ~new_n7486 & ~new_n7706;
  assign new_n7708 = new_n7701 & ~new_n7707;
  assign new_n7709 = ~new_n7701 & new_n7707;
  assign new_n7710 = ~new_n7708 & ~new_n7709;
  assign new_n7711 = ~new_n7700 & new_n7710;
  assign new_n7712 = new_n7701 & new_n7706;
  assign new_n7713 = ~new_n7711 & ~new_n7712;
  assign new_n7714 = new_n7698 & ~new_n7713;
  assign new_n7715 = ~new_n7696 & ~new_n7714;
  assign new_n7716 = new_n7691 & ~new_n7715;
  assign new_n7717 = ~new_n7689 & ~new_n7716;
  assign new_n7718 = new_n7497 & new_n7683;
  assign new_n7719 = ~new_n7684 & ~new_n7718;
  assign new_n7720 = new_n7717 & new_n7719;
  assign new_n7721 = ~new_n7684 & ~new_n7720;
  assign new_n7722 = new_n7312 & new_n7721;
  assign new_n7723 = ~new_n7312 & ~new_n7721;
  assign new_n7724 = ~new_n7722 & ~new_n7723;
  assign new_n7725 = ~new_n7717 & ~new_n7719;
  assign new_n7726 = ~new_n7720 & ~new_n7725;
  assign new_n7727 = ~new_n7691 & new_n7715;
  assign new_n7728 = ~new_n7716 & ~new_n7727;
  assign new_n7729 = new_n7299 & ~new_n7301;
  assign new_n7730 = ~new_n7302 & ~new_n7729;
  assign new_n7731 = new_n7700 & ~new_n7710;
  assign new_n7732 = ~new_n7711 & ~new_n7731;
  assign new_n7733 = ~new_n7289 & ~new_n7291;
  assign new_n7734 = ~new_n7292 & ~new_n7733;
  assign new_n7735 = ~new_n7703 & ~new_n7705;
  assign new_n7736 = ~new_n7706 & ~new_n7735;
  assign new_n7737 = new_n7734 & new_n7736;
  assign new_n7738 = ~new_n7732 & ~new_n7737;
  assign new_n7739 = new_n7292 & ~new_n7294;
  assign new_n7740 = ~new_n7295 & ~new_n7739;
  assign new_n7741 = new_n7732 & new_n7737;
  assign new_n7742 = ~new_n7738 & ~new_n7741;
  assign new_n7743 = new_n7740 & new_n7742;
  assign new_n7744 = ~new_n7738 & ~new_n7743;
  assign new_n7745 = new_n7730 & ~new_n7744;
  assign new_n7746 = ~new_n7698 & new_n7713;
  assign new_n7747 = ~new_n7714 & ~new_n7746;
  assign new_n7748 = ~new_n7730 & new_n7744;
  assign new_n7749 = ~new_n7745 & ~new_n7748;
  assign new_n7750 = ~new_n7747 & new_n7749;
  assign new_n7751 = ~new_n7745 & ~new_n7750;
  assign new_n7752 = new_n7728 & new_n7751;
  assign new_n7753 = new_n7306 & ~new_n7308;
  assign new_n7754 = ~new_n7309 & ~new_n7753;
  assign new_n7755 = ~new_n7728 & ~new_n7751;
  assign new_n7756 = ~new_n7752 & ~new_n7755;
  assign new_n7757 = new_n7754 & new_n7756;
  assign new_n7758 = ~new_n7752 & ~new_n7757;
  assign new_n7759 = ~new_n7726 & ~new_n7758;
  assign new_n7760 = ~new_n7278 & ~new_n7310;
  assign new_n7761 = ~new_n7311 & ~new_n7760;
  assign new_n7762 = new_n7726 & new_n7758;
  assign new_n7763 = ~new_n7759 & ~new_n7762;
  assign new_n7764 = ~new_n7761 & new_n7763;
  assign new_n7765 = ~new_n7759 & ~new_n7764;
  assign new_n7766 = new_n7724 & ~new_n7765;
  assign new_n7767 = ~new_n7722 & ~new_n7766;
  assign new_n7768 = A469 & A470;
  assign new_n7769 = A472 & A473;
  assign new_n7770 = ~new_n7768 & ~new_n7769;
  assign new_n7771 = A471 & A474;
  assign new_n7772 = ~new_n7770 & new_n7771;
  assign new_n7773 = ~A469 & ~A470;
  assign new_n7774 = ~A471 & A474;
  assign new_n7775 = new_n7769 & new_n7774;
  assign new_n7776 = ~A471 & ~new_n7768;
  assign new_n7777 = ~A472 & ~A473;
  assign new_n7778 = ~new_n7769 & ~new_n7777;
  assign new_n7779 = A474 & ~new_n7778;
  assign new_n7780 = ~A474 & ~new_n7769;
  assign new_n7781 = ~new_n7776 & ~new_n7780;
  assign new_n7782 = ~new_n7779 & new_n7781;
  assign new_n7783 = ~new_n7775 & ~new_n7782;
  assign new_n7784 = ~new_n7773 & ~new_n7783;
  assign new_n7785 = A473 & new_n7768;
  assign new_n7786 = new_n7772 & ~new_n7785;
  assign new_n7787 = ~new_n7771 & new_n7773;
  assign new_n7788 = new_n7777 & new_n7787;
  assign new_n7789 = A471 & ~A474;
  assign new_n7790 = new_n7768 & ~new_n7777;
  assign new_n7791 = new_n7789 & new_n7790;
  assign new_n7792 = ~new_n7788 & ~new_n7791;
  assign new_n7793 = ~new_n7786 & new_n7792;
  assign new_n7794 = ~new_n7784 & new_n7793;
  assign new_n7795 = ~new_n7773 & ~new_n7794;
  assign new_n7796 = ~new_n7772 & ~new_n7795;
  assign new_n7797 = A463 & A464;
  assign new_n7798 = A467 & A468;
  assign new_n7799 = ~new_n7797 & new_n7798;
  assign new_n7800 = ~A468 & new_n7797;
  assign new_n7801 = A465 & A466;
  assign new_n7802 = ~new_n7799 & new_n7801;
  assign new_n7803 = ~new_n7800 & new_n7802;
  assign new_n7804 = ~A465 & ~A466;
  assign new_n7805 = ~new_n7797 & new_n7804;
  assign new_n7806 = ~A463 & ~A464;
  assign new_n7807 = new_n7798 & ~new_n7806;
  assign new_n7808 = ~new_n7805 & new_n7807;
  assign new_n7809 = ~new_n7801 & ~new_n7808;
  assign new_n7810 = ~new_n7803 & ~new_n7809;
  assign new_n7811 = ~new_n7797 & ~new_n7801;
  assign new_n7812 = ~A467 & ~A468;
  assign new_n7813 = ~new_n7804 & ~new_n7806;
  assign new_n7814 = ~new_n7812 & new_n7813;
  assign new_n7815 = ~new_n7811 & new_n7814;
  assign new_n7816 = ~new_n7810 & ~new_n7815;
  assign new_n7817 = new_n7796 & new_n7816;
  assign new_n7818 = ~new_n7768 & ~new_n7773;
  assign new_n7819 = ~new_n7774 & ~new_n7789;
  assign new_n7820 = new_n7818 & ~new_n7819;
  assign new_n7821 = ~new_n7818 & new_n7819;
  assign new_n7822 = ~new_n7820 & ~new_n7821;
  assign new_n7823 = new_n7778 & new_n7822;
  assign new_n7824 = ~new_n7778 & ~new_n7822;
  assign new_n7825 = ~new_n7823 & ~new_n7824;
  assign new_n7826 = ~new_n7798 & ~new_n7812;
  assign new_n7827 = ~new_n7801 & ~new_n7804;
  assign new_n7828 = new_n7826 & ~new_n7827;
  assign new_n7829 = ~new_n7826 & new_n7827;
  assign new_n7830 = ~new_n7828 & ~new_n7829;
  assign new_n7831 = ~new_n7797 & ~new_n7806;
  assign new_n7832 = ~new_n7830 & new_n7831;
  assign new_n7833 = new_n7830 & ~new_n7831;
  assign new_n7834 = ~new_n7832 & ~new_n7833;
  assign new_n7835 = new_n7825 & new_n7834;
  assign new_n7836 = ~new_n7801 & new_n7806;
  assign new_n7837 = new_n7812 & new_n7836;
  assign new_n7838 = new_n7805 & ~new_n7832;
  assign new_n7839 = ~new_n7815 & ~new_n7838;
  assign new_n7840 = ~new_n7798 & ~new_n7839;
  assign new_n7841 = ~new_n7810 & ~new_n7837;
  assign new_n7842 = ~new_n7840 & new_n7841;
  assign new_n7843 = ~new_n7835 & ~new_n7842;
  assign new_n7844 = new_n7835 & new_n7842;
  assign new_n7845 = ~new_n7843 & ~new_n7844;
  assign new_n7846 = new_n7776 & new_n7780;
  assign new_n7847 = ~new_n7823 & new_n7846;
  assign new_n7848 = new_n7794 & ~new_n7847;
  assign new_n7849 = new_n7845 & ~new_n7848;
  assign new_n7850 = ~new_n7843 & ~new_n7849;
  assign new_n7851 = ~new_n7796 & ~new_n7816;
  assign new_n7852 = ~new_n7817 & ~new_n7851;
  assign new_n7853 = ~new_n7850 & new_n7852;
  assign new_n7854 = ~new_n7817 & ~new_n7853;
  assign new_n7855 = A475 & A476;
  assign new_n7856 = A478 & A479;
  assign new_n7857 = ~new_n7855 & ~new_n7856;
  assign new_n7858 = A477 & A480;
  assign new_n7859 = ~new_n7857 & new_n7858;
  assign new_n7860 = ~A475 & ~A476;
  assign new_n7861 = ~A477 & A480;
  assign new_n7862 = new_n7856 & new_n7861;
  assign new_n7863 = ~A477 & ~new_n7855;
  assign new_n7864 = ~A478 & ~A479;
  assign new_n7865 = ~new_n7856 & ~new_n7864;
  assign new_n7866 = A480 & ~new_n7865;
  assign new_n7867 = ~A480 & ~new_n7856;
  assign new_n7868 = ~new_n7863 & ~new_n7867;
  assign new_n7869 = ~new_n7866 & new_n7868;
  assign new_n7870 = ~new_n7862 & ~new_n7869;
  assign new_n7871 = ~new_n7860 & ~new_n7870;
  assign new_n7872 = A479 & new_n7855;
  assign new_n7873 = new_n7859 & ~new_n7872;
  assign new_n7874 = ~new_n7858 & new_n7860;
  assign new_n7875 = new_n7864 & new_n7874;
  assign new_n7876 = A477 & ~A480;
  assign new_n7877 = new_n7855 & ~new_n7864;
  assign new_n7878 = new_n7876 & new_n7877;
  assign new_n7879 = ~new_n7875 & ~new_n7878;
  assign new_n7880 = ~new_n7873 & new_n7879;
  assign new_n7881 = ~new_n7871 & new_n7880;
  assign new_n7882 = ~new_n7860 & ~new_n7881;
  assign new_n7883 = ~new_n7859 & ~new_n7882;
  assign new_n7884 = A481 & A482;
  assign new_n7885 = A484 & A485;
  assign new_n7886 = ~new_n7884 & ~new_n7885;
  assign new_n7887 = A483 & A486;
  assign new_n7888 = ~new_n7886 & new_n7887;
  assign new_n7889 = ~A481 & ~A482;
  assign new_n7890 = ~A483 & A486;
  assign new_n7891 = new_n7885 & new_n7890;
  assign new_n7892 = ~A483 & ~new_n7884;
  assign new_n7893 = ~A484 & ~A485;
  assign new_n7894 = ~new_n7885 & ~new_n7893;
  assign new_n7895 = A486 & ~new_n7894;
  assign new_n7896 = ~A486 & ~new_n7885;
  assign new_n7897 = ~new_n7892 & ~new_n7896;
  assign new_n7898 = ~new_n7895 & new_n7897;
  assign new_n7899 = ~new_n7891 & ~new_n7898;
  assign new_n7900 = ~new_n7889 & ~new_n7899;
  assign new_n7901 = A485 & new_n7884;
  assign new_n7902 = new_n7888 & ~new_n7901;
  assign new_n7903 = ~new_n7887 & new_n7889;
  assign new_n7904 = new_n7893 & new_n7903;
  assign new_n7905 = A483 & ~A486;
  assign new_n7906 = new_n7884 & ~new_n7893;
  assign new_n7907 = new_n7905 & new_n7906;
  assign new_n7908 = ~new_n7904 & ~new_n7907;
  assign new_n7909 = ~new_n7902 & new_n7908;
  assign new_n7910 = ~new_n7900 & new_n7909;
  assign new_n7911 = ~new_n7889 & ~new_n7910;
  assign new_n7912 = ~new_n7888 & ~new_n7911;
  assign new_n7913 = new_n7883 & new_n7912;
  assign new_n7914 = ~new_n7855 & ~new_n7860;
  assign new_n7915 = ~new_n7861 & ~new_n7876;
  assign new_n7916 = new_n7914 & ~new_n7915;
  assign new_n7917 = ~new_n7914 & new_n7915;
  assign new_n7918 = ~new_n7916 & ~new_n7917;
  assign new_n7919 = new_n7865 & new_n7918;
  assign new_n7920 = ~new_n7865 & ~new_n7918;
  assign new_n7921 = ~new_n7919 & ~new_n7920;
  assign new_n7922 = ~new_n7884 & ~new_n7889;
  assign new_n7923 = ~new_n7890 & ~new_n7905;
  assign new_n7924 = new_n7922 & ~new_n7923;
  assign new_n7925 = ~new_n7922 & new_n7923;
  assign new_n7926 = ~new_n7924 & ~new_n7925;
  assign new_n7927 = new_n7894 & new_n7926;
  assign new_n7928 = ~new_n7894 & ~new_n7926;
  assign new_n7929 = ~new_n7927 & ~new_n7928;
  assign new_n7930 = new_n7921 & new_n7929;
  assign new_n7931 = new_n7892 & new_n7896;
  assign new_n7932 = ~new_n7927 & new_n7931;
  assign new_n7933 = new_n7910 & ~new_n7932;
  assign new_n7934 = ~new_n7930 & ~new_n7933;
  assign new_n7935 = new_n7930 & new_n7933;
  assign new_n7936 = ~new_n7934 & ~new_n7935;
  assign new_n7937 = new_n7863 & new_n7867;
  assign new_n7938 = ~new_n7919 & new_n7937;
  assign new_n7939 = new_n7881 & ~new_n7938;
  assign new_n7940 = new_n7936 & ~new_n7939;
  assign new_n7941 = ~new_n7934 & ~new_n7940;
  assign new_n7942 = ~new_n7883 & ~new_n7912;
  assign new_n7943 = ~new_n7913 & ~new_n7942;
  assign new_n7944 = ~new_n7941 & new_n7943;
  assign new_n7945 = ~new_n7913 & ~new_n7944;
  assign new_n7946 = new_n7854 & new_n7945;
  assign new_n7947 = new_n7850 & ~new_n7852;
  assign new_n7948 = ~new_n7853 & ~new_n7947;
  assign new_n7949 = ~new_n7936 & new_n7939;
  assign new_n7950 = ~new_n7940 & ~new_n7949;
  assign new_n7951 = ~new_n7845 & new_n7848;
  assign new_n7952 = ~new_n7849 & ~new_n7951;
  assign new_n7953 = ~new_n7950 & ~new_n7952;
  assign new_n7954 = new_n7950 & new_n7952;
  assign new_n7955 = ~new_n7921 & ~new_n7929;
  assign new_n7956 = ~new_n7930 & ~new_n7955;
  assign new_n7957 = ~new_n7825 & ~new_n7834;
  assign new_n7958 = ~new_n7835 & ~new_n7957;
  assign new_n7959 = new_n7956 & new_n7958;
  assign new_n7960 = ~new_n7954 & new_n7959;
  assign new_n7961 = ~new_n7953 & ~new_n7960;
  assign new_n7962 = ~new_n7948 & ~new_n7961;
  assign new_n7963 = new_n7941 & ~new_n7943;
  assign new_n7964 = ~new_n7944 & ~new_n7963;
  assign new_n7965 = new_n7948 & new_n7961;
  assign new_n7966 = ~new_n7962 & ~new_n7965;
  assign new_n7967 = ~new_n7964 & new_n7966;
  assign new_n7968 = ~new_n7962 & ~new_n7967;
  assign new_n7969 = ~new_n7854 & ~new_n7945;
  assign new_n7970 = ~new_n7946 & ~new_n7969;
  assign new_n7971 = ~new_n7968 & new_n7970;
  assign new_n7972 = ~new_n7946 & ~new_n7971;
  assign new_n7973 = A487 & A488;
  assign new_n7974 = A490 & A491;
  assign new_n7975 = ~new_n7973 & ~new_n7974;
  assign new_n7976 = A489 & A492;
  assign new_n7977 = ~new_n7975 & new_n7976;
  assign new_n7978 = ~A487 & ~A488;
  assign new_n7979 = ~A489 & A492;
  assign new_n7980 = new_n7974 & new_n7979;
  assign new_n7981 = ~A489 & ~new_n7973;
  assign new_n7982 = ~A490 & ~A491;
  assign new_n7983 = ~new_n7974 & ~new_n7982;
  assign new_n7984 = A492 & ~new_n7983;
  assign new_n7985 = ~A492 & ~new_n7974;
  assign new_n7986 = ~new_n7981 & ~new_n7985;
  assign new_n7987 = ~new_n7984 & new_n7986;
  assign new_n7988 = ~new_n7980 & ~new_n7987;
  assign new_n7989 = ~new_n7978 & ~new_n7988;
  assign new_n7990 = A491 & new_n7973;
  assign new_n7991 = new_n7977 & ~new_n7990;
  assign new_n7992 = ~new_n7976 & new_n7978;
  assign new_n7993 = new_n7982 & new_n7992;
  assign new_n7994 = A489 & ~A492;
  assign new_n7995 = new_n7973 & ~new_n7982;
  assign new_n7996 = new_n7994 & new_n7995;
  assign new_n7997 = ~new_n7993 & ~new_n7996;
  assign new_n7998 = ~new_n7991 & new_n7997;
  assign new_n7999 = ~new_n7989 & new_n7998;
  assign new_n8000 = ~new_n7978 & ~new_n7999;
  assign new_n8001 = ~new_n7977 & ~new_n8000;
  assign new_n8002 = ~A493 & ~A495;
  assign new_n8003 = A493 & A495;
  assign new_n8004 = ~new_n8002 & ~new_n8003;
  assign new_n8005 = ~A494 & new_n8004;
  assign new_n8006 = ~new_n8002 & ~new_n8005;
  assign new_n8007 = ~A496 & ~A497;
  assign new_n8008 = new_n8006 & ~new_n8007;
  assign new_n8009 = A496 & A497;
  assign new_n8010 = ~A498 & ~new_n8009;
  assign new_n8011 = new_n8008 & ~new_n8010;
  assign new_n8012 = ~A498 & ~new_n8008;
  assign new_n8013 = A494 & ~new_n8004;
  assign new_n8014 = ~new_n8005 & ~new_n8013;
  assign new_n8015 = ~new_n8006 & ~new_n8009;
  assign new_n8016 = new_n8006 & new_n8009;
  assign new_n8017 = ~new_n8015 & ~new_n8016;
  assign new_n8018 = A498 & ~new_n8017;
  assign new_n8019 = ~new_n8012 & ~new_n8014;
  assign new_n8020 = ~new_n8018 & new_n8019;
  assign new_n8021 = ~new_n8011 & ~new_n8020;
  assign new_n8022 = new_n8001 & new_n8021;
  assign new_n8023 = ~new_n7973 & ~new_n7978;
  assign new_n8024 = ~new_n7979 & ~new_n7994;
  assign new_n8025 = new_n8023 & ~new_n8024;
  assign new_n8026 = ~new_n8023 & new_n8024;
  assign new_n8027 = ~new_n8025 & ~new_n8026;
  assign new_n8028 = new_n7983 & new_n8027;
  assign new_n8029 = new_n7981 & new_n7985;
  assign new_n8030 = ~new_n8028 & new_n8029;
  assign new_n8031 = new_n7999 & ~new_n8030;
  assign new_n8032 = A498 & ~new_n8014;
  assign new_n8033 = ~new_n8006 & new_n8007;
  assign new_n8034 = ~new_n8032 & new_n8033;
  assign new_n8035 = ~new_n8006 & new_n8010;
  assign new_n8036 = ~new_n8011 & ~new_n8035;
  assign new_n8037 = new_n8014 & ~new_n8036;
  assign new_n8038 = ~new_n8020 & ~new_n8034;
  assign new_n8039 = ~new_n8037 & new_n8038;
  assign new_n8040 = ~new_n8031 & ~new_n8039;
  assign new_n8041 = ~new_n7983 & ~new_n8027;
  assign new_n8042 = ~new_n8028 & ~new_n8041;
  assign new_n8043 = ~A498 & new_n8014;
  assign new_n8044 = ~new_n8032 & ~new_n8043;
  assign new_n8045 = ~new_n8007 & ~new_n8009;
  assign new_n8046 = ~new_n8044 & new_n8045;
  assign new_n8047 = new_n8044 & ~new_n8045;
  assign new_n8048 = ~new_n8046 & ~new_n8047;
  assign new_n8049 = new_n8042 & ~new_n8048;
  assign new_n8050 = new_n8031 & new_n8039;
  assign new_n8051 = ~new_n8040 & ~new_n8050;
  assign new_n8052 = ~new_n8049 & new_n8051;
  assign new_n8053 = ~new_n8040 & ~new_n8052;
  assign new_n8054 = ~new_n8001 & ~new_n8021;
  assign new_n8055 = ~new_n8022 & ~new_n8054;
  assign new_n8056 = ~new_n8053 & new_n8055;
  assign new_n8057 = ~new_n8022 & ~new_n8056;
  assign new_n8058 = ~A505 & ~A506;
  assign new_n8059 = A505 & A506;
  assign new_n8060 = ~A507 & ~new_n8059;
  assign new_n8061 = ~new_n8058 & ~new_n8060;
  assign new_n8062 = A509 & A510;
  assign new_n8063 = new_n8061 & new_n8062;
  assign new_n8064 = A507 & new_n8059;
  assign new_n8065 = ~A508 & ~new_n8064;
  assign new_n8066 = new_n8061 & ~new_n8065;
  assign new_n8067 = A509 & new_n8066;
  assign new_n8068 = A507 & A508;
  assign new_n8069 = new_n8059 & new_n8068;
  assign new_n8070 = ~new_n8067 & ~new_n8069;
  assign new_n8071 = ~A510 & ~new_n8070;
  assign new_n8072 = ~A509 & ~A510;
  assign new_n8073 = ~new_n8058 & ~new_n8072;
  assign new_n8074 = new_n8060 & ~new_n8062;
  assign new_n8075 = ~new_n8073 & new_n8074;
  assign new_n8076 = ~new_n8063 & ~new_n8075;
  assign new_n8077 = ~A508 & ~new_n8076;
  assign new_n8078 = ~A509 & A510;
  assign new_n8079 = new_n8066 & new_n8078;
  assign new_n8080 = new_n8058 & ~new_n8068;
  assign new_n8081 = A508 & new_n8062;
  assign new_n8082 = ~new_n8064 & new_n8081;
  assign new_n8083 = ~new_n8080 & new_n8082;
  assign new_n8084 = ~new_n8079 & ~new_n8083;
  assign new_n8085 = ~new_n8077 & new_n8084;
  assign new_n8086 = ~new_n8071 & new_n8085;
  assign new_n8087 = ~new_n8065 & ~new_n8086;
  assign new_n8088 = ~new_n8063 & ~new_n8087;
  assign new_n8089 = ~A500 & ~A501;
  assign new_n8090 = A500 & A501;
  assign new_n8091 = ~new_n8089 & ~new_n8090;
  assign new_n8092 = ~A499 & new_n8091;
  assign new_n8093 = ~new_n8089 & ~new_n8092;
  assign new_n8094 = ~A502 & ~A503;
  assign new_n8095 = new_n8093 & ~new_n8094;
  assign new_n8096 = A502 & A503;
  assign new_n8097 = ~A504 & ~new_n8096;
  assign new_n8098 = new_n8095 & ~new_n8097;
  assign new_n8099 = ~A504 & ~new_n8095;
  assign new_n8100 = A499 & ~new_n8091;
  assign new_n8101 = ~new_n8092 & ~new_n8100;
  assign new_n8102 = ~new_n8093 & ~new_n8096;
  assign new_n8103 = new_n8093 & new_n8096;
  assign new_n8104 = ~new_n8102 & ~new_n8103;
  assign new_n8105 = A504 & ~new_n8104;
  assign new_n8106 = ~new_n8099 & ~new_n8101;
  assign new_n8107 = ~new_n8105 & new_n8106;
  assign new_n8108 = ~new_n8098 & ~new_n8107;
  assign new_n8109 = new_n8088 & new_n8108;
  assign new_n8110 = A507 & ~A510;
  assign new_n8111 = ~A507 & A510;
  assign new_n8112 = ~new_n8110 & ~new_n8111;
  assign new_n8113 = ~new_n8058 & ~new_n8059;
  assign new_n8114 = ~A508 & ~A509;
  assign new_n8115 = A508 & A509;
  assign new_n8116 = ~new_n8114 & ~new_n8115;
  assign new_n8117 = new_n8113 & ~new_n8116;
  assign new_n8118 = ~new_n8113 & new_n8116;
  assign new_n8119 = ~new_n8117 & ~new_n8118;
  assign new_n8120 = new_n8112 & new_n8119;
  assign new_n8121 = ~new_n8112 & ~new_n8119;
  assign new_n8122 = ~new_n8120 & ~new_n8121;
  assign new_n8123 = A504 & ~new_n8101;
  assign new_n8124 = ~A504 & new_n8101;
  assign new_n8125 = ~new_n8123 & ~new_n8124;
  assign new_n8126 = ~new_n8094 & ~new_n8096;
  assign new_n8127 = ~new_n8125 & new_n8126;
  assign new_n8128 = new_n8125 & ~new_n8126;
  assign new_n8129 = ~new_n8127 & ~new_n8128;
  assign new_n8130 = new_n8122 & ~new_n8129;
  assign new_n8131 = ~new_n8093 & new_n8094;
  assign new_n8132 = ~new_n8123 & new_n8131;
  assign new_n8133 = ~new_n8093 & new_n8097;
  assign new_n8134 = ~new_n8098 & ~new_n8133;
  assign new_n8135 = new_n8101 & ~new_n8134;
  assign new_n8136 = ~new_n8107 & ~new_n8132;
  assign new_n8137 = ~new_n8135 & new_n8136;
  assign new_n8138 = ~new_n8130 & ~new_n8137;
  assign new_n8139 = new_n8072 & new_n8080;
  assign new_n8140 = new_n8086 & ~new_n8139;
  assign new_n8141 = new_n8130 & new_n8137;
  assign new_n8142 = ~new_n8138 & ~new_n8141;
  assign new_n8143 = ~new_n8140 & new_n8142;
  assign new_n8144 = ~new_n8138 & ~new_n8143;
  assign new_n8145 = ~new_n8088 & ~new_n8108;
  assign new_n8146 = ~new_n8109 & ~new_n8145;
  assign new_n8147 = ~new_n8144 & new_n8146;
  assign new_n8148 = ~new_n8109 & ~new_n8147;
  assign new_n8149 = new_n8057 & new_n8148;
  assign new_n8150 = new_n8053 & ~new_n8055;
  assign new_n8151 = ~new_n8056 & ~new_n8150;
  assign new_n8152 = ~new_n8042 & new_n8048;
  assign new_n8153 = ~new_n8049 & ~new_n8152;
  assign new_n8154 = ~new_n8122 & new_n8129;
  assign new_n8155 = ~new_n8130 & ~new_n8154;
  assign new_n8156 = new_n8153 & new_n8155;
  assign new_n8157 = new_n8051 & new_n8156;
  assign new_n8158 = new_n8140 & ~new_n8142;
  assign new_n8159 = ~new_n8143 & ~new_n8158;
  assign new_n8160 = ~new_n8049 & ~new_n8156;
  assign new_n8161 = new_n8051 & ~new_n8160;
  assign new_n8162 = ~new_n8051 & new_n8160;
  assign new_n8163 = ~new_n8161 & ~new_n8162;
  assign new_n8164 = ~new_n8159 & new_n8163;
  assign new_n8165 = ~new_n8157 & ~new_n8164;
  assign new_n8166 = ~new_n8151 & ~new_n8165;
  assign new_n8167 = new_n8144 & ~new_n8146;
  assign new_n8168 = ~new_n8147 & ~new_n8167;
  assign new_n8169 = new_n8151 & new_n8165;
  assign new_n8170 = ~new_n8166 & ~new_n8169;
  assign new_n8171 = ~new_n8168 & new_n8170;
  assign new_n8172 = ~new_n8166 & ~new_n8171;
  assign new_n8173 = ~new_n8057 & ~new_n8148;
  assign new_n8174 = ~new_n8149 & ~new_n8173;
  assign new_n8175 = ~new_n8172 & new_n8174;
  assign new_n8176 = ~new_n8149 & ~new_n8175;
  assign new_n8177 = ~new_n7972 & ~new_n8176;
  assign new_n8178 = new_n7972 & new_n8176;
  assign new_n8179 = ~new_n8177 & ~new_n8178;
  assign new_n8180 = new_n7968 & ~new_n7970;
  assign new_n8181 = ~new_n7971 & ~new_n8180;
  assign new_n8182 = new_n8159 & ~new_n8163;
  assign new_n8183 = ~new_n8164 & ~new_n8182;
  assign new_n8184 = ~new_n7953 & ~new_n7954;
  assign new_n8185 = ~new_n8153 & ~new_n8155;
  assign new_n8186 = ~new_n8156 & ~new_n8185;
  assign new_n8187 = ~new_n7956 & ~new_n7958;
  assign new_n8188 = ~new_n7959 & ~new_n8187;
  assign new_n8189 = new_n8186 & new_n8188;
  assign new_n8190 = ~new_n7959 & ~new_n8189;
  assign new_n8191 = new_n8184 & ~new_n8190;
  assign new_n8192 = ~new_n8184 & new_n8190;
  assign new_n8193 = ~new_n8191 & ~new_n8192;
  assign new_n8194 = new_n8183 & new_n8193;
  assign new_n8195 = new_n8184 & new_n8189;
  assign new_n8196 = ~new_n8194 & ~new_n8195;
  assign new_n8197 = new_n7964 & ~new_n7966;
  assign new_n8198 = ~new_n7967 & ~new_n8197;
  assign new_n8199 = new_n8196 & ~new_n8198;
  assign new_n8200 = new_n8168 & ~new_n8170;
  assign new_n8201 = ~new_n8171 & ~new_n8200;
  assign new_n8202 = ~new_n8196 & new_n8198;
  assign new_n8203 = ~new_n8199 & ~new_n8202;
  assign new_n8204 = ~new_n8201 & new_n8203;
  assign new_n8205 = ~new_n8199 & ~new_n8204;
  assign new_n8206 = ~new_n8181 & ~new_n8205;
  assign new_n8207 = new_n8172 & ~new_n8174;
  assign new_n8208 = ~new_n8175 & ~new_n8207;
  assign new_n8209 = new_n8181 & new_n8205;
  assign new_n8210 = ~new_n8206 & ~new_n8209;
  assign new_n8211 = ~new_n8208 & new_n8210;
  assign new_n8212 = ~new_n8206 & ~new_n8211;
  assign new_n8213 = new_n8179 & new_n8212;
  assign new_n8214 = ~new_n8177 & ~new_n8213;
  assign new_n8215 = ~A551 & ~A552;
  assign new_n8216 = A551 & A552;
  assign new_n8217 = ~new_n8215 & ~new_n8216;
  assign new_n8218 = A549 & A550;
  assign new_n8219 = A547 & A548;
  assign new_n8220 = new_n8218 & ~new_n8219;
  assign new_n8221 = ~A549 & ~A550;
  assign new_n8222 = ~new_n8218 & ~new_n8221;
  assign new_n8223 = ~A547 & ~A548;
  assign new_n8224 = ~new_n8219 & ~new_n8223;
  assign new_n8225 = ~new_n8222 & new_n8224;
  assign new_n8226 = ~new_n8218 & ~new_n8223;
  assign new_n8227 = ~new_n8225 & new_n8226;
  assign new_n8228 = ~new_n8220 & ~new_n8227;
  assign new_n8229 = new_n8215 & new_n8228;
  assign new_n8230 = ~new_n8217 & ~new_n8229;
  assign new_n8231 = new_n8222 & ~new_n8224;
  assign new_n8232 = ~new_n8218 & ~new_n8231;
  assign new_n8233 = ~new_n8223 & ~new_n8232;
  assign new_n8234 = ~new_n8230 & new_n8233;
  assign new_n8235 = new_n8216 & ~new_n8228;
  assign new_n8236 = ~new_n8234 & ~new_n8235;
  assign new_n8237 = ~new_n8215 & new_n8233;
  assign new_n8238 = new_n8236 & ~new_n8237;
  assign new_n8239 = ~A554 & ~A555;
  assign new_n8240 = A554 & A555;
  assign new_n8241 = ~new_n8239 & ~new_n8240;
  assign new_n8242 = ~A553 & new_n8241;
  assign new_n8243 = ~new_n8239 & ~new_n8242;
  assign new_n8244 = ~A557 & ~A558;
  assign new_n8245 = A557 & A558;
  assign new_n8246 = ~new_n8244 & ~new_n8245;
  assign new_n8247 = ~A556 & new_n8246;
  assign new_n8248 = ~new_n8244 & ~new_n8247;
  assign new_n8249 = ~new_n8243 & ~new_n8248;
  assign new_n8250 = A556 & ~new_n8246;
  assign new_n8251 = ~new_n8247 & ~new_n8250;
  assign new_n8252 = A553 & ~new_n8241;
  assign new_n8253 = ~new_n8242 & ~new_n8252;
  assign new_n8254 = ~new_n8251 & ~new_n8253;
  assign new_n8255 = new_n8243 & new_n8248;
  assign new_n8256 = ~new_n8254 & ~new_n8255;
  assign new_n8257 = ~new_n8249 & ~new_n8256;
  assign new_n8258 = ~new_n8238 & new_n8257;
  assign new_n8259 = new_n8251 & new_n8253;
  assign new_n8260 = ~new_n8254 & ~new_n8259;
  assign new_n8261 = ~new_n8225 & ~new_n8231;
  assign new_n8262 = new_n8217 & ~new_n8261;
  assign new_n8263 = ~new_n8217 & new_n8261;
  assign new_n8264 = ~new_n8262 & ~new_n8263;
  assign new_n8265 = new_n8260 & new_n8264;
  assign new_n8266 = ~new_n8254 & ~new_n8265;
  assign new_n8267 = ~new_n8249 & ~new_n8255;
  assign new_n8268 = ~new_n8266 & new_n8267;
  assign new_n8269 = new_n8266 & ~new_n8267;
  assign new_n8270 = ~new_n8268 & ~new_n8269;
  assign new_n8271 = ~new_n8216 & new_n8221;
  assign new_n8272 = new_n8223 & new_n8271;
  assign new_n8273 = ~new_n8229 & ~new_n8272;
  assign new_n8274 = new_n8236 & new_n8273;
  assign new_n8275 = new_n8270 & new_n8274;
  assign new_n8276 = new_n8265 & new_n8267;
  assign new_n8277 = ~new_n8275 & ~new_n8276;
  assign new_n8278 = new_n8238 & ~new_n8257;
  assign new_n8279 = ~new_n8258 & ~new_n8278;
  assign new_n8280 = ~new_n8277 & new_n8279;
  assign new_n8281 = ~new_n8258 & ~new_n8280;
  assign new_n8282 = A541 & A542;
  assign new_n8283 = A544 & A545;
  assign new_n8284 = ~new_n8282 & ~new_n8283;
  assign new_n8285 = A543 & A546;
  assign new_n8286 = ~new_n8284 & new_n8285;
  assign new_n8287 = ~A541 & ~A542;
  assign new_n8288 = ~A543 & A546;
  assign new_n8289 = new_n8283 & new_n8288;
  assign new_n8290 = ~A543 & ~new_n8282;
  assign new_n8291 = ~A544 & ~A545;
  assign new_n8292 = ~new_n8283 & ~new_n8291;
  assign new_n8293 = A546 & ~new_n8292;
  assign new_n8294 = ~A546 & ~new_n8283;
  assign new_n8295 = ~new_n8290 & ~new_n8294;
  assign new_n8296 = ~new_n8293 & new_n8295;
  assign new_n8297 = ~new_n8289 & ~new_n8296;
  assign new_n8298 = ~new_n8287 & ~new_n8297;
  assign new_n8299 = A545 & new_n8282;
  assign new_n8300 = new_n8286 & ~new_n8299;
  assign new_n8301 = ~new_n8285 & new_n8287;
  assign new_n8302 = new_n8291 & new_n8301;
  assign new_n8303 = A543 & ~A546;
  assign new_n8304 = new_n8282 & ~new_n8291;
  assign new_n8305 = new_n8303 & new_n8304;
  assign new_n8306 = ~new_n8302 & ~new_n8305;
  assign new_n8307 = ~new_n8300 & new_n8306;
  assign new_n8308 = ~new_n8298 & new_n8307;
  assign new_n8309 = ~new_n8287 & ~new_n8308;
  assign new_n8310 = ~new_n8286 & ~new_n8309;
  assign new_n8311 = ~A539 & ~A540;
  assign new_n8312 = A539 & A540;
  assign new_n8313 = ~new_n8311 & ~new_n8312;
  assign new_n8314 = ~A538 & new_n8313;
  assign new_n8315 = ~new_n8311 & ~new_n8314;
  assign new_n8316 = ~A536 & ~A537;
  assign new_n8317 = A536 & A537;
  assign new_n8318 = ~new_n8316 & ~new_n8317;
  assign new_n8319 = ~A535 & new_n8318;
  assign new_n8320 = ~new_n8316 & ~new_n8319;
  assign new_n8321 = new_n8315 & new_n8320;
  assign new_n8322 = A535 & ~new_n8318;
  assign new_n8323 = ~new_n8319 & ~new_n8322;
  assign new_n8324 = A538 & ~new_n8313;
  assign new_n8325 = ~new_n8314 & ~new_n8324;
  assign new_n8326 = ~new_n8323 & ~new_n8325;
  assign new_n8327 = ~new_n8315 & ~new_n8320;
  assign new_n8328 = ~new_n8321 & ~new_n8327;
  assign new_n8329 = new_n8326 & new_n8328;
  assign new_n8330 = ~new_n8321 & ~new_n8329;
  assign new_n8331 = ~new_n8310 & ~new_n8330;
  assign new_n8332 = new_n8310 & new_n8330;
  assign new_n8333 = ~new_n8331 & ~new_n8332;
  assign new_n8334 = new_n8323 & new_n8325;
  assign new_n8335 = ~new_n8282 & ~new_n8287;
  assign new_n8336 = ~new_n8288 & ~new_n8303;
  assign new_n8337 = new_n8335 & ~new_n8336;
  assign new_n8338 = ~new_n8335 & new_n8336;
  assign new_n8339 = ~new_n8337 & ~new_n8338;
  assign new_n8340 = new_n8292 & new_n8339;
  assign new_n8341 = ~new_n8292 & ~new_n8339;
  assign new_n8342 = ~new_n8340 & ~new_n8341;
  assign new_n8343 = ~new_n8326 & ~new_n8334;
  assign new_n8344 = ~new_n8342 & new_n8343;
  assign new_n8345 = ~new_n8334 & ~new_n8344;
  assign new_n8346 = new_n8290 & new_n8294;
  assign new_n8347 = ~new_n8340 & new_n8346;
  assign new_n8348 = new_n8308 & ~new_n8347;
  assign new_n8349 = ~new_n8345 & ~new_n8348;
  assign new_n8350 = new_n8345 & new_n8348;
  assign new_n8351 = ~new_n8349 & ~new_n8350;
  assign new_n8352 = ~new_n8328 & new_n8351;
  assign new_n8353 = ~new_n8329 & ~new_n8349;
  assign new_n8354 = ~new_n8352 & new_n8353;
  assign new_n8355 = new_n8333 & new_n8354;
  assign new_n8356 = ~new_n8331 & ~new_n8355;
  assign new_n8357 = new_n8281 & new_n8356;
  assign new_n8358 = new_n8277 & ~new_n8279;
  assign new_n8359 = ~new_n8280 & ~new_n8358;
  assign new_n8360 = ~new_n8270 & ~new_n8274;
  assign new_n8361 = ~new_n8275 & ~new_n8360;
  assign new_n8362 = new_n8342 & ~new_n8343;
  assign new_n8363 = ~new_n8344 & ~new_n8362;
  assign new_n8364 = ~new_n8260 & ~new_n8264;
  assign new_n8365 = ~new_n8265 & ~new_n8364;
  assign new_n8366 = ~new_n8363 & new_n8365;
  assign new_n8367 = ~new_n8361 & ~new_n8366;
  assign new_n8368 = new_n8328 & ~new_n8351;
  assign new_n8369 = ~new_n8352 & ~new_n8368;
  assign new_n8370 = new_n8361 & new_n8366;
  assign new_n8371 = ~new_n8367 & ~new_n8370;
  assign new_n8372 = new_n8369 & new_n8371;
  assign new_n8373 = ~new_n8367 & ~new_n8372;
  assign new_n8374 = ~new_n8359 & ~new_n8373;
  assign new_n8375 = ~new_n8333 & ~new_n8354;
  assign new_n8376 = ~new_n8355 & ~new_n8375;
  assign new_n8377 = new_n8359 & new_n8373;
  assign new_n8378 = ~new_n8374 & ~new_n8377;
  assign new_n8379 = ~new_n8376 & new_n8378;
  assign new_n8380 = ~new_n8374 & ~new_n8379;
  assign new_n8381 = ~new_n8281 & ~new_n8356;
  assign new_n8382 = ~new_n8357 & ~new_n8381;
  assign new_n8383 = ~new_n8380 & new_n8382;
  assign new_n8384 = ~new_n8357 & ~new_n8383;
  assign new_n8385 = A517 & A518;
  assign new_n8386 = A520 & A521;
  assign new_n8387 = ~new_n8385 & ~new_n8386;
  assign new_n8388 = A519 & A522;
  assign new_n8389 = ~new_n8387 & new_n8388;
  assign new_n8390 = ~A517 & ~A518;
  assign new_n8391 = ~A519 & A522;
  assign new_n8392 = new_n8386 & new_n8391;
  assign new_n8393 = ~A519 & ~new_n8385;
  assign new_n8394 = ~A520 & ~A521;
  assign new_n8395 = ~new_n8386 & ~new_n8394;
  assign new_n8396 = A522 & ~new_n8395;
  assign new_n8397 = ~A522 & ~new_n8386;
  assign new_n8398 = ~new_n8393 & ~new_n8397;
  assign new_n8399 = ~new_n8396 & new_n8398;
  assign new_n8400 = ~new_n8392 & ~new_n8399;
  assign new_n8401 = ~new_n8390 & ~new_n8400;
  assign new_n8402 = A521 & new_n8385;
  assign new_n8403 = new_n8389 & ~new_n8402;
  assign new_n8404 = ~new_n8388 & new_n8390;
  assign new_n8405 = new_n8394 & new_n8404;
  assign new_n8406 = A519 & ~A522;
  assign new_n8407 = new_n8385 & ~new_n8394;
  assign new_n8408 = new_n8406 & new_n8407;
  assign new_n8409 = ~new_n8405 & ~new_n8408;
  assign new_n8410 = ~new_n8403 & new_n8409;
  assign new_n8411 = ~new_n8401 & new_n8410;
  assign new_n8412 = ~new_n8390 & ~new_n8411;
  assign new_n8413 = ~new_n8389 & ~new_n8412;
  assign new_n8414 = ~A512 & ~A513;
  assign new_n8415 = A512 & A513;
  assign new_n8416 = ~new_n8414 & ~new_n8415;
  assign new_n8417 = ~A511 & new_n8416;
  assign new_n8418 = ~new_n8414 & ~new_n8417;
  assign new_n8419 = ~A514 & ~A515;
  assign new_n8420 = new_n8418 & ~new_n8419;
  assign new_n8421 = A514 & A515;
  assign new_n8422 = ~A516 & ~new_n8421;
  assign new_n8423 = new_n8420 & ~new_n8422;
  assign new_n8424 = ~A516 & ~new_n8420;
  assign new_n8425 = A511 & ~new_n8416;
  assign new_n8426 = ~new_n8417 & ~new_n8425;
  assign new_n8427 = ~new_n8418 & ~new_n8421;
  assign new_n8428 = new_n8418 & new_n8421;
  assign new_n8429 = ~new_n8427 & ~new_n8428;
  assign new_n8430 = A516 & ~new_n8429;
  assign new_n8431 = ~new_n8424 & ~new_n8426;
  assign new_n8432 = ~new_n8430 & new_n8431;
  assign new_n8433 = ~new_n8423 & ~new_n8432;
  assign new_n8434 = new_n8413 & new_n8433;
  assign new_n8435 = ~new_n8385 & ~new_n8390;
  assign new_n8436 = ~new_n8391 & ~new_n8406;
  assign new_n8437 = new_n8435 & ~new_n8436;
  assign new_n8438 = ~new_n8435 & new_n8436;
  assign new_n8439 = ~new_n8437 & ~new_n8438;
  assign new_n8440 = new_n8395 & new_n8439;
  assign new_n8441 = new_n8393 & new_n8397;
  assign new_n8442 = ~new_n8440 & new_n8441;
  assign new_n8443 = new_n8411 & ~new_n8442;
  assign new_n8444 = A516 & ~new_n8426;
  assign new_n8445 = ~new_n8418 & new_n8419;
  assign new_n8446 = ~new_n8444 & new_n8445;
  assign new_n8447 = ~new_n8418 & new_n8422;
  assign new_n8448 = ~new_n8423 & ~new_n8447;
  assign new_n8449 = new_n8426 & ~new_n8448;
  assign new_n8450 = ~new_n8432 & ~new_n8446;
  assign new_n8451 = ~new_n8449 & new_n8450;
  assign new_n8452 = ~new_n8443 & ~new_n8451;
  assign new_n8453 = ~new_n8395 & ~new_n8439;
  assign new_n8454 = ~new_n8440 & ~new_n8453;
  assign new_n8455 = ~A516 & new_n8426;
  assign new_n8456 = ~new_n8444 & ~new_n8455;
  assign new_n8457 = ~new_n8419 & ~new_n8421;
  assign new_n8458 = ~new_n8456 & new_n8457;
  assign new_n8459 = new_n8456 & ~new_n8457;
  assign new_n8460 = ~new_n8458 & ~new_n8459;
  assign new_n8461 = new_n8454 & ~new_n8460;
  assign new_n8462 = new_n8443 & new_n8451;
  assign new_n8463 = ~new_n8452 & ~new_n8462;
  assign new_n8464 = ~new_n8461 & new_n8463;
  assign new_n8465 = ~new_n8452 & ~new_n8464;
  assign new_n8466 = ~new_n8413 & ~new_n8433;
  assign new_n8467 = ~new_n8434 & ~new_n8466;
  assign new_n8468 = ~new_n8465 & new_n8467;
  assign new_n8469 = ~new_n8434 & ~new_n8468;
  assign new_n8470 = ~A532 & ~A533;
  assign new_n8471 = A532 & A533;
  assign new_n8472 = ~new_n8470 & ~new_n8471;
  assign new_n8473 = ~A534 & new_n8472;
  assign new_n8474 = ~new_n8470 & ~new_n8473;
  assign new_n8475 = ~A530 & ~A531;
  assign new_n8476 = A530 & A531;
  assign new_n8477 = ~new_n8475 & ~new_n8476;
  assign new_n8478 = ~A529 & new_n8477;
  assign new_n8479 = ~new_n8475 & ~new_n8478;
  assign new_n8480 = ~new_n8474 & ~new_n8479;
  assign new_n8481 = A529 & ~new_n8477;
  assign new_n8482 = ~new_n8478 & ~new_n8481;
  assign new_n8483 = A534 & ~new_n8472;
  assign new_n8484 = ~new_n8473 & ~new_n8483;
  assign new_n8485 = ~new_n8482 & ~new_n8484;
  assign new_n8486 = new_n8474 & new_n8479;
  assign new_n8487 = ~new_n8480 & ~new_n8486;
  assign new_n8488 = ~new_n8485 & new_n8487;
  assign new_n8489 = ~new_n8480 & ~new_n8488;
  assign new_n8490 = A523 & A524;
  assign new_n8491 = ~A527 & ~A528;
  assign new_n8492 = A525 & A526;
  assign new_n8493 = ~new_n8490 & new_n8492;
  assign new_n8494 = ~A525 & ~A526;
  assign new_n8495 = ~new_n8492 & ~new_n8494;
  assign new_n8496 = ~A523 & ~A524;
  assign new_n8497 = ~new_n8490 & ~new_n8496;
  assign new_n8498 = ~new_n8495 & new_n8497;
  assign new_n8499 = ~new_n8492 & ~new_n8496;
  assign new_n8500 = ~new_n8498 & new_n8499;
  assign new_n8501 = ~new_n8493 & ~new_n8500;
  assign new_n8502 = new_n8491 & new_n8501;
  assign new_n8503 = new_n8490 & new_n8502;
  assign new_n8504 = A527 & A528;
  assign new_n8505 = ~new_n8501 & new_n8504;
  assign new_n8506 = ~new_n8503 & ~new_n8505;
  assign new_n8507 = ~new_n8490 & ~new_n8498;
  assign new_n8508 = ~new_n8491 & ~new_n8494;
  assign new_n8509 = ~new_n8507 & new_n8508;
  assign new_n8510 = new_n8506 & ~new_n8509;
  assign new_n8511 = ~new_n8489 & new_n8510;
  assign new_n8512 = new_n8482 & new_n8484;
  assign new_n8513 = ~new_n8485 & ~new_n8512;
  assign new_n8514 = ~new_n8491 & ~new_n8504;
  assign new_n8515 = new_n8495 & ~new_n8497;
  assign new_n8516 = ~new_n8498 & ~new_n8515;
  assign new_n8517 = new_n8514 & ~new_n8516;
  assign new_n8518 = ~new_n8514 & new_n8516;
  assign new_n8519 = ~new_n8517 & ~new_n8518;
  assign new_n8520 = new_n8513 & new_n8519;
  assign new_n8521 = ~new_n8485 & ~new_n8520;
  assign new_n8522 = ~new_n8487 & ~new_n8521;
  assign new_n8523 = ~new_n8488 & ~new_n8522;
  assign new_n8524 = new_n8487 & new_n8520;
  assign new_n8525 = ~new_n8523 & ~new_n8524;
  assign new_n8526 = ~new_n8504 & new_n8509;
  assign new_n8527 = new_n8494 & new_n8496;
  assign new_n8528 = ~new_n8504 & new_n8527;
  assign new_n8529 = ~new_n8502 & ~new_n8528;
  assign new_n8530 = ~new_n8526 & new_n8529;
  assign new_n8531 = new_n8506 & new_n8530;
  assign new_n8532 = new_n8525 & ~new_n8531;
  assign new_n8533 = ~new_n8523 & ~new_n8532;
  assign new_n8534 = new_n8489 & ~new_n8510;
  assign new_n8535 = ~new_n8511 & ~new_n8534;
  assign new_n8536 = ~new_n8533 & new_n8535;
  assign new_n8537 = ~new_n8511 & ~new_n8536;
  assign new_n8538 = new_n8469 & new_n8537;
  assign new_n8539 = new_n8465 & ~new_n8467;
  assign new_n8540 = ~new_n8468 & ~new_n8539;
  assign new_n8541 = ~new_n8454 & new_n8460;
  assign new_n8542 = ~new_n8461 & ~new_n8541;
  assign new_n8543 = ~new_n8513 & ~new_n8519;
  assign new_n8544 = ~new_n8520 & ~new_n8543;
  assign new_n8545 = new_n8542 & new_n8544;
  assign new_n8546 = new_n8463 & new_n8545;
  assign new_n8547 = ~new_n8525 & new_n8531;
  assign new_n8548 = ~new_n8532 & ~new_n8547;
  assign new_n8549 = ~new_n8461 & ~new_n8545;
  assign new_n8550 = new_n8463 & ~new_n8549;
  assign new_n8551 = ~new_n8463 & new_n8549;
  assign new_n8552 = ~new_n8550 & ~new_n8551;
  assign new_n8553 = ~new_n8548 & new_n8552;
  assign new_n8554 = ~new_n8546 & ~new_n8553;
  assign new_n8555 = ~new_n8540 & ~new_n8554;
  assign new_n8556 = new_n8533 & ~new_n8535;
  assign new_n8557 = ~new_n8536 & ~new_n8556;
  assign new_n8558 = new_n8540 & new_n8554;
  assign new_n8559 = ~new_n8555 & ~new_n8558;
  assign new_n8560 = ~new_n8557 & new_n8559;
  assign new_n8561 = ~new_n8555 & ~new_n8560;
  assign new_n8562 = ~new_n8469 & ~new_n8537;
  assign new_n8563 = ~new_n8538 & ~new_n8562;
  assign new_n8564 = ~new_n8561 & new_n8563;
  assign new_n8565 = ~new_n8538 & ~new_n8564;
  assign new_n8566 = ~new_n8384 & new_n8565;
  assign new_n8567 = new_n8380 & ~new_n8382;
  assign new_n8568 = ~new_n8383 & ~new_n8567;
  assign new_n8569 = new_n8557 & ~new_n8559;
  assign new_n8570 = ~new_n8560 & ~new_n8569;
  assign new_n8571 = ~new_n8369 & ~new_n8371;
  assign new_n8572 = ~new_n8372 & ~new_n8571;
  assign new_n8573 = new_n8548 & ~new_n8552;
  assign new_n8574 = ~new_n8553 & ~new_n8573;
  assign new_n8575 = new_n8572 & ~new_n8574;
  assign new_n8576 = ~new_n8572 & new_n8574;
  assign new_n8577 = ~new_n8542 & ~new_n8544;
  assign new_n8578 = ~new_n8545 & ~new_n8577;
  assign new_n8579 = new_n8363 & ~new_n8365;
  assign new_n8580 = ~new_n8366 & ~new_n8579;
  assign new_n8581 = new_n8578 & new_n8580;
  assign new_n8582 = ~new_n8576 & ~new_n8581;
  assign new_n8583 = ~new_n8575 & ~new_n8582;
  assign new_n8584 = new_n8570 & new_n8583;
  assign new_n8585 = new_n8376 & ~new_n8378;
  assign new_n8586 = ~new_n8379 & ~new_n8585;
  assign new_n8587 = ~new_n8570 & ~new_n8583;
  assign new_n8588 = ~new_n8584 & ~new_n8587;
  assign new_n8589 = ~new_n8586 & new_n8588;
  assign new_n8590 = ~new_n8584 & ~new_n8589;
  assign new_n8591 = ~new_n8568 & ~new_n8590;
  assign new_n8592 = new_n8561 & ~new_n8563;
  assign new_n8593 = ~new_n8564 & ~new_n8592;
  assign new_n8594 = new_n8568 & new_n8590;
  assign new_n8595 = ~new_n8591 & ~new_n8594;
  assign new_n8596 = new_n8593 & new_n8595;
  assign new_n8597 = ~new_n8591 & ~new_n8596;
  assign new_n8598 = new_n8384 & ~new_n8565;
  assign new_n8599 = ~new_n8566 & ~new_n8598;
  assign new_n8600 = new_n8597 & new_n8599;
  assign new_n8601 = ~new_n8566 & ~new_n8600;
  assign new_n8602 = ~new_n8214 & new_n8601;
  assign new_n8603 = new_n8214 & ~new_n8601;
  assign new_n8604 = ~new_n8602 & ~new_n8603;
  assign new_n8605 = ~new_n8179 & ~new_n8212;
  assign new_n8606 = ~new_n8213 & ~new_n8605;
  assign new_n8607 = ~new_n8597 & ~new_n8599;
  assign new_n8608 = ~new_n8600 & ~new_n8607;
  assign new_n8609 = ~new_n8606 & new_n8608;
  assign new_n8610 = new_n8606 & ~new_n8608;
  assign new_n8611 = ~new_n8609 & ~new_n8610;
  assign new_n8612 = new_n8201 & ~new_n8203;
  assign new_n8613 = ~new_n8204 & ~new_n8612;
  assign new_n8614 = ~new_n8183 & ~new_n8193;
  assign new_n8615 = ~new_n8194 & ~new_n8614;
  assign new_n8616 = ~new_n8575 & ~new_n8576;
  assign new_n8617 = ~new_n8578 & ~new_n8580;
  assign new_n8618 = ~new_n8581 & ~new_n8617;
  assign new_n8619 = ~new_n8186 & ~new_n8188;
  assign new_n8620 = ~new_n8189 & ~new_n8619;
  assign new_n8621 = new_n8618 & new_n8620;
  assign new_n8622 = ~new_n8581 & ~new_n8621;
  assign new_n8623 = new_n8616 & ~new_n8622;
  assign new_n8624 = ~new_n8616 & new_n8622;
  assign new_n8625 = ~new_n8623 & ~new_n8624;
  assign new_n8626 = ~new_n8615 & new_n8625;
  assign new_n8627 = ~new_n8621 & ~new_n8625;
  assign new_n8628 = ~new_n8626 & ~new_n8627;
  assign new_n8629 = new_n8613 & ~new_n8628;
  assign new_n8630 = new_n8586 & ~new_n8588;
  assign new_n8631 = ~new_n8589 & ~new_n8630;
  assign new_n8632 = ~new_n8613 & new_n8628;
  assign new_n8633 = ~new_n8629 & ~new_n8632;
  assign new_n8634 = ~new_n8631 & new_n8633;
  assign new_n8635 = ~new_n8629 & ~new_n8634;
  assign new_n8636 = ~new_n8593 & ~new_n8595;
  assign new_n8637 = ~new_n8596 & ~new_n8636;
  assign new_n8638 = new_n8635 & new_n8637;
  assign new_n8639 = new_n8208 & ~new_n8210;
  assign new_n8640 = ~new_n8211 & ~new_n8639;
  assign new_n8641 = ~new_n8635 & ~new_n8637;
  assign new_n8642 = ~new_n8638 & ~new_n8641;
  assign new_n8643 = ~new_n8640 & new_n8642;
  assign new_n8644 = ~new_n8638 & ~new_n8643;
  assign new_n8645 = new_n8611 & new_n8644;
  assign new_n8646 = ~new_n8609 & ~new_n8645;
  assign new_n8647 = new_n8604 & new_n8646;
  assign new_n8648 = ~new_n8602 & ~new_n8647;
  assign new_n8649 = ~new_n7767 & ~new_n8648;
  assign new_n8650 = new_n7767 & new_n8648;
  assign new_n8651 = ~new_n8649 & ~new_n8650;
  assign new_n8652 = ~new_n7724 & new_n7765;
  assign new_n8653 = ~new_n7766 & ~new_n8652;
  assign new_n8654 = ~new_n8611 & ~new_n8644;
  assign new_n8655 = ~new_n8645 & ~new_n8654;
  assign new_n8656 = new_n8640 & ~new_n8642;
  assign new_n8657 = ~new_n8643 & ~new_n8656;
  assign new_n8658 = ~new_n7754 & ~new_n7756;
  assign new_n8659 = ~new_n7757 & ~new_n8658;
  assign new_n8660 = new_n8657 & new_n8659;
  assign new_n8661 = new_n7747 & ~new_n7749;
  assign new_n8662 = ~new_n7750 & ~new_n8661;
  assign new_n8663 = ~new_n7740 & ~new_n7742;
  assign new_n8664 = ~new_n7743 & ~new_n8663;
  assign new_n8665 = ~new_n8618 & ~new_n8620;
  assign new_n8666 = ~new_n8621 & ~new_n8665;
  assign new_n8667 = ~new_n7734 & ~new_n7736;
  assign new_n8668 = ~new_n7737 & ~new_n8667;
  assign new_n8669 = new_n8666 & new_n8668;
  assign new_n8670 = ~new_n8664 & new_n8669;
  assign new_n8671 = new_n8615 & ~new_n8625;
  assign new_n8672 = ~new_n8626 & ~new_n8671;
  assign new_n8673 = new_n8664 & ~new_n8669;
  assign new_n8674 = ~new_n8670 & ~new_n8673;
  assign new_n8675 = ~new_n8672 & new_n8674;
  assign new_n8676 = ~new_n8670 & ~new_n8675;
  assign new_n8677 = ~new_n8662 & ~new_n8676;
  assign new_n8678 = new_n8631 & ~new_n8633;
  assign new_n8679 = ~new_n8634 & ~new_n8678;
  assign new_n8680 = new_n8662 & new_n8676;
  assign new_n8681 = ~new_n8677 & ~new_n8680;
  assign new_n8682 = ~new_n8679 & new_n8681;
  assign new_n8683 = ~new_n8677 & ~new_n8682;
  assign new_n8684 = ~new_n8657 & ~new_n8659;
  assign new_n8685 = ~new_n8660 & ~new_n8684;
  assign new_n8686 = ~new_n8683 & new_n8685;
  assign new_n8687 = ~new_n8660 & ~new_n8686;
  assign new_n8688 = ~new_n8655 & ~new_n8687;
  assign new_n8689 = new_n7761 & ~new_n7763;
  assign new_n8690 = ~new_n7764 & ~new_n8689;
  assign new_n8691 = new_n8655 & new_n8687;
  assign new_n8692 = ~new_n8688 & ~new_n8691;
  assign new_n8693 = new_n8690 & new_n8692;
  assign new_n8694 = ~new_n8688 & ~new_n8693;
  assign new_n8695 = ~new_n8653 & new_n8694;
  assign new_n8696 = ~new_n8604 & ~new_n8646;
  assign new_n8697 = ~new_n8647 & ~new_n8696;
  assign new_n8698 = new_n8653 & ~new_n8694;
  assign new_n8699 = ~new_n8695 & ~new_n8698;
  assign new_n8700 = ~new_n8697 & new_n8699;
  assign new_n8701 = ~new_n8695 & ~new_n8700;
  assign new_n8702 = new_n8651 & new_n8701;
  assign new_n8703 = ~new_n8649 & ~new_n8702;
  assign new_n8704 = A757 & A758;
  assign new_n8705 = A760 & A761;
  assign new_n8706 = ~new_n8704 & ~new_n8705;
  assign new_n8707 = A759 & A762;
  assign new_n8708 = ~new_n8706 & new_n8707;
  assign new_n8709 = ~A757 & ~A758;
  assign new_n8710 = ~A759 & A762;
  assign new_n8711 = new_n8705 & new_n8710;
  assign new_n8712 = ~A759 & ~new_n8704;
  assign new_n8713 = ~A760 & ~A761;
  assign new_n8714 = ~new_n8705 & ~new_n8713;
  assign new_n8715 = A762 & ~new_n8714;
  assign new_n8716 = ~A762 & ~new_n8705;
  assign new_n8717 = ~new_n8712 & ~new_n8716;
  assign new_n8718 = ~new_n8715 & new_n8717;
  assign new_n8719 = ~new_n8711 & ~new_n8718;
  assign new_n8720 = ~new_n8709 & ~new_n8719;
  assign new_n8721 = A761 & new_n8704;
  assign new_n8722 = new_n8708 & ~new_n8721;
  assign new_n8723 = ~new_n8707 & new_n8709;
  assign new_n8724 = new_n8713 & new_n8723;
  assign new_n8725 = A759 & ~A762;
  assign new_n8726 = new_n8704 & ~new_n8713;
  assign new_n8727 = new_n8725 & new_n8726;
  assign new_n8728 = ~new_n8724 & ~new_n8727;
  assign new_n8729 = ~new_n8722 & new_n8728;
  assign new_n8730 = ~new_n8720 & new_n8729;
  assign new_n8731 = ~new_n8709 & ~new_n8730;
  assign new_n8732 = ~new_n8708 & ~new_n8731;
  assign new_n8733 = A751 & A752;
  assign new_n8734 = A754 & A755;
  assign new_n8735 = ~new_n8733 & ~new_n8734;
  assign new_n8736 = A753 & A756;
  assign new_n8737 = ~new_n8735 & new_n8736;
  assign new_n8738 = ~A751 & ~A752;
  assign new_n8739 = ~A753 & A756;
  assign new_n8740 = new_n8734 & new_n8739;
  assign new_n8741 = ~A753 & ~new_n8733;
  assign new_n8742 = ~A754 & ~A755;
  assign new_n8743 = ~new_n8734 & ~new_n8742;
  assign new_n8744 = A756 & ~new_n8743;
  assign new_n8745 = ~A756 & ~new_n8734;
  assign new_n8746 = ~new_n8741 & ~new_n8745;
  assign new_n8747 = ~new_n8744 & new_n8746;
  assign new_n8748 = ~new_n8740 & ~new_n8747;
  assign new_n8749 = ~new_n8738 & ~new_n8748;
  assign new_n8750 = A755 & new_n8733;
  assign new_n8751 = new_n8737 & ~new_n8750;
  assign new_n8752 = ~new_n8736 & new_n8738;
  assign new_n8753 = new_n8742 & new_n8752;
  assign new_n8754 = A753 & ~A756;
  assign new_n8755 = new_n8733 & ~new_n8742;
  assign new_n8756 = new_n8754 & new_n8755;
  assign new_n8757 = ~new_n8753 & ~new_n8756;
  assign new_n8758 = ~new_n8751 & new_n8757;
  assign new_n8759 = ~new_n8749 & new_n8758;
  assign new_n8760 = ~new_n8738 & ~new_n8759;
  assign new_n8761 = ~new_n8737 & ~new_n8760;
  assign new_n8762 = new_n8732 & new_n8761;
  assign new_n8763 = ~new_n8733 & ~new_n8738;
  assign new_n8764 = ~new_n8739 & ~new_n8754;
  assign new_n8765 = new_n8763 & ~new_n8764;
  assign new_n8766 = ~new_n8763 & new_n8764;
  assign new_n8767 = ~new_n8765 & ~new_n8766;
  assign new_n8768 = new_n8743 & new_n8767;
  assign new_n8769 = ~new_n8743 & ~new_n8767;
  assign new_n8770 = ~new_n8768 & ~new_n8769;
  assign new_n8771 = ~new_n8704 & ~new_n8709;
  assign new_n8772 = ~new_n8710 & ~new_n8725;
  assign new_n8773 = new_n8771 & ~new_n8772;
  assign new_n8774 = ~new_n8771 & new_n8772;
  assign new_n8775 = ~new_n8773 & ~new_n8774;
  assign new_n8776 = new_n8714 & new_n8775;
  assign new_n8777 = ~new_n8714 & ~new_n8775;
  assign new_n8778 = ~new_n8776 & ~new_n8777;
  assign new_n8779 = new_n8770 & new_n8778;
  assign new_n8780 = new_n8712 & new_n8716;
  assign new_n8781 = ~new_n8776 & new_n8780;
  assign new_n8782 = new_n8730 & ~new_n8781;
  assign new_n8783 = ~new_n8779 & ~new_n8782;
  assign new_n8784 = new_n8779 & new_n8782;
  assign new_n8785 = ~new_n8783 & ~new_n8784;
  assign new_n8786 = new_n8741 & new_n8745;
  assign new_n8787 = ~new_n8768 & new_n8786;
  assign new_n8788 = new_n8759 & ~new_n8787;
  assign new_n8789 = new_n8785 & ~new_n8788;
  assign new_n8790 = ~new_n8783 & ~new_n8789;
  assign new_n8791 = ~new_n8732 & ~new_n8761;
  assign new_n8792 = ~new_n8762 & ~new_n8791;
  assign new_n8793 = ~new_n8790 & new_n8792;
  assign new_n8794 = ~new_n8762 & ~new_n8793;
  assign new_n8795 = ~A773 & ~A774;
  assign new_n8796 = A773 & A774;
  assign new_n8797 = ~new_n8795 & ~new_n8796;
  assign new_n8798 = ~A772 & new_n8797;
  assign new_n8799 = ~new_n8795 & ~new_n8798;
  assign new_n8800 = ~A770 & ~A771;
  assign new_n8801 = A770 & A771;
  assign new_n8802 = ~new_n8800 & ~new_n8801;
  assign new_n8803 = ~A769 & new_n8802;
  assign new_n8804 = ~new_n8800 & ~new_n8803;
  assign new_n8805 = ~new_n8799 & ~new_n8804;
  assign new_n8806 = A769 & ~new_n8802;
  assign new_n8807 = ~new_n8803 & ~new_n8806;
  assign new_n8808 = A772 & ~new_n8797;
  assign new_n8809 = ~new_n8798 & ~new_n8808;
  assign new_n8810 = ~new_n8807 & ~new_n8809;
  assign new_n8811 = new_n8799 & new_n8804;
  assign new_n8812 = ~new_n8805 & ~new_n8811;
  assign new_n8813 = ~new_n8810 & new_n8812;
  assign new_n8814 = ~new_n8805 & ~new_n8813;
  assign new_n8815 = A763 & A764;
  assign new_n8816 = ~A767 & ~A768;
  assign new_n8817 = A765 & A766;
  assign new_n8818 = ~new_n8815 & new_n8817;
  assign new_n8819 = ~A765 & ~A766;
  assign new_n8820 = ~new_n8817 & ~new_n8819;
  assign new_n8821 = ~A763 & ~A764;
  assign new_n8822 = ~new_n8815 & ~new_n8821;
  assign new_n8823 = ~new_n8820 & new_n8822;
  assign new_n8824 = ~new_n8817 & ~new_n8821;
  assign new_n8825 = ~new_n8823 & new_n8824;
  assign new_n8826 = ~new_n8818 & ~new_n8825;
  assign new_n8827 = new_n8816 & new_n8826;
  assign new_n8828 = new_n8815 & new_n8827;
  assign new_n8829 = A767 & A768;
  assign new_n8830 = ~new_n8826 & new_n8829;
  assign new_n8831 = ~new_n8828 & ~new_n8830;
  assign new_n8832 = ~new_n8815 & ~new_n8823;
  assign new_n8833 = ~new_n8816 & ~new_n8819;
  assign new_n8834 = ~new_n8832 & new_n8833;
  assign new_n8835 = new_n8831 & ~new_n8834;
  assign new_n8836 = ~new_n8814 & new_n8835;
  assign new_n8837 = new_n8807 & new_n8809;
  assign new_n8838 = ~new_n8810 & ~new_n8837;
  assign new_n8839 = ~new_n8816 & ~new_n8829;
  assign new_n8840 = new_n8820 & ~new_n8822;
  assign new_n8841 = ~new_n8823 & ~new_n8840;
  assign new_n8842 = new_n8839 & ~new_n8841;
  assign new_n8843 = ~new_n8839 & new_n8841;
  assign new_n8844 = ~new_n8842 & ~new_n8843;
  assign new_n8845 = new_n8838 & ~new_n8844;
  assign new_n8846 = ~new_n8837 & ~new_n8845;
  assign new_n8847 = ~new_n8812 & new_n8846;
  assign new_n8848 = new_n8812 & ~new_n8846;
  assign new_n8849 = ~new_n8847 & ~new_n8848;
  assign new_n8850 = ~new_n8829 & new_n8834;
  assign new_n8851 = new_n8819 & new_n8821;
  assign new_n8852 = ~new_n8829 & new_n8851;
  assign new_n8853 = ~new_n8827 & ~new_n8852;
  assign new_n8854 = ~new_n8850 & new_n8853;
  assign new_n8855 = new_n8831 & new_n8854;
  assign new_n8856 = ~new_n8849 & ~new_n8855;
  assign new_n8857 = ~new_n8813 & ~new_n8847;
  assign new_n8858 = ~new_n8856 & ~new_n8857;
  assign new_n8859 = new_n8814 & ~new_n8835;
  assign new_n8860 = ~new_n8836 & ~new_n8859;
  assign new_n8861 = ~new_n8858 & new_n8860;
  assign new_n8862 = ~new_n8836 & ~new_n8861;
  assign new_n8863 = ~new_n8794 & ~new_n8862;
  assign new_n8864 = new_n8794 & new_n8862;
  assign new_n8865 = ~new_n8863 & ~new_n8864;
  assign new_n8866 = new_n8790 & ~new_n8792;
  assign new_n8867 = ~new_n8793 & ~new_n8866;
  assign new_n8868 = ~new_n8785 & new_n8788;
  assign new_n8869 = ~new_n8789 & ~new_n8868;
  assign new_n8870 = ~new_n8770 & ~new_n8778;
  assign new_n8871 = ~new_n8779 & ~new_n8870;
  assign new_n8872 = ~new_n8838 & new_n8844;
  assign new_n8873 = ~new_n8845 & ~new_n8872;
  assign new_n8874 = new_n8871 & ~new_n8873;
  assign new_n8875 = ~new_n8869 & new_n8874;
  assign new_n8876 = new_n8849 & new_n8855;
  assign new_n8877 = ~new_n8856 & ~new_n8876;
  assign new_n8878 = new_n8869 & ~new_n8874;
  assign new_n8879 = ~new_n8875 & ~new_n8878;
  assign new_n8880 = ~new_n8877 & new_n8879;
  assign new_n8881 = ~new_n8875 & ~new_n8880;
  assign new_n8882 = ~new_n8867 & ~new_n8881;
  assign new_n8883 = new_n8858 & ~new_n8860;
  assign new_n8884 = ~new_n8861 & ~new_n8883;
  assign new_n8885 = new_n8867 & new_n8881;
  assign new_n8886 = ~new_n8882 & ~new_n8885;
  assign new_n8887 = ~new_n8884 & new_n8886;
  assign new_n8888 = ~new_n8882 & ~new_n8887;
  assign new_n8889 = new_n8865 & new_n8888;
  assign new_n8890 = ~new_n8863 & ~new_n8889;
  assign new_n8891 = ~A793 & ~A794;
  assign new_n8892 = A793 & A794;
  assign new_n8893 = ~A795 & ~new_n8892;
  assign new_n8894 = ~new_n8891 & ~new_n8893;
  assign new_n8895 = A797 & A798;
  assign new_n8896 = new_n8894 & new_n8895;
  assign new_n8897 = A795 & new_n8892;
  assign new_n8898 = ~A796 & ~new_n8897;
  assign new_n8899 = new_n8894 & ~new_n8898;
  assign new_n8900 = A797 & new_n8899;
  assign new_n8901 = A795 & A796;
  assign new_n8902 = new_n8892 & new_n8901;
  assign new_n8903 = ~new_n8900 & ~new_n8902;
  assign new_n8904 = ~A798 & ~new_n8903;
  assign new_n8905 = ~A797 & ~A798;
  assign new_n8906 = ~new_n8891 & ~new_n8905;
  assign new_n8907 = new_n8893 & ~new_n8895;
  assign new_n8908 = ~new_n8906 & new_n8907;
  assign new_n8909 = ~new_n8896 & ~new_n8908;
  assign new_n8910 = ~A796 & ~new_n8909;
  assign new_n8911 = ~A797 & A798;
  assign new_n8912 = new_n8899 & new_n8911;
  assign new_n8913 = new_n8891 & ~new_n8901;
  assign new_n8914 = A796 & new_n8895;
  assign new_n8915 = ~new_n8897 & new_n8914;
  assign new_n8916 = ~new_n8913 & new_n8915;
  assign new_n8917 = ~new_n8912 & ~new_n8916;
  assign new_n8918 = ~new_n8910 & new_n8917;
  assign new_n8919 = ~new_n8904 & new_n8918;
  assign new_n8920 = ~new_n8898 & ~new_n8919;
  assign new_n8921 = ~new_n8896 & ~new_n8920;
  assign new_n8922 = ~A788 & ~A789;
  assign new_n8923 = A788 & A789;
  assign new_n8924 = ~new_n8922 & ~new_n8923;
  assign new_n8925 = ~A787 & new_n8924;
  assign new_n8926 = ~new_n8922 & ~new_n8925;
  assign new_n8927 = ~A790 & ~A791;
  assign new_n8928 = new_n8926 & ~new_n8927;
  assign new_n8929 = A790 & A791;
  assign new_n8930 = ~A792 & ~new_n8929;
  assign new_n8931 = new_n8928 & ~new_n8930;
  assign new_n8932 = ~A792 & ~new_n8928;
  assign new_n8933 = A787 & ~new_n8924;
  assign new_n8934 = ~new_n8925 & ~new_n8933;
  assign new_n8935 = ~new_n8926 & ~new_n8929;
  assign new_n8936 = new_n8926 & new_n8929;
  assign new_n8937 = ~new_n8935 & ~new_n8936;
  assign new_n8938 = A792 & ~new_n8937;
  assign new_n8939 = ~new_n8932 & ~new_n8934;
  assign new_n8940 = ~new_n8938 & new_n8939;
  assign new_n8941 = ~new_n8931 & ~new_n8940;
  assign new_n8942 = ~new_n8921 & ~new_n8941;
  assign new_n8943 = new_n8921 & new_n8941;
  assign new_n8944 = ~new_n8942 & ~new_n8943;
  assign new_n8945 = A795 & ~A798;
  assign new_n8946 = ~A795 & A798;
  assign new_n8947 = ~new_n8945 & ~new_n8946;
  assign new_n8948 = ~new_n8891 & ~new_n8892;
  assign new_n8949 = ~A796 & ~A797;
  assign new_n8950 = A796 & A797;
  assign new_n8951 = ~new_n8949 & ~new_n8950;
  assign new_n8952 = new_n8948 & ~new_n8951;
  assign new_n8953 = ~new_n8948 & new_n8951;
  assign new_n8954 = ~new_n8952 & ~new_n8953;
  assign new_n8955 = new_n8947 & new_n8954;
  assign new_n8956 = ~new_n8947 & ~new_n8954;
  assign new_n8957 = ~new_n8955 & ~new_n8956;
  assign new_n8958 = A792 & ~new_n8934;
  assign new_n8959 = ~A792 & new_n8934;
  assign new_n8960 = ~new_n8958 & ~new_n8959;
  assign new_n8961 = ~new_n8927 & ~new_n8929;
  assign new_n8962 = ~new_n8960 & new_n8961;
  assign new_n8963 = new_n8960 & ~new_n8961;
  assign new_n8964 = ~new_n8962 & ~new_n8963;
  assign new_n8965 = new_n8957 & ~new_n8964;
  assign new_n8966 = ~new_n8926 & new_n8927;
  assign new_n8967 = ~new_n8958 & new_n8966;
  assign new_n8968 = ~new_n8926 & new_n8930;
  assign new_n8969 = ~new_n8931 & ~new_n8968;
  assign new_n8970 = new_n8934 & ~new_n8969;
  assign new_n8971 = ~new_n8940 & ~new_n8967;
  assign new_n8972 = ~new_n8970 & new_n8971;
  assign new_n8973 = ~new_n8965 & ~new_n8972;
  assign new_n8974 = new_n8905 & new_n8913;
  assign new_n8975 = new_n8919 & ~new_n8974;
  assign new_n8976 = new_n8965 & new_n8972;
  assign new_n8977 = ~new_n8973 & ~new_n8976;
  assign new_n8978 = ~new_n8975 & new_n8977;
  assign new_n8979 = ~new_n8973 & ~new_n8978;
  assign new_n8980 = new_n8944 & new_n8979;
  assign new_n8981 = ~new_n8942 & ~new_n8980;
  assign new_n8982 = A775 & A776;
  assign new_n8983 = A778 & A779;
  assign new_n8984 = ~new_n8982 & ~new_n8983;
  assign new_n8985 = A777 & A780;
  assign new_n8986 = ~new_n8984 & new_n8985;
  assign new_n8987 = ~A775 & ~A776;
  assign new_n8988 = ~A777 & A780;
  assign new_n8989 = new_n8983 & new_n8988;
  assign new_n8990 = ~A777 & ~new_n8982;
  assign new_n8991 = ~A778 & ~A779;
  assign new_n8992 = ~new_n8983 & ~new_n8991;
  assign new_n8993 = A780 & ~new_n8992;
  assign new_n8994 = ~A780 & ~new_n8983;
  assign new_n8995 = ~new_n8990 & ~new_n8994;
  assign new_n8996 = ~new_n8993 & new_n8995;
  assign new_n8997 = ~new_n8989 & ~new_n8996;
  assign new_n8998 = ~new_n8987 & ~new_n8997;
  assign new_n8999 = A779 & new_n8982;
  assign new_n9000 = new_n8986 & ~new_n8999;
  assign new_n9001 = A777 & ~A780;
  assign new_n9002 = new_n8982 & ~new_n8991;
  assign new_n9003 = new_n9001 & new_n9002;
  assign new_n9004 = ~new_n8985 & new_n8987;
  assign new_n9005 = new_n8991 & new_n9004;
  assign new_n9006 = ~new_n9003 & ~new_n9005;
  assign new_n9007 = ~new_n9000 & new_n9006;
  assign new_n9008 = ~new_n8998 & new_n9007;
  assign new_n9009 = ~new_n8987 & ~new_n9008;
  assign new_n9010 = ~new_n8986 & ~new_n9009;
  assign new_n9011 = A781 & A782;
  assign new_n9012 = A784 & A785;
  assign new_n9013 = ~new_n9011 & ~new_n9012;
  assign new_n9014 = A783 & A786;
  assign new_n9015 = ~new_n9013 & new_n9014;
  assign new_n9016 = ~A781 & ~A782;
  assign new_n9017 = ~A783 & A786;
  assign new_n9018 = new_n9012 & new_n9017;
  assign new_n9019 = ~A783 & ~new_n9011;
  assign new_n9020 = ~A784 & ~A785;
  assign new_n9021 = ~new_n9012 & ~new_n9020;
  assign new_n9022 = A786 & ~new_n9021;
  assign new_n9023 = ~A786 & ~new_n9012;
  assign new_n9024 = ~new_n9019 & ~new_n9023;
  assign new_n9025 = ~new_n9022 & new_n9024;
  assign new_n9026 = ~new_n9018 & ~new_n9025;
  assign new_n9027 = ~new_n9016 & ~new_n9026;
  assign new_n9028 = A785 & new_n9011;
  assign new_n9029 = new_n9015 & ~new_n9028;
  assign new_n9030 = A783 & ~A786;
  assign new_n9031 = new_n9011 & ~new_n9020;
  assign new_n9032 = new_n9030 & new_n9031;
  assign new_n9033 = ~new_n9014 & new_n9016;
  assign new_n9034 = new_n9020 & new_n9033;
  assign new_n9035 = ~new_n9032 & ~new_n9034;
  assign new_n9036 = ~new_n9029 & new_n9035;
  assign new_n9037 = ~new_n9027 & new_n9036;
  assign new_n9038 = ~new_n9016 & ~new_n9037;
  assign new_n9039 = ~new_n9015 & ~new_n9038;
  assign new_n9040 = new_n9010 & new_n9039;
  assign new_n9041 = ~new_n9011 & ~new_n9016;
  assign new_n9042 = ~new_n9017 & ~new_n9030;
  assign new_n9043 = new_n9041 & ~new_n9042;
  assign new_n9044 = ~new_n9041 & new_n9042;
  assign new_n9045 = ~new_n9043 & ~new_n9044;
  assign new_n9046 = new_n9021 & new_n9045;
  assign new_n9047 = new_n9019 & new_n9023;
  assign new_n9048 = ~new_n9046 & new_n9047;
  assign new_n9049 = new_n9037 & ~new_n9048;
  assign new_n9050 = ~new_n8982 & ~new_n8987;
  assign new_n9051 = ~new_n8988 & ~new_n9001;
  assign new_n9052 = new_n9050 & ~new_n9051;
  assign new_n9053 = ~new_n9050 & new_n9051;
  assign new_n9054 = ~new_n9052 & ~new_n9053;
  assign new_n9055 = new_n8992 & new_n9054;
  assign new_n9056 = new_n8990 & new_n8994;
  assign new_n9057 = ~new_n9055 & new_n9056;
  assign new_n9058 = new_n9008 & ~new_n9057;
  assign new_n9059 = ~new_n9049 & ~new_n9058;
  assign new_n9060 = new_n9049 & new_n9058;
  assign new_n9061 = ~new_n9021 & ~new_n9045;
  assign new_n9062 = ~new_n9046 & ~new_n9061;
  assign new_n9063 = ~new_n8992 & ~new_n9054;
  assign new_n9064 = ~new_n9055 & ~new_n9063;
  assign new_n9065 = new_n9062 & new_n9064;
  assign new_n9066 = ~new_n9060 & ~new_n9065;
  assign new_n9067 = ~new_n9059 & ~new_n9066;
  assign new_n9068 = ~new_n9010 & ~new_n9039;
  assign new_n9069 = ~new_n9040 & ~new_n9068;
  assign new_n9070 = ~new_n9067 & new_n9069;
  assign new_n9071 = ~new_n9040 & ~new_n9070;
  assign new_n9072 = ~new_n8981 & new_n9071;
  assign new_n9073 = ~new_n8944 & ~new_n8979;
  assign new_n9074 = ~new_n8980 & ~new_n9073;
  assign new_n9075 = new_n9067 & ~new_n9069;
  assign new_n9076 = ~new_n9070 & ~new_n9075;
  assign new_n9077 = new_n9074 & ~new_n9076;
  assign new_n9078 = ~new_n9074 & new_n9076;
  assign new_n9079 = ~new_n9077 & ~new_n9078;
  assign new_n9080 = new_n8975 & ~new_n8977;
  assign new_n9081 = ~new_n8978 & ~new_n9080;
  assign new_n9082 = ~new_n9062 & ~new_n9064;
  assign new_n9083 = ~new_n9065 & ~new_n9082;
  assign new_n9084 = ~new_n8957 & new_n8964;
  assign new_n9085 = ~new_n8965 & ~new_n9084;
  assign new_n9086 = new_n9083 & new_n9085;
  assign new_n9087 = new_n9081 & ~new_n9086;
  assign new_n9088 = ~new_n9081 & new_n9086;
  assign new_n9089 = ~new_n9065 & ~new_n9086;
  assign new_n9090 = ~new_n9059 & ~new_n9060;
  assign new_n9091 = new_n9081 & ~new_n9090;
  assign new_n9092 = ~new_n9081 & new_n9090;
  assign new_n9093 = ~new_n9091 & ~new_n9092;
  assign new_n9094 = new_n9089 & new_n9093;
  assign new_n9095 = ~new_n9089 & ~new_n9093;
  assign new_n9096 = ~new_n9094 & ~new_n9095;
  assign new_n9097 = ~new_n9088 & ~new_n9096;
  assign new_n9098 = ~new_n9087 & ~new_n9097;
  assign new_n9099 = new_n9079 & new_n9098;
  assign new_n9100 = ~new_n9077 & ~new_n9099;
  assign new_n9101 = new_n8981 & ~new_n9071;
  assign new_n9102 = ~new_n9072 & ~new_n9101;
  assign new_n9103 = ~new_n9100 & new_n9102;
  assign new_n9104 = ~new_n9072 & ~new_n9103;
  assign new_n9105 = ~new_n8890 & new_n9104;
  assign new_n9106 = new_n8890 & ~new_n9104;
  assign new_n9107 = ~new_n9105 & ~new_n9106;
  assign new_n9108 = ~new_n8865 & ~new_n8888;
  assign new_n9109 = ~new_n8889 & ~new_n9108;
  assign new_n9110 = new_n8884 & ~new_n8886;
  assign new_n9111 = ~new_n8887 & ~new_n9110;
  assign new_n9112 = new_n8877 & ~new_n8879;
  assign new_n9113 = ~new_n8880 & ~new_n9112;
  assign new_n9114 = ~new_n9096 & new_n9113;
  assign new_n9115 = new_n9096 & ~new_n9113;
  assign new_n9116 = ~new_n9083 & ~new_n9085;
  assign new_n9117 = ~new_n9086 & ~new_n9116;
  assign new_n9118 = ~new_n8871 & new_n8873;
  assign new_n9119 = ~new_n8874 & ~new_n9118;
  assign new_n9120 = new_n9117 & new_n9119;
  assign new_n9121 = ~new_n9115 & new_n9120;
  assign new_n9122 = ~new_n9114 & ~new_n9121;
  assign new_n9123 = ~new_n9111 & new_n9122;
  assign new_n9124 = ~new_n9079 & ~new_n9098;
  assign new_n9125 = ~new_n9099 & ~new_n9124;
  assign new_n9126 = new_n9111 & ~new_n9122;
  assign new_n9127 = ~new_n9123 & ~new_n9126;
  assign new_n9128 = ~new_n9125 & new_n9127;
  assign new_n9129 = ~new_n9123 & ~new_n9128;
  assign new_n9130 = new_n9109 & ~new_n9129;
  assign new_n9131 = new_n9100 & ~new_n9102;
  assign new_n9132 = ~new_n9103 & ~new_n9131;
  assign new_n9133 = ~new_n9109 & new_n9129;
  assign new_n9134 = ~new_n9130 & ~new_n9133;
  assign new_n9135 = ~new_n9132 & new_n9134;
  assign new_n9136 = ~new_n9130 & ~new_n9135;
  assign new_n9137 = new_n9107 & ~new_n9136;
  assign new_n9138 = ~new_n9105 & ~new_n9137;
  assign new_n9139 = ~A824 & ~A825;
  assign new_n9140 = A824 & A825;
  assign new_n9141 = ~new_n9139 & ~new_n9140;
  assign new_n9142 = ~A823 & new_n9141;
  assign new_n9143 = ~new_n9139 & ~new_n9142;
  assign new_n9144 = ~A826 & ~A827;
  assign new_n9145 = new_n9143 & ~new_n9144;
  assign new_n9146 = A826 & A827;
  assign new_n9147 = ~A828 & ~new_n9146;
  assign new_n9148 = new_n9145 & ~new_n9147;
  assign new_n9149 = ~A828 & ~new_n9145;
  assign new_n9150 = A823 & ~new_n9141;
  assign new_n9151 = ~new_n9142 & ~new_n9150;
  assign new_n9152 = ~new_n9143 & ~new_n9146;
  assign new_n9153 = new_n9143 & new_n9146;
  assign new_n9154 = ~new_n9152 & ~new_n9153;
  assign new_n9155 = A828 & ~new_n9154;
  assign new_n9156 = ~new_n9149 & ~new_n9151;
  assign new_n9157 = ~new_n9155 & new_n9156;
  assign new_n9158 = ~new_n9148 & ~new_n9157;
  assign new_n9159 = ~A833 & ~A834;
  assign new_n9160 = A829 & A830;
  assign new_n9161 = A831 & A832;
  assign new_n9162 = ~new_n9160 & ~new_n9161;
  assign new_n9163 = ~A829 & ~A830;
  assign new_n9164 = ~A831 & ~A832;
  assign new_n9165 = ~new_n9163 & ~new_n9164;
  assign new_n9166 = ~new_n9159 & ~new_n9162;
  assign new_n9167 = new_n9165 & new_n9166;
  assign new_n9168 = new_n9162 & ~new_n9165;
  assign new_n9169 = new_n9160 & new_n9161;
  assign new_n9170 = ~new_n9168 & ~new_n9169;
  assign new_n9171 = ~new_n9159 & ~new_n9170;
  assign new_n9172 = A833 & A834;
  assign new_n9173 = ~new_n9169 & ~new_n9172;
  assign new_n9174 = ~new_n9171 & ~new_n9173;
  assign new_n9175 = ~new_n9167 & ~new_n9174;
  assign new_n9176 = new_n9158 & new_n9175;
  assign new_n9177 = new_n9163 & new_n9164;
  assign new_n9178 = ~new_n9167 & ~new_n9177;
  assign new_n9179 = ~new_n9172 & ~new_n9178;
  assign new_n9180 = new_n9159 & ~new_n9170;
  assign new_n9181 = ~new_n9174 & ~new_n9180;
  assign new_n9182 = ~new_n9179 & new_n9181;
  assign new_n9183 = A828 & ~new_n9151;
  assign new_n9184 = ~new_n9143 & new_n9144;
  assign new_n9185 = ~new_n9183 & new_n9184;
  assign new_n9186 = ~new_n9143 & new_n9147;
  assign new_n9187 = ~new_n9148 & ~new_n9186;
  assign new_n9188 = new_n9151 & ~new_n9187;
  assign new_n9189 = ~new_n9157 & ~new_n9185;
  assign new_n9190 = ~new_n9188 & new_n9189;
  assign new_n9191 = ~new_n9182 & ~new_n9190;
  assign new_n9192 = ~new_n9159 & ~new_n9172;
  assign new_n9193 = ~new_n9161 & ~new_n9164;
  assign new_n9194 = ~new_n9192 & new_n9193;
  assign new_n9195 = new_n9192 & ~new_n9193;
  assign new_n9196 = ~new_n9194 & ~new_n9195;
  assign new_n9197 = ~new_n9160 & ~new_n9163;
  assign new_n9198 = ~new_n9196 & new_n9197;
  assign new_n9199 = new_n9196 & ~new_n9197;
  assign new_n9200 = ~new_n9198 & ~new_n9199;
  assign new_n9201 = ~new_n9144 & ~new_n9146;
  assign new_n9202 = ~A828 & new_n9151;
  assign new_n9203 = ~new_n9183 & ~new_n9202;
  assign new_n9204 = new_n9201 & new_n9203;
  assign new_n9205 = ~new_n9201 & ~new_n9203;
  assign new_n9206 = ~new_n9204 & ~new_n9205;
  assign new_n9207 = new_n9200 & new_n9206;
  assign new_n9208 = new_n9182 & new_n9190;
  assign new_n9209 = ~new_n9191 & ~new_n9208;
  assign new_n9210 = ~new_n9207 & new_n9209;
  assign new_n9211 = ~new_n9191 & ~new_n9210;
  assign new_n9212 = ~new_n9158 & ~new_n9175;
  assign new_n9213 = ~new_n9176 & ~new_n9212;
  assign new_n9214 = ~new_n9211 & new_n9213;
  assign new_n9215 = ~new_n9176 & ~new_n9214;
  assign new_n9216 = ~A842 & ~A843;
  assign new_n9217 = A842 & A843;
  assign new_n9218 = ~new_n9216 & ~new_n9217;
  assign new_n9219 = ~A841 & new_n9218;
  assign new_n9220 = ~new_n9216 & ~new_n9219;
  assign new_n9221 = ~A844 & ~A846;
  assign new_n9222 = A844 & A846;
  assign new_n9223 = ~new_n9221 & ~new_n9222;
  assign new_n9224 = ~A845 & new_n9223;
  assign new_n9225 = ~new_n9221 & ~new_n9224;
  assign new_n9226 = ~new_n9220 & ~new_n9225;
  assign new_n9227 = A845 & ~new_n9223;
  assign new_n9228 = ~new_n9224 & ~new_n9227;
  assign new_n9229 = A841 & ~new_n9218;
  assign new_n9230 = ~new_n9219 & ~new_n9229;
  assign new_n9231 = ~new_n9228 & ~new_n9230;
  assign new_n9232 = new_n9220 & new_n9225;
  assign new_n9233 = ~new_n9226 & ~new_n9232;
  assign new_n9234 = ~new_n9231 & new_n9233;
  assign new_n9235 = ~new_n9226 & ~new_n9234;
  assign new_n9236 = A835 & A836;
  assign new_n9237 = ~A839 & ~A840;
  assign new_n9238 = ~A835 & ~A836;
  assign new_n9239 = A837 & A838;
  assign new_n9240 = ~A837 & ~A838;
  assign new_n9241 = ~new_n9239 & ~new_n9240;
  assign new_n9242 = ~new_n9238 & new_n9241;
  assign new_n9243 = ~new_n9236 & ~new_n9239;
  assign new_n9244 = A838 & new_n9236;
  assign new_n9245 = ~new_n9243 & ~new_n9244;
  assign new_n9246 = ~new_n9242 & ~new_n9245;
  assign new_n9247 = new_n9237 & new_n9246;
  assign new_n9248 = new_n9236 & new_n9247;
  assign new_n9249 = A839 & A840;
  assign new_n9250 = ~new_n9246 & new_n9249;
  assign new_n9251 = ~new_n9248 & ~new_n9250;
  assign new_n9252 = ~new_n9237 & ~new_n9238;
  assign new_n9253 = ~new_n9240 & new_n9252;
  assign new_n9254 = ~new_n9243 & new_n9253;
  assign new_n9255 = new_n9251 & ~new_n9254;
  assign new_n9256 = ~new_n9235 & new_n9255;
  assign new_n9257 = ~new_n9249 & new_n9254;
  assign new_n9258 = new_n9238 & new_n9240;
  assign new_n9259 = ~new_n9249 & new_n9258;
  assign new_n9260 = ~new_n9247 & ~new_n9259;
  assign new_n9261 = ~new_n9257 & new_n9260;
  assign new_n9262 = new_n9251 & new_n9261;
  assign new_n9263 = ~new_n9233 & new_n9262;
  assign new_n9264 = new_n9233 & ~new_n9262;
  assign new_n9265 = ~new_n9263 & ~new_n9264;
  assign new_n9266 = new_n9228 & new_n9230;
  assign new_n9267 = ~new_n9231 & ~new_n9266;
  assign new_n9268 = ~new_n9237 & ~new_n9249;
  assign new_n9269 = new_n9241 & ~new_n9268;
  assign new_n9270 = ~new_n9241 & new_n9268;
  assign new_n9271 = ~new_n9269 & ~new_n9270;
  assign new_n9272 = ~new_n9236 & ~new_n9238;
  assign new_n9273 = ~new_n9271 & new_n9272;
  assign new_n9274 = new_n9271 & ~new_n9272;
  assign new_n9275 = ~new_n9273 & ~new_n9274;
  assign new_n9276 = new_n9267 & ~new_n9275;
  assign new_n9277 = ~new_n9266 & ~new_n9276;
  assign new_n9278 = ~new_n9265 & ~new_n9277;
  assign new_n9279 = ~new_n9234 & ~new_n9263;
  assign new_n9280 = ~new_n9278 & ~new_n9279;
  assign new_n9281 = new_n9235 & ~new_n9255;
  assign new_n9282 = ~new_n9256 & ~new_n9281;
  assign new_n9283 = ~new_n9280 & new_n9282;
  assign new_n9284 = ~new_n9256 & ~new_n9283;
  assign new_n9285 = new_n9215 & new_n9284;
  assign new_n9286 = ~new_n9215 & ~new_n9284;
  assign new_n9287 = ~new_n9285 & ~new_n9286;
  assign new_n9288 = new_n9265 & new_n9277;
  assign new_n9289 = ~new_n9278 & ~new_n9288;
  assign new_n9290 = new_n9207 & ~new_n9209;
  assign new_n9291 = ~new_n9210 & ~new_n9290;
  assign new_n9292 = ~new_n9289 & ~new_n9291;
  assign new_n9293 = ~new_n9267 & new_n9275;
  assign new_n9294 = ~new_n9276 & ~new_n9293;
  assign new_n9295 = ~new_n9200 & ~new_n9206;
  assign new_n9296 = ~new_n9207 & ~new_n9295;
  assign new_n9297 = ~new_n9294 & new_n9296;
  assign new_n9298 = ~new_n9209 & new_n9289;
  assign new_n9299 = new_n9297 & ~new_n9298;
  assign new_n9300 = ~new_n9292 & ~new_n9299;
  assign new_n9301 = new_n9211 & ~new_n9213;
  assign new_n9302 = ~new_n9214 & ~new_n9301;
  assign new_n9303 = ~new_n9300 & ~new_n9302;
  assign new_n9304 = new_n9280 & ~new_n9282;
  assign new_n9305 = ~new_n9283 & ~new_n9304;
  assign new_n9306 = new_n9300 & new_n9302;
  assign new_n9307 = ~new_n9303 & ~new_n9306;
  assign new_n9308 = ~new_n9305 & new_n9307;
  assign new_n9309 = ~new_n9303 & ~new_n9308;
  assign new_n9310 = new_n9287 & ~new_n9309;
  assign new_n9311 = ~new_n9285 & ~new_n9310;
  assign new_n9312 = A801 & A804;
  assign new_n9313 = A799 & A800;
  assign new_n9314 = A802 & A803;
  assign new_n9315 = ~new_n9313 & ~new_n9314;
  assign new_n9316 = new_n9312 & ~new_n9315;
  assign new_n9317 = ~A799 & ~A800;
  assign new_n9318 = ~A801 & A804;
  assign new_n9319 = new_n9314 & new_n9318;
  assign new_n9320 = ~A801 & ~new_n9313;
  assign new_n9321 = ~A802 & ~A803;
  assign new_n9322 = ~new_n9314 & ~new_n9321;
  assign new_n9323 = A804 & ~new_n9322;
  assign new_n9324 = ~A804 & ~new_n9314;
  assign new_n9325 = ~new_n9320 & ~new_n9324;
  assign new_n9326 = ~new_n9323 & new_n9325;
  assign new_n9327 = ~new_n9319 & ~new_n9326;
  assign new_n9328 = ~new_n9317 & ~new_n9327;
  assign new_n9329 = A803 & new_n9313;
  assign new_n9330 = new_n9316 & ~new_n9329;
  assign new_n9331 = A801 & ~A804;
  assign new_n9332 = new_n9313 & ~new_n9321;
  assign new_n9333 = new_n9331 & new_n9332;
  assign new_n9334 = ~new_n9312 & new_n9317;
  assign new_n9335 = new_n9321 & new_n9334;
  assign new_n9336 = ~new_n9333 & ~new_n9335;
  assign new_n9337 = ~new_n9330 & new_n9336;
  assign new_n9338 = ~new_n9328 & new_n9337;
  assign new_n9339 = ~new_n9317 & ~new_n9338;
  assign new_n9340 = ~new_n9316 & ~new_n9339;
  assign new_n9341 = ~A806 & ~A807;
  assign new_n9342 = A806 & A807;
  assign new_n9343 = ~new_n9341 & ~new_n9342;
  assign new_n9344 = ~A805 & new_n9343;
  assign new_n9345 = ~new_n9341 & ~new_n9344;
  assign new_n9346 = ~A808 & ~A809;
  assign new_n9347 = new_n9345 & ~new_n9346;
  assign new_n9348 = A808 & A809;
  assign new_n9349 = ~A810 & ~new_n9348;
  assign new_n9350 = new_n9347 & ~new_n9349;
  assign new_n9351 = ~A810 & ~new_n9347;
  assign new_n9352 = A805 & ~new_n9343;
  assign new_n9353 = ~new_n9344 & ~new_n9352;
  assign new_n9354 = ~new_n9345 & ~new_n9348;
  assign new_n9355 = new_n9345 & new_n9348;
  assign new_n9356 = ~new_n9354 & ~new_n9355;
  assign new_n9357 = A810 & ~new_n9356;
  assign new_n9358 = ~new_n9351 & ~new_n9353;
  assign new_n9359 = ~new_n9357 & new_n9358;
  assign new_n9360 = ~new_n9350 & ~new_n9359;
  assign new_n9361 = new_n9340 & new_n9360;
  assign new_n9362 = ~new_n9313 & ~new_n9317;
  assign new_n9363 = ~new_n9318 & ~new_n9331;
  assign new_n9364 = new_n9362 & ~new_n9363;
  assign new_n9365 = ~new_n9362 & new_n9363;
  assign new_n9366 = ~new_n9364 & ~new_n9365;
  assign new_n9367 = new_n9322 & new_n9366;
  assign new_n9368 = new_n9320 & new_n9324;
  assign new_n9369 = ~new_n9367 & new_n9368;
  assign new_n9370 = new_n9338 & ~new_n9369;
  assign new_n9371 = A810 & ~new_n9353;
  assign new_n9372 = ~new_n9345 & new_n9346;
  assign new_n9373 = ~new_n9371 & new_n9372;
  assign new_n9374 = ~new_n9345 & new_n9349;
  assign new_n9375 = ~new_n9350 & ~new_n9374;
  assign new_n9376 = new_n9353 & ~new_n9375;
  assign new_n9377 = ~new_n9359 & ~new_n9373;
  assign new_n9378 = ~new_n9376 & new_n9377;
  assign new_n9379 = ~new_n9370 & ~new_n9378;
  assign new_n9380 = ~new_n9322 & ~new_n9366;
  assign new_n9381 = ~new_n9367 & ~new_n9380;
  assign new_n9382 = ~A810 & new_n9353;
  assign new_n9383 = ~new_n9371 & ~new_n9382;
  assign new_n9384 = ~new_n9346 & ~new_n9348;
  assign new_n9385 = ~new_n9383 & new_n9384;
  assign new_n9386 = new_n9383 & ~new_n9384;
  assign new_n9387 = ~new_n9385 & ~new_n9386;
  assign new_n9388 = new_n9381 & ~new_n9387;
  assign new_n9389 = new_n9370 & new_n9378;
  assign new_n9390 = ~new_n9379 & ~new_n9389;
  assign new_n9391 = ~new_n9388 & new_n9390;
  assign new_n9392 = ~new_n9379 & ~new_n9391;
  assign new_n9393 = ~new_n9340 & ~new_n9360;
  assign new_n9394 = ~new_n9361 & ~new_n9393;
  assign new_n9395 = ~new_n9392 & new_n9394;
  assign new_n9396 = ~new_n9361 & ~new_n9395;
  assign new_n9397 = ~A818 & ~A819;
  assign new_n9398 = A818 & A819;
  assign new_n9399 = ~new_n9397 & ~new_n9398;
  assign new_n9400 = ~A817 & new_n9399;
  assign new_n9401 = ~new_n9397 & ~new_n9400;
  assign new_n9402 = ~A821 & ~A822;
  assign new_n9403 = A821 & A822;
  assign new_n9404 = ~new_n9402 & ~new_n9403;
  assign new_n9405 = ~A820 & new_n9404;
  assign new_n9406 = ~new_n9402 & ~new_n9405;
  assign new_n9407 = ~new_n9401 & ~new_n9406;
  assign new_n9408 = A820 & ~new_n9404;
  assign new_n9409 = ~new_n9405 & ~new_n9408;
  assign new_n9410 = A817 & ~new_n9399;
  assign new_n9411 = ~new_n9400 & ~new_n9410;
  assign new_n9412 = ~new_n9409 & ~new_n9411;
  assign new_n9413 = new_n9401 & new_n9406;
  assign new_n9414 = ~new_n9407 & ~new_n9413;
  assign new_n9415 = ~new_n9412 & new_n9414;
  assign new_n9416 = ~new_n9407 & ~new_n9415;
  assign new_n9417 = A811 & A812;
  assign new_n9418 = ~A815 & ~A816;
  assign new_n9419 = A813 & A814;
  assign new_n9420 = ~new_n9417 & new_n9419;
  assign new_n9421 = ~A813 & ~A814;
  assign new_n9422 = ~new_n9419 & ~new_n9421;
  assign new_n9423 = ~A811 & ~A812;
  assign new_n9424 = ~new_n9417 & ~new_n9423;
  assign new_n9425 = ~new_n9422 & new_n9424;
  assign new_n9426 = ~new_n9419 & ~new_n9423;
  assign new_n9427 = ~new_n9425 & new_n9426;
  assign new_n9428 = ~new_n9420 & ~new_n9427;
  assign new_n9429 = new_n9418 & new_n9428;
  assign new_n9430 = new_n9417 & new_n9429;
  assign new_n9431 = A815 & A816;
  assign new_n9432 = ~new_n9428 & new_n9431;
  assign new_n9433 = ~new_n9430 & ~new_n9432;
  assign new_n9434 = ~new_n9417 & ~new_n9425;
  assign new_n9435 = ~new_n9418 & ~new_n9421;
  assign new_n9436 = ~new_n9434 & new_n9435;
  assign new_n9437 = new_n9433 & ~new_n9436;
  assign new_n9438 = ~new_n9416 & new_n9437;
  assign new_n9439 = new_n9409 & new_n9411;
  assign new_n9440 = ~new_n9412 & ~new_n9439;
  assign new_n9441 = ~new_n9418 & ~new_n9431;
  assign new_n9442 = new_n9422 & ~new_n9424;
  assign new_n9443 = ~new_n9425 & ~new_n9442;
  assign new_n9444 = new_n9441 & ~new_n9443;
  assign new_n9445 = ~new_n9441 & new_n9443;
  assign new_n9446 = ~new_n9444 & ~new_n9445;
  assign new_n9447 = new_n9440 & ~new_n9446;
  assign new_n9448 = ~new_n9439 & ~new_n9447;
  assign new_n9449 = ~new_n9414 & new_n9448;
  assign new_n9450 = new_n9414 & ~new_n9448;
  assign new_n9451 = ~new_n9449 & ~new_n9450;
  assign new_n9452 = ~new_n9431 & new_n9436;
  assign new_n9453 = new_n9421 & new_n9423;
  assign new_n9454 = ~new_n9431 & new_n9453;
  assign new_n9455 = ~new_n9429 & ~new_n9454;
  assign new_n9456 = ~new_n9452 & new_n9455;
  assign new_n9457 = new_n9433 & new_n9456;
  assign new_n9458 = ~new_n9451 & ~new_n9457;
  assign new_n9459 = ~new_n9415 & ~new_n9449;
  assign new_n9460 = ~new_n9458 & ~new_n9459;
  assign new_n9461 = new_n9416 & ~new_n9437;
  assign new_n9462 = ~new_n9438 & ~new_n9461;
  assign new_n9463 = ~new_n9460 & new_n9462;
  assign new_n9464 = ~new_n9438 & ~new_n9463;
  assign new_n9465 = new_n9396 & new_n9464;
  assign new_n9466 = new_n9392 & ~new_n9394;
  assign new_n9467 = ~new_n9395 & ~new_n9466;
  assign new_n9468 = ~new_n9381 & new_n9387;
  assign new_n9469 = ~new_n9388 & ~new_n9468;
  assign new_n9470 = ~new_n9440 & new_n9446;
  assign new_n9471 = ~new_n9447 & ~new_n9470;
  assign new_n9472 = new_n9469 & ~new_n9471;
  assign new_n9473 = new_n9390 & new_n9472;
  assign new_n9474 = new_n9451 & new_n9457;
  assign new_n9475 = ~new_n9458 & ~new_n9474;
  assign new_n9476 = ~new_n9388 & ~new_n9472;
  assign new_n9477 = new_n9390 & ~new_n9476;
  assign new_n9478 = ~new_n9390 & new_n9476;
  assign new_n9479 = ~new_n9477 & ~new_n9478;
  assign new_n9480 = ~new_n9475 & new_n9479;
  assign new_n9481 = ~new_n9473 & ~new_n9480;
  assign new_n9482 = ~new_n9467 & ~new_n9481;
  assign new_n9483 = new_n9460 & ~new_n9462;
  assign new_n9484 = ~new_n9463 & ~new_n9483;
  assign new_n9485 = new_n9467 & new_n9481;
  assign new_n9486 = ~new_n9482 & ~new_n9485;
  assign new_n9487 = ~new_n9484 & new_n9486;
  assign new_n9488 = ~new_n9482 & ~new_n9487;
  assign new_n9489 = ~new_n9396 & ~new_n9464;
  assign new_n9490 = ~new_n9465 & ~new_n9489;
  assign new_n9491 = ~new_n9488 & new_n9490;
  assign new_n9492 = ~new_n9465 & ~new_n9491;
  assign new_n9493 = ~new_n9311 & ~new_n9492;
  assign new_n9494 = new_n9311 & new_n9492;
  assign new_n9495 = ~new_n9493 & ~new_n9494;
  assign new_n9496 = new_n9488 & ~new_n9490;
  assign new_n9497 = ~new_n9491 & ~new_n9496;
  assign new_n9498 = new_n9305 & ~new_n9307;
  assign new_n9499 = ~new_n9308 & ~new_n9498;
  assign new_n9500 = ~new_n9469 & new_n9471;
  assign new_n9501 = ~new_n9472 & ~new_n9500;
  assign new_n9502 = new_n9294 & ~new_n9296;
  assign new_n9503 = ~new_n9297 & ~new_n9502;
  assign new_n9504 = new_n9501 & new_n9503;
  assign new_n9505 = ~new_n9207 & ~new_n9297;
  assign new_n9506 = new_n9209 & ~new_n9289;
  assign new_n9507 = ~new_n9298 & ~new_n9506;
  assign new_n9508 = new_n9505 & ~new_n9507;
  assign new_n9509 = ~new_n9505 & new_n9507;
  assign new_n9510 = ~new_n9508 & ~new_n9509;
  assign new_n9511 = new_n9504 & new_n9510;
  assign new_n9512 = new_n9475 & ~new_n9479;
  assign new_n9513 = ~new_n9480 & ~new_n9512;
  assign new_n9514 = ~new_n9504 & ~new_n9510;
  assign new_n9515 = ~new_n9511 & ~new_n9514;
  assign new_n9516 = new_n9513 & new_n9515;
  assign new_n9517 = ~new_n9511 & ~new_n9516;
  assign new_n9518 = ~new_n9499 & new_n9517;
  assign new_n9519 = new_n9484 & ~new_n9486;
  assign new_n9520 = ~new_n9487 & ~new_n9519;
  assign new_n9521 = new_n9499 & ~new_n9517;
  assign new_n9522 = ~new_n9518 & ~new_n9521;
  assign new_n9523 = ~new_n9520 & new_n9522;
  assign new_n9524 = ~new_n9518 & ~new_n9523;
  assign new_n9525 = ~new_n9497 & ~new_n9524;
  assign new_n9526 = ~new_n9287 & new_n9309;
  assign new_n9527 = ~new_n9310 & ~new_n9526;
  assign new_n9528 = new_n9497 & new_n9524;
  assign new_n9529 = ~new_n9525 & ~new_n9528;
  assign new_n9530 = ~new_n9527 & new_n9529;
  assign new_n9531 = ~new_n9525 & ~new_n9530;
  assign new_n9532 = new_n9495 & new_n9531;
  assign new_n9533 = ~new_n9493 & ~new_n9532;
  assign new_n9534 = new_n9138 & ~new_n9533;
  assign new_n9535 = ~new_n9495 & ~new_n9531;
  assign new_n9536 = ~new_n9532 & ~new_n9535;
  assign new_n9537 = new_n9527 & ~new_n9529;
  assign new_n9538 = ~new_n9530 & ~new_n9537;
  assign new_n9539 = new_n9520 & ~new_n9522;
  assign new_n9540 = ~new_n9523 & ~new_n9539;
  assign new_n9541 = ~new_n9513 & ~new_n9515;
  assign new_n9542 = ~new_n9516 & ~new_n9541;
  assign new_n9543 = ~new_n9114 & ~new_n9115;
  assign new_n9544 = ~new_n9501 & ~new_n9503;
  assign new_n9545 = ~new_n9504 & ~new_n9544;
  assign new_n9546 = ~new_n9117 & ~new_n9119;
  assign new_n9547 = ~new_n9120 & ~new_n9546;
  assign new_n9548 = new_n9545 & new_n9547;
  assign new_n9549 = ~new_n9120 & ~new_n9548;
  assign new_n9550 = new_n9543 & ~new_n9549;
  assign new_n9551 = ~new_n9543 & new_n9549;
  assign new_n9552 = ~new_n9550 & ~new_n9551;
  assign new_n9553 = ~new_n9542 & new_n9552;
  assign new_n9554 = ~new_n9548 & ~new_n9552;
  assign new_n9555 = ~new_n9553 & ~new_n9554;
  assign new_n9556 = ~new_n9540 & new_n9555;
  assign new_n9557 = new_n9125 & ~new_n9127;
  assign new_n9558 = ~new_n9128 & ~new_n9557;
  assign new_n9559 = new_n9540 & ~new_n9555;
  assign new_n9560 = ~new_n9556 & ~new_n9559;
  assign new_n9561 = ~new_n9558 & new_n9560;
  assign new_n9562 = ~new_n9556 & ~new_n9561;
  assign new_n9563 = new_n9538 & new_n9562;
  assign new_n9564 = new_n9132 & ~new_n9134;
  assign new_n9565 = ~new_n9135 & ~new_n9564;
  assign new_n9566 = ~new_n9538 & ~new_n9562;
  assign new_n9567 = ~new_n9563 & ~new_n9566;
  assign new_n9568 = new_n9565 & new_n9567;
  assign new_n9569 = ~new_n9563 & ~new_n9568;
  assign new_n9570 = new_n9536 & new_n9569;
  assign new_n9571 = ~new_n9107 & new_n9136;
  assign new_n9572 = ~new_n9137 & ~new_n9571;
  assign new_n9573 = ~new_n9536 & ~new_n9569;
  assign new_n9574 = ~new_n9570 & ~new_n9573;
  assign new_n9575 = ~new_n9572 & new_n9574;
  assign new_n9576 = ~new_n9570 & ~new_n9575;
  assign new_n9577 = ~new_n9138 & new_n9533;
  assign new_n9578 = ~new_n9534 & ~new_n9577;
  assign new_n9579 = ~new_n9576 & new_n9578;
  assign new_n9580 = ~new_n9534 & ~new_n9579;
  assign new_n9581 = A691 & A692;
  assign new_n9582 = A694 & A695;
  assign new_n9583 = ~new_n9581 & ~new_n9582;
  assign new_n9584 = A693 & A696;
  assign new_n9585 = ~new_n9583 & new_n9584;
  assign new_n9586 = ~A691 & ~A692;
  assign new_n9587 = ~A693 & A696;
  assign new_n9588 = new_n9582 & new_n9587;
  assign new_n9589 = ~A693 & ~new_n9581;
  assign new_n9590 = ~A694 & ~A695;
  assign new_n9591 = ~new_n9582 & ~new_n9590;
  assign new_n9592 = A696 & ~new_n9591;
  assign new_n9593 = ~A696 & ~new_n9582;
  assign new_n9594 = ~new_n9589 & ~new_n9593;
  assign new_n9595 = ~new_n9592 & new_n9594;
  assign new_n9596 = ~new_n9588 & ~new_n9595;
  assign new_n9597 = ~new_n9586 & ~new_n9596;
  assign new_n9598 = A695 & new_n9581;
  assign new_n9599 = new_n9585 & ~new_n9598;
  assign new_n9600 = ~new_n9584 & new_n9586;
  assign new_n9601 = new_n9590 & new_n9600;
  assign new_n9602 = A693 & ~A696;
  assign new_n9603 = new_n9581 & ~new_n9590;
  assign new_n9604 = new_n9602 & new_n9603;
  assign new_n9605 = ~new_n9601 & ~new_n9604;
  assign new_n9606 = ~new_n9599 & new_n9605;
  assign new_n9607 = ~new_n9597 & new_n9606;
  assign new_n9608 = ~new_n9586 & ~new_n9607;
  assign new_n9609 = ~new_n9585 & ~new_n9608;
  assign new_n9610 = ~A701 & ~A702;
  assign new_n9611 = A701 & A702;
  assign new_n9612 = ~new_n9610 & ~new_n9611;
  assign new_n9613 = ~A700 & new_n9612;
  assign new_n9614 = ~new_n9610 & ~new_n9613;
  assign new_n9615 = ~A698 & ~A699;
  assign new_n9616 = A698 & A699;
  assign new_n9617 = ~new_n9615 & ~new_n9616;
  assign new_n9618 = ~A697 & new_n9617;
  assign new_n9619 = ~new_n9615 & ~new_n9618;
  assign new_n9620 = ~new_n9614 & ~new_n9619;
  assign new_n9621 = A697 & ~new_n9617;
  assign new_n9622 = ~new_n9618 & ~new_n9621;
  assign new_n9623 = A700 & ~new_n9612;
  assign new_n9624 = ~new_n9613 & ~new_n9623;
  assign new_n9625 = ~new_n9622 & ~new_n9624;
  assign new_n9626 = new_n9614 & new_n9619;
  assign new_n9627 = ~new_n9620 & ~new_n9626;
  assign new_n9628 = ~new_n9625 & new_n9627;
  assign new_n9629 = ~new_n9620 & ~new_n9628;
  assign new_n9630 = new_n9609 & ~new_n9629;
  assign new_n9631 = ~new_n9581 & ~new_n9586;
  assign new_n9632 = ~new_n9587 & ~new_n9602;
  assign new_n9633 = new_n9631 & ~new_n9632;
  assign new_n9634 = ~new_n9631 & new_n9632;
  assign new_n9635 = ~new_n9633 & ~new_n9634;
  assign new_n9636 = new_n9591 & new_n9635;
  assign new_n9637 = new_n9589 & new_n9593;
  assign new_n9638 = ~new_n9636 & new_n9637;
  assign new_n9639 = new_n9607 & ~new_n9638;
  assign new_n9640 = ~new_n9627 & new_n9639;
  assign new_n9641 = new_n9627 & ~new_n9639;
  assign new_n9642 = ~new_n9640 & ~new_n9641;
  assign new_n9643 = new_n9622 & new_n9624;
  assign new_n9644 = ~new_n9591 & ~new_n9635;
  assign new_n9645 = ~new_n9636 & ~new_n9644;
  assign new_n9646 = ~new_n9625 & ~new_n9643;
  assign new_n9647 = ~new_n9645 & new_n9646;
  assign new_n9648 = ~new_n9643 & ~new_n9647;
  assign new_n9649 = ~new_n9642 & ~new_n9648;
  assign new_n9650 = ~new_n9628 & ~new_n9640;
  assign new_n9651 = ~new_n9649 & ~new_n9650;
  assign new_n9652 = ~new_n9609 & new_n9629;
  assign new_n9653 = ~new_n9630 & ~new_n9652;
  assign new_n9654 = ~new_n9651 & new_n9653;
  assign new_n9655 = ~new_n9630 & ~new_n9654;
  assign new_n9656 = A685 & A686;
  assign new_n9657 = A688 & A689;
  assign new_n9658 = ~new_n9656 & ~new_n9657;
  assign new_n9659 = A687 & A690;
  assign new_n9660 = ~new_n9658 & new_n9659;
  assign new_n9661 = ~A685 & ~A686;
  assign new_n9662 = ~A687 & A690;
  assign new_n9663 = new_n9657 & new_n9662;
  assign new_n9664 = ~A687 & ~new_n9656;
  assign new_n9665 = ~A688 & ~A689;
  assign new_n9666 = ~new_n9657 & ~new_n9665;
  assign new_n9667 = A690 & ~new_n9666;
  assign new_n9668 = ~A690 & ~new_n9657;
  assign new_n9669 = ~new_n9664 & ~new_n9668;
  assign new_n9670 = ~new_n9667 & new_n9669;
  assign new_n9671 = ~new_n9663 & ~new_n9670;
  assign new_n9672 = ~new_n9661 & ~new_n9671;
  assign new_n9673 = A689 & new_n9656;
  assign new_n9674 = new_n9660 & ~new_n9673;
  assign new_n9675 = ~new_n9659 & new_n9661;
  assign new_n9676 = new_n9665 & new_n9675;
  assign new_n9677 = A687 & ~A690;
  assign new_n9678 = new_n9656 & ~new_n9665;
  assign new_n9679 = new_n9677 & new_n9678;
  assign new_n9680 = ~new_n9676 & ~new_n9679;
  assign new_n9681 = ~new_n9674 & new_n9680;
  assign new_n9682 = ~new_n9672 & new_n9681;
  assign new_n9683 = ~new_n9661 & ~new_n9682;
  assign new_n9684 = ~new_n9660 & ~new_n9683;
  assign new_n9685 = A679 & A680;
  assign new_n9686 = A682 & A683;
  assign new_n9687 = ~new_n9685 & ~new_n9686;
  assign new_n9688 = A681 & A684;
  assign new_n9689 = ~new_n9687 & new_n9688;
  assign new_n9690 = ~A679 & ~A680;
  assign new_n9691 = ~A681 & A684;
  assign new_n9692 = new_n9686 & new_n9691;
  assign new_n9693 = ~A681 & ~new_n9685;
  assign new_n9694 = ~A682 & ~A683;
  assign new_n9695 = ~new_n9686 & ~new_n9694;
  assign new_n9696 = A684 & ~new_n9695;
  assign new_n9697 = ~A684 & ~new_n9686;
  assign new_n9698 = ~new_n9693 & ~new_n9697;
  assign new_n9699 = ~new_n9696 & new_n9698;
  assign new_n9700 = ~new_n9692 & ~new_n9699;
  assign new_n9701 = ~new_n9690 & ~new_n9700;
  assign new_n9702 = A683 & new_n9685;
  assign new_n9703 = new_n9689 & ~new_n9702;
  assign new_n9704 = ~new_n9688 & new_n9690;
  assign new_n9705 = new_n9694 & new_n9704;
  assign new_n9706 = A681 & ~A684;
  assign new_n9707 = new_n9685 & ~new_n9694;
  assign new_n9708 = new_n9706 & new_n9707;
  assign new_n9709 = ~new_n9705 & ~new_n9708;
  assign new_n9710 = ~new_n9703 & new_n9709;
  assign new_n9711 = ~new_n9701 & new_n9710;
  assign new_n9712 = ~new_n9690 & ~new_n9711;
  assign new_n9713 = ~new_n9689 & ~new_n9712;
  assign new_n9714 = ~new_n9684 & ~new_n9713;
  assign new_n9715 = new_n9684 & new_n9713;
  assign new_n9716 = ~new_n9714 & ~new_n9715;
  assign new_n9717 = ~new_n9685 & ~new_n9690;
  assign new_n9718 = ~new_n9691 & ~new_n9706;
  assign new_n9719 = new_n9717 & ~new_n9718;
  assign new_n9720 = ~new_n9717 & new_n9718;
  assign new_n9721 = ~new_n9719 & ~new_n9720;
  assign new_n9722 = new_n9695 & new_n9721;
  assign new_n9723 = new_n9693 & new_n9697;
  assign new_n9724 = ~new_n9722 & new_n9723;
  assign new_n9725 = new_n9711 & ~new_n9724;
  assign new_n9726 = ~new_n9656 & ~new_n9661;
  assign new_n9727 = ~new_n9662 & ~new_n9677;
  assign new_n9728 = new_n9726 & ~new_n9727;
  assign new_n9729 = ~new_n9726 & new_n9727;
  assign new_n9730 = ~new_n9728 & ~new_n9729;
  assign new_n9731 = new_n9666 & new_n9730;
  assign new_n9732 = new_n9664 & new_n9668;
  assign new_n9733 = ~new_n9731 & new_n9732;
  assign new_n9734 = new_n9682 & ~new_n9733;
  assign new_n9735 = new_n9725 & new_n9734;
  assign new_n9736 = ~new_n9695 & ~new_n9721;
  assign new_n9737 = ~new_n9722 & ~new_n9736;
  assign new_n9738 = ~new_n9666 & ~new_n9730;
  assign new_n9739 = ~new_n9731 & ~new_n9738;
  assign new_n9740 = new_n9737 & new_n9739;
  assign new_n9741 = ~new_n9725 & ~new_n9734;
  assign new_n9742 = ~new_n9735 & ~new_n9741;
  assign new_n9743 = new_n9740 & new_n9742;
  assign new_n9744 = ~new_n9735 & ~new_n9743;
  assign new_n9745 = new_n9716 & ~new_n9744;
  assign new_n9746 = ~new_n9714 & ~new_n9745;
  assign new_n9747 = ~new_n9655 & new_n9746;
  assign new_n9748 = new_n9655 & ~new_n9746;
  assign new_n9749 = ~new_n9747 & ~new_n9748;
  assign new_n9750 = new_n9651 & ~new_n9653;
  assign new_n9751 = ~new_n9654 & ~new_n9750;
  assign new_n9752 = ~new_n9716 & new_n9744;
  assign new_n9753 = ~new_n9745 & ~new_n9752;
  assign new_n9754 = new_n9751 & ~new_n9753;
  assign new_n9755 = ~new_n9751 & new_n9753;
  assign new_n9756 = ~new_n9754 & ~new_n9755;
  assign new_n9757 = new_n9642 & new_n9648;
  assign new_n9758 = ~new_n9649 & ~new_n9757;
  assign new_n9759 = new_n9742 & ~new_n9758;
  assign new_n9760 = new_n9645 & ~new_n9646;
  assign new_n9761 = ~new_n9647 & ~new_n9760;
  assign new_n9762 = ~new_n9737 & ~new_n9739;
  assign new_n9763 = ~new_n9740 & ~new_n9762;
  assign new_n9764 = ~new_n9761 & new_n9763;
  assign new_n9765 = ~new_n9740 & ~new_n9764;
  assign new_n9766 = ~new_n9742 & new_n9758;
  assign new_n9767 = ~new_n9759 & ~new_n9766;
  assign new_n9768 = ~new_n9765 & new_n9767;
  assign new_n9769 = ~new_n9759 & ~new_n9768;
  assign new_n9770 = ~new_n9743 & ~new_n9769;
  assign new_n9771 = new_n9756 & ~new_n9770;
  assign new_n9772 = ~new_n9754 & ~new_n9771;
  assign new_n9773 = new_n9749 & ~new_n9772;
  assign new_n9774 = ~new_n9747 & ~new_n9773;
  assign new_n9775 = ~A661 & ~A662;
  assign new_n9776 = A661 & A662;
  assign new_n9777 = ~A663 & ~new_n9776;
  assign new_n9778 = ~new_n9775 & ~new_n9777;
  assign new_n9779 = A665 & A666;
  assign new_n9780 = new_n9778 & new_n9779;
  assign new_n9781 = A663 & new_n9776;
  assign new_n9782 = ~A664 & ~new_n9781;
  assign new_n9783 = new_n9778 & ~new_n9782;
  assign new_n9784 = A665 & new_n9783;
  assign new_n9785 = A663 & A664;
  assign new_n9786 = new_n9776 & new_n9785;
  assign new_n9787 = ~new_n9784 & ~new_n9786;
  assign new_n9788 = ~A666 & ~new_n9787;
  assign new_n9789 = ~A665 & ~A666;
  assign new_n9790 = ~new_n9775 & ~new_n9789;
  assign new_n9791 = new_n9777 & ~new_n9779;
  assign new_n9792 = ~new_n9790 & new_n9791;
  assign new_n9793 = ~new_n9780 & ~new_n9792;
  assign new_n9794 = ~A664 & ~new_n9793;
  assign new_n9795 = ~A665 & A666;
  assign new_n9796 = new_n9783 & new_n9795;
  assign new_n9797 = new_n9775 & ~new_n9785;
  assign new_n9798 = A664 & new_n9779;
  assign new_n9799 = ~new_n9781 & new_n9798;
  assign new_n9800 = ~new_n9797 & new_n9799;
  assign new_n9801 = ~new_n9796 & ~new_n9800;
  assign new_n9802 = ~new_n9794 & new_n9801;
  assign new_n9803 = ~new_n9788 & new_n9802;
  assign new_n9804 = ~new_n9782 & ~new_n9803;
  assign new_n9805 = ~new_n9780 & ~new_n9804;
  assign new_n9806 = A657 & A660;
  assign new_n9807 = A658 & A659;
  assign new_n9808 = A655 & A656;
  assign new_n9809 = ~new_n9807 & ~new_n9808;
  assign new_n9810 = new_n9806 & ~new_n9809;
  assign new_n9811 = ~A655 & ~A656;
  assign new_n9812 = ~A657 & A660;
  assign new_n9813 = new_n9807 & new_n9812;
  assign new_n9814 = ~A657 & ~new_n9808;
  assign new_n9815 = ~A658 & ~A659;
  assign new_n9816 = ~new_n9807 & ~new_n9815;
  assign new_n9817 = A660 & ~new_n9816;
  assign new_n9818 = ~A660 & ~new_n9807;
  assign new_n9819 = ~new_n9814 & ~new_n9818;
  assign new_n9820 = ~new_n9817 & new_n9819;
  assign new_n9821 = ~new_n9813 & ~new_n9820;
  assign new_n9822 = ~new_n9811 & ~new_n9821;
  assign new_n9823 = A659 & new_n9808;
  assign new_n9824 = new_n9810 & ~new_n9823;
  assign new_n9825 = ~new_n9806 & new_n9811;
  assign new_n9826 = new_n9815 & new_n9825;
  assign new_n9827 = A657 & ~A660;
  assign new_n9828 = new_n9808 & ~new_n9815;
  assign new_n9829 = new_n9827 & new_n9828;
  assign new_n9830 = ~new_n9826 & ~new_n9829;
  assign new_n9831 = ~new_n9824 & new_n9830;
  assign new_n9832 = ~new_n9822 & new_n9831;
  assign new_n9833 = ~new_n9811 & ~new_n9832;
  assign new_n9834 = ~new_n9810 & ~new_n9833;
  assign new_n9835 = new_n9805 & new_n9834;
  assign new_n9836 = ~new_n9808 & ~new_n9811;
  assign new_n9837 = ~new_n9812 & ~new_n9827;
  assign new_n9838 = new_n9836 & ~new_n9837;
  assign new_n9839 = ~new_n9836 & new_n9837;
  assign new_n9840 = ~new_n9838 & ~new_n9839;
  assign new_n9841 = new_n9816 & new_n9840;
  assign new_n9842 = ~new_n9816 & ~new_n9840;
  assign new_n9843 = ~new_n9841 & ~new_n9842;
  assign new_n9844 = A663 & ~A666;
  assign new_n9845 = ~A663 & A666;
  assign new_n9846 = ~new_n9844 & ~new_n9845;
  assign new_n9847 = ~new_n9775 & ~new_n9776;
  assign new_n9848 = ~A664 & ~A665;
  assign new_n9849 = A664 & A665;
  assign new_n9850 = ~new_n9848 & ~new_n9849;
  assign new_n9851 = new_n9847 & ~new_n9850;
  assign new_n9852 = ~new_n9847 & new_n9850;
  assign new_n9853 = ~new_n9851 & ~new_n9852;
  assign new_n9854 = new_n9846 & new_n9853;
  assign new_n9855 = ~new_n9846 & ~new_n9853;
  assign new_n9856 = ~new_n9854 & ~new_n9855;
  assign new_n9857 = new_n9843 & new_n9856;
  assign new_n9858 = new_n9814 & new_n9818;
  assign new_n9859 = ~new_n9841 & new_n9858;
  assign new_n9860 = new_n9832 & ~new_n9859;
  assign new_n9861 = ~new_n9857 & ~new_n9860;
  assign new_n9862 = new_n9789 & new_n9797;
  assign new_n9863 = new_n9803 & ~new_n9862;
  assign new_n9864 = new_n9857 & new_n9860;
  assign new_n9865 = ~new_n9861 & ~new_n9864;
  assign new_n9866 = ~new_n9863 & new_n9865;
  assign new_n9867 = ~new_n9861 & ~new_n9866;
  assign new_n9868 = ~new_n9805 & ~new_n9834;
  assign new_n9869 = ~new_n9835 & ~new_n9868;
  assign new_n9870 = ~new_n9867 & new_n9869;
  assign new_n9871 = ~new_n9835 & ~new_n9870;
  assign new_n9872 = A667 & A668;
  assign new_n9873 = A670 & A671;
  assign new_n9874 = ~new_n9872 & ~new_n9873;
  assign new_n9875 = A669 & A672;
  assign new_n9876 = ~new_n9874 & new_n9875;
  assign new_n9877 = ~A667 & ~A668;
  assign new_n9878 = ~A669 & A672;
  assign new_n9879 = new_n9873 & new_n9878;
  assign new_n9880 = ~A669 & ~new_n9872;
  assign new_n9881 = ~A670 & ~A671;
  assign new_n9882 = ~new_n9873 & ~new_n9881;
  assign new_n9883 = A672 & ~new_n9882;
  assign new_n9884 = ~A672 & ~new_n9873;
  assign new_n9885 = ~new_n9880 & ~new_n9884;
  assign new_n9886 = ~new_n9883 & new_n9885;
  assign new_n9887 = ~new_n9879 & ~new_n9886;
  assign new_n9888 = ~new_n9877 & ~new_n9887;
  assign new_n9889 = A671 & new_n9872;
  assign new_n9890 = new_n9876 & ~new_n9889;
  assign new_n9891 = A669 & ~A672;
  assign new_n9892 = new_n9872 & ~new_n9881;
  assign new_n9893 = new_n9891 & new_n9892;
  assign new_n9894 = ~new_n9875 & new_n9877;
  assign new_n9895 = new_n9881 & new_n9894;
  assign new_n9896 = ~new_n9893 & ~new_n9895;
  assign new_n9897 = ~new_n9890 & new_n9896;
  assign new_n9898 = ~new_n9888 & new_n9897;
  assign new_n9899 = ~new_n9877 & ~new_n9898;
  assign new_n9900 = ~new_n9876 & ~new_n9899;
  assign new_n9901 = A673 & A674;
  assign new_n9902 = A676 & A677;
  assign new_n9903 = ~new_n9901 & ~new_n9902;
  assign new_n9904 = A675 & A678;
  assign new_n9905 = ~new_n9903 & new_n9904;
  assign new_n9906 = ~A673 & ~A674;
  assign new_n9907 = ~A675 & A678;
  assign new_n9908 = new_n9902 & new_n9907;
  assign new_n9909 = ~A675 & ~new_n9901;
  assign new_n9910 = ~A676 & ~A677;
  assign new_n9911 = ~new_n9902 & ~new_n9910;
  assign new_n9912 = A678 & ~new_n9911;
  assign new_n9913 = ~A678 & ~new_n9902;
  assign new_n9914 = ~new_n9909 & ~new_n9913;
  assign new_n9915 = ~new_n9912 & new_n9914;
  assign new_n9916 = ~new_n9908 & ~new_n9915;
  assign new_n9917 = ~new_n9906 & ~new_n9916;
  assign new_n9918 = A677 & new_n9901;
  assign new_n9919 = new_n9905 & ~new_n9918;
  assign new_n9920 = ~new_n9904 & new_n9906;
  assign new_n9921 = new_n9910 & new_n9920;
  assign new_n9922 = A675 & ~A678;
  assign new_n9923 = new_n9901 & ~new_n9910;
  assign new_n9924 = new_n9922 & new_n9923;
  assign new_n9925 = ~new_n9921 & ~new_n9924;
  assign new_n9926 = ~new_n9919 & new_n9925;
  assign new_n9927 = ~new_n9917 & new_n9926;
  assign new_n9928 = ~new_n9906 & ~new_n9927;
  assign new_n9929 = ~new_n9905 & ~new_n9928;
  assign new_n9930 = new_n9900 & new_n9929;
  assign new_n9931 = ~new_n9872 & ~new_n9877;
  assign new_n9932 = ~new_n9878 & ~new_n9891;
  assign new_n9933 = new_n9931 & ~new_n9932;
  assign new_n9934 = ~new_n9931 & new_n9932;
  assign new_n9935 = ~new_n9933 & ~new_n9934;
  assign new_n9936 = new_n9882 & new_n9935;
  assign new_n9937 = new_n9880 & new_n9884;
  assign new_n9938 = ~new_n9936 & new_n9937;
  assign new_n9939 = new_n9898 & ~new_n9938;
  assign new_n9940 = ~new_n9901 & ~new_n9906;
  assign new_n9941 = ~new_n9907 & ~new_n9922;
  assign new_n9942 = new_n9940 & ~new_n9941;
  assign new_n9943 = ~new_n9940 & new_n9941;
  assign new_n9944 = ~new_n9942 & ~new_n9943;
  assign new_n9945 = new_n9911 & new_n9944;
  assign new_n9946 = new_n9909 & new_n9913;
  assign new_n9947 = ~new_n9945 & new_n9946;
  assign new_n9948 = new_n9927 & ~new_n9947;
  assign new_n9949 = ~new_n9939 & ~new_n9948;
  assign new_n9950 = ~new_n9882 & ~new_n9935;
  assign new_n9951 = ~new_n9936 & ~new_n9950;
  assign new_n9952 = ~new_n9911 & ~new_n9944;
  assign new_n9953 = ~new_n9945 & ~new_n9952;
  assign new_n9954 = new_n9951 & new_n9953;
  assign new_n9955 = new_n9939 & new_n9948;
  assign new_n9956 = ~new_n9949 & ~new_n9955;
  assign new_n9957 = ~new_n9954 & new_n9956;
  assign new_n9958 = ~new_n9949 & ~new_n9957;
  assign new_n9959 = ~new_n9900 & ~new_n9929;
  assign new_n9960 = ~new_n9930 & ~new_n9959;
  assign new_n9961 = ~new_n9958 & new_n9960;
  assign new_n9962 = ~new_n9930 & ~new_n9961;
  assign new_n9963 = new_n9871 & new_n9962;
  assign new_n9964 = new_n9958 & ~new_n9960;
  assign new_n9965 = ~new_n9961 & ~new_n9964;
  assign new_n9966 = ~new_n9951 & ~new_n9953;
  assign new_n9967 = ~new_n9954 & ~new_n9966;
  assign new_n9968 = ~new_n9843 & ~new_n9856;
  assign new_n9969 = ~new_n9857 & ~new_n9968;
  assign new_n9970 = new_n9967 & new_n9969;
  assign new_n9971 = new_n9956 & new_n9970;
  assign new_n9972 = new_n9863 & ~new_n9865;
  assign new_n9973 = ~new_n9866 & ~new_n9972;
  assign new_n9974 = new_n9954 & ~new_n9956;
  assign new_n9975 = ~new_n9957 & ~new_n9970;
  assign new_n9976 = ~new_n9974 & new_n9975;
  assign new_n9977 = ~new_n9971 & ~new_n9976;
  assign new_n9978 = ~new_n9973 & new_n9977;
  assign new_n9979 = ~new_n9971 & ~new_n9978;
  assign new_n9980 = ~new_n9965 & ~new_n9979;
  assign new_n9981 = new_n9867 & ~new_n9869;
  assign new_n9982 = ~new_n9870 & ~new_n9981;
  assign new_n9983 = new_n9965 & new_n9979;
  assign new_n9984 = ~new_n9980 & ~new_n9983;
  assign new_n9985 = ~new_n9982 & new_n9984;
  assign new_n9986 = ~new_n9980 & ~new_n9985;
  assign new_n9987 = ~new_n9871 & ~new_n9962;
  assign new_n9988 = ~new_n9963 & ~new_n9987;
  assign new_n9989 = ~new_n9986 & new_n9988;
  assign new_n9990 = ~new_n9963 & ~new_n9989;
  assign new_n9991 = ~new_n9774 & new_n9990;
  assign new_n9992 = ~new_n9749 & new_n9772;
  assign new_n9993 = ~new_n9773 & ~new_n9992;
  assign new_n9994 = new_n9986 & ~new_n9988;
  assign new_n9995 = ~new_n9989 & ~new_n9994;
  assign new_n9996 = new_n9993 & ~new_n9995;
  assign new_n9997 = ~new_n9993 & new_n9995;
  assign new_n9998 = ~new_n9996 & ~new_n9997;
  assign new_n9999 = new_n9982 & ~new_n9984;
  assign new_n10000 = ~new_n9985 & ~new_n9999;
  assign new_n10001 = new_n9765 & ~new_n9767;
  assign new_n10002 = ~new_n9768 & ~new_n10001;
  assign new_n10003 = new_n9973 & ~new_n9977;
  assign new_n10004 = ~new_n9978 & ~new_n10003;
  assign new_n10005 = new_n10002 & new_n10004;
  assign new_n10006 = new_n9761 & ~new_n9763;
  assign new_n10007 = ~new_n9764 & ~new_n10006;
  assign new_n10008 = ~new_n9967 & ~new_n9969;
  assign new_n10009 = ~new_n9970 & ~new_n10008;
  assign new_n10010 = new_n10007 & new_n10009;
  assign new_n10011 = ~new_n10002 & ~new_n10004;
  assign new_n10012 = ~new_n10005 & ~new_n10011;
  assign new_n10013 = new_n10010 & new_n10012;
  assign new_n10014 = ~new_n10005 & ~new_n10013;
  assign new_n10015 = new_n10000 & ~new_n10014;
  assign new_n10016 = ~new_n9756 & new_n9770;
  assign new_n10017 = ~new_n9771 & ~new_n10016;
  assign new_n10018 = ~new_n10000 & new_n10014;
  assign new_n10019 = ~new_n10015 & ~new_n10018;
  assign new_n10020 = ~new_n10017 & new_n10019;
  assign new_n10021 = ~new_n10015 & ~new_n10020;
  assign new_n10022 = new_n9998 & new_n10021;
  assign new_n10023 = ~new_n9996 & ~new_n10022;
  assign new_n10024 = new_n9774 & ~new_n9990;
  assign new_n10025 = ~new_n9991 & ~new_n10024;
  assign new_n10026 = ~new_n10023 & new_n10025;
  assign new_n10027 = ~new_n9991 & ~new_n10026;
  assign new_n10028 = A723 & A726;
  assign new_n10029 = A724 & A725;
  assign new_n10030 = A721 & A722;
  assign new_n10031 = ~new_n10029 & ~new_n10030;
  assign new_n10032 = new_n10028 & ~new_n10031;
  assign new_n10033 = ~A721 & ~A722;
  assign new_n10034 = ~A723 & A726;
  assign new_n10035 = new_n10029 & new_n10034;
  assign new_n10036 = ~A723 & ~new_n10030;
  assign new_n10037 = ~A724 & ~A725;
  assign new_n10038 = ~new_n10029 & ~new_n10037;
  assign new_n10039 = A726 & ~new_n10038;
  assign new_n10040 = ~A726 & ~new_n10029;
  assign new_n10041 = ~new_n10036 & ~new_n10040;
  assign new_n10042 = ~new_n10039 & new_n10041;
  assign new_n10043 = ~new_n10035 & ~new_n10042;
  assign new_n10044 = ~new_n10033 & ~new_n10043;
  assign new_n10045 = A725 & new_n10030;
  assign new_n10046 = new_n10032 & ~new_n10045;
  assign new_n10047 = ~new_n10028 & new_n10033;
  assign new_n10048 = new_n10037 & new_n10047;
  assign new_n10049 = A723 & ~A726;
  assign new_n10050 = new_n10030 & ~new_n10037;
  assign new_n10051 = new_n10049 & new_n10050;
  assign new_n10052 = ~new_n10048 & ~new_n10051;
  assign new_n10053 = ~new_n10046 & new_n10052;
  assign new_n10054 = ~new_n10044 & new_n10053;
  assign new_n10055 = ~new_n10033 & ~new_n10054;
  assign new_n10056 = ~new_n10032 & ~new_n10055;
  assign new_n10057 = ~A718 & ~A719;
  assign new_n10058 = ~A716 & ~A717;
  assign new_n10059 = A716 & A717;
  assign new_n10060 = ~new_n10058 & ~new_n10059;
  assign new_n10061 = ~A715 & new_n10060;
  assign new_n10062 = ~new_n10058 & ~new_n10061;
  assign new_n10063 = ~new_n10057 & new_n10062;
  assign new_n10064 = A718 & A719;
  assign new_n10065 = ~A720 & ~new_n10064;
  assign new_n10066 = new_n10063 & ~new_n10065;
  assign new_n10067 = ~A720 & ~new_n10063;
  assign new_n10068 = A715 & ~new_n10060;
  assign new_n10069 = ~new_n10061 & ~new_n10068;
  assign new_n10070 = ~new_n10062 & ~new_n10064;
  assign new_n10071 = new_n10062 & new_n10064;
  assign new_n10072 = ~new_n10070 & ~new_n10071;
  assign new_n10073 = A720 & ~new_n10072;
  assign new_n10074 = ~new_n10067 & ~new_n10069;
  assign new_n10075 = ~new_n10073 & new_n10074;
  assign new_n10076 = ~new_n10066 & ~new_n10075;
  assign new_n10077 = ~new_n10056 & ~new_n10076;
  assign new_n10078 = new_n10056 & new_n10076;
  assign new_n10079 = ~new_n10077 & ~new_n10078;
  assign new_n10080 = ~new_n10030 & ~new_n10033;
  assign new_n10081 = ~new_n10034 & ~new_n10049;
  assign new_n10082 = new_n10080 & ~new_n10081;
  assign new_n10083 = ~new_n10080 & new_n10081;
  assign new_n10084 = ~new_n10082 & ~new_n10083;
  assign new_n10085 = new_n10038 & new_n10084;
  assign new_n10086 = new_n10036 & new_n10040;
  assign new_n10087 = ~new_n10085 & new_n10086;
  assign new_n10088 = new_n10054 & ~new_n10087;
  assign new_n10089 = A720 & ~new_n10069;
  assign new_n10090 = new_n10057 & ~new_n10062;
  assign new_n10091 = ~new_n10089 & new_n10090;
  assign new_n10092 = ~new_n10062 & new_n10065;
  assign new_n10093 = ~new_n10066 & ~new_n10092;
  assign new_n10094 = new_n10069 & ~new_n10093;
  assign new_n10095 = ~new_n10075 & ~new_n10091;
  assign new_n10096 = ~new_n10094 & new_n10095;
  assign new_n10097 = ~new_n10088 & ~new_n10096;
  assign new_n10098 = ~new_n10038 & ~new_n10084;
  assign new_n10099 = ~new_n10085 & ~new_n10098;
  assign new_n10100 = ~A720 & new_n10069;
  assign new_n10101 = ~new_n10089 & ~new_n10100;
  assign new_n10102 = ~new_n10057 & ~new_n10064;
  assign new_n10103 = ~new_n10101 & new_n10102;
  assign new_n10104 = new_n10101 & ~new_n10102;
  assign new_n10105 = ~new_n10103 & ~new_n10104;
  assign new_n10106 = new_n10099 & ~new_n10105;
  assign new_n10107 = new_n10088 & new_n10096;
  assign new_n10108 = ~new_n10097 & ~new_n10107;
  assign new_n10109 = ~new_n10106 & new_n10108;
  assign new_n10110 = ~new_n10097 & ~new_n10109;
  assign new_n10111 = new_n10079 & new_n10110;
  assign new_n10112 = ~new_n10077 & ~new_n10111;
  assign new_n10113 = A705 & A708;
  assign new_n10114 = A706 & A707;
  assign new_n10115 = A703 & A704;
  assign new_n10116 = ~new_n10114 & ~new_n10115;
  assign new_n10117 = new_n10113 & ~new_n10116;
  assign new_n10118 = ~A703 & ~A704;
  assign new_n10119 = ~A705 & A708;
  assign new_n10120 = new_n10114 & new_n10119;
  assign new_n10121 = ~A705 & ~new_n10115;
  assign new_n10122 = ~A706 & ~A707;
  assign new_n10123 = ~new_n10114 & ~new_n10122;
  assign new_n10124 = A708 & ~new_n10123;
  assign new_n10125 = ~A708 & ~new_n10114;
  assign new_n10126 = ~new_n10121 & ~new_n10125;
  assign new_n10127 = ~new_n10124 & new_n10126;
  assign new_n10128 = ~new_n10120 & ~new_n10127;
  assign new_n10129 = ~new_n10118 & ~new_n10128;
  assign new_n10130 = A707 & new_n10115;
  assign new_n10131 = new_n10117 & ~new_n10130;
  assign new_n10132 = A705 & ~A708;
  assign new_n10133 = new_n10115 & ~new_n10122;
  assign new_n10134 = new_n10132 & new_n10133;
  assign new_n10135 = ~new_n10113 & new_n10118;
  assign new_n10136 = new_n10122 & new_n10135;
  assign new_n10137 = ~new_n10134 & ~new_n10136;
  assign new_n10138 = ~new_n10131 & new_n10137;
  assign new_n10139 = ~new_n10129 & new_n10138;
  assign new_n10140 = ~new_n10118 & ~new_n10139;
  assign new_n10141 = ~new_n10117 & ~new_n10140;
  assign new_n10142 = ~A712 & ~A713;
  assign new_n10143 = ~A709 & ~A711;
  assign new_n10144 = A709 & A711;
  assign new_n10145 = ~new_n10143 & ~new_n10144;
  assign new_n10146 = ~A710 & new_n10145;
  assign new_n10147 = ~new_n10143 & ~new_n10146;
  assign new_n10148 = ~new_n10142 & new_n10147;
  assign new_n10149 = A712 & A713;
  assign new_n10150 = ~A714 & ~new_n10149;
  assign new_n10151 = new_n10148 & ~new_n10150;
  assign new_n10152 = ~A714 & ~new_n10148;
  assign new_n10153 = A710 & ~new_n10145;
  assign new_n10154 = ~new_n10146 & ~new_n10153;
  assign new_n10155 = ~new_n10147 & ~new_n10149;
  assign new_n10156 = new_n10147 & new_n10149;
  assign new_n10157 = ~new_n10155 & ~new_n10156;
  assign new_n10158 = A714 & ~new_n10157;
  assign new_n10159 = ~new_n10152 & ~new_n10154;
  assign new_n10160 = ~new_n10158 & new_n10159;
  assign new_n10161 = ~new_n10151 & ~new_n10160;
  assign new_n10162 = new_n10141 & new_n10161;
  assign new_n10163 = ~new_n10115 & ~new_n10118;
  assign new_n10164 = ~new_n10119 & ~new_n10132;
  assign new_n10165 = new_n10163 & ~new_n10164;
  assign new_n10166 = ~new_n10163 & new_n10164;
  assign new_n10167 = ~new_n10165 & ~new_n10166;
  assign new_n10168 = new_n10123 & new_n10167;
  assign new_n10169 = new_n10121 & new_n10125;
  assign new_n10170 = ~new_n10168 & new_n10169;
  assign new_n10171 = new_n10139 & ~new_n10170;
  assign new_n10172 = A714 & ~new_n10154;
  assign new_n10173 = new_n10142 & ~new_n10147;
  assign new_n10174 = ~new_n10172 & new_n10173;
  assign new_n10175 = ~new_n10147 & new_n10150;
  assign new_n10176 = ~new_n10151 & ~new_n10175;
  assign new_n10177 = new_n10154 & ~new_n10176;
  assign new_n10178 = ~new_n10160 & ~new_n10174;
  assign new_n10179 = ~new_n10177 & new_n10178;
  assign new_n10180 = ~new_n10171 & ~new_n10179;
  assign new_n10181 = ~new_n10123 & ~new_n10167;
  assign new_n10182 = ~new_n10168 & ~new_n10181;
  assign new_n10183 = ~A714 & new_n10154;
  assign new_n10184 = ~new_n10172 & ~new_n10183;
  assign new_n10185 = ~new_n10142 & ~new_n10149;
  assign new_n10186 = ~new_n10184 & new_n10185;
  assign new_n10187 = new_n10184 & ~new_n10185;
  assign new_n10188 = ~new_n10186 & ~new_n10187;
  assign new_n10189 = new_n10182 & ~new_n10188;
  assign new_n10190 = new_n10171 & new_n10179;
  assign new_n10191 = ~new_n10180 & ~new_n10190;
  assign new_n10192 = ~new_n10189 & new_n10191;
  assign new_n10193 = ~new_n10180 & ~new_n10192;
  assign new_n10194 = ~new_n10141 & ~new_n10161;
  assign new_n10195 = ~new_n10162 & ~new_n10194;
  assign new_n10196 = ~new_n10193 & new_n10195;
  assign new_n10197 = ~new_n10162 & ~new_n10196;
  assign new_n10198 = ~new_n10112 & new_n10197;
  assign new_n10199 = new_n10112 & ~new_n10197;
  assign new_n10200 = ~new_n10198 & ~new_n10199;
  assign new_n10201 = new_n10193 & ~new_n10195;
  assign new_n10202 = ~new_n10196 & ~new_n10201;
  assign new_n10203 = ~new_n10079 & ~new_n10110;
  assign new_n10204 = ~new_n10111 & ~new_n10203;
  assign new_n10205 = ~new_n10202 & new_n10204;
  assign new_n10206 = new_n10106 & ~new_n10108;
  assign new_n10207 = ~new_n10109 & ~new_n10206;
  assign new_n10208 = new_n10189 & ~new_n10191;
  assign new_n10209 = ~new_n10192 & ~new_n10208;
  assign new_n10210 = ~new_n10207 & ~new_n10209;
  assign new_n10211 = ~new_n10099 & new_n10105;
  assign new_n10212 = ~new_n10106 & ~new_n10211;
  assign new_n10213 = ~new_n10182 & new_n10188;
  assign new_n10214 = ~new_n10189 & ~new_n10213;
  assign new_n10215 = new_n10212 & new_n10214;
  assign new_n10216 = ~new_n10191 & new_n10207;
  assign new_n10217 = new_n10215 & ~new_n10216;
  assign new_n10218 = ~new_n10210 & ~new_n10217;
  assign new_n10219 = new_n10202 & ~new_n10204;
  assign new_n10220 = ~new_n10205 & ~new_n10219;
  assign new_n10221 = ~new_n10218 & new_n10220;
  assign new_n10222 = ~new_n10205 & ~new_n10221;
  assign new_n10223 = new_n10200 & ~new_n10222;
  assign new_n10224 = ~new_n10198 & ~new_n10223;
  assign new_n10225 = A742 & A743;
  assign new_n10226 = ~A740 & ~A741;
  assign new_n10227 = A740 & A741;
  assign new_n10228 = ~new_n10226 & ~new_n10227;
  assign new_n10229 = ~A739 & new_n10228;
  assign new_n10230 = ~new_n10226 & ~new_n10229;
  assign new_n10231 = new_n10225 & new_n10230;
  assign new_n10232 = ~A742 & ~A743;
  assign new_n10233 = A739 & ~new_n10228;
  assign new_n10234 = ~new_n10229 & ~new_n10233;
  assign new_n10235 = ~A744 & new_n10234;
  assign new_n10236 = A744 & ~new_n10234;
  assign new_n10237 = ~new_n10235 & ~new_n10236;
  assign new_n10238 = new_n10230 & ~new_n10232;
  assign new_n10239 = new_n10237 & new_n10238;
  assign new_n10240 = ~new_n10225 & ~new_n10230;
  assign new_n10241 = ~new_n10231 & new_n10236;
  assign new_n10242 = ~new_n10240 & new_n10241;
  assign new_n10243 = ~new_n10239 & ~new_n10242;
  assign new_n10244 = ~new_n10231 & new_n10243;
  assign new_n10245 = ~A746 & ~A747;
  assign new_n10246 = A746 & A747;
  assign new_n10247 = ~new_n10245 & ~new_n10246;
  assign new_n10248 = ~A745 & new_n10247;
  assign new_n10249 = ~new_n10245 & ~new_n10248;
  assign new_n10250 = ~A749 & ~A750;
  assign new_n10251 = A749 & A750;
  assign new_n10252 = ~new_n10250 & ~new_n10251;
  assign new_n10253 = ~A748 & new_n10252;
  assign new_n10254 = ~new_n10250 & ~new_n10253;
  assign new_n10255 = ~new_n10249 & ~new_n10254;
  assign new_n10256 = new_n10249 & new_n10254;
  assign new_n10257 = A748 & ~new_n10252;
  assign new_n10258 = ~new_n10253 & ~new_n10257;
  assign new_n10259 = A745 & ~new_n10247;
  assign new_n10260 = ~new_n10248 & ~new_n10259;
  assign new_n10261 = ~new_n10258 & ~new_n10260;
  assign new_n10262 = ~new_n10256 & ~new_n10261;
  assign new_n10263 = ~new_n10255 & ~new_n10262;
  assign new_n10264 = ~new_n10244 & new_n10263;
  assign new_n10265 = ~new_n10255 & ~new_n10256;
  assign new_n10266 = ~new_n10225 & ~new_n10232;
  assign new_n10267 = new_n10237 & ~new_n10266;
  assign new_n10268 = ~new_n10237 & new_n10266;
  assign new_n10269 = ~new_n10267 & ~new_n10268;
  assign new_n10270 = new_n10258 & new_n10260;
  assign new_n10271 = ~new_n10261 & ~new_n10270;
  assign new_n10272 = ~new_n10269 & new_n10271;
  assign new_n10273 = ~new_n10261 & ~new_n10272;
  assign new_n10274 = new_n10265 & ~new_n10273;
  assign new_n10275 = ~new_n10265 & new_n10273;
  assign new_n10276 = ~new_n10274 & ~new_n10275;
  assign new_n10277 = new_n10231 & ~new_n10233;
  assign new_n10278 = ~new_n10235 & ~new_n10267;
  assign new_n10279 = new_n10240 & ~new_n10278;
  assign new_n10280 = new_n10243 & ~new_n10277;
  assign new_n10281 = ~new_n10279 & new_n10280;
  assign new_n10282 = new_n10276 & new_n10281;
  assign new_n10283 = new_n10265 & new_n10272;
  assign new_n10284 = ~new_n10282 & ~new_n10283;
  assign new_n10285 = new_n10244 & ~new_n10263;
  assign new_n10286 = ~new_n10264 & ~new_n10285;
  assign new_n10287 = ~new_n10284 & new_n10286;
  assign new_n10288 = ~new_n10264 & ~new_n10287;
  assign new_n10289 = A735 & A738;
  assign new_n10290 = A736 & A737;
  assign new_n10291 = A733 & A734;
  assign new_n10292 = ~new_n10290 & ~new_n10291;
  assign new_n10293 = new_n10289 & ~new_n10292;
  assign new_n10294 = ~A733 & ~A734;
  assign new_n10295 = ~A735 & A738;
  assign new_n10296 = new_n10290 & new_n10295;
  assign new_n10297 = ~A735 & ~new_n10291;
  assign new_n10298 = ~A736 & ~A737;
  assign new_n10299 = ~new_n10290 & ~new_n10298;
  assign new_n10300 = A738 & ~new_n10299;
  assign new_n10301 = ~A738 & ~new_n10290;
  assign new_n10302 = ~new_n10297 & ~new_n10301;
  assign new_n10303 = ~new_n10300 & new_n10302;
  assign new_n10304 = ~new_n10296 & ~new_n10303;
  assign new_n10305 = ~new_n10294 & ~new_n10304;
  assign new_n10306 = A737 & new_n10291;
  assign new_n10307 = new_n10293 & ~new_n10306;
  assign new_n10308 = A735 & ~A738;
  assign new_n10309 = new_n10291 & ~new_n10298;
  assign new_n10310 = new_n10308 & new_n10309;
  assign new_n10311 = ~new_n10289 & new_n10294;
  assign new_n10312 = new_n10298 & new_n10311;
  assign new_n10313 = ~new_n10310 & ~new_n10312;
  assign new_n10314 = ~new_n10307 & new_n10313;
  assign new_n10315 = ~new_n10305 & new_n10314;
  assign new_n10316 = ~new_n10294 & ~new_n10315;
  assign new_n10317 = ~new_n10293 & ~new_n10316;
  assign new_n10318 = A729 & A732;
  assign new_n10319 = A730 & A731;
  assign new_n10320 = A727 & A728;
  assign new_n10321 = ~new_n10319 & ~new_n10320;
  assign new_n10322 = new_n10318 & ~new_n10321;
  assign new_n10323 = ~A727 & ~A728;
  assign new_n10324 = ~A729 & A732;
  assign new_n10325 = new_n10319 & new_n10324;
  assign new_n10326 = ~A729 & ~new_n10320;
  assign new_n10327 = ~A730 & ~A731;
  assign new_n10328 = ~new_n10319 & ~new_n10327;
  assign new_n10329 = A732 & ~new_n10328;
  assign new_n10330 = ~A732 & ~new_n10319;
  assign new_n10331 = ~new_n10326 & ~new_n10330;
  assign new_n10332 = ~new_n10329 & new_n10331;
  assign new_n10333 = ~new_n10325 & ~new_n10332;
  assign new_n10334 = ~new_n10323 & ~new_n10333;
  assign new_n10335 = A731 & new_n10320;
  assign new_n10336 = new_n10322 & ~new_n10335;
  assign new_n10337 = ~new_n10318 & new_n10323;
  assign new_n10338 = new_n10327 & new_n10337;
  assign new_n10339 = A729 & ~A732;
  assign new_n10340 = new_n10320 & ~new_n10327;
  assign new_n10341 = new_n10339 & new_n10340;
  assign new_n10342 = ~new_n10338 & ~new_n10341;
  assign new_n10343 = ~new_n10336 & new_n10342;
  assign new_n10344 = ~new_n10334 & new_n10343;
  assign new_n10345 = ~new_n10323 & ~new_n10344;
  assign new_n10346 = ~new_n10322 & ~new_n10345;
  assign new_n10347 = new_n10317 & new_n10346;
  assign new_n10348 = ~new_n10320 & ~new_n10323;
  assign new_n10349 = ~new_n10324 & ~new_n10339;
  assign new_n10350 = new_n10348 & ~new_n10349;
  assign new_n10351 = ~new_n10348 & new_n10349;
  assign new_n10352 = ~new_n10350 & ~new_n10351;
  assign new_n10353 = new_n10328 & new_n10352;
  assign new_n10354 = ~new_n10328 & ~new_n10352;
  assign new_n10355 = ~new_n10353 & ~new_n10354;
  assign new_n10356 = ~new_n10291 & ~new_n10294;
  assign new_n10357 = ~new_n10295 & ~new_n10308;
  assign new_n10358 = new_n10356 & ~new_n10357;
  assign new_n10359 = ~new_n10356 & new_n10357;
  assign new_n10360 = ~new_n10358 & ~new_n10359;
  assign new_n10361 = new_n10299 & new_n10360;
  assign new_n10362 = ~new_n10299 & ~new_n10360;
  assign new_n10363 = ~new_n10361 & ~new_n10362;
  assign new_n10364 = new_n10355 & new_n10363;
  assign new_n10365 = new_n10326 & new_n10330;
  assign new_n10366 = ~new_n10353 & new_n10365;
  assign new_n10367 = new_n10344 & ~new_n10366;
  assign new_n10368 = ~new_n10364 & ~new_n10367;
  assign new_n10369 = new_n10364 & new_n10367;
  assign new_n10370 = ~new_n10368 & ~new_n10369;
  assign new_n10371 = new_n10297 & new_n10301;
  assign new_n10372 = ~new_n10361 & new_n10371;
  assign new_n10373 = new_n10315 & ~new_n10372;
  assign new_n10374 = new_n10370 & ~new_n10373;
  assign new_n10375 = ~new_n10368 & ~new_n10374;
  assign new_n10376 = ~new_n10317 & ~new_n10346;
  assign new_n10377 = ~new_n10347 & ~new_n10376;
  assign new_n10378 = ~new_n10375 & new_n10377;
  assign new_n10379 = ~new_n10347 & ~new_n10378;
  assign new_n10380 = ~new_n10288 & new_n10379;
  assign new_n10381 = new_n10288 & ~new_n10379;
  assign new_n10382 = ~new_n10380 & ~new_n10381;
  assign new_n10383 = new_n10284 & ~new_n10286;
  assign new_n10384 = ~new_n10287 & ~new_n10383;
  assign new_n10385 = ~new_n10370 & new_n10373;
  assign new_n10386 = ~new_n10374 & ~new_n10385;
  assign new_n10387 = ~new_n10276 & ~new_n10281;
  assign new_n10388 = ~new_n10282 & ~new_n10387;
  assign new_n10389 = new_n10386 & ~new_n10388;
  assign new_n10390 = ~new_n10355 & ~new_n10363;
  assign new_n10391 = ~new_n10364 & ~new_n10390;
  assign new_n10392 = new_n10269 & ~new_n10271;
  assign new_n10393 = ~new_n10272 & ~new_n10392;
  assign new_n10394 = new_n10391 & new_n10393;
  assign new_n10395 = ~new_n10386 & new_n10388;
  assign new_n10396 = ~new_n10389 & ~new_n10395;
  assign new_n10397 = ~new_n10394 & new_n10396;
  assign new_n10398 = ~new_n10389 & ~new_n10397;
  assign new_n10399 = new_n10384 & new_n10398;
  assign new_n10400 = new_n10375 & ~new_n10377;
  assign new_n10401 = ~new_n10378 & ~new_n10400;
  assign new_n10402 = ~new_n10384 & ~new_n10398;
  assign new_n10403 = ~new_n10399 & ~new_n10402;
  assign new_n10404 = ~new_n10401 & new_n10403;
  assign new_n10405 = ~new_n10399 & ~new_n10404;
  assign new_n10406 = new_n10382 & ~new_n10405;
  assign new_n10407 = ~new_n10380 & ~new_n10406;
  assign new_n10408 = new_n10224 & new_n10407;
  assign new_n10409 = ~new_n10382 & new_n10405;
  assign new_n10410 = ~new_n10406 & ~new_n10409;
  assign new_n10411 = new_n10218 & ~new_n10220;
  assign new_n10412 = ~new_n10221 & ~new_n10411;
  assign new_n10413 = new_n10401 & ~new_n10403;
  assign new_n10414 = ~new_n10404 & ~new_n10413;
  assign new_n10415 = new_n10412 & new_n10414;
  assign new_n10416 = ~new_n10412 & ~new_n10414;
  assign new_n10417 = ~new_n10415 & ~new_n10416;
  assign new_n10418 = new_n10394 & ~new_n10396;
  assign new_n10419 = ~new_n10397 & ~new_n10418;
  assign new_n10420 = ~new_n10189 & ~new_n10215;
  assign new_n10421 = new_n10191 & ~new_n10207;
  assign new_n10422 = ~new_n10216 & ~new_n10421;
  assign new_n10423 = new_n10420 & new_n10422;
  assign new_n10424 = ~new_n10420 & ~new_n10422;
  assign new_n10425 = ~new_n10423 & ~new_n10424;
  assign new_n10426 = ~new_n10419 & ~new_n10425;
  assign new_n10427 = ~new_n10212 & ~new_n10214;
  assign new_n10428 = ~new_n10215 & ~new_n10427;
  assign new_n10429 = ~new_n10391 & ~new_n10393;
  assign new_n10430 = ~new_n10394 & ~new_n10429;
  assign new_n10431 = new_n10428 & new_n10430;
  assign new_n10432 = new_n10419 & new_n10425;
  assign new_n10433 = ~new_n10426 & ~new_n10432;
  assign new_n10434 = new_n10431 & new_n10433;
  assign new_n10435 = ~new_n10426 & ~new_n10434;
  assign new_n10436 = new_n10417 & ~new_n10435;
  assign new_n10437 = ~new_n10415 & ~new_n10436;
  assign new_n10438 = ~new_n10410 & new_n10437;
  assign new_n10439 = ~new_n10200 & new_n10222;
  assign new_n10440 = ~new_n10223 & ~new_n10439;
  assign new_n10441 = new_n10410 & ~new_n10437;
  assign new_n10442 = ~new_n10438 & ~new_n10441;
  assign new_n10443 = ~new_n10440 & new_n10442;
  assign new_n10444 = ~new_n10438 & ~new_n10443;
  assign new_n10445 = ~new_n10224 & ~new_n10407;
  assign new_n10446 = ~new_n10408 & ~new_n10445;
  assign new_n10447 = ~new_n10444 & new_n10446;
  assign new_n10448 = ~new_n10408 & ~new_n10447;
  assign new_n10449 = ~new_n10027 & ~new_n10448;
  assign new_n10450 = new_n10027 & new_n10448;
  assign new_n10451 = new_n10023 & ~new_n10025;
  assign new_n10452 = ~new_n10026 & ~new_n10451;
  assign new_n10453 = new_n10444 & ~new_n10446;
  assign new_n10454 = ~new_n10447 & ~new_n10453;
  assign new_n10455 = ~new_n10452 & ~new_n10454;
  assign new_n10456 = ~new_n9998 & ~new_n10021;
  assign new_n10457 = ~new_n10022 & ~new_n10456;
  assign new_n10458 = ~new_n10417 & new_n10435;
  assign new_n10459 = ~new_n10436 & ~new_n10458;
  assign new_n10460 = ~new_n10431 & ~new_n10433;
  assign new_n10461 = ~new_n10434 & ~new_n10460;
  assign new_n10462 = new_n10012 & new_n10461;
  assign new_n10463 = ~new_n10428 & ~new_n10430;
  assign new_n10464 = ~new_n10431 & ~new_n10463;
  assign new_n10465 = ~new_n10007 & ~new_n10009;
  assign new_n10466 = ~new_n10010 & ~new_n10465;
  assign new_n10467 = new_n10464 & new_n10466;
  assign new_n10468 = ~new_n10010 & ~new_n10467;
  assign new_n10469 = ~new_n10012 & ~new_n10461;
  assign new_n10470 = ~new_n10462 & ~new_n10469;
  assign new_n10471 = ~new_n10468 & new_n10470;
  assign new_n10472 = ~new_n10462 & ~new_n10471;
  assign new_n10473 = ~new_n10013 & ~new_n10472;
  assign new_n10474 = ~new_n10459 & ~new_n10473;
  assign new_n10475 = new_n10017 & ~new_n10019;
  assign new_n10476 = ~new_n10020 & ~new_n10475;
  assign new_n10477 = new_n10459 & new_n10473;
  assign new_n10478 = ~new_n10474 & ~new_n10477;
  assign new_n10479 = ~new_n10476 & new_n10478;
  assign new_n10480 = ~new_n10474 & ~new_n10479;
  assign new_n10481 = ~new_n10457 & new_n10480;
  assign new_n10482 = new_n10440 & ~new_n10442;
  assign new_n10483 = ~new_n10443 & ~new_n10482;
  assign new_n10484 = new_n10457 & ~new_n10480;
  assign new_n10485 = ~new_n10481 & ~new_n10484;
  assign new_n10486 = ~new_n10483 & new_n10485;
  assign new_n10487 = ~new_n10481 & ~new_n10486;
  assign new_n10488 = new_n10452 & new_n10454;
  assign new_n10489 = ~new_n10455 & ~new_n10488;
  assign new_n10490 = ~new_n10487 & new_n10489;
  assign new_n10491 = ~new_n10455 & ~new_n10490;
  assign new_n10492 = ~new_n10450 & new_n10491;
  assign new_n10493 = ~new_n10449 & ~new_n10492;
  assign new_n10494 = new_n9580 & ~new_n10493;
  assign new_n10495 = new_n10487 & ~new_n10489;
  assign new_n10496 = ~new_n10490 & ~new_n10495;
  assign new_n10497 = ~new_n9565 & ~new_n9567;
  assign new_n10498 = ~new_n9568 & ~new_n10497;
  assign new_n10499 = new_n10483 & ~new_n10485;
  assign new_n10500 = ~new_n10486 & ~new_n10499;
  assign new_n10501 = ~new_n10498 & new_n10500;
  assign new_n10502 = new_n10476 & ~new_n10478;
  assign new_n10503 = ~new_n10479 & ~new_n10502;
  assign new_n10504 = ~new_n10464 & ~new_n10466;
  assign new_n10505 = ~new_n10467 & ~new_n10504;
  assign new_n10506 = ~new_n9545 & ~new_n9547;
  assign new_n10507 = ~new_n9548 & ~new_n10506;
  assign new_n10508 = new_n10505 & new_n10507;
  assign new_n10509 = new_n10468 & ~new_n10470;
  assign new_n10510 = ~new_n10471 & ~new_n10509;
  assign new_n10511 = ~new_n10508 & ~new_n10510;
  assign new_n10512 = new_n9542 & ~new_n9552;
  assign new_n10513 = ~new_n9553 & ~new_n10512;
  assign new_n10514 = new_n10508 & new_n10510;
  assign new_n10515 = ~new_n10511 & ~new_n10514;
  assign new_n10516 = new_n10513 & new_n10515;
  assign new_n10517 = ~new_n10511 & ~new_n10516;
  assign new_n10518 = new_n10503 & ~new_n10517;
  assign new_n10519 = new_n9558 & ~new_n9560;
  assign new_n10520 = ~new_n9561 & ~new_n10519;
  assign new_n10521 = ~new_n10503 & new_n10517;
  assign new_n10522 = ~new_n10518 & ~new_n10521;
  assign new_n10523 = ~new_n10520 & new_n10522;
  assign new_n10524 = ~new_n10518 & ~new_n10523;
  assign new_n10525 = new_n10498 & ~new_n10500;
  assign new_n10526 = ~new_n10501 & ~new_n10525;
  assign new_n10527 = new_n10524 & new_n10526;
  assign new_n10528 = ~new_n10501 & ~new_n10527;
  assign new_n10529 = ~new_n10496 & new_n10528;
  assign new_n10530 = new_n9572 & ~new_n9574;
  assign new_n10531 = ~new_n9575 & ~new_n10530;
  assign new_n10532 = new_n10496 & ~new_n10528;
  assign new_n10533 = ~new_n10529 & ~new_n10532;
  assign new_n10534 = ~new_n10531 & new_n10533;
  assign new_n10535 = ~new_n10529 & ~new_n10534;
  assign new_n10536 = ~new_n10449 & ~new_n10450;
  assign new_n10537 = new_n10491 & ~new_n10536;
  assign new_n10538 = ~new_n10491 & new_n10536;
  assign new_n10539 = ~new_n10537 & ~new_n10538;
  assign new_n10540 = new_n10535 & new_n10539;
  assign new_n10541 = new_n9576 & ~new_n9578;
  assign new_n10542 = ~new_n9579 & ~new_n10541;
  assign new_n10543 = ~new_n10535 & ~new_n10539;
  assign new_n10544 = ~new_n10540 & ~new_n10543;
  assign new_n10545 = new_n10542 & new_n10544;
  assign new_n10546 = ~new_n10540 & ~new_n10545;
  assign new_n10547 = ~new_n9580 & new_n10493;
  assign new_n10548 = ~new_n10494 & ~new_n10547;
  assign new_n10549 = new_n10546 & new_n10548;
  assign new_n10550 = ~new_n10494 & ~new_n10549;
  assign new_n10551 = new_n8703 & ~new_n10550;
  assign new_n10552 = ~new_n8703 & new_n10550;
  assign new_n10553 = ~new_n10551 & ~new_n10552;
  assign new_n10554 = ~new_n8651 & ~new_n8701;
  assign new_n10555 = ~new_n8702 & ~new_n10554;
  assign new_n10556 = ~new_n10542 & ~new_n10544;
  assign new_n10557 = ~new_n10545 & ~new_n10556;
  assign new_n10558 = new_n8697 & ~new_n8699;
  assign new_n10559 = ~new_n8700 & ~new_n10558;
  assign new_n10560 = ~new_n10557 & new_n10559;
  assign new_n10561 = ~new_n8690 & ~new_n8692;
  assign new_n10562 = ~new_n8693 & ~new_n10561;
  assign new_n10563 = new_n8683 & ~new_n8685;
  assign new_n10564 = ~new_n8686 & ~new_n10563;
  assign new_n10565 = new_n8679 & ~new_n8681;
  assign new_n10566 = ~new_n8682 & ~new_n10565;
  assign new_n10567 = new_n8672 & ~new_n8674;
  assign new_n10568 = ~new_n8675 & ~new_n10567;
  assign new_n10569 = ~new_n10513 & ~new_n10515;
  assign new_n10570 = ~new_n10516 & ~new_n10569;
  assign new_n10571 = ~new_n10568 & new_n10570;
  assign new_n10572 = ~new_n8666 & ~new_n8668;
  assign new_n10573 = ~new_n8669 & ~new_n10572;
  assign new_n10574 = ~new_n10505 & ~new_n10507;
  assign new_n10575 = ~new_n10508 & ~new_n10574;
  assign new_n10576 = new_n10573 & new_n10575;
  assign new_n10577 = new_n10568 & ~new_n10570;
  assign new_n10578 = ~new_n10571 & ~new_n10577;
  assign new_n10579 = ~new_n10576 & new_n10578;
  assign new_n10580 = ~new_n10571 & ~new_n10579;
  assign new_n10581 = ~new_n10566 & ~new_n10580;
  assign new_n10582 = new_n10520 & ~new_n10522;
  assign new_n10583 = ~new_n10523 & ~new_n10582;
  assign new_n10584 = new_n10566 & new_n10580;
  assign new_n10585 = ~new_n10581 & ~new_n10584;
  assign new_n10586 = new_n10583 & new_n10585;
  assign new_n10587 = ~new_n10581 & ~new_n10586;
  assign new_n10588 = ~new_n10564 & ~new_n10587;
  assign new_n10589 = ~new_n10524 & ~new_n10526;
  assign new_n10590 = ~new_n10527 & ~new_n10589;
  assign new_n10591 = new_n10564 & new_n10587;
  assign new_n10592 = ~new_n10588 & ~new_n10591;
  assign new_n10593 = ~new_n10590 & new_n10592;
  assign new_n10594 = ~new_n10588 & ~new_n10593;
  assign new_n10595 = new_n10562 & new_n10594;
  assign new_n10596 = new_n10531 & ~new_n10533;
  assign new_n10597 = ~new_n10534 & ~new_n10596;
  assign new_n10598 = ~new_n10562 & ~new_n10594;
  assign new_n10599 = ~new_n10595 & ~new_n10598;
  assign new_n10600 = ~new_n10597 & new_n10599;
  assign new_n10601 = ~new_n10595 & ~new_n10600;
  assign new_n10602 = new_n10557 & ~new_n10559;
  assign new_n10603 = ~new_n10560 & ~new_n10602;
  assign new_n10604 = new_n10601 & new_n10603;
  assign new_n10605 = ~new_n10560 & ~new_n10604;
  assign new_n10606 = new_n10555 & new_n10605;
  assign new_n10607 = ~new_n10546 & ~new_n10548;
  assign new_n10608 = ~new_n10549 & ~new_n10607;
  assign new_n10609 = ~new_n10555 & ~new_n10605;
  assign new_n10610 = ~new_n10606 & ~new_n10609;
  assign new_n10611 = ~new_n10608 & new_n10610;
  assign new_n10612 = ~new_n10606 & ~new_n10611;
  assign new_n10613 = new_n10553 & new_n10612;
  assign new_n10614 = ~new_n10553 & ~new_n10612;
  assign new_n10615 = ~new_n10613 & ~new_n10614;
  assign new_n10616 = ~new_n6931 & ~new_n10615;
  assign new_n10617 = new_n6931 & new_n10615;
  assign new_n10618 = new_n10608 & ~new_n10610;
  assign new_n10619 = ~new_n10611 & ~new_n10618;
  assign new_n10620 = new_n6916 & ~new_n6918;
  assign new_n10621 = ~new_n6919 & ~new_n10620;
  assign new_n10622 = ~new_n10601 & ~new_n10603;
  assign new_n10623 = ~new_n10604 & ~new_n10622;
  assign new_n10624 = ~new_n10621 & new_n10623;
  assign new_n10625 = ~new_n6878 & new_n6911;
  assign new_n10626 = ~new_n6912 & ~new_n10625;
  assign new_n10627 = new_n10597 & ~new_n10599;
  assign new_n10628 = ~new_n10600 & ~new_n10627;
  assign new_n10629 = ~new_n10626 & ~new_n10628;
  assign new_n10630 = new_n6907 & ~new_n6909;
  assign new_n10631 = ~new_n6910 & ~new_n10630;
  assign new_n10632 = new_n10590 & ~new_n10592;
  assign new_n10633 = ~new_n10593 & ~new_n10632;
  assign new_n10634 = new_n10631 & ~new_n10633;
  assign new_n10635 = ~new_n10631 & new_n10633;
  assign new_n10636 = ~new_n10634 & ~new_n10635;
  assign new_n10637 = ~new_n6887 & ~new_n6902;
  assign new_n10638 = ~new_n6903 & ~new_n10637;
  assign new_n10639 = ~new_n10583 & ~new_n10585;
  assign new_n10640 = ~new_n10586 & ~new_n10639;
  assign new_n10641 = ~new_n10638 & ~new_n10640;
  assign new_n10642 = new_n6889 & ~new_n6899;
  assign new_n10643 = ~new_n6900 & ~new_n10642;
  assign new_n10644 = new_n10576 & ~new_n10578;
  assign new_n10645 = ~new_n10579 & ~new_n10644;
  assign new_n10646 = new_n10643 & ~new_n10645;
  assign new_n10647 = ~new_n10573 & ~new_n10575;
  assign new_n10648 = ~new_n10576 & ~new_n10647;
  assign new_n10649 = ~new_n10578 & ~new_n10643;
  assign new_n10650 = ~new_n6892 & new_n6894;
  assign new_n10651 = ~new_n6895 & ~new_n10650;
  assign new_n10652 = new_n10648 & new_n10651;
  assign new_n10653 = ~new_n10649 & new_n10652;
  assign new_n10654 = ~new_n10646 & ~new_n10653;
  assign new_n10655 = new_n10638 & new_n10640;
  assign new_n10656 = ~new_n10641 & ~new_n10655;
  assign new_n10657 = ~new_n10654 & new_n10656;
  assign new_n10658 = ~new_n10641 & ~new_n10657;
  assign new_n10659 = new_n10636 & ~new_n10658;
  assign new_n10660 = ~new_n10634 & ~new_n10659;
  assign new_n10661 = ~new_n10629 & ~new_n10660;
  assign new_n10662 = new_n10621 & ~new_n10623;
  assign new_n10663 = new_n10626 & new_n10628;
  assign new_n10664 = ~new_n10661 & ~new_n10663;
  assign new_n10665 = ~new_n10662 & new_n10664;
  assign new_n10666 = ~new_n10624 & ~new_n10665;
  assign new_n10667 = ~new_n10619 & ~new_n10666;
  assign new_n10668 = new_n6923 & ~new_n6925;
  assign new_n10669 = ~new_n6926 & ~new_n10668;
  assign new_n10670 = new_n10619 & new_n10666;
  assign new_n10671 = ~new_n10669 & ~new_n10670;
  assign new_n10672 = ~new_n10667 & ~new_n10671;
  assign new_n10673 = ~new_n10617 & new_n10672;
  assign new_n10674 = ~new_n10616 & ~new_n10673;
  assign new_n10675 = new_n6929 & ~new_n10674;
  assign new_n10676 = ~new_n10551 & ~new_n10613;
  assign new_n10677 = ~new_n6859 & ~new_n6862;
  assign new_n10678 = ~new_n10676 & ~new_n10677;
  assign new_n10679 = ~new_n10616 & ~new_n10617;
  assign new_n10680 = new_n10667 & ~new_n10669;
  assign new_n10681 = ~new_n10672 & ~new_n10680;
  assign new_n10682 = new_n10679 & new_n10681;
  assign new_n10683 = new_n10669 & new_n10670;
  assign new_n10684 = ~new_n10679 & new_n10683;
  assign new_n10685 = ~new_n10682 & ~new_n10684;
  assign new_n10686 = ~new_n10636 & new_n10658;
  assign new_n10687 = ~new_n10659 & ~new_n10686;
  assign new_n10688 = new_n10578 & new_n10643;
  assign new_n10689 = new_n10653 & ~new_n10688;
  assign new_n10690 = ~new_n10643 & new_n10645;
  assign new_n10691 = ~new_n10646 & ~new_n10690;
  assign new_n10692 = ~new_n10648 & ~new_n10651;
  assign new_n10693 = ~new_n10691 & new_n10692;
  assign new_n10694 = ~new_n10689 & ~new_n10693;
  assign new_n10695 = ~A1000 & ~new_n10694;
  assign new_n10696 = new_n10654 & ~new_n10656;
  assign new_n10697 = ~new_n10657 & ~new_n10695;
  assign new_n10698 = ~new_n10696 & new_n10697;
  assign new_n10699 = ~new_n10687 & ~new_n10698;
  assign new_n10700 = ~new_n10624 & ~new_n10662;
  assign new_n10701 = new_n10661 & new_n10700;
  assign new_n10702 = ~new_n10663 & ~new_n10700;
  assign new_n10703 = ~new_n10629 & ~new_n10663;
  assign new_n10704 = new_n10660 & ~new_n10703;
  assign new_n10705 = ~new_n10699 & ~new_n10704;
  assign new_n10706 = ~new_n10701 & new_n10705;
  assign new_n10707 = ~new_n10702 & new_n10706;
  assign new_n10708 = ~new_n10685 & new_n10707;
  assign new_n10709 = new_n10676 & new_n10677;
  assign new_n10710 = ~new_n6929 & ~new_n10709;
  assign new_n10711 = new_n10674 & new_n10710;
  assign new_n10712 = ~new_n10708 & new_n10711;
  assign new_n10713 = ~new_n10678 & ~new_n10712;
  assign new_n10714 = new_n10708 & ~new_n10711;
  assign new_n10715 = ~new_n10675 & ~new_n10714;
  assign maj = new_n10713 | ~new_n10715;
endmodule


