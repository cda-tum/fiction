module top ( 
    \1 , 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124, 125,
    128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223, 226,
    232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317, 322,
    326, 329, 330, 343, 349, 350,
    1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002,
    5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361  );
  input  \1 , 13, 20, 33, 41, 45, 50, 58, 68, 77, 87, 97, 107, 116, 124,
    125, 128, 132, 137, 143, 150, 159, 169, 179, 190, 200, 213, 222, 223,
    226, 232, 238, 244, 250, 257, 264, 270, 274, 283, 294, 303, 311, 317,
    322, 326, 329, 330, 343, 349, 350;
  output 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944,
    5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361;
  wire n73, n74, n76, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1058, n1059, n1060, n1061, n1062, n1063, n1065,
    n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109;
  assign n73 = ~50 & ~58;
  assign n74 = ~68 & n73;
  assign 1713 = ~77 & n74;
  assign n76 = ~97 & ~107;
  assign 1947 = ~87 | n76;
  assign n78 = ~58 & ~68;
  assign n79 = 50 & ~n78;
  assign n80 = \1  & 13;
  assign n81 = 20 & n80;
  assign n82 = n79 & n81;
  assign n83 = ~257 & ~264;
  assign n84 = 250 & ~n83;
  assign n85 = \1  & ~13;
  assign n86 = 20 & n85;
  assign n87 = n84 & n86;
  assign n88 = 50 & 226;
  assign n89 = 58 & 232;
  assign n90 = 68 & 238;
  assign n91 = 77 & 244;
  assign n92 = ~n88 & ~n89;
  assign n93 = ~n90 & n92;
  assign n94 = ~n91 & n93;
  assign n95 = 87 & 250;
  assign n96 = 97 & 257;
  assign n97 = 107 & 264;
  assign n98 = 116 & 270;
  assign n99 = ~n95 & ~n96;
  assign n100 = ~n97 & n99;
  assign n101 = ~n98 & n100;
  assign n102 = n94 & n101;
  assign n103 = ~n81 & ~n86;
  assign n104 = ~n102 & n103;
  assign n105 = ~n82 & ~n87;
  assign 3195 = ~n104 & n105;
  assign n107 = ~264 & 270;
  assign n108 = 264 & ~270;
  assign n109 = ~n107 & ~n108;
  assign n110 = ~250 & 257;
  assign n111 = 250 & ~257;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~n109 & n112;
  assign n114 = n109 & ~n112;
  assign n115 = ~n113 & ~n114;
  assign n116 = ~238 & 244;
  assign n117 = 238 & ~244;
  assign n118 = ~n116 & ~n117;
  assign n119 = ~226 & 232;
  assign n120 = 226 & ~232;
  assign n121 = ~n119 & ~n120;
  assign n122 = ~n118 & n121;
  assign n123 = n118 & ~n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = ~n115 & n124;
  assign n126 = n115 & ~n124;
  assign 3833 = ~n125 & ~n126;
  assign n128 = 107 & ~116;
  assign n129 = ~107 & 116;
  assign n130 = ~n128 & ~n129;
  assign n131 = 87 & ~97;
  assign n132 = ~87 & 97;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n130 & n133;
  assign n135 = n130 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = 68 & ~77;
  assign n138 = ~68 & 77;
  assign n139 = ~n137 & ~n138;
  assign n140 = 50 & 58;
  assign n141 = ~n73 & ~n140;
  assign n142 = ~n139 & n141;
  assign n143 = n139 & ~n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = ~n136 & n144;
  assign n146 = n136 & ~n144;
  assign 3987 = n145 | n146;
  assign n148 = ~87 & ~97;
  assign n149 = ~107 & n148;
  assign n150 = 20 & ~n149;
  assign n151 = ~20 & 33;
  assign n152 = 97 & n151;
  assign n153 = ~20 & ~n151;
  assign n154 = 68 & n153;
  assign n155 = ~n150 & ~n152;
  assign n156 = ~n154 & n155;
  assign n157 = \1  & 20;
  assign n158 = 33 & n157;
  assign n159 = ~n80 & ~n158;
  assign n160 = ~n156 & ~n159;
  assign n161 = 13 & 20;
  assign n162 = ~\1  & n161;
  assign n163 = ~87 & n162;
  assign n164 = ~\1  & 33;
  assign n165 = n159 & ~n162;
  assign n166 = 87 & ~n164;
  assign n167 = n165 & n166;
  assign n168 = ~n160 & ~n163;
  assign n169 = ~n167 & n168;
  assign n170 = 33 & 41;
  assign n171 = n80 & ~n170;
  assign n172 = ~\1  & 45;
  assign n173 = 250 & ~n171;
  assign n174 = ~n172 & n173;
  assign n175 = 274 & ~n171;
  assign n176 = n172 & n175;
  assign n177 = 33 & 116;
  assign n178 = ~33 & ~349;
  assign n179 = 238 & n178;
  assign n180 = ~33 & ~n178;
  assign n181 = 244 & n180;
  assign n182 = ~n177 & ~n179;
  assign n183 = ~n181 & n182;
  assign n184 = n171 & ~n183;
  assign n185 = ~n174 & ~n176;
  assign n186 = ~n184 & n185;
  assign n187 = 169 & ~n169;
  assign n188 = ~n186 & n187;
  assign n189 = 179 & ~n169;
  assign n190 = n186 & n189;
  assign n191 = ~n188 & ~n190;
  assign n192 = 190 & n169;
  assign n193 = n186 & n192;
  assign n194 = 200 & n169;
  assign n195 = ~n186 & n194;
  assign n196 = ~n193 & ~n195;
  assign n197 = n169 & n196;
  assign n198 = n191 & ~n197;
  assign n199 = ~97 & 107;
  assign n200 = 97 & ~107;
  assign n201 = ~n199 & ~n200;
  assign n202 = 20 & n201;
  assign n203 = 107 & n151;
  assign n204 = 77 & n153;
  assign n205 = ~n202 & ~n203;
  assign n206 = ~n204 & n205;
  assign n207 = ~n159 & ~n206;
  assign n208 = ~97 & n162;
  assign n209 = 97 & ~n164;
  assign n210 = n165 & n209;
  assign n211 = ~n207 & ~n208;
  assign n212 = ~n210 & n211;
  assign n213 = ~41 & n172;
  assign n214 = 257 & ~n171;
  assign n215 = ~n213 & n214;
  assign n216 = n175 & n213;
  assign n217 = 33 & 283;
  assign n218 = 244 & n178;
  assign n219 = 250 & n180;
  assign n220 = ~n217 & ~n218;
  assign n221 = ~n219 & n220;
  assign n222 = n171 & ~n221;
  assign n223 = ~n215 & ~n216;
  assign n224 = ~n222 & n223;
  assign n225 = 169 & ~n212;
  assign n226 = ~n224 & n225;
  assign n227 = 179 & ~n212;
  assign n228 = n224 & n227;
  assign n229 = ~n226 & ~n228;
  assign n230 = 190 & n212;
  assign n231 = n224 & n230;
  assign n232 = 200 & n212;
  assign n233 = ~n224 & n232;
  assign n234 = ~n231 & ~n233;
  assign n235 = n212 & n234;
  assign n236 = n229 & ~n235;
  assign n237 = 20 & ~107;
  assign n238 = 116 & n151;
  assign n239 = 87 & n153;
  assign n240 = ~n237 & ~n238;
  assign n241 = ~n239 & n240;
  assign n242 = ~n159 & ~n241;
  assign n243 = ~107 & n162;
  assign n244 = 107 & ~n164;
  assign n245 = n165 & n244;
  assign n246 = ~n242 & ~n243;
  assign n247 = ~n245 & n246;
  assign n248 = 264 & ~n171;
  assign n249 = ~n213 & n248;
  assign n250 = 33 & 294;
  assign n251 = 250 & n178;
  assign n252 = 257 & n180;
  assign n253 = ~n250 & ~n251;
  assign n254 = ~n252 & n253;
  assign n255 = n171 & ~n254;
  assign n256 = ~n216 & ~n249;
  assign n257 = ~n255 & n256;
  assign n258 = 169 & ~n247;
  assign n259 = ~n257 & n258;
  assign n260 = 179 & ~n247;
  assign n261 = n257 & n260;
  assign n262 = ~n259 & ~n261;
  assign n263 = 190 & n247;
  assign n264 = n257 & n263;
  assign n265 = 200 & n247;
  assign n266 = ~n257 & n265;
  assign n267 = ~n264 & ~n266;
  assign n268 = n247 & n267;
  assign n269 = n262 & ~n268;
  assign n270 = 20 & 116;
  assign n271 = 283 & n151;
  assign n272 = 97 & n153;
  assign n273 = ~n270 & ~n271;
  assign n274 = ~n272 & n273;
  assign n275 = ~n159 & ~n274;
  assign n276 = ~116 & n162;
  assign n277 = 116 & ~n164;
  assign n278 = n165 & n277;
  assign n279 = ~n275 & ~n276;
  assign n280 = ~n278 & n279;
  assign n281 = 270 & ~n171;
  assign n282 = ~n213 & n281;
  assign n283 = 33 & 303;
  assign n284 = 257 & n178;
  assign n285 = 264 & n180;
  assign n286 = ~n283 & ~n284;
  assign n287 = ~n285 & n286;
  assign n288 = n171 & ~n287;
  assign n289 = ~n216 & ~n282;
  assign n290 = ~n288 & n289;
  assign n291 = 169 & ~n280;
  assign n292 = ~n290 & n291;
  assign n293 = 179 & ~n280;
  assign n294 = n290 & n293;
  assign n295 = ~n292 & ~n294;
  assign n296 = 190 & n280;
  assign n297 = n290 & n296;
  assign n298 = 200 & n280;
  assign n299 = ~n290 & n298;
  assign n300 = ~n297 & ~n299;
  assign n301 = n280 & n300;
  assign n302 = n295 & ~n301;
  assign n303 = n198 & n236;
  assign n304 = n269 & n303;
  assign n305 = n302 & n304;
  assign n306 = 20 & ~n74;
  assign n307 = 58 & n151;
  assign n308 = 150 & n153;
  assign n309 = ~n306 & ~n307;
  assign n310 = ~n308 & n309;
  assign n311 = ~n159 & ~n310;
  assign n312 = ~50 & n162;
  assign n313 = ~\1  & 20;
  assign n314 = 50 & ~n313;
  assign n315 = n165 & n314;
  assign n316 = ~n311 & ~n312;
  assign n317 = ~n315 & n316;
  assign n318 = ~41 & ~45;
  assign n319 = ~\1  & ~n318;
  assign n320 = 226 & ~n171;
  assign n321 = ~n319 & n320;
  assign n322 = n175 & n319;
  assign n323 = 33 & 77;
  assign n324 = 222 & n178;
  assign n325 = 223 & n180;
  assign n326 = ~n323 & ~n324;
  assign n327 = ~n325 & n326;
  assign n328 = n171 & ~n327;
  assign n329 = ~n321 & ~n322;
  assign n330 = ~n328 & n329;
  assign n331 = 169 & ~n317;
  assign n332 = ~n330 & n331;
  assign n333 = 179 & ~n317;
  assign n334 = n330 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = 190 & n317;
  assign n337 = n330 & n336;
  assign n338 = 200 & n317;
  assign n339 = ~n330 & n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = n317 & n340;
  assign n342 = n335 & ~n341;
  assign n343 = ~58 & 68;
  assign n344 = 58 & ~68;
  assign n345 = ~n343 & ~n344;
  assign n346 = 20 & n345;
  assign n347 = 68 & n151;
  assign n348 = 159 & n153;
  assign n349 = ~n346 & ~n347;
  assign n350 = ~n348 & n349;
  assign n351 = ~n159 & ~n350;
  assign n352 = ~58 & n162;
  assign n353 = 58 & ~n313;
  assign n354 = n165 & n353;
  assign n355 = ~n351 & ~n352;
  assign n356 = ~n354 & n355;
  assign n357 = 232 & ~n171;
  assign n358 = ~n319 & n357;
  assign n359 = 33 & 87;
  assign n360 = 223 & n178;
  assign n361 = 226 & n180;
  assign n362 = ~n359 & ~n360;
  assign n363 = ~n361 & n362;
  assign n364 = n171 & ~n363;
  assign n365 = ~n322 & ~n358;
  assign n366 = ~n364 & n365;
  assign n367 = 169 & ~n356;
  assign n368 = ~n366 & n367;
  assign n369 = 179 & ~n356;
  assign n370 = n366 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = 190 & n356;
  assign n373 = n366 & n372;
  assign n374 = 200 & n356;
  assign n375 = ~n366 & n374;
  assign n376 = ~n373 & ~n375;
  assign n377 = n356 & n376;
  assign n378 = n371 & ~n377;
  assign n379 = 20 & ~68;
  assign n380 = 77 & n151;
  assign n381 = 50 & n153;
  assign n382 = ~n379 & ~n380;
  assign n383 = ~n381 & n382;
  assign n384 = ~n159 & ~n383;
  assign n385 = ~68 & n162;
  assign n386 = 68 & ~n313;
  assign n387 = n165 & n386;
  assign n388 = ~n384 & ~n385;
  assign n389 = ~n387 & n388;
  assign n390 = 238 & ~n171;
  assign n391 = ~n319 & n390;
  assign n392 = 33 & 97;
  assign n393 = 226 & n178;
  assign n394 = 232 & n180;
  assign n395 = ~n392 & ~n393;
  assign n396 = ~n394 & n395;
  assign n397 = n171 & ~n396;
  assign n398 = ~n322 & ~n391;
  assign n399 = ~n397 & n398;
  assign n400 = 169 & ~n389;
  assign n401 = ~n399 & n400;
  assign n402 = 179 & ~n389;
  assign n403 = n399 & n402;
  assign n404 = ~n401 & ~n403;
  assign n405 = 190 & n389;
  assign n406 = n399 & n405;
  assign n407 = 200 & n389;
  assign n408 = ~n399 & n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = n389 & n409;
  assign n411 = n404 & ~n410;
  assign n412 = 20 & 77;
  assign n413 = 87 & n151;
  assign n414 = 58 & n153;
  assign n415 = ~n412 & ~n413;
  assign n416 = ~n414 & n415;
  assign n417 = ~n159 & ~n416;
  assign n418 = ~77 & n162;
  assign n419 = 77 & ~n313;
  assign n420 = n165 & n419;
  assign n421 = ~n417 & ~n418;
  assign n422 = ~n420 & n421;
  assign n423 = 244 & ~n171;
  assign n424 = ~n319 & n423;
  assign n425 = 33 & 107;
  assign n426 = 232 & n178;
  assign n427 = 238 & n180;
  assign n428 = ~n425 & ~n426;
  assign n429 = ~n427 & n428;
  assign n430 = n171 & ~n429;
  assign n431 = ~n322 & ~n424;
  assign n432 = ~n430 & n431;
  assign n433 = 169 & ~n422;
  assign n434 = ~n432 & n433;
  assign n435 = 179 & ~n422;
  assign n436 = n432 & n435;
  assign n437 = ~n434 & ~n436;
  assign n438 = 190 & n422;
  assign n439 = n432 & n438;
  assign n440 = 200 & n422;
  assign n441 = ~n432 & n440;
  assign n442 = ~n439 & ~n441;
  assign n443 = n422 & n442;
  assign n444 = n437 & ~n443;
  assign n445 = n342 & n378;
  assign n446 = n411 & n445;
  assign n447 = n444 & n446;
  assign 4028 = n305 & n447;
  assign n449 = n198 & ~n229;
  assign n450 = ~n262 & n303;
  assign n451 = n236 & ~n295;
  assign n452 = n269 & n451;
  assign n453 = n198 & n452;
  assign n454 = n191 & ~n449;
  assign n455 = ~n450 & n454;
  assign n456 = ~n453 & n455;
  assign n457 = n447 & ~n456;
  assign n458 = n342 & ~n371;
  assign n459 = ~n404 & n445;
  assign n460 = n378 & ~n437;
  assign n461 = n411 & n460;
  assign n462 = n342 & n461;
  assign n463 = n335 & ~n458;
  assign n464 = ~n459 & n463;
  assign n465 = ~n462 & n464;
  assign 4145 = n457 | ~n465;
  assign n467 = ~\1  & 13;
  assign n468 = ~20 & n467;
  assign n469 = 213 & n468;
  assign n470 = 343 & n469;
  assign n471 = ~n280 & n470;
  assign n472 = ~n302 & n471;
  assign n473 = n302 & ~n471;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n247 & n470;
  assign n476 = ~n269 & n475;
  assign n477 = n269 & ~n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n474 & ~n478;
  assign n480 = ~n262 & ~n470;
  assign n481 = ~n295 & ~n470;
  assign n482 = ~n478 & n481;
  assign n483 = ~n480 & ~n482;
  assign n484 = 330 & n479;
  assign n485 = n483 & n484;
  assign 4589 = ~n483 | n485;
  assign n487 = ~41 & n86;
  assign n488 = n79 & n487;
  assign n489 = ~n186 & ~n224;
  assign n490 = ~n257 & n489;
  assign n491 = ~n290 & n490;
  assign n492 = ~179 & n491;
  assign n493 = n186 & n224;
  assign n494 = n257 & n493;
  assign n495 = n290 & n494;
  assign n496 = 179 & n495;
  assign n497 = ~n492 & ~n496;
  assign n498 = n470 & ~n497;
  assign n499 = n305 & ~n470;
  assign n500 = ~n498 & ~n499;
  assign n501 = ~n456 & ~n470;
  assign n502 = 330 & ~n500;
  assign n503 = ~n501 & n502;
  assign n504 = ~n501 & ~n503;
  assign n505 = ~\1  & ~n504;
  assign n506 = ~116 & n149;
  assign n507 = \1  & ~n487;
  assign n508 = n506 & n507;
  assign n509 = ~n488 & ~n505;
  assign 4667 = n508 | ~n509;
  assign n511 = ~330 & ~n474;
  assign n512 = 330 & n474;
  assign n513 = ~n511 & ~n512;
  assign n514 = 13 & ~20;
  assign n515 = 45 & n514;
  assign n516 = \1  & ~n515;
  assign n517 = ~n513 & ~n516;
  assign n518 = n487 & ~n513;
  assign n519 = 20 & ~190;
  assign n520 = 20 & 200;
  assign n521 = 20 & 179;
  assign n522 = ~n520 & ~n521;
  assign n523 = n519 & n522;
  assign n524 = 159 & n523;
  assign n525 = n520 & ~n521;
  assign n526 = n519 & n525;
  assign n527 = 107 & n526;
  assign n528 = ~n519 & n522;
  assign n529 = 97 & n528;
  assign n530 = ~n519 & n525;
  assign n531 = 87 & n530;
  assign n532 = ~200 & n521;
  assign n533 = n519 & n532;
  assign n534 = 77 & n533;
  assign n535 = 200 & n521;
  assign n536 = n519 & n535;
  assign n537 = 68 & n536;
  assign n538 = ~n519 & n532;
  assign n539 = 58 & n538;
  assign n540 = ~n519 & n535;
  assign n541 = 50 & n540;
  assign n542 = ~n524 & ~n527;
  assign n543 = ~n529 & n542;
  assign n544 = ~n531 & n543;
  assign n545 = ~n534 & n544;
  assign n546 = ~n537 & n545;
  assign n547 = ~n539 & n546;
  assign n548 = ~n541 & n547;
  assign n549 = ~33 & n548;
  assign n550 = 329 & n523;
  assign n551 = 283 & n526;
  assign n552 = 294 & n528;
  assign n553 = 303 & n530;
  assign n554 = 311 & n533;
  assign n555 = 317 & n536;
  assign n556 = 322 & n538;
  assign n557 = 326 & n540;
  assign n558 = ~n550 & ~n551;
  assign n559 = ~n552 & n558;
  assign n560 = ~n553 & n559;
  assign n561 = ~n554 & n560;
  assign n562 = ~n555 & n561;
  assign n563 = ~n556 & n562;
  assign n564 = ~n557 & n563;
  assign n565 = 33 & n564;
  assign n566 = ~n549 & ~n565;
  assign n567 = 20 & ~169;
  assign n568 = n80 & ~n567;
  assign n569 = ~n566 & n568;
  assign n570 = ~13 & ~20;
  assign n571 = ~33 & n570;
  assign n572 = n474 & n571;
  assign n573 = 45 & ~n144;
  assign n574 = ~45 & n79;
  assign n575 = ~n573 & ~n574;
  assign n576 = 33 & n86;
  assign n577 = n575 & n576;
  assign n578 = ~33 & n86;
  assign n579 = 1947 & n578;
  assign n580 = ~n576 & ~n578;
  assign n581 = ~116 & n580;
  assign n582 = ~n577 & ~n579;
  assign n583 = ~n581 & n582;
  assign n584 = ~n568 & ~n571;
  assign n585 = ~n583 & n584;
  assign n586 = ~n569 & ~n572;
  assign n587 = ~n585 & n586;
  assign n588 = ~n487 & n516;
  assign n589 = n587 & n588;
  assign n590 = ~n517 & ~n518;
  assign 4815 = n589 | ~n590;
  assign n592 = ~n422 & n470;
  assign n593 = ~n444 & n592;
  assign n594 = n444 & ~n592;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n501 & ~n595;
  assign n597 = n501 & n595;
  assign n598 = ~n596 & ~n597;
  assign n599 = n502 & n598;
  assign n600 = ~n502 & ~n598;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n516 & ~n601;
  assign n603 = n487 & ~n601;
  assign n604 = 132 & n523;
  assign n605 = 68 & n526;
  assign n606 = 58 & n528;
  assign n607 = 50 & n530;
  assign n608 = 159 & n533;
  assign n609 = 150 & n536;
  assign n610 = 143 & n538;
  assign n611 = 137 & n540;
  assign n612 = ~n604 & ~n605;
  assign n613 = ~n606 & n612;
  assign n614 = ~n607 & n613;
  assign n615 = ~n608 & n614;
  assign n616 = ~n609 & n615;
  assign n617 = ~n610 & n616;
  assign n618 = ~n611 & n617;
  assign n619 = ~33 & n618;
  assign n620 = 311 & n523;
  assign n621 = 87 & n526;
  assign n622 = 107 & n530;
  assign n623 = 116 & n533;
  assign n624 = 283 & n536;
  assign n625 = 294 & n538;
  assign n626 = 303 & n540;
  assign n627 = ~n620 & ~n621;
  assign n628 = ~n529 & n627;
  assign n629 = ~n622 & n628;
  assign n630 = ~n623 & n629;
  assign n631 = ~n624 & n630;
  assign n632 = ~n625 & n631;
  assign n633 = ~n626 & n632;
  assign n634 = 33 & n633;
  assign n635 = ~n619 & ~n634;
  assign n636 = n568 & ~n635;
  assign n637 = ~13 & ~33;
  assign n638 = n595 & n637;
  assign n639 = ~n568 & ~n637;
  assign n640 = ~77 & n639;
  assign n641 = ~n636 & ~n638;
  assign n642 = ~n640 & n641;
  assign n643 = n588 & n642;
  assign n644 = ~n602 & ~n603;
  assign 4944 = n643 | ~n644;
  assign n646 = 77 & ~n345;
  assign n647 = 50 & n646;
  assign n648 = ~50 & 68;
  assign n649 = ~n647 & ~n648;
  assign n650 = n85 & ~n649;
  assign n651 = 116 & ~n201;
  assign n652 = n81 & n651;
  assign n653 = ~n356 & n469;
  assign n654 = ~n378 & n653;
  assign n655 = n378 & ~n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n389 & n470;
  assign n658 = ~n411 & n657;
  assign n659 = n411 & ~n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n500 & ~n656;
  assign n662 = ~n660 & n661;
  assign n663 = ~n595 & n662;
  assign n664 = n447 & ~n500;
  assign n665 = n663 & ~n664;
  assign n666 = ~n663 & n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = 330 & ~n667;
  assign n669 = n447 & n501;
  assign n670 = n465 & ~n669;
  assign n671 = ~n371 & ~n469;
  assign n672 = ~n404 & ~n470;
  assign n673 = ~n656 & n672;
  assign n674 = ~n437 & ~n470;
  assign n675 = ~n656 & ~n660;
  assign n676 = n674 & n675;
  assign n677 = ~n595 & n675;
  assign n678 = n501 & n677;
  assign n679 = ~n671 & ~n673;
  assign n680 = ~n676 & n679;
  assign n681 = ~n678 & n680;
  assign n682 = ~n670 & n681;
  assign n683 = n670 & ~n681;
  assign n684 = ~n682 & ~n683;
  assign n685 = n668 & n684;
  assign n686 = ~n668 & ~n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n81 & ~n85;
  assign n689 = ~n687 & n688;
  assign n690 = ~n650 & ~n652;
  assign 5002 = n689 | ~n690;
  assign n692 = ~n212 & n470;
  assign n693 = ~n236 & n692;
  assign n694 = n236 & ~n692;
  assign n695 = ~n693 & ~n694;
  assign n696 = n479 & ~n695;
  assign n697 = 330 & n696;
  assign n698 = ~n169 & n470;
  assign n699 = ~n198 & n698;
  assign n700 = n198 & ~n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n229 & ~n470;
  assign n703 = n480 & ~n695;
  assign n704 = ~n478 & ~n695;
  assign n705 = n481 & n704;
  assign n706 = ~n702 & ~n703;
  assign n707 = ~n705 & n706;
  assign n708 = ~n701 & n707;
  assign n709 = n701 & ~n707;
  assign n710 = ~n708 & ~n709;
  assign n711 = n697 & n710;
  assign n712 = ~n697 & ~n710;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n516 & ~n713;
  assign n715 = ~n504 & ~n713;
  assign n716 = 330 & ~n474;
  assign n717 = ~n478 & ~n481;
  assign n718 = n478 & n481;
  assign n719 = ~n717 & ~n718;
  assign n720 = n716 & n719;
  assign n721 = ~n716 & ~n719;
  assign n722 = ~n720 & ~n721;
  assign n723 = n483 & ~n695;
  assign n724 = ~n483 & n695;
  assign n725 = ~n723 & ~n724;
  assign n726 = n484 & n725;
  assign n727 = ~n484 & ~n725;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n722 & ~n728;
  assign n730 = ~n713 & n729;
  assign n731 = n504 & n730;
  assign n732 = ~n715 & ~n731;
  assign n733 = n487 & ~n732;
  assign n734 = 137 & n523;
  assign n735 = 77 & n526;
  assign n736 = 68 & n528;
  assign n737 = 58 & n530;
  assign n738 = 50 & n533;
  assign n739 = 159 & n536;
  assign n740 = 150 & n538;
  assign n741 = 143 & n540;
  assign n742 = ~n734 & ~n735;
  assign n743 = ~n736 & n742;
  assign n744 = ~n737 & n743;
  assign n745 = ~n738 & n744;
  assign n746 = ~n739 & n745;
  assign n747 = ~n740 & n746;
  assign n748 = ~n741 & n747;
  assign n749 = ~33 & n748;
  assign n750 = 317 & n523;
  assign n751 = 97 & n526;
  assign n752 = 107 & n528;
  assign n753 = 116 & n530;
  assign n754 = 283 & n533;
  assign n755 = 294 & n536;
  assign n756 = 303 & n538;
  assign n757 = 311 & n540;
  assign n758 = ~n750 & ~n751;
  assign n759 = ~n752 & n758;
  assign n760 = ~n753 & n759;
  assign n761 = ~n754 & n760;
  assign n762 = ~n755 & n761;
  assign n763 = ~n756 & n762;
  assign n764 = ~n757 & n763;
  assign n765 = 33 & n764;
  assign n766 = ~n749 & ~n765;
  assign n767 = n568 & ~n766;
  assign n768 = n571 & n701;
  assign n769 = ~n115 & n576;
  assign n770 = ~87 & n580;
  assign n771 = ~n578 & ~n769;
  assign n772 = ~n770 & n771;
  assign n773 = n584 & ~n772;
  assign n774 = ~n767 & ~n768;
  assign n775 = ~n773 & n774;
  assign n776 = n588 & n775;
  assign n777 = ~n714 & ~n733;
  assign 5045 = n776 | ~n777;
  assign n779 = ~n516 & ~n722;
  assign n780 = n504 & ~n722;
  assign n781 = ~n504 & n722;
  assign n782 = ~n780 & ~n781;
  assign n783 = n487 & n782;
  assign n784 = 150 & n523;
  assign n785 = 87 & n528;
  assign n786 = 77 & n530;
  assign n787 = 68 & n533;
  assign n788 = 58 & n536;
  assign n789 = 50 & n538;
  assign n790 = 159 & n540;
  assign n791 = ~n751 & ~n784;
  assign n792 = ~n785 & n791;
  assign n793 = ~n786 & n792;
  assign n794 = ~n787 & n793;
  assign n795 = ~n788 & n794;
  assign n796 = ~n789 & n795;
  assign n797 = ~n790 & n796;
  assign n798 = ~33 & n797;
  assign n799 = 326 & n523;
  assign n800 = 116 & n526;
  assign n801 = 283 & n528;
  assign n802 = 294 & n530;
  assign n803 = 303 & n533;
  assign n804 = 311 & n536;
  assign n805 = 317 & n538;
  assign n806 = 322 & n540;
  assign n807 = ~n799 & ~n800;
  assign n808 = ~n801 & n807;
  assign n809 = ~n802 & n808;
  assign n810 = ~n803 & n809;
  assign n811 = ~n804 & n810;
  assign n812 = ~n805 & n811;
  assign n813 = ~n806 & n812;
  assign n814 = 33 & n813;
  assign n815 = ~n798 & ~n814;
  assign n816 = n568 & ~n815;
  assign n817 = n478 & n571;
  assign n818 = 45 & n124;
  assign n819 = 68 & 77;
  assign n820 = n506 & ~n819;
  assign n821 = ~50 & n820;
  assign n822 = 58 & n821;
  assign n823 = ~45 & n822;
  assign n824 = ~n818 & ~n823;
  assign n825 = n576 & n824;
  assign n826 = ~n506 & n578;
  assign n827 = ~107 & n580;
  assign n828 = ~n825 & ~n826;
  assign n829 = ~n827 & n828;
  assign n830 = n584 & ~n829;
  assign n831 = ~n816 & ~n817;
  assign n832 = ~n830 & n831;
  assign n833 = n588 & n832;
  assign n834 = ~n779 & ~n783;
  assign 5047 = n833 | ~n834;
  assign n836 = ~n516 & ~n728;
  assign n837 = n728 & n780;
  assign n838 = ~n728 & ~n780;
  assign n839 = ~n837 & ~n838;
  assign n840 = n487 & ~n839;
  assign n841 = 143 & n523;
  assign n842 = 77 & n528;
  assign n843 = 68 & n530;
  assign n844 = 58 & n533;
  assign n845 = 50 & n536;
  assign n846 = 159 & n538;
  assign n847 = 150 & n540;
  assign n848 = ~n621 & ~n841;
  assign n849 = ~n842 & n848;
  assign n850 = ~n843 & n849;
  assign n851 = ~n844 & n850;
  assign n852 = ~n845 & n851;
  assign n853 = ~n846 & n852;
  assign n854 = ~n847 & n853;
  assign n855 = ~33 & n854;
  assign n856 = 322 & n523;
  assign n857 = 116 & n528;
  assign n858 = 283 & n530;
  assign n859 = 294 & n533;
  assign n860 = 303 & n536;
  assign n861 = 311 & n538;
  assign n862 = 317 & n540;
  assign n863 = ~n527 & ~n856;
  assign n864 = ~n857 & n863;
  assign n865 = ~n858 & n864;
  assign n866 = ~n859 & n865;
  assign n867 = ~n860 & n866;
  assign n868 = ~n861 & n867;
  assign n869 = ~n862 & n868;
  assign n870 = 33 & n869;
  assign n871 = ~n855 & ~n870;
  assign n872 = n568 & ~n871;
  assign n873 = n571 & n695;
  assign n874 = ~n136 & n576;
  assign n875 = ~97 & n580;
  assign n876 = ~n578 & ~n874;
  assign n877 = ~n875 & n876;
  assign n878 = n584 & ~n877;
  assign n879 = ~n872 & ~n873;
  assign n880 = ~n878 & n879;
  assign n881 = n588 & n880;
  assign n882 = ~n836 & ~n840;
  assign 5078 = n881 | ~n882;
  assign n884 = ~n500 & ~n595;
  assign n885 = ~n660 & n884;
  assign n886 = 330 & n885;
  assign n887 = ~n660 & n674;
  assign n888 = ~n595 & ~n660;
  assign n889 = n501 & n888;
  assign n890 = ~n672 & ~n887;
  assign n891 = ~n889 & n890;
  assign n892 = ~n656 & n891;
  assign n893 = n656 & ~n891;
  assign n894 = ~n892 & ~n893;
  assign n895 = n886 & n894;
  assign n896 = ~n886 & ~n894;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n516 & ~n897;
  assign n899 = 330 & n884;
  assign n900 = n501 & ~n595;
  assign n901 = ~n674 & ~n900;
  assign n902 = ~n660 & n901;
  assign n903 = n660 & ~n901;
  assign n904 = ~n902 & ~n903;
  assign n905 = n899 & n904;
  assign n906 = ~n899 & ~n904;
  assign n907 = ~n905 & ~n906;
  assign n908 = 330 & n664;
  assign n909 = n670 & n908;
  assign n910 = n670 & ~n909;
  assign n911 = ~n907 & n910;
  assign n912 = n897 & n911;
  assign n913 = ~n897 & ~n911;
  assign n914 = ~n912 & ~n913;
  assign n915 = n487 & ~n914;
  assign n916 = 125 & n523;
  assign n917 = 50 & n526;
  assign n918 = 159 & n528;
  assign n919 = 150 & n530;
  assign n920 = 143 & n533;
  assign n921 = 137 & n536;
  assign n922 = 132 & n538;
  assign n923 = 128 & n540;
  assign n924 = ~n916 & ~n917;
  assign n925 = ~n918 & n924;
  assign n926 = ~n919 & n925;
  assign n927 = ~n920 & n926;
  assign n928 = ~n921 & n927;
  assign n929 = ~n922 & n928;
  assign n930 = ~n923 & n929;
  assign n931 = ~33 & n930;
  assign n932 = 294 & n523;
  assign n933 = 97 & n533;
  assign n934 = 107 & n536;
  assign n935 = 116 & n538;
  assign n936 = 283 & n540;
  assign n937 = ~n605 & ~n932;
  assign n938 = ~n842 & n937;
  assign n939 = ~n531 & n938;
  assign n940 = ~n933 & n939;
  assign n941 = ~n934 & n940;
  assign n942 = ~n935 & n941;
  assign n943 = ~n936 & n942;
  assign n944 = 33 & n943;
  assign n945 = ~n931 & ~n944;
  assign n946 = n568 & ~n945;
  assign n947 = n637 & n656;
  assign n948 = ~58 & n639;
  assign n949 = ~n946 & ~n947;
  assign n950 = ~n948 & n949;
  assign n951 = n588 & n950;
  assign n952 = ~n898 & ~n915;
  assign 5102 = n951 | ~n952;
  assign n954 = 330 & n663;
  assign n955 = ~n317 & n469;
  assign n956 = ~n342 & n955;
  assign n957 = n342 & ~n955;
  assign n958 = ~n956 & ~n957;
  assign n959 = n681 & ~n958;
  assign n960 = ~n681 & n958;
  assign n961 = ~n959 & ~n960;
  assign n962 = n954 & n961;
  assign n963 = ~n954 & ~n961;
  assign n964 = ~n962 & ~n963;
  assign n965 = ~n516 & ~n964;
  assign n966 = ~n910 & ~n964;
  assign n967 = ~n897 & ~n907;
  assign n968 = ~n964 & n967;
  assign n969 = n910 & n968;
  assign n970 = ~n966 & ~n969;
  assign n971 = n487 & ~n970;
  assign n972 = 124 & n523;
  assign n973 = 159 & n526;
  assign n974 = 150 & n528;
  assign n975 = 143 & n530;
  assign n976 = 137 & n533;
  assign n977 = 132 & n536;
  assign n978 = 128 & n538;
  assign n979 = 125 & n540;
  assign n980 = ~n972 & ~n973;
  assign n981 = ~n974 & n980;
  assign n982 = ~n975 & n981;
  assign n983 = ~n976 & n982;
  assign n984 = ~n977 & n983;
  assign n985 = ~n978 & n984;
  assign n986 = ~n979 & n985;
  assign n987 = ~33 & ~41;
  assign n988 = n986 & n987;
  assign n989 = 283 & n523;
  assign n990 = 58 & n526;
  assign n991 = 87 & n533;
  assign n992 = 97 & n536;
  assign n993 = 107 & n538;
  assign n994 = 116 & n540;
  assign n995 = ~n989 & ~n990;
  assign n996 = ~n736 & n995;
  assign n997 = ~n786 & n996;
  assign n998 = ~n991 & n997;
  assign n999 = ~n992 & n998;
  assign n1000 = ~n993 & n999;
  assign n1001 = ~n994 & n1000;
  assign n1002 = 33 & ~41;
  assign n1003 = n1001 & n1002;
  assign n1004 = ~n987 & ~n1002;
  assign n1005 = ~50 & n1004;
  assign n1006 = ~n988 & ~n1003;
  assign n1007 = ~n1005 & n1006;
  assign n1008 = n568 & ~n1007;
  assign n1009 = n637 & n958;
  assign n1010 = ~50 & n639;
  assign n1011 = ~n1008 & ~n1009;
  assign n1012 = ~n1010 & n1011;
  assign n1013 = n588 & n1012;
  assign n1014 = ~n965 & ~n971;
  assign 5120 = n1013 | ~n1014;
  assign n1016 = ~n516 & ~n907;
  assign n1017 = n907 & ~n910;
  assign n1018 = ~n911 & ~n1017;
  assign n1019 = n487 & n1018;
  assign n1020 = 128 & n523;
  assign n1021 = 50 & n528;
  assign n1022 = 159 & n530;
  assign n1023 = 150 & n533;
  assign n1024 = 143 & n536;
  assign n1025 = 137 & n538;
  assign n1026 = 132 & n540;
  assign n1027 = ~n990 & ~n1020;
  assign n1028 = ~n1021 & n1027;
  assign n1029 = ~n1022 & n1028;
  assign n1030 = ~n1023 & n1029;
  assign n1031 = ~n1024 & n1030;
  assign n1032 = ~n1025 & n1031;
  assign n1033 = ~n1026 & n1032;
  assign n1034 = ~33 & n1033;
  assign n1035 = 303 & n523;
  assign n1036 = 97 & n530;
  assign n1037 = 107 & n533;
  assign n1038 = 116 & n536;
  assign n1039 = 283 & n538;
  assign n1040 = 294 & n540;
  assign n1041 = ~n735 & ~n1035;
  assign n1042 = ~n785 & n1041;
  assign n1043 = ~n1036 & n1042;
  assign n1044 = ~n1037 & n1043;
  assign n1045 = ~n1038 & n1044;
  assign n1046 = ~n1039 & n1045;
  assign n1047 = ~n1040 & n1046;
  assign n1048 = 33 & n1047;
  assign n1049 = ~n1034 & ~n1048;
  assign n1050 = n568 & ~n1049;
  assign n1051 = n637 & n660;
  assign n1052 = ~68 & n639;
  assign n1053 = ~n1050 & ~n1051;
  assign n1054 = ~n1052 & n1053;
  assign n1055 = n588 & n1054;
  assign n1056 = ~n1016 & ~n1019;
  assign 5121 = n1055 | ~n1056;
  assign n1058 = ~4815 & ~5047;
  assign n1059 = ~5078 & n1058;
  assign n1060 = ~5045 & n1059;
  assign n1061 = ~4944 & ~5121;
  assign n1062 = ~5102 & n1061;
  assign n1063 = ~5120 & n1062;
  assign 5192 = ~n1060 | ~n1063;
  assign n1065 = 213 & ~343;
  assign n1066 = ~5102 & ~5120;
  assign n1067 = n1065 & n1066;
  assign n1068 = 5192 & ~n1067;
  assign 5231 = ~213 | ~n1068;
  assign n1070 = 5045 & ~5078;
  assign n1071 = ~5045 & 5078;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = ~4815 & 5047;
  assign n1074 = 4815 & ~5047;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = ~n1072 & n1075;
  assign n1077 = n1072 & ~n1075;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~4944 & 5121;
  assign n1080 = 4944 & ~5121;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = 5102 & ~n1065;
  assign n1083 = 5120 & ~n1065;
  assign n1084 = n1082 & ~n1083;
  assign n1085 = ~n1082 & n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = 350 & n1065;
  assign n1088 = ~n1081 & ~n1086;
  assign n1089 = n1087 & n1088;
  assign n1090 = ~n1081 & n1086;
  assign n1091 = ~n1087 & n1090;
  assign n1092 = n1081 & ~n1086;
  assign n1093 = ~n1087 & n1092;
  assign n1094 = n1081 & n1086;
  assign n1095 = n1087 & n1094;
  assign n1096 = ~n1089 & ~n1091;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = ~n1095 & n1097;
  assign n1099 = n1078 & n1098;
  assign n1100 = ~n1078 & ~n1098;
  assign 5360 = n1099 | n1100;
  assign n1102 = ~5102 & 5120;
  assign n1103 = 5102 & ~5120;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = n1081 & ~n1104;
  assign n1106 = ~n1081 & n1104;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = n1078 & ~n1107;
  assign n1109 = ~n1078 & n1107;
  assign 5361 = ~n1108 & ~n1109;
endmodule


