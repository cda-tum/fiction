// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    p_4_1_, p_26_9_, p_130_58_, p_53_19_, p_64_22_, p_67_23_, p_91_35_,
    p_94_36_, p_136_62_, p_173_76_, p_293_112_, p_545_150_, p_2174_161_,
    p_3717_169_, p_25_8_, p_106_40_, p_14_3_, p_52_18_, p_113_43_,
    p_117_47_, p_534_149_, p_24_7_, p_272_105_, p_302_114_, p_4091_175_,
    p_61_21_, p_100_38_, p_170_75_, p_210_89_, p_226_93_, p_373_133_,
    p_23_6_, p_167_74_, p_206_87_, p_400_137_, p_457_142_, p_1694_160_,
    p_4090_174_, p_11_2_, p_123_53_, p_315_117_, p_514_147_, p_1690_158_,
    p_4115_177_, p_109_41_, p_257_102_, p_323_119_, p_435_140_, p_559_154_,
    p_31_11_, p_34_12_, p_114_44_, p_118_48_, p_120_50_, p_176_77_,
    p_324_120_, p_552_152_, p_20_5_, p_40_14_, p_140_64_, p_549_151_,
    p_4092_176_, p_146_67_, p_242_97_, p_374_134_, p_4089_173_, p_203_86_,
    p_254_101_, p_308_116_, p_331_121_, p_37_13_, p_97_37_, p_127_55_,
    p_179_78_, p_468_143_, p_3552_168_, p_4088_172_, p_1_0_, p_182_79_,
    p_200_85_, p_233_94_, p_273_106_, p_490_145_, p_3550_167_, p_17_4_,
    p_137_63_, p_2824_163_, p_4087_171_, p_49_17_, p_70_24_, p_86_32_,
    p_87_33_, p_88_34_, p_217_90_, p_251_100_, p_351_127_, p_358_128_,
    p_369_131_, p_3173_164_, p_145_66_, p_241_96_, p_341_125_, p_348_126_,
    p_411_138_, p_46_16_, p_73_25_, p_83_31_, p_141_65_, p_152_69_,
    p_191_82_, p_234_95_, p_338_124_, p_121_51_, p_158_71_, p_248_99_,
    p_264_103_, p_361_129_, p_389_136_, p_446_141_, p_43_15_, p_76_26_,
    p_164_73_, p_556_153_, p_3548_166_, p_280_107_, p_82_30_, p_307_115_,
    p_335_123_, p_115_45_, p_128_56_, p_149_68_, p_245_98_, p_386_135_,
    p_3546_165_, p_131_59_, p_209_88_, p_218_91_, p_422_139_, p_1497_156_,
    p_1689_157_, p_27_10_, p_103_39_, p_112_42_, p_116_46_, p_122_52_,
    p_185_80_, p_265_104_, p_562_155_, p_1691_159_, p_79_27_, p_197_84_,
    p_299_113_, p_332_122_, p_503_146_, p_126_54_, p_135_61_, p_292_111_,
    p_194_83_, p_289_110_, p_366_130_, p_479_144_, p_2358_162_, p_80_28_,
    p_129_57_, p_188_81_, p_316_118_, p_54_20_, p_161_72_, p_523_148_,
    p_81_29_, p_119_49_, p_132_60_, p_155_70_, p_225_92_, p_281_108_,
    p_288_109_, p_372_132_, p_3724_170_,
    p_591_1894_, p_604_223_, p_664_2223_, p_690_2484_, p_699_2227_,
    p_618_1925_, p_588_1696_, p_615_1750_, p_688_2317_, p_704_1281_,
    p_818_2273_, p_869_2181_, p_973_202_, p_593_733_, p_600_259_,
    p_611_275_, p_648_2295_, p_822_1933_, p_757_2190_, p_722_2131_,
    p_802_2183_, p_1000_2168_, p_606_407_, p_682_2296_, p_792_2188_,
    p_838_2064_, p_603_225_, p_921_664_, p_629_1926_, p_892_408_,
    p_949_852_, p_612_263_, p_772_2299_, p_797_2191_, p_661_2178_,
    p_727_2298_, p_849_219_, p_939_853_, p_598_1623_, p_634_665_,
    p_636_1280_, p_742_2238_, p_767_2479_, p_836_2128_, p_693_2179_,
    p_702_2228_, p_807_2480_, p_594_224_, p_654_2315_, p_658_2483_,
    p_820_1283_, p_861_2070_, p_875_2125_, p_978_851_, p_685_2316_,
    p_815_627_, p_834_2123_, p_882_2456_, p_926_624_, p_621_1893_,
    p_676_2229_, p_667_2224_, p_696_2226_, p_787_2186_, p_877_2126_,
    p_1002_1920_, p_1004_1977_, p_670_2225_, p_712_2297_, p_298_299_,
    p_715_1278_, p_809_655_, p_843_2455_, p_867_2237_, p_602_222_,
    p_859_2132_, p_863_2276_, p_623_2152_, p_810_356_, p_642_2222_,
    p_777_2278_, p_830_2182_, p_626_1752_, p_632_1692_, p_645_2271_,
    p_679_2272_, p_707_1277_, p_737_2279_, p_782_2239_, p_850_217_,
    p_717_1282_, p_747_2187_, p_826_2275_, p_845_845_, p_871_2127_,
    p_585_2236_, p_865_2277_, p_673_1276_, p_887_528_, p_923_619_,
    p_144_354_, p_732_2300_, p_854_2268_, p_873_2124_, p_889_734_,
    p_599_269_, p_752_2189_, p_610_1519_, p_824_2274_, p_851_218_,
    p_813_2260_, p_832_2133_, p_848_330_, p_993_850_, p_575_2240_,
    p_601_220_, p_639_1275_, p_651_2314_, p_656_621_, p_762_2184_,
    p_828_2233_, p_847_465_, p_998_2163_  );
  input  p_4_1_, p_26_9_, p_130_58_, p_53_19_, p_64_22_, p_67_23_,
    p_91_35_, p_94_36_, p_136_62_, p_173_76_, p_293_112_, p_545_150_,
    p_2174_161_, p_3717_169_, p_25_8_, p_106_40_, p_14_3_, p_52_18_,
    p_113_43_, p_117_47_, p_534_149_, p_24_7_, p_272_105_, p_302_114_,
    p_4091_175_, p_61_21_, p_100_38_, p_170_75_, p_210_89_, p_226_93_,
    p_373_133_, p_23_6_, p_167_74_, p_206_87_, p_400_137_, p_457_142_,
    p_1694_160_, p_4090_174_, p_11_2_, p_123_53_, p_315_117_, p_514_147_,
    p_1690_158_, p_4115_177_, p_109_41_, p_257_102_, p_323_119_,
    p_435_140_, p_559_154_, p_31_11_, p_34_12_, p_114_44_, p_118_48_,
    p_120_50_, p_176_77_, p_324_120_, p_552_152_, p_20_5_, p_40_14_,
    p_140_64_, p_549_151_, p_4092_176_, p_146_67_, p_242_97_, p_374_134_,
    p_4089_173_, p_203_86_, p_254_101_, p_308_116_, p_331_121_, p_37_13_,
    p_97_37_, p_127_55_, p_179_78_, p_468_143_, p_3552_168_, p_4088_172_,
    p_1_0_, p_182_79_, p_200_85_, p_233_94_, p_273_106_, p_490_145_,
    p_3550_167_, p_17_4_, p_137_63_, p_2824_163_, p_4087_171_, p_49_17_,
    p_70_24_, p_86_32_, p_87_33_, p_88_34_, p_217_90_, p_251_100_,
    p_351_127_, p_358_128_, p_369_131_, p_3173_164_, p_145_66_, p_241_96_,
    p_341_125_, p_348_126_, p_411_138_, p_46_16_, p_73_25_, p_83_31_,
    p_141_65_, p_152_69_, p_191_82_, p_234_95_, p_338_124_, p_121_51_,
    p_158_71_, p_248_99_, p_264_103_, p_361_129_, p_389_136_, p_446_141_,
    p_43_15_, p_76_26_, p_164_73_, p_556_153_, p_3548_166_, p_280_107_,
    p_82_30_, p_307_115_, p_335_123_, p_115_45_, p_128_56_, p_149_68_,
    p_245_98_, p_386_135_, p_3546_165_, p_131_59_, p_209_88_, p_218_91_,
    p_422_139_, p_1497_156_, p_1689_157_, p_27_10_, p_103_39_, p_112_42_,
    p_116_46_, p_122_52_, p_185_80_, p_265_104_, p_562_155_, p_1691_159_,
    p_79_27_, p_197_84_, p_299_113_, p_332_122_, p_503_146_, p_126_54_,
    p_135_61_, p_292_111_, p_194_83_, p_289_110_, p_366_130_, p_479_144_,
    p_2358_162_, p_80_28_, p_129_57_, p_188_81_, p_316_118_, p_54_20_,
    p_161_72_, p_523_148_, p_81_29_, p_119_49_, p_132_60_, p_155_70_,
    p_225_92_, p_281_108_, p_288_109_, p_372_132_, p_3724_170_;
  output p_591_1894_, p_604_223_, p_664_2223_, p_690_2484_, p_699_2227_,
    p_618_1925_, p_588_1696_, p_615_1750_, p_688_2317_, p_704_1281_,
    p_818_2273_, p_869_2181_, p_973_202_, p_593_733_, p_600_259_,
    p_611_275_, p_648_2295_, p_822_1933_, p_757_2190_, p_722_2131_,
    p_802_2183_, p_1000_2168_, p_606_407_, p_682_2296_, p_792_2188_,
    p_838_2064_, p_603_225_, p_921_664_, p_629_1926_, p_892_408_,
    p_949_852_, p_612_263_, p_772_2299_, p_797_2191_, p_661_2178_,
    p_727_2298_, p_849_219_, p_939_853_, p_598_1623_, p_634_665_,
    p_636_1280_, p_742_2238_, p_767_2479_, p_836_2128_, p_693_2179_,
    p_702_2228_, p_807_2480_, p_594_224_, p_654_2315_, p_658_2483_,
    p_820_1283_, p_861_2070_, p_875_2125_, p_978_851_, p_685_2316_,
    p_815_627_, p_834_2123_, p_882_2456_, p_926_624_, p_621_1893_,
    p_676_2229_, p_667_2224_, p_696_2226_, p_787_2186_, p_877_2126_,
    p_1002_1920_, p_1004_1977_, p_670_2225_, p_712_2297_, p_298_299_,
    p_715_1278_, p_809_655_, p_843_2455_, p_867_2237_, p_602_222_,
    p_859_2132_, p_863_2276_, p_623_2152_, p_810_356_, p_642_2222_,
    p_777_2278_, p_830_2182_, p_626_1752_, p_632_1692_, p_645_2271_,
    p_679_2272_, p_707_1277_, p_737_2279_, p_782_2239_, p_850_217_,
    p_717_1282_, p_747_2187_, p_826_2275_, p_845_845_, p_871_2127_,
    p_585_2236_, p_865_2277_, p_673_1276_, p_887_528_, p_923_619_,
    p_144_354_, p_732_2300_, p_854_2268_, p_873_2124_, p_889_734_,
    p_599_269_, p_752_2189_, p_610_1519_, p_824_2274_, p_851_218_,
    p_813_2260_, p_832_2133_, p_848_330_, p_993_850_, p_575_2240_,
    p_601_220_, p_639_1275_, p_651_2314_, p_656_621_, p_762_2184_,
    p_828_2233_, p_847_465_, p_998_2163_;
  wire new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1378,
    new_n1380, new_n1381, new_n1382, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1433, new_n1434, new_n1435, new_n1437, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1477, new_n1478, new_n1479,
    new_n1481, new_n1482, new_n1483, new_n1484, new_n1485, new_n1486,
    new_n1487, new_n1488, new_n1489, new_n1490, new_n1492, new_n1493,
    new_n1494, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1526, new_n1527, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1539, new_n1540, new_n1542,
    new_n1543, new_n1544, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1611, new_n1612, new_n1613, new_n1614, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1639, new_n1640, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1731, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1855, new_n1856, new_n1857, new_n1858,
    new_n1859, new_n1860, new_n1861, new_n1862, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1879,
    new_n1880, new_n1881, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1896, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912;
  assign new_n302 = p_264_103_ & p_335_123_;
  assign new_n303 = p_257_102_ & ~p_335_123_;
  assign new_n304 = ~new_n302 & ~new_n303;
  assign new_n305 = p_389_136_ & new_n304;
  assign new_n306 = ~p_389_136_ & ~new_n304;
  assign new_n307 = ~new_n305 & ~new_n306;
  assign new_n308 = p_241_96_ & p_335_123_;
  assign new_n309 = p_234_95_ & ~p_335_123_;
  assign new_n310 = ~new_n308 & ~new_n309;
  assign new_n311 = p_435_140_ & new_n310;
  assign new_n312 = ~p_435_140_ & ~new_n310;
  assign new_n313 = ~new_n311 & ~new_n312;
  assign new_n314 = p_280_107_ & p_335_123_;
  assign new_n315 = p_273_106_ & ~p_335_123_;
  assign new_n316 = ~new_n314 & ~new_n315;
  assign new_n317 = p_411_138_ & ~new_n316;
  assign new_n318 = p_272_105_ & p_335_123_;
  assign new_n319 = ~p_335_123_ & p_265_104_;
  assign new_n320 = ~new_n318 & ~new_n319;
  assign new_n321 = p_400_137_ & new_n320;
  assign new_n322 = ~p_400_137_ & ~new_n320;
  assign new_n323 = ~new_n321 & ~new_n322;
  assign new_n324 = ~new_n307 & ~new_n313;
  assign new_n325 = new_n317 & new_n324;
  assign new_n326 = ~new_n323 & new_n325;
  assign new_n327 = p_335_123_ & p_288_109_;
  assign new_n328 = ~p_335_123_ & p_281_108_;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = p_374_134_ & ~new_n329;
  assign new_n331 = p_411_138_ & new_n316;
  assign new_n332 = ~p_411_138_ & ~new_n316;
  assign new_n333 = ~new_n331 & ~new_n332;
  assign new_n334 = ~new_n307 & new_n330;
  assign new_n335 = ~new_n323 & new_n334;
  assign new_n336 = ~new_n313 & new_n335;
  assign new_n337 = ~new_n333 & new_n336;
  assign new_n338 = p_389_136_ & ~new_n304;
  assign new_n339 = ~new_n313 & new_n338;
  assign new_n340 = p_400_137_ & ~new_n320;
  assign new_n341 = ~new_n313 & new_n340;
  assign new_n342 = ~new_n307 & new_n341;
  assign new_n343 = p_435_140_ & ~new_n310;
  assign new_n344 = ~new_n326 & ~new_n337;
  assign new_n345 = ~new_n339 & new_n344;
  assign new_n346 = ~new_n342 & new_n345;
  assign new_n347 = ~new_n343 & new_n346;
  assign new_n348 = p_335_123_ & p_209_88_;
  assign new_n349 = p_206_87_ & ~p_335_123_;
  assign new_n350 = ~new_n348 & ~new_n349;
  assign new_n351 = p_446_141_ & new_n350;
  assign new_n352 = ~p_446_141_ & ~new_n350;
  assign new_n353 = ~new_n351 & ~new_n352;
  assign new_n354 = p_335_123_ & p_225_92_;
  assign new_n355 = ~p_335_123_ & p_218_91_;
  assign new_n356 = ~new_n354 & ~new_n355;
  assign new_n357 = p_468_143_ & new_n356;
  assign new_n358 = ~p_468_143_ & ~new_n356;
  assign new_n359 = ~new_n357 & ~new_n358;
  assign new_n360 = p_217_90_ & p_335_123_;
  assign new_n361 = p_210_89_ & ~p_335_123_;
  assign new_n362 = ~new_n360 & ~new_n361;
  assign new_n363 = p_457_142_ & new_n362;
  assign new_n364 = ~p_457_142_ & ~new_n362;
  assign new_n365 = ~new_n363 & ~new_n364;
  assign new_n366 = p_233_94_ & p_335_123_;
  assign new_n367 = p_226_93_ & ~p_335_123_;
  assign new_n368 = ~new_n366 & ~new_n367;
  assign new_n369 = p_422_139_ & new_n368;
  assign new_n370 = ~p_422_139_ & ~new_n368;
  assign new_n371 = ~new_n369 & ~new_n370;
  assign new_n372 = ~new_n353 & ~new_n359;
  assign new_n373 = ~new_n365 & new_n372;
  assign new_n374 = ~new_n371 & new_n373;
  assign new_n375 = ~new_n347 & new_n374;
  assign new_n376 = p_422_139_ & ~new_n368;
  assign new_n377 = ~new_n353 & ~new_n365;
  assign new_n378 = new_n376 & new_n377;
  assign new_n379 = ~new_n359 & new_n378;
  assign new_n380 = p_457_142_ & ~new_n362;
  assign new_n381 = ~new_n353 & new_n380;
  assign new_n382 = p_468_143_ & ~new_n356;
  assign new_n383 = ~new_n353 & new_n382;
  assign new_n384 = ~new_n365 & new_n383;
  assign new_n385 = p_446_141_ & ~new_n350;
  assign new_n386 = ~new_n379 & ~new_n381;
  assign new_n387 = ~new_n384 & new_n386;
  assign new_n388 = ~new_n385 & new_n387;
  assign p_591_1894_ = new_n375 | ~new_n388;
  assign new_n390 = p_1690_158_ & p_1689_157_;
  assign new_n391 = p_158_71_ & new_n390;
  assign new_n392 = ~p_374_134_ & ~new_n329;
  assign new_n393 = p_374_134_ & new_n329;
  assign new_n394 = ~new_n392 & ~new_n393;
  assign new_n395 = p_4_1_ & ~new_n394;
  assign new_n396 = ~new_n330 & ~new_n395;
  assign new_n397 = new_n333 & ~new_n396;
  assign new_n398 = ~new_n333 & new_n396;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = p_4091_175_ & ~p_4092_176_;
  assign new_n401 = ~new_n399 & new_n400;
  assign new_n402 = ~p_4091_175_ & p_4092_176_;
  assign new_n403 = p_126_54_ & new_n402;
  assign new_n404 = ~p_273_106_ & ~p_3548_166_;
  assign new_n405 = p_273_106_ & ~p_3546_165_;
  assign new_n406 = ~p_411_138_ & ~new_n404;
  assign new_n407 = ~new_n405 & new_n406;
  assign new_n408 = ~p_273_106_ & ~p_3550_167_;
  assign new_n409 = p_411_138_ & new_n408;
  assign new_n410 = p_273_106_ & p_411_138_;
  assign new_n411 = ~p_3552_168_ & new_n410;
  assign new_n412 = ~new_n409 & ~new_n411;
  assign new_n413 = ~new_n407 & new_n412;
  assign new_n414 = ~p_4091_175_ & ~p_4092_176_;
  assign new_n415 = new_n413 & new_n414;
  assign new_n416 = ~new_n401 & ~new_n403;
  assign p_877_2126_ = ~new_n415 & new_n416;
  assign new_n418 = ~p_1690_158_ & p_1689_157_;
  assign new_n419 = ~p_877_2126_ & new_n418;
  assign new_n420 = p_1690_158_ & ~p_1689_157_;
  assign new_n421 = p_188_81_ & new_n420;
  assign new_n422 = p_358_128_ & p_332_122_;
  assign new_n423 = p_351_127_ & ~p_332_122_;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = ~p_534_149_ & ~new_n424;
  assign new_n426 = p_534_149_ & new_n424;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = p_332_122_ & p_366_130_;
  assign new_n429 = p_361_129_ & ~p_332_122_;
  assign new_n430 = ~new_n428 & ~new_n429;
  assign new_n431 = p_54_20_ & new_n430;
  assign new_n432 = new_n430 & ~new_n431;
  assign new_n433 = new_n427 & ~new_n432;
  assign new_n434 = ~new_n427 & new_n432;
  assign new_n435 = ~new_n433 & ~new_n434;
  assign new_n436 = new_n400 & ~new_n435;
  assign new_n437 = p_129_57_ & new_n402;
  assign new_n438 = ~p_351_127_ & ~p_3548_166_;
  assign new_n439 = p_351_127_ & ~p_3546_165_;
  assign new_n440 = ~p_534_149_ & ~new_n438;
  assign new_n441 = ~new_n439 & new_n440;
  assign new_n442 = ~p_3550_167_ & ~p_351_127_;
  assign new_n443 = p_534_149_ & new_n442;
  assign new_n444 = p_534_149_ & p_351_127_;
  assign new_n445 = ~p_3552_168_ & new_n444;
  assign new_n446 = ~new_n443 & ~new_n445;
  assign new_n447 = ~new_n441 & new_n446;
  assign new_n448 = new_n414 & new_n447;
  assign new_n449 = ~new_n436 & ~new_n437;
  assign p_838_2064_ = ~new_n448 & new_n449;
  assign new_n451 = ~p_1690_158_ & ~p_1689_157_;
  assign new_n452 = ~p_838_2064_ & new_n451;
  assign new_n453 = ~new_n391 & ~new_n419;
  assign new_n454 = ~new_n421 & new_n453;
  assign new_n455 = ~new_n452 & new_n454;
  assign p_664_2223_ = p_137_63_ & ~new_n455;
  assign new_n457 = p_1694_160_ & p_1691_159_;
  assign new_n458 = p_179_78_ & new_n457;
  assign new_n459 = p_4092_176_ & p_97_37_;
  assign new_n460 = ~new_n307 & ~new_n323;
  assign new_n461 = new_n330 & new_n460;
  assign new_n462 = ~new_n333 & new_n461;
  assign new_n463 = ~new_n323 & ~new_n333;
  assign new_n464 = ~new_n307 & new_n463;
  assign new_n465 = ~new_n394 & new_n464;
  assign new_n466 = ~new_n307 & new_n340;
  assign new_n467 = ~new_n307 & new_n317;
  assign new_n468 = ~new_n323 & new_n467;
  assign new_n469 = ~new_n462 & ~new_n465;
  assign new_n470 = ~new_n466 & new_n469;
  assign new_n471 = ~new_n468 & new_n470;
  assign new_n472 = ~new_n338 & new_n471;
  assign new_n473 = ~new_n333 & ~new_n394;
  assign new_n474 = new_n330 & ~new_n333;
  assign new_n475 = ~new_n317 & ~new_n474;
  assign new_n476 = ~new_n473 & new_n475;
  assign new_n477 = ~new_n394 & new_n463;
  assign new_n478 = new_n317 & ~new_n323;
  assign new_n479 = ~new_n323 & new_n330;
  assign new_n480 = ~new_n333 & new_n479;
  assign new_n481 = ~new_n477 & ~new_n478;
  assign new_n482 = ~new_n480 & new_n481;
  assign new_n483 = ~new_n340 & new_n482;
  assign new_n484 = ~p_374_134_ & new_n329;
  assign new_n485 = new_n483 & new_n484;
  assign new_n486 = ~new_n483 & ~new_n484;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = new_n476 & ~new_n487;
  assign new_n489 = ~new_n476 & new_n487;
  assign new_n490 = ~new_n488 & ~new_n489;
  assign new_n491 = new_n472 & ~new_n490;
  assign new_n492 = ~new_n472 & new_n490;
  assign new_n493 = ~new_n491 & ~new_n492;
  assign new_n494 = new_n394 & ~new_n493;
  assign new_n495 = ~new_n394 & new_n493;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = new_n333 & ~new_n496;
  assign new_n498 = ~new_n333 & new_n496;
  assign new_n499 = ~new_n497 & ~new_n498;
  assign new_n500 = new_n313 & ~new_n499;
  assign new_n501 = ~new_n313 & new_n499;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = new_n323 & ~new_n502;
  assign new_n504 = ~new_n323 & new_n502;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = new_n307 & ~new_n505;
  assign new_n507 = ~new_n307 & new_n505;
  assign new_n508 = ~new_n506 & ~new_n507;
  assign new_n509 = p_1497_156_ & ~new_n508;
  assign new_n510 = ~new_n462 & ~new_n466;
  assign new_n511 = ~new_n468 & new_n510;
  assign new_n512 = ~new_n338 & new_n511;
  assign new_n513 = ~new_n478 & ~new_n480;
  assign new_n514 = ~new_n340 & new_n513;
  assign new_n515 = new_n330 & ~new_n514;
  assign new_n516 = ~new_n330 & new_n514;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = ~new_n475 & ~new_n517;
  assign new_n519 = new_n475 & new_n517;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = ~new_n512 & ~new_n520;
  assign new_n522 = new_n512 & new_n520;
  assign new_n523 = ~new_n521 & ~new_n522;
  assign new_n524 = new_n394 & ~new_n523;
  assign new_n525 = ~new_n394 & new_n523;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = new_n333 & ~new_n526;
  assign new_n528 = ~new_n333 & new_n526;
  assign new_n529 = ~new_n527 & ~new_n528;
  assign new_n530 = new_n313 & ~new_n529;
  assign new_n531 = ~new_n313 & new_n529;
  assign new_n532 = ~new_n530 & ~new_n531;
  assign new_n533 = new_n323 & ~new_n532;
  assign new_n534 = ~new_n323 & new_n532;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536 = new_n307 & ~new_n535;
  assign new_n537 = ~new_n307 & new_n535;
  assign new_n538 = ~new_n536 & ~new_n537;
  assign new_n539 = ~p_1497_156_ & new_n538;
  assign new_n540 = ~new_n509 & ~new_n539;
  assign new_n541 = new_n324 & ~new_n333;
  assign new_n542 = ~new_n323 & new_n541;
  assign new_n543 = ~new_n394 & new_n542;
  assign new_n544 = new_n347 & ~new_n543;
  assign new_n545 = ~new_n359 & ~new_n365;
  assign new_n546 = ~new_n371 & new_n545;
  assign new_n547 = ~new_n365 & new_n382;
  assign new_n548 = ~new_n365 & new_n376;
  assign new_n549 = ~new_n359 & new_n548;
  assign new_n550 = ~new_n546 & ~new_n547;
  assign new_n551 = ~new_n549 & new_n550;
  assign new_n552 = ~new_n380 & new_n551;
  assign new_n553 = ~new_n359 & ~new_n371;
  assign new_n554 = ~new_n359 & new_n376;
  assign new_n555 = ~new_n382 & ~new_n554;
  assign new_n556 = ~new_n553 & new_n555;
  assign new_n557 = ~p_422_139_ & new_n368;
  assign new_n558 = new_n556 & new_n557;
  assign new_n559 = ~new_n556 & ~new_n557;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = new_n552 & ~new_n560;
  assign new_n562 = ~new_n552 & new_n560;
  assign new_n563 = ~new_n561 & ~new_n562;
  assign new_n564 = new_n371 & ~new_n563;
  assign new_n565 = ~new_n371 & new_n563;
  assign new_n566 = ~new_n564 & ~new_n565;
  assign new_n567 = new_n359 & ~new_n566;
  assign new_n568 = ~new_n359 & new_n566;
  assign new_n569 = ~new_n567 & ~new_n568;
  assign new_n570 = new_n353 & ~new_n569;
  assign new_n571 = ~new_n353 & new_n569;
  assign new_n572 = ~new_n570 & ~new_n571;
  assign new_n573 = new_n365 & ~new_n572;
  assign new_n574 = ~new_n365 & new_n572;
  assign new_n575 = ~new_n573 & ~new_n574;
  assign new_n576 = p_1497_156_ & ~new_n544;
  assign new_n577 = ~new_n575 & new_n576;
  assign new_n578 = ~p_1497_156_ & ~new_n347;
  assign new_n579 = ~new_n575 & new_n578;
  assign new_n580 = ~new_n547 & ~new_n549;
  assign new_n581 = ~new_n380 & new_n580;
  assign new_n582 = new_n376 & ~new_n555;
  assign new_n583 = ~new_n376 & new_n555;
  assign new_n584 = ~new_n582 & ~new_n583;
  assign new_n585 = ~new_n581 & ~new_n584;
  assign new_n586 = new_n581 & new_n584;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = new_n371 & ~new_n587;
  assign new_n589 = ~new_n371 & new_n587;
  assign new_n590 = ~new_n588 & ~new_n589;
  assign new_n591 = new_n359 & ~new_n590;
  assign new_n592 = ~new_n359 & new_n590;
  assign new_n593 = ~new_n591 & ~new_n592;
  assign new_n594 = new_n353 & ~new_n593;
  assign new_n595 = ~new_n353 & new_n593;
  assign new_n596 = ~new_n594 & ~new_n595;
  assign new_n597 = new_n365 & ~new_n596;
  assign new_n598 = ~new_n365 & new_n596;
  assign new_n599 = ~new_n597 & ~new_n598;
  assign new_n600 = p_1497_156_ & new_n544;
  assign new_n601 = ~new_n599 & new_n600;
  assign new_n602 = ~p_1497_156_ & new_n347;
  assign new_n603 = ~new_n599 & new_n602;
  assign new_n604 = ~new_n577 & ~new_n579;
  assign new_n605 = ~new_n601 & new_n604;
  assign new_n606 = ~new_n603 & new_n605;
  assign new_n607 = new_n540 & ~new_n606;
  assign new_n608 = ~new_n540 & new_n606;
  assign new_n609 = ~new_n607 & ~new_n608;
  assign new_n610 = p_4091_175_ & new_n609;
  assign new_n611 = ~p_226_93_ & p_254_101_;
  assign new_n612 = p_226_93_ & p_242_97_;
  assign new_n613 = ~p_422_139_ & ~new_n611;
  assign new_n614 = ~new_n612 & new_n613;
  assign new_n615 = ~p_226_93_ & p_251_100_;
  assign new_n616 = p_422_139_ & new_n615;
  assign new_n617 = p_226_93_ & p_422_139_;
  assign new_n618 = p_248_99_ & new_n617;
  assign new_n619 = ~new_n616 & ~new_n618;
  assign new_n620 = ~new_n614 & new_n619;
  assign new_n621 = p_254_101_ & ~p_218_91_;
  assign new_n622 = p_242_97_ & p_218_91_;
  assign new_n623 = ~p_468_143_ & ~new_n621;
  assign new_n624 = ~new_n622 & new_n623;
  assign new_n625 = p_251_100_ & ~p_218_91_;
  assign new_n626 = p_468_143_ & new_n625;
  assign new_n627 = p_468_143_ & p_218_91_;
  assign new_n628 = p_248_99_ & new_n627;
  assign new_n629 = ~new_n626 & ~new_n628;
  assign new_n630 = ~new_n624 & new_n629;
  assign new_n631 = ~new_n620 & new_n630;
  assign new_n632 = new_n620 & ~new_n630;
  assign new_n633 = ~new_n631 & ~new_n632;
  assign new_n634 = ~p_210_89_ & p_254_101_;
  assign new_n635 = p_210_89_ & p_242_97_;
  assign new_n636 = ~p_457_142_ & ~new_n634;
  assign new_n637 = ~new_n635 & new_n636;
  assign new_n638 = ~p_210_89_ & p_251_100_;
  assign new_n639 = p_457_142_ & new_n638;
  assign new_n640 = p_210_89_ & p_457_142_;
  assign new_n641 = p_248_99_ & new_n640;
  assign new_n642 = ~new_n639 & ~new_n641;
  assign new_n643 = ~new_n637 & new_n642;
  assign new_n644 = ~p_206_87_ & p_254_101_;
  assign new_n645 = p_206_87_ & p_242_97_;
  assign new_n646 = ~p_446_141_ & ~new_n644;
  assign new_n647 = ~new_n645 & new_n646;
  assign new_n648 = ~p_206_87_ & p_251_100_;
  assign new_n649 = p_446_141_ & new_n648;
  assign new_n650 = p_206_87_ & p_446_141_;
  assign new_n651 = p_248_99_ & new_n650;
  assign new_n652 = ~new_n649 & ~new_n651;
  assign new_n653 = ~new_n647 & new_n652;
  assign new_n654 = ~new_n643 & new_n653;
  assign new_n655 = new_n643 & ~new_n653;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = new_n633 & ~new_n656;
  assign new_n658 = ~new_n633 & new_n656;
  assign new_n659 = ~new_n657 & ~new_n658;
  assign new_n660 = p_254_101_ & ~p_281_108_;
  assign new_n661 = p_242_97_ & p_281_108_;
  assign new_n662 = ~p_374_134_ & ~new_n660;
  assign new_n663 = ~new_n661 & new_n662;
  assign new_n664 = p_251_100_ & ~p_281_108_;
  assign new_n665 = p_374_134_ & new_n664;
  assign new_n666 = p_374_134_ & p_281_108_;
  assign new_n667 = p_248_99_ & new_n666;
  assign new_n668 = ~new_n665 & ~new_n667;
  assign new_n669 = ~new_n663 & new_n668;
  assign new_n670 = ~p_257_102_ & p_254_101_;
  assign new_n671 = p_257_102_ & p_242_97_;
  assign new_n672 = ~p_389_136_ & ~new_n670;
  assign new_n673 = ~new_n671 & new_n672;
  assign new_n674 = ~p_257_102_ & p_251_100_;
  assign new_n675 = p_389_136_ & new_n674;
  assign new_n676 = p_257_102_ & p_389_136_;
  assign new_n677 = p_248_99_ & new_n676;
  assign new_n678 = ~new_n675 & ~new_n677;
  assign new_n679 = ~new_n673 & new_n678;
  assign new_n680 = p_254_101_ & ~p_234_95_;
  assign new_n681 = p_242_97_ & p_234_95_;
  assign new_n682 = ~p_435_140_ & ~new_n680;
  assign new_n683 = ~new_n681 & new_n682;
  assign new_n684 = p_251_100_ & ~p_234_95_;
  assign new_n685 = p_435_140_ & new_n684;
  assign new_n686 = p_435_140_ & p_234_95_;
  assign new_n687 = p_248_99_ & new_n686;
  assign new_n688 = ~new_n685 & ~new_n687;
  assign new_n689 = ~new_n683 & new_n688;
  assign new_n690 = ~new_n679 & new_n689;
  assign new_n691 = new_n679 & ~new_n689;
  assign new_n692 = ~new_n690 & ~new_n691;
  assign new_n693 = p_254_101_ & ~p_273_106_;
  assign new_n694 = p_242_97_ & p_273_106_;
  assign new_n695 = ~p_411_138_ & ~new_n693;
  assign new_n696 = ~new_n694 & new_n695;
  assign new_n697 = ~p_273_106_ & p_251_100_;
  assign new_n698 = p_411_138_ & new_n697;
  assign new_n699 = p_248_99_ & new_n410;
  assign new_n700 = ~new_n698 & ~new_n699;
  assign new_n701 = ~new_n696 & new_n700;
  assign new_n702 = p_254_101_ & ~p_265_104_;
  assign new_n703 = p_242_97_ & p_265_104_;
  assign new_n704 = ~p_400_137_ & ~new_n702;
  assign new_n705 = ~new_n703 & new_n704;
  assign new_n706 = p_251_100_ & ~p_265_104_;
  assign new_n707 = p_400_137_ & new_n706;
  assign new_n708 = p_400_137_ & p_265_104_;
  assign new_n709 = p_248_99_ & new_n708;
  assign new_n710 = ~new_n707 & ~new_n709;
  assign new_n711 = ~new_n705 & new_n710;
  assign new_n712 = ~new_n701 & new_n711;
  assign new_n713 = new_n701 & ~new_n711;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = ~new_n669 & ~new_n692;
  assign new_n716 = ~new_n714 & new_n715;
  assign new_n717 = new_n692 & ~new_n714;
  assign new_n718 = new_n669 & new_n717;
  assign new_n719 = ~new_n716 & ~new_n718;
  assign new_n720 = new_n669 & ~new_n692;
  assign new_n721 = new_n714 & new_n720;
  assign new_n722 = new_n692 & new_n714;
  assign new_n723 = ~new_n669 & new_n722;
  assign new_n724 = ~new_n721 & ~new_n723;
  assign new_n725 = new_n719 & new_n724;
  assign new_n726 = new_n659 & ~new_n725;
  assign new_n727 = ~new_n659 & new_n725;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = ~p_4091_175_ & ~new_n728;
  assign new_n730 = ~new_n610 & ~new_n729;
  assign new_n731 = ~p_4092_176_ & ~new_n730;
  assign new_n732 = ~new_n459 & ~new_n731;
  assign new_n733 = ~p_1694_160_ & p_1691_159_;
  assign new_n734 = ~new_n732 & new_n733;
  assign new_n735 = p_1694_160_ & ~p_1691_159_;
  assign new_n736 = p_176_77_ & new_n735;
  assign new_n737 = p_94_36_ & p_4092_176_;
  assign new_n738 = p_338_124_ & p_332_122_;
  assign new_n739 = p_332_122_ & ~new_n738;
  assign new_n740 = p_514_147_ & new_n739;
  assign new_n741 = ~p_514_147_ & ~new_n739;
  assign new_n742 = ~new_n740 & ~new_n741;
  assign new_n743 = p_348_126_ & p_332_122_;
  assign new_n744 = p_341_125_ & ~p_332_122_;
  assign new_n745 = ~new_n743 & ~new_n744;
  assign new_n746 = p_523_148_ & new_n745;
  assign new_n747 = ~p_523_148_ & ~new_n745;
  assign new_n748 = ~new_n746 & ~new_n747;
  assign new_n749 = p_331_121_ & p_332_122_;
  assign new_n750 = p_324_120_ & ~p_332_122_;
  assign new_n751 = ~new_n749 & ~new_n750;
  assign new_n752 = p_503_146_ & new_n751;
  assign new_n753 = ~p_503_146_ & ~new_n751;
  assign new_n754 = ~new_n752 & ~new_n753;
  assign new_n755 = ~new_n742 & ~new_n748;
  assign new_n756 = ~new_n430 & new_n755;
  assign new_n757 = ~new_n427 & new_n756;
  assign new_n758 = ~new_n427 & ~new_n748;
  assign new_n759 = ~new_n742 & new_n758;
  assign new_n760 = new_n430 & new_n759;
  assign new_n761 = p_523_148_ & ~new_n745;
  assign new_n762 = ~new_n742 & new_n761;
  assign new_n763 = p_534_149_ & ~new_n424;
  assign new_n764 = ~new_n742 & new_n763;
  assign new_n765 = ~new_n748 & new_n764;
  assign new_n766 = p_514_147_ & ~new_n739;
  assign new_n767 = ~new_n757 & ~new_n760;
  assign new_n768 = ~new_n762 & new_n767;
  assign new_n769 = ~new_n765 & new_n768;
  assign new_n770 = ~new_n766 & new_n769;
  assign new_n771 = ~new_n427 & new_n430;
  assign new_n772 = ~new_n427 & ~new_n430;
  assign new_n773 = ~new_n763 & ~new_n772;
  assign new_n774 = ~new_n771 & new_n773;
  assign new_n775 = new_n430 & new_n758;
  assign new_n776 = ~new_n748 & new_n763;
  assign new_n777 = ~new_n430 & ~new_n748;
  assign new_n778 = ~new_n427 & new_n777;
  assign new_n779 = ~new_n775 & ~new_n776;
  assign new_n780 = ~new_n778 & new_n779;
  assign new_n781 = ~new_n761 & new_n780;
  assign new_n782 = new_n774 & ~new_n781;
  assign new_n783 = ~new_n774 & new_n781;
  assign new_n784 = ~new_n782 & ~new_n783;
  assign new_n785 = new_n770 & ~new_n784;
  assign new_n786 = ~new_n770 & new_n784;
  assign new_n787 = ~new_n785 & ~new_n786;
  assign new_n788 = ~new_n430 & ~new_n787;
  assign new_n789 = new_n430 & new_n787;
  assign new_n790 = ~new_n788 & ~new_n789;
  assign new_n791 = new_n427 & ~new_n790;
  assign new_n792 = ~new_n427 & new_n790;
  assign new_n793 = ~new_n791 & ~new_n792;
  assign new_n794 = new_n754 & ~new_n793;
  assign new_n795 = ~new_n754 & new_n793;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = new_n748 & ~new_n796;
  assign new_n798 = ~new_n748 & new_n796;
  assign new_n799 = ~new_n797 & ~new_n798;
  assign new_n800 = new_n742 & ~new_n799;
  assign new_n801 = ~new_n742 & new_n799;
  assign new_n802 = ~new_n800 & ~new_n801;
  assign new_n803 = p_2174_161_ & ~new_n802;
  assign new_n804 = ~new_n757 & ~new_n762;
  assign new_n805 = ~new_n765 & new_n804;
  assign new_n806 = ~new_n766 & new_n805;
  assign new_n807 = ~new_n776 & ~new_n778;
  assign new_n808 = ~new_n761 & new_n807;
  assign new_n809 = ~new_n430 & ~new_n808;
  assign new_n810 = new_n430 & new_n808;
  assign new_n811 = ~new_n809 & ~new_n810;
  assign new_n812 = ~new_n773 & ~new_n811;
  assign new_n813 = new_n773 & new_n811;
  assign new_n814 = ~new_n812 & ~new_n813;
  assign new_n815 = ~new_n806 & ~new_n814;
  assign new_n816 = new_n806 & new_n814;
  assign new_n817 = ~new_n815 & ~new_n816;
  assign new_n818 = ~new_n430 & ~new_n817;
  assign new_n819 = new_n430 & new_n817;
  assign new_n820 = ~new_n818 & ~new_n819;
  assign new_n821 = new_n427 & ~new_n820;
  assign new_n822 = ~new_n427 & new_n820;
  assign new_n823 = ~new_n821 & ~new_n822;
  assign new_n824 = new_n754 & ~new_n823;
  assign new_n825 = ~new_n754 & new_n823;
  assign new_n826 = ~new_n824 & ~new_n825;
  assign new_n827 = new_n748 & ~new_n826;
  assign new_n828 = ~new_n748 & new_n826;
  assign new_n829 = ~new_n827 & ~new_n828;
  assign new_n830 = new_n742 & ~new_n829;
  assign new_n831 = ~new_n742 & new_n829;
  assign new_n832 = ~new_n830 & ~new_n831;
  assign new_n833 = ~p_2174_161_ & new_n832;
  assign new_n834 = ~new_n803 & ~new_n833;
  assign new_n835 = ~new_n742 & ~new_n754;
  assign new_n836 = ~new_n427 & new_n835;
  assign new_n837 = ~new_n748 & new_n836;
  assign new_n838 = new_n430 & new_n837;
  assign new_n839 = new_n763 & new_n835;
  assign new_n840 = ~new_n748 & new_n839;
  assign new_n841 = ~new_n430 & ~new_n742;
  assign new_n842 = ~new_n748 & new_n841;
  assign new_n843 = ~new_n754 & new_n842;
  assign new_n844 = ~new_n427 & new_n843;
  assign new_n845 = ~new_n754 & new_n766;
  assign new_n846 = ~new_n754 & new_n761;
  assign new_n847 = ~new_n742 & new_n846;
  assign new_n848 = p_503_146_ & ~new_n751;
  assign new_n849 = ~new_n840 & ~new_n844;
  assign new_n850 = ~new_n845 & new_n849;
  assign new_n851 = ~new_n847 & new_n850;
  assign new_n852 = ~new_n848 & new_n851;
  assign new_n853 = ~new_n838 & new_n852;
  assign new_n854 = p_307_115_ & p_332_122_;
  assign new_n855 = p_302_114_ & ~p_332_122_;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = p_299_113_ & p_332_122_;
  assign new_n858 = p_293_112_ & ~p_332_122_;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = p_315_117_ & p_332_122_;
  assign new_n861 = p_308_116_ & ~p_332_122_;
  assign new_n862 = ~new_n860 & ~new_n861;
  assign new_n863 = p_479_144_ & new_n862;
  assign new_n864 = ~p_479_144_ & ~new_n862;
  assign new_n865 = ~new_n863 & ~new_n864;
  assign new_n866 = p_323_119_ & p_332_122_;
  assign new_n867 = ~p_332_122_ & p_316_118_;
  assign new_n868 = ~new_n866 & ~new_n867;
  assign new_n869 = p_490_145_ & new_n868;
  assign new_n870 = ~p_490_145_ & ~new_n868;
  assign new_n871 = ~new_n869 & ~new_n870;
  assign new_n872 = new_n856 & ~new_n865;
  assign new_n873 = ~new_n871 & new_n872;
  assign new_n874 = p_479_144_ & ~new_n862;
  assign new_n875 = new_n856 & new_n874;
  assign new_n876 = p_490_145_ & ~new_n868;
  assign new_n877 = new_n856 & new_n876;
  assign new_n878 = ~new_n865 & new_n877;
  assign new_n879 = ~new_n873 & ~new_n875;
  assign new_n880 = ~new_n878 & new_n879;
  assign new_n881 = new_n856 & new_n880;
  assign new_n882 = ~new_n865 & ~new_n871;
  assign new_n883 = ~new_n865 & new_n876;
  assign new_n884 = ~new_n874 & ~new_n883;
  assign new_n885 = ~new_n882 & new_n884;
  assign new_n886 = ~p_490_145_ & new_n868;
  assign new_n887 = new_n885 & new_n886;
  assign new_n888 = ~new_n885 & ~new_n886;
  assign new_n889 = ~new_n887 & ~new_n888;
  assign new_n890 = new_n881 & ~new_n889;
  assign new_n891 = ~new_n881 & new_n889;
  assign new_n892 = ~new_n890 & ~new_n891;
  assign new_n893 = new_n871 & ~new_n892;
  assign new_n894 = ~new_n871 & new_n892;
  assign new_n895 = ~new_n893 & ~new_n894;
  assign new_n896 = new_n865 & ~new_n895;
  assign new_n897 = ~new_n865 & new_n895;
  assign new_n898 = ~new_n896 & ~new_n897;
  assign new_n899 = ~new_n859 & ~new_n898;
  assign new_n900 = new_n859 & new_n898;
  assign new_n901 = ~new_n899 & ~new_n900;
  assign new_n902 = ~new_n856 & ~new_n901;
  assign new_n903 = new_n856 & new_n901;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = p_2174_161_ & ~new_n853;
  assign new_n906 = ~new_n904 & new_n905;
  assign new_n907 = ~p_2174_161_ & ~new_n852;
  assign new_n908 = ~new_n904 & new_n907;
  assign new_n909 = ~new_n875 & ~new_n878;
  assign new_n910 = new_n856 & new_n909;
  assign new_n911 = new_n876 & ~new_n884;
  assign new_n912 = ~new_n876 & new_n884;
  assign new_n913 = ~new_n911 & ~new_n912;
  assign new_n914 = ~new_n910 & ~new_n913;
  assign new_n915 = new_n910 & new_n913;
  assign new_n916 = ~new_n914 & ~new_n915;
  assign new_n917 = new_n871 & ~new_n916;
  assign new_n918 = ~new_n871 & new_n916;
  assign new_n919 = ~new_n917 & ~new_n918;
  assign new_n920 = new_n865 & ~new_n919;
  assign new_n921 = ~new_n865 & new_n919;
  assign new_n922 = ~new_n920 & ~new_n921;
  assign new_n923 = ~new_n859 & ~new_n922;
  assign new_n924 = new_n859 & new_n922;
  assign new_n925 = ~new_n923 & ~new_n924;
  assign new_n926 = ~new_n856 & ~new_n925;
  assign new_n927 = new_n856 & new_n925;
  assign new_n928 = ~new_n926 & ~new_n927;
  assign new_n929 = p_2174_161_ & new_n853;
  assign new_n930 = ~new_n928 & new_n929;
  assign new_n931 = ~p_2174_161_ & new_n852;
  assign new_n932 = ~new_n928 & new_n931;
  assign new_n933 = ~new_n906 & ~new_n908;
  assign new_n934 = ~new_n930 & new_n933;
  assign new_n935 = ~new_n932 & new_n934;
  assign new_n936 = new_n834 & ~new_n935;
  assign new_n937 = ~new_n834 & new_n935;
  assign new_n938 = ~new_n936 & ~new_n937;
  assign new_n939 = p_4091_175_ & new_n938;
  assign new_n940 = p_254_101_ & ~p_316_118_;
  assign new_n941 = p_242_97_ & p_316_118_;
  assign new_n942 = ~p_490_145_ & ~new_n940;
  assign new_n943 = ~new_n941 & new_n942;
  assign new_n944 = p_251_100_ & ~p_316_118_;
  assign new_n945 = p_490_145_ & new_n944;
  assign new_n946 = p_490_145_ & p_316_118_;
  assign new_n947 = p_248_99_ & new_n946;
  assign new_n948 = ~new_n945 & ~new_n947;
  assign new_n949 = ~new_n943 & new_n948;
  assign new_n950 = p_254_101_ & ~p_308_116_;
  assign new_n951 = p_242_97_ & p_308_116_;
  assign new_n952 = ~p_479_144_ & ~new_n950;
  assign new_n953 = ~new_n951 & new_n952;
  assign new_n954 = ~p_308_116_ & p_251_100_;
  assign new_n955 = p_479_144_ & new_n954;
  assign new_n956 = p_308_116_ & p_479_144_;
  assign new_n957 = p_248_99_ & new_n956;
  assign new_n958 = ~new_n955 & ~new_n957;
  assign new_n959 = ~new_n953 & new_n958;
  assign new_n960 = ~new_n949 & new_n959;
  assign new_n961 = new_n949 & ~new_n959;
  assign new_n962 = ~new_n960 & ~new_n961;
  assign new_n963 = ~p_302_114_ & p_251_100_;
  assign new_n964 = p_302_114_ & p_248_99_;
  assign new_n965 = ~new_n963 & ~new_n964;
  assign new_n966 = ~p_293_112_ & p_254_101_;
  assign new_n967 = p_293_112_ & p_242_97_;
  assign new_n968 = ~new_n966 & ~new_n967;
  assign new_n969 = ~new_n965 & ~new_n968;
  assign new_n970 = new_n965 & new_n968;
  assign new_n971 = ~new_n969 & ~new_n970;
  assign new_n972 = new_n962 & ~new_n971;
  assign new_n973 = ~new_n962 & new_n971;
  assign new_n974 = ~new_n972 & ~new_n973;
  assign new_n975 = p_251_100_ & ~p_361_129_;
  assign new_n976 = p_248_99_ & p_361_129_;
  assign new_n977 = ~new_n975 & ~new_n976;
  assign new_n978 = ~p_514_147_ & ~p_242_97_;
  assign new_n979 = p_514_147_ & p_248_99_;
  assign new_n980 = ~new_n978 & ~new_n979;
  assign new_n981 = ~p_324_120_ & p_254_101_;
  assign new_n982 = p_324_120_ & p_242_97_;
  assign new_n983 = ~p_503_146_ & ~new_n981;
  assign new_n984 = ~new_n982 & new_n983;
  assign new_n985 = ~p_324_120_ & p_251_100_;
  assign new_n986 = p_503_146_ & new_n985;
  assign new_n987 = p_324_120_ & p_503_146_;
  assign new_n988 = p_248_99_ & new_n987;
  assign new_n989 = ~new_n986 & ~new_n988;
  assign new_n990 = ~new_n984 & new_n989;
  assign new_n991 = ~new_n980 & new_n990;
  assign new_n992 = new_n980 & ~new_n990;
  assign new_n993 = ~new_n991 & ~new_n992;
  assign new_n994 = p_254_101_ & ~p_351_127_;
  assign new_n995 = p_242_97_ & p_351_127_;
  assign new_n996 = ~p_534_149_ & ~new_n994;
  assign new_n997 = ~new_n995 & new_n996;
  assign new_n998 = p_251_100_ & ~p_351_127_;
  assign new_n999 = p_534_149_ & new_n998;
  assign new_n1000 = p_248_99_ & new_n444;
  assign new_n1001 = ~new_n999 & ~new_n1000;
  assign new_n1002 = ~new_n997 & new_n1001;
  assign new_n1003 = p_254_101_ & ~p_341_125_;
  assign new_n1004 = p_242_97_ & p_341_125_;
  assign new_n1005 = ~p_523_148_ & ~new_n1003;
  assign new_n1006 = ~new_n1004 & new_n1005;
  assign new_n1007 = p_251_100_ & ~p_341_125_;
  assign new_n1008 = p_523_148_ & new_n1007;
  assign new_n1009 = p_341_125_ & p_523_148_;
  assign new_n1010 = p_248_99_ & new_n1009;
  assign new_n1011 = ~new_n1008 & ~new_n1010;
  assign new_n1012 = ~new_n1006 & new_n1011;
  assign new_n1013 = ~new_n1002 & new_n1012;
  assign new_n1014 = new_n1002 & ~new_n1012;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = ~new_n977 & ~new_n993;
  assign new_n1017 = ~new_n1015 & new_n1016;
  assign new_n1018 = new_n993 & ~new_n1015;
  assign new_n1019 = new_n977 & new_n1018;
  assign new_n1020 = ~new_n1017 & ~new_n1019;
  assign new_n1021 = new_n977 & ~new_n993;
  assign new_n1022 = new_n1015 & new_n1021;
  assign new_n1023 = new_n993 & new_n1015;
  assign new_n1024 = ~new_n977 & new_n1023;
  assign new_n1025 = ~new_n1022 & ~new_n1024;
  assign new_n1026 = new_n1020 & new_n1025;
  assign new_n1027 = new_n974 & ~new_n1026;
  assign new_n1028 = ~new_n974 & new_n1026;
  assign new_n1029 = ~new_n1027 & ~new_n1028;
  assign new_n1030 = ~p_4091_175_ & ~new_n1029;
  assign new_n1031 = ~new_n939 & ~new_n1030;
  assign new_n1032 = ~p_4092_176_ & ~new_n1031;
  assign new_n1033 = ~new_n737 & ~new_n1032;
  assign new_n1034 = ~p_1694_160_ & ~p_1691_159_;
  assign new_n1035 = ~new_n1033 & new_n1034;
  assign new_n1036 = ~new_n458 & ~new_n734;
  assign new_n1037 = ~new_n736 & new_n1036;
  assign new_n1038 = ~new_n1035 & new_n1037;
  assign p_690_2484_ = ~p_137_63_ | new_n1038;
  assign new_n1040 = p_152_69_ & new_n457;
  assign new_n1041 = p_4_1_ & new_n473;
  assign new_n1042 = ~new_n474 & ~new_n1041;
  assign new_n1043 = ~new_n317 & new_n1042;
  assign new_n1044 = new_n323 & ~new_n1043;
  assign new_n1045 = ~new_n323 & new_n1043;
  assign new_n1046 = ~new_n1044 & ~new_n1045;
  assign new_n1047 = new_n400 & ~new_n1046;
  assign new_n1048 = p_127_55_ & new_n402;
  assign new_n1049 = ~p_3548_166_ & ~p_265_104_;
  assign new_n1050 = ~p_3546_165_ & p_265_104_;
  assign new_n1051 = ~p_400_137_ & ~new_n1049;
  assign new_n1052 = ~new_n1050 & new_n1051;
  assign new_n1053 = ~p_3550_167_ & ~p_265_104_;
  assign new_n1054 = p_400_137_ & new_n1053;
  assign new_n1055 = ~p_3552_168_ & new_n708;
  assign new_n1056 = ~new_n1054 & ~new_n1055;
  assign new_n1057 = ~new_n1052 & new_n1056;
  assign new_n1058 = new_n414 & new_n1057;
  assign new_n1059 = ~new_n1047 & ~new_n1048;
  assign p_875_2125_ = ~new_n1058 & new_n1059;
  assign new_n1061 = new_n733 & ~p_875_2125_;
  assign new_n1062 = p_155_70_ & new_n735;
  assign new_n1063 = p_54_20_ & new_n771;
  assign new_n1064 = ~new_n772 & ~new_n1063;
  assign new_n1065 = ~new_n763 & new_n1064;
  assign new_n1066 = new_n748 & ~new_n1065;
  assign new_n1067 = ~new_n748 & new_n1065;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n400 & ~new_n1068;
  assign new_n1070 = p_119_49_ & new_n402;
  assign new_n1071 = ~p_341_125_ & ~p_3548_166_;
  assign new_n1072 = p_341_125_ & ~p_3546_165_;
  assign new_n1073 = ~p_523_148_ & ~new_n1071;
  assign new_n1074 = ~new_n1072 & new_n1073;
  assign new_n1075 = ~p_3550_167_ & ~p_341_125_;
  assign new_n1076 = p_523_148_ & new_n1075;
  assign new_n1077 = ~p_3552_168_ & new_n1009;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = ~new_n1074 & new_n1078;
  assign new_n1080 = new_n414 & new_n1079;
  assign new_n1081 = ~new_n1069 & ~new_n1070;
  assign p_836_2128_ = ~new_n1080 & new_n1081;
  assign new_n1083 = new_n1034 & ~p_836_2128_;
  assign new_n1084 = ~new_n1040 & ~new_n1061;
  assign new_n1085 = ~new_n1062 & new_n1084;
  assign new_n1086 = ~new_n1083 & new_n1085;
  assign p_699_2227_ = p_137_63_ & ~new_n1086;
  assign new_n1088 = new_n859 & ~new_n871;
  assign new_n1089 = ~new_n865 & new_n1088;
  assign new_n1090 = new_n856 & new_n1089;
  assign new_n1091 = ~new_n852 & new_n1090;
  assign new_n1092 = new_n856 & new_n859;
  assign new_n1093 = new_n876 & new_n1092;
  assign new_n1094 = ~new_n865 & new_n1093;
  assign new_n1095 = ~new_n856 & new_n859;
  assign new_n1096 = new_n859 & new_n874;
  assign new_n1097 = new_n856 & new_n1096;
  assign new_n1098 = ~new_n1094 & ~new_n1095;
  assign new_n1099 = ~new_n1097 & new_n1098;
  assign new_n1100 = new_n859 & new_n1099;
  assign p_618_1925_ = new_n1091 | ~new_n1100;
  assign p_588_1696_ = new_n374 & new_n543;
  assign new_n1103 = ~new_n427 & ~new_n754;
  assign new_n1104 = new_n430 & new_n1103;
  assign new_n1105 = ~new_n748 & new_n1104;
  assign new_n1106 = ~new_n742 & new_n1105;
  assign p_615_1750_ = new_n1090 & new_n1106;
  assign new_n1108 = p_161_72_ & new_n457;
  assign new_n1109 = new_n353 & ~new_n552;
  assign new_n1110 = ~new_n353 & new_n552;
  assign new_n1111 = ~new_n1109 & ~new_n1110;
  assign new_n1112 = ~new_n313 & ~new_n333;
  assign new_n1113 = ~new_n394 & new_n1112;
  assign new_n1114 = ~new_n323 & new_n1113;
  assign new_n1115 = ~new_n307 & new_n1114;
  assign new_n1116 = p_4_1_ & new_n1115;
  assign new_n1117 = new_n347 & ~new_n1116;
  assign new_n1118 = ~new_n1111 & ~new_n1117;
  assign new_n1119 = new_n376 & new_n545;
  assign new_n1120 = ~new_n547 & ~new_n1119;
  assign new_n1121 = ~new_n380 & new_n1120;
  assign new_n1122 = new_n353 & new_n1121;
  assign new_n1123 = ~new_n353 & ~new_n1121;
  assign new_n1124 = ~new_n1122 & ~new_n1123;
  assign new_n1125 = new_n1117 & new_n1124;
  assign new_n1126 = ~new_n1118 & ~new_n1125;
  assign new_n1127 = new_n400 & ~new_n1126;
  assign new_n1128 = p_115_45_ & new_n402;
  assign new_n1129 = new_n414 & new_n653;
  assign new_n1130 = ~new_n1127 & ~new_n1128;
  assign p_863_2276_ = ~new_n1129 & new_n1130;
  assign new_n1132 = new_n733 & ~p_863_2276_;
  assign new_n1133 = p_191_82_ & new_n735;
  assign new_n1134 = ~new_n859 & ~new_n881;
  assign new_n1135 = new_n859 & new_n881;
  assign new_n1136 = ~new_n1134 & ~new_n1135;
  assign new_n1137 = p_54_20_ & new_n1106;
  assign new_n1138 = new_n852 & ~new_n1137;
  assign new_n1139 = ~new_n1136 & ~new_n1138;
  assign new_n1140 = new_n872 & new_n876;
  assign new_n1141 = ~new_n875 & ~new_n1140;
  assign new_n1142 = new_n856 & new_n1141;
  assign new_n1143 = ~new_n859 & new_n1142;
  assign new_n1144 = new_n859 & ~new_n1142;
  assign new_n1145 = ~new_n1143 & ~new_n1144;
  assign new_n1146 = new_n1138 & new_n1145;
  assign p_623_2152_ = ~new_n1139 & ~new_n1146;
  assign new_n1148 = new_n400 & ~p_623_2152_;
  assign new_n1149 = p_123_53_ & new_n402;
  assign new_n1150 = new_n414 & ~new_n968;
  assign new_n1151 = ~new_n1148 & ~new_n1149;
  assign p_824_2274_ = ~new_n1150 & new_n1151;
  assign new_n1153 = new_n1034 & ~p_824_2274_;
  assign new_n1154 = ~new_n1108 & ~new_n1132;
  assign new_n1155 = ~new_n1133 & new_n1154;
  assign new_n1156 = ~new_n1153 & new_n1155;
  assign p_688_2317_ = p_137_63_ & ~new_n1156;
  assign p_809_655_ = ~p_31_11_ | ~p_27_10_;
  assign new_n1159 = p_88_34_ & ~p_2358_162_;
  assign new_n1160 = p_34_12_ & p_2358_162_;
  assign new_n1161 = ~new_n1159 & ~new_n1160;
  assign p_704_1281_ = p_809_655_ | new_n1161;
  assign new_n1163 = p_3717_169_ & p_3724_170_;
  assign new_n1164 = ~p_623_2152_ & new_n1163;
  assign new_n1165 = p_132_60_ & new_n859;
  assign new_n1166 = p_132_60_ & ~new_n1165;
  assign new_n1167 = new_n859 & ~new_n1165;
  assign new_n1168 = ~new_n1166 & ~new_n1167;
  assign new_n1169 = ~p_3717_169_ & p_3724_170_;
  assign new_n1170 = ~new_n1168 & new_n1169;
  assign new_n1171 = p_3717_169_ & ~p_3724_170_;
  assign new_n1172 = p_123_53_ & new_n1171;
  assign new_n1173 = ~p_3717_169_ & ~p_3724_170_;
  assign new_n1174 = ~new_n968 & new_n1173;
  assign new_n1175 = ~new_n1164 & ~new_n1170;
  assign new_n1176 = ~new_n1172 & new_n1175;
  assign new_n1177 = ~new_n1174 & new_n1176;
  assign new_n1178 = p_4115_177_ & p_135_61_;
  assign p_818_2273_ = ~new_n1177 & ~new_n1178;
  assign new_n1180 = new_n371 & ~new_n1117;
  assign new_n1181 = ~new_n371 & new_n1117;
  assign new_n1182 = ~new_n1180 & ~new_n1181;
  assign new_n1183 = new_n400 & ~new_n1182;
  assign new_n1184 = p_113_43_ & new_n402;
  assign new_n1185 = ~p_226_93_ & ~p_3548_166_;
  assign new_n1186 = p_226_93_ & ~p_3546_165_;
  assign new_n1187 = ~p_422_139_ & ~new_n1185;
  assign new_n1188 = ~new_n1186 & new_n1187;
  assign new_n1189 = ~p_226_93_ & ~p_3550_167_;
  assign new_n1190 = p_422_139_ & new_n1189;
  assign new_n1191 = ~p_3552_168_ & new_n617;
  assign new_n1192 = ~new_n1190 & ~new_n1191;
  assign new_n1193 = ~new_n1188 & new_n1192;
  assign new_n1194 = new_n414 & new_n1193;
  assign new_n1195 = ~new_n1183 & ~new_n1184;
  assign p_869_2181_ = ~new_n1194 & new_n1195;
  assign new_n1197 = p_167_74_ & new_n390;
  assign new_n1198 = new_n359 & new_n557;
  assign new_n1199 = ~new_n359 & ~new_n557;
  assign new_n1200 = ~new_n1198 & ~new_n1199;
  assign new_n1201 = ~new_n1117 & new_n1200;
  assign new_n1202 = new_n359 & new_n376;
  assign new_n1203 = ~new_n359 & ~new_n376;
  assign new_n1204 = ~new_n1202 & ~new_n1203;
  assign new_n1205 = new_n1117 & ~new_n1204;
  assign new_n1206 = ~new_n1201 & ~new_n1205;
  assign new_n1207 = new_n400 & ~new_n1206;
  assign new_n1208 = p_53_19_ & new_n402;
  assign new_n1209 = ~p_3548_166_ & ~p_218_91_;
  assign new_n1210 = ~p_3546_165_ & p_218_91_;
  assign new_n1211 = ~p_468_143_ & ~new_n1209;
  assign new_n1212 = ~new_n1210 & new_n1211;
  assign new_n1213 = ~p_3550_167_ & ~p_218_91_;
  assign new_n1214 = p_468_143_ & new_n1213;
  assign new_n1215 = ~p_3552_168_ & new_n627;
  assign new_n1216 = ~new_n1214 & ~new_n1215;
  assign new_n1217 = ~new_n1212 & new_n1216;
  assign new_n1218 = new_n414 & new_n1217;
  assign new_n1219 = ~new_n1207 & ~new_n1208;
  assign p_867_2237_ = ~new_n1218 & new_n1219;
  assign new_n1221 = new_n418 & ~p_867_2237_;
  assign new_n1222 = p_197_84_ & new_n420;
  assign new_n1223 = new_n865 & new_n886;
  assign new_n1224 = ~new_n865 & ~new_n886;
  assign new_n1225 = ~new_n1223 & ~new_n1224;
  assign new_n1226 = ~new_n1138 & new_n1225;
  assign new_n1227 = new_n865 & new_n876;
  assign new_n1228 = ~new_n865 & ~new_n876;
  assign new_n1229 = ~new_n1227 & ~new_n1228;
  assign new_n1230 = new_n1138 & ~new_n1229;
  assign new_n1231 = ~new_n1226 & ~new_n1230;
  assign new_n1232 = new_n400 & ~new_n1231;
  assign new_n1233 = p_116_46_ & new_n402;
  assign new_n1234 = new_n414 & new_n959;
  assign new_n1235 = ~new_n1232 & ~new_n1233;
  assign p_828_2233_ = ~new_n1234 & new_n1235;
  assign new_n1237 = new_n451 & ~p_828_2233_;
  assign new_n1238 = ~new_n1197 & ~new_n1221;
  assign new_n1239 = ~new_n1222 & new_n1238;
  assign new_n1240 = ~new_n1237 & new_n1239;
  assign p_648_2295_ = p_137_63_ & ~new_n1240;
  assign new_n1242 = p_54_20_ & ~new_n430;
  assign new_n1243 = ~p_54_20_ & new_n430;
  assign new_n1244 = ~new_n1242 & ~new_n1243;
  assign new_n1245 = new_n400 & ~new_n1244;
  assign new_n1246 = p_131_59_ & new_n402;
  assign new_n1247 = new_n414 & new_n977;
  assign new_n1248 = ~new_n1245 & ~new_n1246;
  assign p_822_1933_ = ~new_n1247 & new_n1248;
  assign new_n1250 = p_4088_172_ & p_4087_171_;
  assign new_n1251 = p_17_4_ & new_n1250;
  assign new_n1252 = p_4088_172_ & ~p_4087_171_;
  assign new_n1253 = ~p_875_2125_ & new_n1252;
  assign new_n1254 = ~p_4088_172_ & p_4087_171_;
  assign new_n1255 = p_73_25_ & new_n1254;
  assign new_n1256 = ~p_4088_172_ & ~p_4087_171_;
  assign new_n1257 = ~p_836_2128_ & new_n1256;
  assign new_n1258 = ~new_n1251 & ~new_n1253;
  assign new_n1259 = ~new_n1255 & new_n1258;
  assign p_757_2190_ = new_n1257 | ~new_n1259;
  assign new_n1261 = p_61_21_ & new_n1250;
  assign new_n1262 = p_4_1_ & new_n394;
  assign new_n1263 = ~p_4_1_ & ~new_n394;
  assign new_n1264 = ~new_n1262 & ~new_n1263;
  assign new_n1265 = new_n400 & ~new_n1264;
  assign new_n1266 = p_117_47_ & new_n402;
  assign new_n1267 = ~p_3548_166_ & ~p_281_108_;
  assign new_n1268 = ~p_3546_165_ & p_281_108_;
  assign new_n1269 = ~p_374_134_ & ~new_n1267;
  assign new_n1270 = ~new_n1268 & new_n1269;
  assign new_n1271 = ~p_3550_167_ & ~p_281_108_;
  assign new_n1272 = p_374_134_ & new_n1271;
  assign new_n1273 = ~p_3552_168_ & new_n666;
  assign new_n1274 = ~new_n1272 & ~new_n1273;
  assign new_n1275 = ~new_n1270 & new_n1274;
  assign new_n1276 = new_n414 & new_n1275;
  assign new_n1277 = ~new_n1265 & ~new_n1266;
  assign p_861_2070_ = ~new_n1276 & new_n1277;
  assign new_n1279 = new_n1252 & ~p_861_2070_;
  assign new_n1280 = p_11_2_ & new_n1254;
  assign new_n1281 = ~p_822_1933_ & new_n1256;
  assign new_n1282 = ~new_n1261 & ~new_n1279;
  assign new_n1283 = ~new_n1280 & new_n1282;
  assign p_722_2131_ = new_n1281 | ~new_n1283;
  assign new_n1285 = p_4090_174_ & p_4089_173_;
  assign new_n1286 = p_70_24_ & new_n1285;
  assign new_n1287 = ~p_4090_174_ & p_4089_173_;
  assign new_n1288 = ~p_877_2126_ & new_n1287;
  assign new_n1289 = p_4090_174_ & ~p_4089_173_;
  assign new_n1290 = p_67_23_ & new_n1289;
  assign new_n1291 = ~p_4090_174_ & ~p_4089_173_;
  assign new_n1292 = ~p_838_2064_ & new_n1291;
  assign new_n1293 = ~new_n1286 & ~new_n1288;
  assign new_n1294 = ~new_n1290 & new_n1293;
  assign p_802_2183_ = new_n1292 | ~new_n1294;
  assign new_n1296 = ~new_n316 & new_n329;
  assign new_n1297 = new_n316 & ~new_n329;
  assign new_n1298 = ~new_n1296 & ~new_n1297;
  assign new_n1299 = ~new_n304 & new_n320;
  assign new_n1300 = new_n304 & ~new_n320;
  assign new_n1301 = ~new_n1299 & ~new_n1300;
  assign new_n1302 = new_n1298 & ~new_n1301;
  assign new_n1303 = ~new_n1298 & new_n1301;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = new_n310 & ~new_n368;
  assign new_n1306 = ~new_n310 & new_n368;
  assign new_n1307 = ~new_n1305 & ~new_n1306;
  assign new_n1308 = p_335_123_ & p_292_111_;
  assign new_n1309 = ~p_335_123_ & p_289_110_;
  assign new_n1310 = ~new_n1308 & ~new_n1309;
  assign new_n1311 = new_n350 & ~new_n1310;
  assign new_n1312 = ~new_n350 & new_n1310;
  assign new_n1313 = ~new_n1311 & ~new_n1312;
  assign new_n1314 = new_n356 & ~new_n362;
  assign new_n1315 = ~new_n356 & new_n362;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = ~new_n1307 & ~new_n1313;
  assign new_n1318 = ~new_n1316 & new_n1317;
  assign new_n1319 = new_n1313 & ~new_n1316;
  assign new_n1320 = new_n1307 & new_n1319;
  assign new_n1321 = ~new_n1318 & ~new_n1320;
  assign new_n1322 = new_n1307 & ~new_n1313;
  assign new_n1323 = new_n1316 & new_n1322;
  assign new_n1324 = new_n1313 & new_n1316;
  assign new_n1325 = ~new_n1307 & new_n1324;
  assign new_n1326 = ~new_n1323 & ~new_n1325;
  assign new_n1327 = new_n1321 & new_n1326;
  assign new_n1328 = new_n1304 & ~new_n1327;
  assign new_n1329 = ~new_n1304 & new_n1327;
  assign p_1000_2168_ = new_n1328 | new_n1329;
  assign new_n1331 = p_167_74_ & new_n457;
  assign new_n1332 = new_n733 & ~p_867_2237_;
  assign new_n1333 = p_197_84_ & new_n735;
  assign new_n1334 = new_n1034 & ~p_828_2233_;
  assign new_n1335 = ~new_n1331 & ~new_n1332;
  assign new_n1336 = ~new_n1333 & new_n1335;
  assign new_n1337 = ~new_n1334 & new_n1336;
  assign p_682_2296_ = p_137_63_ & ~new_n1337;
  assign new_n1339 = p_20_5_ & new_n1285;
  assign new_n1340 = ~new_n323 & new_n473;
  assign new_n1341 = p_4_1_ & new_n1340;
  assign new_n1342 = ~new_n478 & ~new_n1341;
  assign new_n1343 = ~new_n480 & new_n1342;
  assign new_n1344 = ~new_n340 & new_n1343;
  assign new_n1345 = new_n307 & ~new_n1344;
  assign new_n1346 = ~new_n307 & new_n1344;
  assign new_n1347 = ~new_n1345 & ~new_n1346;
  assign new_n1348 = new_n400 & ~new_n1347;
  assign new_n1349 = p_128_56_ & new_n402;
  assign new_n1350 = ~p_257_102_ & ~p_3548_166_;
  assign new_n1351 = p_257_102_ & ~p_3546_165_;
  assign new_n1352 = ~p_389_136_ & ~new_n1350;
  assign new_n1353 = ~new_n1351 & new_n1352;
  assign new_n1354 = ~p_257_102_ & ~p_3550_167_;
  assign new_n1355 = p_389_136_ & new_n1354;
  assign new_n1356 = ~p_3552_168_ & new_n676;
  assign new_n1357 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = ~new_n1353 & new_n1357;
  assign new_n1359 = new_n414 & new_n1358;
  assign new_n1360 = ~new_n1348 & ~new_n1349;
  assign p_873_2124_ = ~new_n1359 & new_n1360;
  assign new_n1362 = new_n1287 & ~p_873_2124_;
  assign new_n1363 = p_76_26_ & new_n1289;
  assign new_n1364 = ~new_n748 & new_n771;
  assign new_n1365 = p_54_20_ & new_n1364;
  assign new_n1366 = ~new_n776 & ~new_n1365;
  assign new_n1367 = ~new_n778 & new_n1366;
  assign new_n1368 = ~new_n761 & new_n1367;
  assign new_n1369 = new_n742 & ~new_n1368;
  assign new_n1370 = ~new_n742 & new_n1368;
  assign new_n1371 = ~new_n1369 & ~new_n1370;
  assign new_n1372 = new_n400 & ~new_n1371;
  assign new_n1373 = p_130_58_ & new_n402;
  assign new_n1374 = ~p_514_147_ & p_3546_165_;
  assign new_n1375 = p_514_147_ & ~p_3552_168_;
  assign new_n1376 = ~new_n1374 & ~new_n1375;
  assign new_n1377 = new_n414 & new_n1376;
  assign new_n1378 = ~new_n1372 & ~new_n1373;
  assign p_834_2123_ = ~new_n1377 & new_n1378;
  assign new_n1380 = new_n1291 & ~p_834_2123_;
  assign new_n1381 = ~new_n1339 & ~new_n1362;
  assign new_n1382 = ~new_n1363 & new_n1381;
  assign p_792_2188_ = new_n1380 | ~new_n1382;
  assign new_n1384 = new_n859 & ~new_n865;
  assign new_n1385 = new_n856 & new_n1384;
  assign new_n1386 = ~new_n871 & new_n1385;
  assign new_n1387 = ~new_n852 & new_n1386;
  assign p_629_1926_ = ~new_n1100 | new_n1387;
  assign new_n1389 = p_49_17_ & new_n1285;
  assign new_n1390 = ~new_n553 & ~new_n554;
  assign new_n1391 = ~new_n382 & new_n1390;
  assign new_n1392 = new_n365 & ~new_n1391;
  assign new_n1393 = ~new_n365 & new_n1391;
  assign new_n1394 = ~new_n1392 & ~new_n1393;
  assign new_n1395 = ~new_n1117 & ~new_n1394;
  assign new_n1396 = new_n365 & new_n555;
  assign new_n1397 = ~new_n365 & ~new_n555;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = new_n1117 & new_n1398;
  assign new_n1400 = ~new_n1395 & ~new_n1399;
  assign new_n1401 = new_n400 & ~new_n1400;
  assign new_n1402 = p_114_44_ & new_n402;
  assign new_n1403 = ~p_210_89_ & ~p_3548_166_;
  assign new_n1404 = p_210_89_ & ~p_3546_165_;
  assign new_n1405 = ~p_457_142_ & ~new_n1403;
  assign new_n1406 = ~new_n1404 & new_n1405;
  assign new_n1407 = ~p_210_89_ & ~p_3550_167_;
  assign new_n1408 = p_457_142_ & new_n1407;
  assign new_n1409 = ~p_3552_168_ & new_n640;
  assign new_n1410 = ~new_n1408 & ~new_n1409;
  assign new_n1411 = ~new_n1406 & new_n1410;
  assign new_n1412 = new_n414 & new_n1411;
  assign new_n1413 = ~new_n1401 & ~new_n1402;
  assign p_865_2277_ = ~new_n1412 & new_n1413;
  assign new_n1415 = new_n1287 & ~p_865_2277_;
  assign new_n1416 = p_46_16_ & new_n1289;
  assign new_n1417 = ~new_n882 & ~new_n883;
  assign new_n1418 = ~new_n874 & new_n1417;
  assign new_n1419 = ~new_n856 & ~new_n1418;
  assign new_n1420 = new_n856 & new_n1418;
  assign new_n1421 = ~new_n1419 & ~new_n1420;
  assign new_n1422 = ~new_n1138 & ~new_n1421;
  assign new_n1423 = ~new_n856 & new_n884;
  assign new_n1424 = new_n856 & ~new_n884;
  assign new_n1425 = ~new_n1423 & ~new_n1424;
  assign new_n1426 = new_n1138 & new_n1425;
  assign new_n1427 = ~new_n1422 & ~new_n1426;
  assign new_n1428 = new_n400 & ~new_n1427;
  assign new_n1429 = p_121_51_ & new_n402;
  assign new_n1430 = new_n414 & new_n965;
  assign new_n1431 = ~new_n1428 & ~new_n1429;
  assign p_826_2275_ = ~new_n1430 & new_n1431;
  assign new_n1433 = new_n1291 & ~p_826_2275_;
  assign new_n1434 = ~new_n1389 & ~new_n1415;
  assign new_n1435 = ~new_n1416 & new_n1434;
  assign p_772_2299_ = new_n1433 | ~new_n1435;
  assign new_n1437 = p_17_4_ & new_n1285;
  assign new_n1438 = ~p_875_2125_ & new_n1287;
  assign new_n1439 = p_73_25_ & new_n1289;
  assign new_n1440 = ~p_836_2128_ & new_n1291;
  assign new_n1441 = ~new_n1437 & ~new_n1438;
  assign new_n1442 = ~new_n1439 & new_n1441;
  assign p_797_2191_ = new_n1440 | ~new_n1442;
  assign new_n1444 = p_185_80_ & new_n390;
  assign new_n1445 = new_n418 & ~p_861_2070_;
  assign new_n1446 = p_182_79_ & new_n420;
  assign new_n1447 = new_n451 & ~p_822_1933_;
  assign new_n1448 = ~new_n1444 & ~new_n1445;
  assign new_n1449 = ~new_n1446 & new_n1448;
  assign new_n1450 = ~new_n1447 & new_n1449;
  assign p_661_2178_ = p_137_63_ & ~new_n1450;
  assign new_n1452 = p_106_40_ & new_n1250;
  assign new_n1453 = ~p_863_2276_ & new_n1252;
  assign new_n1454 = p_109_41_ & new_n1254;
  assign new_n1455 = ~p_824_2274_ & new_n1256;
  assign new_n1456 = ~new_n1452 & ~new_n1453;
  assign new_n1457 = ~new_n1454 & new_n1456;
  assign p_727_2298_ = new_n1455 | ~new_n1457;
  assign new_n1459 = ~p_324_120_ & ~p_3548_166_;
  assign new_n1460 = p_324_120_ & ~p_3546_165_;
  assign new_n1461 = ~p_503_146_ & ~new_n1459;
  assign new_n1462 = ~new_n1460 & new_n1461;
  assign new_n1463 = ~p_324_120_ & ~p_3550_167_;
  assign new_n1464 = p_503_146_ & new_n1463;
  assign new_n1465 = ~p_3552_168_ & new_n987;
  assign new_n1466 = ~new_n1464 & ~new_n1465;
  assign new_n1467 = ~new_n1462 & new_n1466;
  assign new_n1468 = ~new_n1079 & ~new_n1467;
  assign new_n1469 = ~new_n1376 & new_n1468;
  assign new_n1470 = ~new_n447 & new_n1469;
  assign new_n1471 = ~new_n959 & new_n968;
  assign new_n1472 = ~new_n965 & new_n1471;
  assign new_n1473 = ~new_n949 & new_n1472;
  assign new_n1474 = ~new_n977 & new_n1470;
  assign p_598_1623_ = new_n1473 & new_n1474;
  assign p_634_665_ = p_373_133_ & p_1_0_;
  assign new_n1477 = p_86_32_ & ~p_2358_162_;
  assign new_n1478 = p_87_33_ & p_2358_162_;
  assign new_n1479 = ~new_n1477 & ~new_n1478;
  assign p_636_1280_ = p_809_655_ | new_n1479;
  assign new_n1481 = p_40_14_ & new_n1250;
  assign new_n1482 = ~p_869_2181_ & new_n1252;
  assign new_n1483 = p_91_35_ & new_n1254;
  assign new_n1484 = new_n871 & ~new_n1138;
  assign new_n1485 = ~new_n871 & new_n1138;
  assign new_n1486 = ~new_n1484 & ~new_n1485;
  assign new_n1487 = new_n400 & ~new_n1486;
  assign new_n1488 = p_112_42_ & new_n402;
  assign new_n1489 = new_n414 & new_n949;
  assign new_n1490 = ~new_n1487 & ~new_n1488;
  assign p_830_2182_ = ~new_n1489 & new_n1490;
  assign new_n1492 = new_n1256 & ~p_830_2182_;
  assign new_n1493 = ~new_n1481 & ~new_n1482;
  assign new_n1494 = ~new_n1483 & new_n1493;
  assign p_742_2238_ = new_n1492 | ~new_n1494;
  assign new_n1496 = p_64_22_ & new_n1250;
  assign new_n1497 = ~new_n732 & new_n1252;
  assign new_n1498 = p_14_3_ & new_n1254;
  assign new_n1499 = ~new_n1033 & new_n1256;
  assign new_n1500 = ~new_n1496 & ~new_n1497;
  assign new_n1501 = ~new_n1498 & new_n1500;
  assign p_767_2479_ = new_n1499 | ~new_n1501;
  assign new_n1503 = p_185_80_ & new_n457;
  assign new_n1504 = new_n733 & ~p_861_2070_;
  assign new_n1505 = p_182_79_ & new_n735;
  assign new_n1506 = new_n1034 & ~p_822_1933_;
  assign new_n1507 = ~new_n1503 & ~new_n1504;
  assign new_n1508 = ~new_n1505 & new_n1507;
  assign new_n1509 = ~new_n1506 & new_n1508;
  assign p_693_2179_ = p_137_63_ & ~new_n1509;
  assign new_n1511 = p_146_67_ & new_n457;
  assign new_n1512 = new_n733 & ~p_873_2124_;
  assign new_n1513 = p_149_68_ & new_n735;
  assign new_n1514 = new_n1034 & ~p_834_2123_;
  assign new_n1515 = ~new_n1511 & ~new_n1512;
  assign new_n1516 = ~new_n1513 & new_n1515;
  assign new_n1517 = ~new_n1514 & new_n1516;
  assign p_702_2228_ = p_137_63_ & ~new_n1517;
  assign new_n1519 = p_64_22_ & new_n1285;
  assign new_n1520 = ~new_n732 & new_n1287;
  assign new_n1521 = p_14_3_ & new_n1289;
  assign new_n1522 = ~new_n1033 & new_n1291;
  assign new_n1523 = ~new_n1519 & ~new_n1520;
  assign new_n1524 = ~new_n1521 & new_n1523;
  assign p_807_2480_ = new_n1522 | ~new_n1524;
  assign new_n1526 = p_161_72_ & new_n390;
  assign new_n1527 = new_n418 & ~p_863_2276_;
  assign new_n1528 = p_191_82_ & new_n420;
  assign new_n1529 = new_n451 & ~p_824_2274_;
  assign new_n1530 = ~new_n1526 & ~new_n1527;
  assign new_n1531 = ~new_n1528 & new_n1530;
  assign new_n1532 = ~new_n1529 & new_n1531;
  assign p_654_2315_ = p_137_63_ & ~new_n1532;
  assign new_n1534 = p_179_78_ & new_n390;
  assign new_n1535 = new_n418 & ~new_n732;
  assign new_n1536 = p_176_77_ & new_n420;
  assign new_n1537 = new_n451 & ~new_n1033;
  assign new_n1538 = ~new_n1534 & ~new_n1535;
  assign new_n1539 = ~new_n1536 & new_n1538;
  assign new_n1540 = ~new_n1537 & new_n1539;
  assign p_658_2483_ = ~p_137_63_ | new_n1540;
  assign new_n1542 = p_83_31_ & ~p_2358_162_;
  assign new_n1543 = p_83_31_ & p_2358_162_;
  assign new_n1544 = ~new_n1542 & ~new_n1543;
  assign p_820_1283_ = p_809_655_ | new_n1544;
  assign new_n1546 = p_164_73_ & new_n457;
  assign new_n1547 = new_n733 & ~p_865_2277_;
  assign new_n1548 = p_194_83_ & new_n735;
  assign new_n1549 = new_n1034 & ~p_826_2275_;
  assign new_n1550 = ~new_n1546 & ~new_n1547;
  assign new_n1551 = ~new_n1548 & new_n1550;
  assign new_n1552 = ~new_n1549 & new_n1551;
  assign p_685_2316_ = p_137_63_ & ~new_n1552;
  assign p_815_627_ = p_136_62_ & ~p_3173_164_;
  assign new_n1555 = p_4091_175_ & p_4092_176_;
  assign new_n1556 = new_n400 & ~new_n609;
  assign new_n1557 = p_118_48_ & new_n402;
  assign new_n1558 = new_n414 & new_n728;
  assign new_n1559 = ~new_n1555 & ~new_n1556;
  assign new_n1560 = ~new_n1557 & new_n1559;
  assign p_882_2456_ = new_n1558 | ~new_n1560;
  assign new_n1562 = ~new_n353 & ~new_n371;
  assign new_n1563 = ~new_n359 & new_n1562;
  assign new_n1564 = ~new_n365 & new_n1563;
  assign new_n1565 = ~new_n347 & new_n1564;
  assign p_621_1893_ = ~new_n388 | new_n1565;
  assign new_n1567 = p_170_75_ & new_n457;
  assign new_n1568 = ~new_n307 & ~new_n333;
  assign new_n1569 = ~new_n394 & new_n1568;
  assign new_n1570 = ~new_n323 & new_n1569;
  assign new_n1571 = p_4_1_ & new_n1570;
  assign new_n1572 = ~new_n462 & ~new_n1571;
  assign new_n1573 = ~new_n466 & new_n1572;
  assign new_n1574 = ~new_n468 & new_n1573;
  assign new_n1575 = ~new_n338 & new_n1574;
  assign new_n1576 = new_n313 & ~new_n1575;
  assign new_n1577 = ~new_n313 & new_n1575;
  assign new_n1578 = ~new_n1576 & ~new_n1577;
  assign new_n1579 = new_n400 & ~new_n1578;
  assign new_n1580 = p_122_52_ & new_n402;
  assign new_n1581 = ~p_234_95_ & ~p_3548_166_;
  assign new_n1582 = p_234_95_ & ~p_3546_165_;
  assign new_n1583 = ~p_435_140_ & ~new_n1581;
  assign new_n1584 = ~new_n1582 & new_n1583;
  assign new_n1585 = ~p_3550_167_ & ~p_234_95_;
  assign new_n1586 = p_435_140_ & new_n1585;
  assign new_n1587 = ~p_3552_168_ & new_n686;
  assign new_n1588 = ~new_n1586 & ~new_n1587;
  assign new_n1589 = ~new_n1584 & new_n1588;
  assign new_n1590 = new_n414 & new_n1589;
  assign new_n1591 = ~new_n1579 & ~new_n1580;
  assign p_871_2127_ = ~new_n1590 & new_n1591;
  assign new_n1593 = new_n733 & ~p_871_2127_;
  assign new_n1594 = p_200_85_ & new_n735;
  assign new_n1595 = ~new_n427 & ~new_n742;
  assign new_n1596 = new_n430 & new_n1595;
  assign new_n1597 = ~new_n748 & new_n1596;
  assign new_n1598 = p_54_20_ & new_n1597;
  assign new_n1599 = ~new_n757 & ~new_n1598;
  assign new_n1600 = ~new_n762 & new_n1599;
  assign new_n1601 = ~new_n765 & new_n1600;
  assign new_n1602 = ~new_n766 & new_n1601;
  assign new_n1603 = new_n754 & ~new_n1602;
  assign new_n1604 = ~new_n754 & new_n1602;
  assign new_n1605 = ~new_n1603 & ~new_n1604;
  assign new_n1606 = new_n400 & ~new_n1605;
  assign new_n1607 = p_52_18_ & new_n402;
  assign new_n1608 = new_n414 & new_n1467;
  assign new_n1609 = ~new_n1606 & ~new_n1607;
  assign p_832_2133_ = ~new_n1608 & new_n1609;
  assign new_n1611 = new_n1034 & ~p_832_2133_;
  assign new_n1612 = ~new_n1567 & ~new_n1593;
  assign new_n1613 = ~new_n1594 & new_n1612;
  assign new_n1614 = ~new_n1611 & new_n1613;
  assign p_676_2229_ = p_137_63_ & ~new_n1614;
  assign new_n1616 = p_152_69_ & new_n390;
  assign new_n1617 = new_n418 & ~p_875_2125_;
  assign new_n1618 = p_155_70_ & new_n420;
  assign new_n1619 = new_n451 & ~p_836_2128_;
  assign new_n1620 = ~new_n1616 & ~new_n1617;
  assign new_n1621 = ~new_n1618 & new_n1620;
  assign new_n1622 = ~new_n1619 & new_n1621;
  assign p_667_2224_ = p_137_63_ & ~new_n1622;
  assign new_n1624 = p_158_71_ & new_n457;
  assign new_n1625 = ~p_877_2126_ & new_n733;
  assign new_n1626 = p_188_81_ & new_n735;
  assign new_n1627 = ~p_838_2064_ & new_n1034;
  assign new_n1628 = ~new_n1624 & ~new_n1625;
  assign new_n1629 = ~new_n1626 & new_n1628;
  assign new_n1630 = ~new_n1627 & new_n1629;
  assign p_696_2226_ = p_137_63_ & ~new_n1630;
  assign new_n1632 = p_37_13_ & new_n1285;
  assign new_n1633 = new_n1287 & ~p_871_2127_;
  assign new_n1634 = p_43_15_ & new_n1289;
  assign new_n1635 = new_n1291 & ~p_832_2133_;
  assign new_n1636 = ~new_n1632 & ~new_n1633;
  assign new_n1637 = ~new_n1634 & new_n1636;
  assign p_787_2186_ = new_n1635 | ~new_n1637;
  assign new_n1639 = p_308_116_ & ~p_316_118_;
  assign new_n1640 = ~p_308_116_ & p_316_118_;
  assign new_n1641 = ~new_n1639 & ~new_n1640;
  assign new_n1642 = p_293_112_ & ~p_302_114_;
  assign new_n1643 = ~p_293_112_ & p_302_114_;
  assign new_n1644 = ~new_n1642 & ~new_n1643;
  assign new_n1645 = new_n1641 & ~new_n1644;
  assign new_n1646 = ~new_n1641 & new_n1644;
  assign new_n1647 = ~new_n1645 & ~new_n1646;
  assign new_n1648 = ~p_369_131_ & p_361_129_;
  assign new_n1649 = p_369_131_ & ~p_361_129_;
  assign new_n1650 = ~new_n1648 & ~new_n1649;
  assign new_n1651 = ~p_351_127_ & p_341_125_;
  assign new_n1652 = p_351_127_ & ~p_341_125_;
  assign new_n1653 = ~new_n1651 & ~new_n1652;
  assign new_n1654 = ~p_324_120_ & ~new_n1650;
  assign new_n1655 = ~new_n1653 & new_n1654;
  assign new_n1656 = p_324_120_ & ~new_n1653;
  assign new_n1657 = new_n1650 & new_n1656;
  assign new_n1658 = ~new_n1655 & ~new_n1657;
  assign new_n1659 = ~p_324_120_ & new_n1650;
  assign new_n1660 = new_n1653 & new_n1659;
  assign new_n1661 = p_324_120_ & new_n1653;
  assign new_n1662 = ~new_n1650 & new_n1661;
  assign new_n1663 = ~new_n1660 & ~new_n1662;
  assign new_n1664 = new_n1658 & new_n1663;
  assign new_n1665 = new_n1647 & ~new_n1664;
  assign new_n1666 = ~new_n1647 & new_n1664;
  assign p_1002_1920_ = new_n1665 | new_n1666;
  assign new_n1668 = ~p_226_93_ & p_218_91_;
  assign new_n1669 = p_226_93_ & ~p_218_91_;
  assign new_n1670 = ~new_n1668 & ~new_n1669;
  assign new_n1671 = ~p_210_89_ & p_206_87_;
  assign new_n1672 = p_210_89_ & ~p_206_87_;
  assign new_n1673 = ~new_n1671 & ~new_n1672;
  assign new_n1674 = new_n1670 & ~new_n1673;
  assign new_n1675 = ~new_n1670 & new_n1673;
  assign new_n1676 = ~new_n1674 & ~new_n1675;
  assign new_n1677 = ~p_289_110_ & p_281_108_;
  assign new_n1678 = p_289_110_ & ~p_281_108_;
  assign new_n1679 = ~new_n1677 & ~new_n1678;
  assign new_n1680 = ~p_257_102_ & p_234_95_;
  assign new_n1681 = p_257_102_ & ~p_234_95_;
  assign new_n1682 = ~new_n1680 & ~new_n1681;
  assign new_n1683 = ~p_273_106_ & p_265_104_;
  assign new_n1684 = p_273_106_ & ~p_265_104_;
  assign new_n1685 = ~new_n1683 & ~new_n1684;
  assign new_n1686 = ~new_n1679 & ~new_n1682;
  assign new_n1687 = ~new_n1685 & new_n1686;
  assign new_n1688 = new_n1682 & ~new_n1685;
  assign new_n1689 = new_n1679 & new_n1688;
  assign new_n1690 = ~new_n1687 & ~new_n1689;
  assign new_n1691 = new_n1679 & ~new_n1682;
  assign new_n1692 = new_n1685 & new_n1691;
  assign new_n1693 = new_n1682 & new_n1685;
  assign new_n1694 = ~new_n1679 & new_n1693;
  assign new_n1695 = ~new_n1692 & ~new_n1694;
  assign new_n1696 = new_n1690 & new_n1695;
  assign new_n1697 = new_n1676 & ~new_n1696;
  assign new_n1698 = ~new_n1676 & new_n1696;
  assign p_1004_1977_ = new_n1697 | new_n1698;
  assign new_n1700 = p_146_67_ & new_n390;
  assign new_n1701 = new_n418 & ~p_873_2124_;
  assign new_n1702 = p_149_68_ & new_n420;
  assign new_n1703 = new_n451 & ~p_834_2123_;
  assign new_n1704 = ~new_n1700 & ~new_n1701;
  assign new_n1705 = ~new_n1702 & new_n1704;
  assign new_n1706 = ~new_n1703 & new_n1705;
  assign p_670_2225_ = p_137_63_ & ~new_n1706;
  assign new_n1708 = p_106_40_ & new_n1285;
  assign new_n1709 = ~p_863_2276_ & new_n1287;
  assign new_n1710 = p_109_41_ & new_n1289;
  assign new_n1711 = ~p_824_2274_ & new_n1291;
  assign new_n1712 = ~new_n1708 & ~new_n1709;
  assign new_n1713 = ~new_n1710 & new_n1712;
  assign p_712_2297_ = new_n1711 | ~new_n1713;
  assign new_n1715 = p_2358_162_ & p_809_655_;
  assign new_n1716 = p_2358_162_ & ~p_809_655_;
  assign new_n1717 = p_80_28_ & new_n1716;
  assign new_n1718 = ~p_2358_162_ & p_809_655_;
  assign new_n1719 = ~p_2358_162_ & ~p_809_655_;
  assign new_n1720 = p_82_30_ & new_n1719;
  assign new_n1721 = ~new_n1715 & ~new_n1717;
  assign new_n1722 = ~new_n1718 & new_n1721;
  assign new_n1723 = ~new_n1720 & new_n1722;
  assign p_715_1278_ = p_141_65_ & ~new_n1723;
  assign new_n1725 = new_n400 & ~new_n938;
  assign new_n1726 = p_120_50_ & new_n402;
  assign new_n1727 = new_n414 & new_n1029;
  assign new_n1728 = ~new_n1555 & ~new_n1725;
  assign new_n1729 = ~new_n1726 & new_n1728;
  assign p_843_2455_ = new_n1727 | ~new_n1729;
  assign new_n1731 = p_61_21_ & new_n1285;
  assign new_n1732 = ~p_861_2070_ & new_n1287;
  assign new_n1733 = p_11_2_ & new_n1289;
  assign new_n1734 = ~p_822_1933_ & new_n1291;
  assign new_n1735 = ~new_n1731 & ~new_n1732;
  assign new_n1736 = ~new_n1733 & new_n1735;
  assign p_859_2132_ = new_n1734 | ~new_n1736;
  assign p_810_356_ = p_145_66_ & p_141_65_;
  assign new_n1739 = p_170_75_ & new_n390;
  assign new_n1740 = new_n418 & ~p_871_2127_;
  assign new_n1741 = p_200_85_ & new_n420;
  assign new_n1742 = new_n451 & ~p_832_2133_;
  assign new_n1743 = ~new_n1739 & ~new_n1740;
  assign new_n1744 = ~new_n1741 & new_n1743;
  assign new_n1745 = ~new_n1742 & new_n1744;
  assign p_642_2222_ = p_137_63_ & ~new_n1745;
  assign new_n1747 = p_103_39_ & new_n1285;
  assign new_n1748 = ~p_867_2237_ & new_n1287;
  assign new_n1749 = p_100_38_ & new_n1289;
  assign new_n1750 = ~p_828_2233_ & new_n1291;
  assign new_n1751 = ~new_n1747 & ~new_n1748;
  assign new_n1752 = ~new_n1749 & new_n1751;
  assign p_777_2278_ = new_n1750 | ~new_n1752;
  assign p_626_1752_ = new_n838 & new_n1386;
  assign p_632_1692_ = new_n1115 & new_n1564;
  assign new_n1756 = p_173_76_ & new_n390;
  assign new_n1757 = new_n418 & ~p_869_2181_;
  assign new_n1758 = p_203_86_ & new_n420;
  assign new_n1759 = new_n451 & ~p_830_2182_;
  assign new_n1760 = ~new_n1756 & ~new_n1757;
  assign new_n1761 = ~new_n1758 & new_n1760;
  assign new_n1762 = ~new_n1759 & new_n1761;
  assign p_645_2271_ = p_137_63_ & ~new_n1762;
  assign new_n1764 = p_173_76_ & new_n457;
  assign new_n1765 = new_n733 & ~p_869_2181_;
  assign new_n1766 = p_203_86_ & new_n735;
  assign new_n1767 = new_n1034 & ~p_830_2182_;
  assign new_n1768 = ~new_n1764 & ~new_n1765;
  assign new_n1769 = ~new_n1766 & new_n1768;
  assign new_n1770 = ~new_n1767 & new_n1769;
  assign p_679_2272_ = p_137_63_ & ~new_n1770;
  assign new_n1772 = p_23_6_ & new_n1716;
  assign new_n1773 = p_79_27_ & new_n1719;
  assign new_n1774 = ~new_n1715 & ~new_n1772;
  assign new_n1775 = ~new_n1718 & new_n1774;
  assign new_n1776 = ~new_n1773 & new_n1775;
  assign p_707_1277_ = p_141_65_ & ~new_n1776;
  assign new_n1778 = p_103_39_ & new_n1250;
  assign new_n1779 = ~p_867_2237_ & new_n1252;
  assign new_n1780 = p_100_38_ & new_n1254;
  assign new_n1781 = ~p_828_2233_ & new_n1256;
  assign new_n1782 = ~new_n1778 & ~new_n1779;
  assign new_n1783 = ~new_n1780 & new_n1782;
  assign p_737_2279_ = new_n1781 | ~new_n1783;
  assign new_n1785 = p_40_14_ & new_n1285;
  assign new_n1786 = ~p_869_2181_ & new_n1287;
  assign new_n1787 = p_91_35_ & new_n1289;
  assign new_n1788 = new_n1291 & ~p_830_2182_;
  assign new_n1789 = ~new_n1785 & ~new_n1786;
  assign new_n1790 = ~new_n1787 & new_n1789;
  assign p_782_2239_ = new_n1788 | ~new_n1790;
  assign new_n1792 = p_37_13_ & new_n1250;
  assign new_n1793 = new_n1252 & ~p_871_2127_;
  assign new_n1794 = p_43_15_ & new_n1254;
  assign new_n1795 = new_n1256 & ~p_832_2133_;
  assign new_n1796 = ~new_n1792 & ~new_n1793;
  assign new_n1797 = ~new_n1794 & new_n1796;
  assign p_747_2187_ = new_n1795 | ~new_n1797;
  assign p_845_845_ = p_2824_163_ | ~p_27_10_;
  assign new_n1800 = new_n1371 & new_n1605;
  assign new_n1801 = new_n435 & new_n1800;
  assign new_n1802 = new_n1068 & new_n1801;
  assign new_n1803 = new_n1244 & new_n1802;
  assign new_n1804 = new_n1427 & new_n1803;
  assign new_n1805 = p_623_2152_ & new_n1804;
  assign new_n1806 = new_n1486 & new_n1805;
  assign p_585_2236_ = new_n1231 & new_n1806;
  assign new_n1808 = p_81_29_ & new_n1716;
  assign new_n1809 = p_26_9_ & new_n1719;
  assign new_n1810 = ~new_n1715 & ~new_n1808;
  assign new_n1811 = ~new_n1718 & new_n1810;
  assign new_n1812 = ~new_n1809 & new_n1811;
  assign p_673_1276_ = p_141_65_ & ~new_n1812;
  assign new_n1814 = p_49_17_ & new_n1250;
  assign new_n1815 = new_n1252 & ~p_865_2277_;
  assign new_n1816 = p_46_16_ & new_n1254;
  assign new_n1817 = new_n1256 & ~p_826_2275_;
  assign new_n1818 = ~new_n1814 & ~new_n1815;
  assign new_n1819 = ~new_n1816 & new_n1818;
  assign p_732_2300_ = new_n1817 | ~new_n1819;
  assign new_n1821 = ~new_n862 & new_n868;
  assign new_n1822 = new_n862 & ~new_n868;
  assign new_n1823 = ~new_n1821 & ~new_n1822;
  assign new_n1824 = new_n856 & ~new_n859;
  assign new_n1825 = ~new_n1095 & ~new_n1824;
  assign new_n1826 = new_n1823 & ~new_n1825;
  assign new_n1827 = ~new_n1823 & new_n1825;
  assign new_n1828 = ~new_n1826 & ~new_n1827;
  assign new_n1829 = ~new_n424 & new_n745;
  assign new_n1830 = new_n424 & ~new_n745;
  assign new_n1831 = ~new_n1829 & ~new_n1830;
  assign new_n1832 = new_n739 & ~new_n751;
  assign new_n1833 = ~new_n739 & new_n751;
  assign new_n1834 = ~new_n1832 & ~new_n1833;
  assign new_n1835 = p_332_122_ & p_372_132_;
  assign new_n1836 = p_369_131_ & ~p_332_122_;
  assign new_n1837 = ~new_n1835 & ~new_n1836;
  assign new_n1838 = new_n430 & ~new_n1837;
  assign new_n1839 = ~new_n430 & new_n1837;
  assign new_n1840 = ~new_n1838 & ~new_n1839;
  assign new_n1841 = ~new_n1831 & ~new_n1834;
  assign new_n1842 = ~new_n1840 & new_n1841;
  assign new_n1843 = new_n1834 & ~new_n1840;
  assign new_n1844 = new_n1831 & new_n1843;
  assign new_n1845 = ~new_n1842 & ~new_n1844;
  assign new_n1846 = new_n1831 & ~new_n1834;
  assign new_n1847 = new_n1840 & new_n1846;
  assign new_n1848 = new_n1834 & new_n1840;
  assign new_n1849 = ~new_n1831 & new_n1848;
  assign new_n1850 = ~new_n1847 & ~new_n1849;
  assign new_n1851 = new_n1845 & new_n1850;
  assign new_n1852 = new_n1828 & ~new_n1851;
  assign new_n1853 = ~new_n1828 & new_n1851;
  assign p_998_2163_ = new_n1852 | new_n1853;
  assign new_n1855 = ~p_1002_1920_ & ~p_1004_1977_;
  assign new_n1856 = ~p_998_2163_ & new_n1855;
  assign new_n1857 = ~p_1000_2168_ & new_n1856;
  assign new_n1858 = p_562_155_ & new_n1857;
  assign new_n1859 = p_559_154_ & p_552_152_;
  assign new_n1860 = p_556_153_ & new_n1859;
  assign new_n1861 = p_386_135_ & new_n1860;
  assign new_n1862 = p_245_98_ & new_n1858;
  assign p_854_2268_ = new_n1861 & new_n1862;
  assign new_n1864 = p_20_5_ & new_n1250;
  assign new_n1865 = new_n1252 & ~p_873_2124_;
  assign new_n1866 = p_76_26_ & new_n1254;
  assign new_n1867 = new_n1256 & ~p_834_2123_;
  assign new_n1868 = ~new_n1864 & ~new_n1865;
  assign new_n1869 = ~new_n1866 & new_n1868;
  assign p_752_2189_ = new_n1867 | ~new_n1869;
  assign new_n1871 = ~new_n413 & ~new_n1358;
  assign new_n1872 = ~new_n1057 & new_n1871;
  assign new_n1873 = ~new_n1275 & new_n1872;
  assign new_n1874 = ~new_n1193 & ~new_n1411;
  assign new_n1875 = ~new_n1217 & new_n1874;
  assign new_n1876 = ~new_n1589 & new_n1875;
  assign new_n1877 = ~new_n653 & new_n1873;
  assign p_610_1519_ = new_n1876 & new_n1877;
  assign new_n1879 = ~p_623_2152_ & ~new_n1168;
  assign new_n1880 = ~p_623_2152_ & ~new_n1879;
  assign new_n1881 = ~new_n1168 & ~new_n1879;
  assign p_813_2260_ = new_n1880 | new_n1881;
  assign new_n1883 = new_n1347 & new_n1578;
  assign new_n1884 = new_n399 & new_n1883;
  assign new_n1885 = new_n1046 & new_n1884;
  assign new_n1886 = new_n1264 & new_n1885;
  assign new_n1887 = new_n1400 & new_n1886;
  assign new_n1888 = new_n1126 & new_n1887;
  assign new_n1889 = new_n1182 & new_n1888;
  assign p_575_2240_ = new_n1206 & new_n1889;
  assign p_601_220_ = p_552_152_ & p_562_155_;
  assign new_n1892 = p_25_8_ & new_n1716;
  assign new_n1893 = p_24_7_ & new_n1719;
  assign new_n1894 = ~new_n1715 & ~new_n1892;
  assign new_n1895 = ~new_n1718 & new_n1894;
  assign new_n1896 = ~new_n1893 & new_n1895;
  assign p_639_1275_ = p_141_65_ & ~new_n1896;
  assign new_n1898 = p_164_73_ & new_n390;
  assign new_n1899 = new_n418 & ~p_865_2277_;
  assign new_n1900 = p_194_83_ & new_n420;
  assign new_n1901 = new_n451 & ~p_826_2275_;
  assign new_n1902 = ~new_n1898 & ~new_n1899;
  assign new_n1903 = ~new_n1900 & new_n1902;
  assign new_n1904 = ~new_n1901 & new_n1903;
  assign p_651_2314_ = p_137_63_ & ~new_n1904;
  assign p_656_621_ = ~p_140_64_ | p_809_655_;
  assign new_n1907 = p_70_24_ & new_n1250;
  assign new_n1908 = ~p_877_2126_ & new_n1252;
  assign new_n1909 = p_67_23_ & new_n1254;
  assign new_n1910 = ~p_838_2064_ & new_n1256;
  assign new_n1911 = ~new_n1907 & ~new_n1908;
  assign new_n1912 = ~new_n1909 & new_n1911;
  assign p_762_2184_ = new_n1910 | ~new_n1912;
  assign p_847_465_ = ~p_556_153_ | ~p_386_135_;
  assign p_604_223_ = ~p_545_150_;
  assign p_593_733_ = ~p_299_113_;
  assign p_600_259_ = ~p_366_130_;
  assign p_611_275_ = ~p_338_124_;
  assign p_606_407_ = ~p_549_151_;
  assign p_612_263_ = ~p_358_128_;
  assign p_849_219_ = ~p_552_152_;
  assign p_850_217_ = ~p_562_155_;
  assign p_599_269_ = ~p_348_126_;
  assign p_851_218_ = ~p_559_154_;
  assign p_848_330_ = ~p_245_98_;
  assign p_973_202_ = p_3173_164_;
  assign p_603_225_ = p_604_223_;
  assign p_921_664_ = p_1_0_;
  assign p_892_408_ = p_549_151_;
  assign p_949_852_ = p_1_0_;
  assign p_939_853_ = p_1_0_;
  assign p_594_224_ = p_604_223_;
  assign p_978_851_ = p_1_0_;
  assign p_926_624_ = p_137_63_;
  assign p_298_299_ = p_293_112_;
  assign p_602_222_ = p_606_407_;
  assign p_717_1282_ = p_704_1281_;
  assign p_887_528_ = p_299_113_;
  assign p_923_619_ = p_141_65_;
  assign p_144_354_ = p_141_65_;
  assign p_889_734_ = p_299_113_;
  assign p_993_850_ = p_1_0_;
endmodule


