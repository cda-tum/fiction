// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_, pv96_20_,
    pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_, pv32_18_,
    pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_, pv32_19_,
    pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_, pv131_1_,
    pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_, pv64_5_,
    pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_,
    pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_  );
  input  pv96_30_, pv96_31_, pv96_10_, pv96_21_, pv138_4_, pv96_11_,
    pv96_20_, pv138_3_, pv138_2_, pv131_18_, pv138_0_, pv131_19_, pv32_7_,
    pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv131_3_, pv131_29_, pv32_6_,
    pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv131_2_, pv131_28_, pv32_5_,
    pv131_1_, pv32_4_, pv131_0_, pv32_3_, pv64_4_, pv96_5_, pv32_2_,
    pv64_5_, pv96_4_, pv32_1_, pv64_2_, pv96_7_, pv32_0_, pv64_3_, pv96_6_,
    pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_, pv97_0_,
    pv131_21_, pv32_11_, pv32_20_, pv64_9_, pv64_18_, pv64_27_, pv96_0_,
    pv131_20_, pv32_12_, pv32_23_, pv32_30_, pv64_6_, pv64_15_, pv64_26_,
    pv96_3_, pv99_0_, pv131_9_, pv131_23_, pv134_0_, pv32_13_, pv32_22_,
    pv32_31_, pv64_7_, pv64_16_, pv64_25_, pv96_2_, pv98_0_, pv131_8_,
    pv131_22_, pv32_14_, pv32_25_, pv131_7_, pv131_25_, pv131_30_,
    pv133_1_, pv32_15_, pv32_24_, pv131_6_, pv131_24_, pv131_31_, pv133_0_,
    pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv131_5_, pv131_27_, pv32_8_,
    pv32_17_, pv32_26_, pv64_29_, pv131_4_, pv131_26_, pv64_20_, pv64_31_,
    pv96_16_, pv96_27_, pv131_16_, pv64_10_, pv96_17_, pv96_26_, pv131_17_,
    pv96_18_, pv96_29_, pv131_14_, pv96_19_, pv96_28_, pv131_15_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv131_12_, pv64_14_, pv64_23_, pv96_13_,
    pv96_22_, pv131_13_, pv64_11_, pv64_22_, pv96_14_, pv96_25_, pv131_10_,
    pv64_12_, pv64_21_, pv64_30_, pv96_15_, pv96_24_, pv131_11_;
  output pv198_17_, pv205_3_, pv198_16_, pv205_4_, pv198_19_, pv205_5_,
    pv198_18_, pv205_6_, pv198_8_, pv198_13_, pv198_7_, pv198_12_,
    pv205_0_, pv198_15_, pv205_1_, pv198_9_, pv198_14_, pv205_2_, pv166_7_,
    pv166_10_, pv166_23_, pv198_4_, pv198_22_, pv166_8_, pv166_24_,
    pv198_3_, pv198_23_, pv166_5_, pv166_21_, pv198_6_, pv198_24_,
    pv166_6_, pv166_22_, pv198_5_, pv198_25_, pv166_14_, pv198_0_,
    pv198_26_, pv166_13_, pv166_20_, pv198_27_, pv166_9_, pv166_12_,
    pv198_2_, pv198_28_, pv166_11_, pv198_1_, pv198_29_, pv166_18_,
    pv166_0_, pv166_17_, pv166_16_, pv166_15_, pv166_3_, pv166_27_,
    pv198_31_, pv166_4_, pv198_30_, pv166_1_, pv166_25_, pv198_20_,
    pv166_2_, pv166_19_, pv166_26_, pv198_21_, pv198_11_, pv198_10_;
  wire new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n230, new_n231, new_n232, new_n233, new_n234, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n289, new_n290, new_n291, new_n292, new_n293, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n333, new_n334, new_n335, new_n336,
    new_n338, new_n339, new_n340, new_n341, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n355, new_n356, new_n357, new_n358, new_n360, new_n361, new_n362,
    new_n363, new_n365, new_n366, new_n367, new_n368, new_n369, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n377, new_n378, new_n379,
    new_n380, new_n382, new_n383, new_n384, new_n385, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n399, new_n400, new_n401, new_n402, new_n404, new_n405,
    new_n406, new_n407, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n421, new_n422,
    new_n423, new_n424, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n438, new_n439,
    new_n440, new_n441, new_n443, new_n444, new_n445, new_n446, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n454, new_n455, new_n456,
    new_n457, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n476, new_n477, new_n478, new_n479, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n493, new_n494, new_n495, new_n496, new_n498, new_n499,
    new_n500, new_n501, new_n503, new_n504, new_n505, new_n506, new_n508,
    new_n509, new_n510, new_n511, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592;
  assign new_n206 = pv138_4_ & ~pv138_0_;
  assign new_n207 = ~pv138_2_ & new_n206;
  assign new_n208 = pv96_13_ & new_n207;
  assign new_n209 = pv138_4_ & pv138_0_;
  assign new_n210 = pv138_2_ & new_n209;
  assign new_n211 = ~pv131_13_ & new_n210;
  assign new_n212 = ~pv138_2_ & new_n209;
  assign new_n213 = pv131_13_ & new_n212;
  assign new_n214 = ~pv138_4_ & pv138_2_;
  assign new_n215 = ~new_n208 & ~new_n211;
  assign new_n216 = ~new_n213 & ~new_n214;
  assign pv198_17_ = ~new_n215 | ~new_n216;
  assign new_n218 = pv138_3_ & ~pv138_0_;
  assign new_n219 = ~pv138_2_ & new_n218;
  assign new_n220 = pv96_31_ & new_n219;
  assign new_n221 = pv138_3_ & pv138_0_;
  assign new_n222 = pv138_2_ & new_n221;
  assign new_n223 = ~pv131_31_ & new_n222;
  assign new_n224 = ~pv138_2_ & new_n221;
  assign new_n225 = pv131_31_ & new_n224;
  assign new_n226 = ~pv138_3_ & pv138_2_;
  assign new_n227 = ~new_n220 & ~new_n223;
  assign new_n228 = ~new_n225 & ~new_n226;
  assign pv205_3_ = ~new_n227 | ~new_n228;
  assign new_n230 = pv96_12_ & new_n207;
  assign new_n231 = ~pv131_12_ & new_n210;
  assign new_n232 = pv131_12_ & new_n212;
  assign new_n233 = ~new_n230 & ~new_n231;
  assign new_n234 = ~new_n214 & ~new_n232;
  assign pv198_16_ = ~new_n233 | ~new_n234;
  assign new_n236 = pv97_0_ & new_n219;
  assign new_n237 = ~pv133_0_ & new_n222;
  assign new_n238 = pv133_0_ & new_n224;
  assign new_n239 = ~new_n236 & ~new_n237;
  assign new_n240 = ~new_n226 & ~new_n238;
  assign pv205_4_ = ~new_n239 | ~new_n240;
  assign new_n242 = pv96_15_ & new_n207;
  assign new_n243 = ~pv131_15_ & new_n210;
  assign new_n244 = pv131_15_ & new_n212;
  assign new_n245 = ~new_n242 & ~new_n243;
  assign new_n246 = ~new_n214 & ~new_n244;
  assign pv198_19_ = ~new_n245 | ~new_n246;
  assign new_n248 = pv98_0_ & new_n219;
  assign new_n249 = ~pv133_1_ & new_n222;
  assign new_n250 = pv133_1_ & new_n224;
  assign new_n251 = ~new_n248 & ~new_n249;
  assign new_n252 = ~new_n226 & ~new_n250;
  assign pv205_5_ = ~new_n251 | ~new_n252;
  assign new_n254 = pv96_14_ & new_n207;
  assign new_n255 = ~pv131_14_ & new_n210;
  assign new_n256 = pv131_14_ & new_n212;
  assign new_n257 = ~new_n254 & ~new_n255;
  assign new_n258 = ~new_n214 & ~new_n256;
  assign pv198_18_ = ~new_n257 | ~new_n258;
  assign new_n260 = pv134_0_ & new_n224;
  assign new_n261 = pv99_0_ & new_n219;
  assign new_n262 = pv134_0_ & new_n222;
  assign new_n263 = ~new_n260 & ~new_n261;
  assign pv205_6_ = new_n262 | ~new_n263;
  assign new_n265 = pv96_4_ & new_n207;
  assign new_n266 = ~pv131_4_ & new_n210;
  assign new_n267 = pv131_4_ & new_n212;
  assign new_n268 = ~new_n265 & ~new_n266;
  assign new_n269 = ~new_n214 & ~new_n267;
  assign pv198_8_ = ~new_n268 | ~new_n269;
  assign new_n271 = pv96_9_ & new_n207;
  assign new_n272 = ~pv131_9_ & new_n210;
  assign new_n273 = pv131_9_ & new_n212;
  assign new_n274 = ~new_n271 & ~new_n272;
  assign new_n275 = ~new_n214 & ~new_n273;
  assign pv198_13_ = ~new_n274 | ~new_n275;
  assign new_n277 = pv96_3_ & new_n207;
  assign new_n278 = ~pv131_3_ & new_n210;
  assign new_n279 = pv131_3_ & new_n212;
  assign new_n280 = ~new_n277 & ~new_n278;
  assign new_n281 = ~new_n214 & ~new_n279;
  assign pv198_7_ = ~new_n280 | ~new_n281;
  assign new_n283 = pv96_8_ & new_n207;
  assign new_n284 = ~pv131_8_ & new_n210;
  assign new_n285 = pv131_8_ & new_n212;
  assign new_n286 = ~new_n283 & ~new_n284;
  assign new_n287 = ~new_n214 & ~new_n285;
  assign pv198_12_ = ~new_n286 | ~new_n287;
  assign new_n289 = pv96_28_ & new_n219;
  assign new_n290 = ~pv131_28_ & new_n222;
  assign new_n291 = pv131_28_ & new_n224;
  assign new_n292 = ~new_n289 & ~new_n290;
  assign new_n293 = ~new_n226 & ~new_n291;
  assign pv205_0_ = ~new_n292 | ~new_n293;
  assign new_n295 = pv96_11_ & new_n207;
  assign new_n296 = ~pv131_11_ & new_n210;
  assign new_n297 = pv131_11_ & new_n212;
  assign new_n298 = ~new_n295 & ~new_n296;
  assign new_n299 = ~new_n214 & ~new_n297;
  assign pv198_15_ = ~new_n298 | ~new_n299;
  assign new_n301 = pv96_29_ & new_n219;
  assign new_n302 = ~pv131_29_ & new_n222;
  assign new_n303 = pv131_29_ & new_n224;
  assign new_n304 = ~new_n301 & ~new_n302;
  assign new_n305 = ~new_n226 & ~new_n303;
  assign pv205_1_ = ~new_n304 | ~new_n305;
  assign new_n307 = pv96_5_ & new_n207;
  assign new_n308 = ~pv131_5_ & new_n210;
  assign new_n309 = pv131_5_ & new_n212;
  assign new_n310 = ~new_n307 & ~new_n308;
  assign new_n311 = ~new_n214 & ~new_n309;
  assign pv198_9_ = ~new_n310 | ~new_n311;
  assign new_n313 = pv96_10_ & new_n207;
  assign new_n314 = ~pv131_10_ & new_n210;
  assign new_n315 = pv131_10_ & new_n212;
  assign new_n316 = ~new_n313 & ~new_n314;
  assign new_n317 = ~new_n214 & ~new_n315;
  assign pv198_14_ = ~new_n316 | ~new_n317;
  assign new_n319 = pv96_30_ & new_n219;
  assign new_n320 = ~pv131_30_ & new_n222;
  assign new_n321 = pv131_30_ & new_n224;
  assign new_n322 = ~new_n319 & ~new_n320;
  assign new_n323 = ~new_n226 & ~new_n321;
  assign pv205_2_ = ~new_n322 | ~new_n323;
  assign new_n325 = ~pv138_2_ & pv138_0_;
  assign new_n326 = pv64_7_ & new_n325;
  assign new_n327 = ~pv138_2_ & ~pv138_0_;
  assign new_n328 = pv32_7_ & new_n327;
  assign new_n329 = pv138_2_ & pv138_0_;
  assign new_n330 = ~pv64_7_ & new_n329;
  assign new_n331 = ~new_n326 & ~new_n328;
  assign pv166_7_ = new_n330 | ~new_n331;
  assign new_n333 = pv64_10_ & new_n325;
  assign new_n334 = pv32_10_ & new_n327;
  assign new_n335 = ~pv64_10_ & new_n329;
  assign new_n336 = ~new_n333 & ~new_n334;
  assign pv166_10_ = new_n335 | ~new_n336;
  assign new_n338 = pv64_23_ & new_n325;
  assign new_n339 = pv32_23_ & new_n327;
  assign new_n340 = ~pv64_23_ & new_n329;
  assign new_n341 = ~new_n338 & ~new_n339;
  assign pv166_23_ = new_n340 | ~new_n341;
  assign new_n343 = pv96_0_ & new_n207;
  assign new_n344 = ~pv131_0_ & new_n210;
  assign new_n345 = pv131_0_ & new_n212;
  assign new_n346 = ~new_n343 & ~new_n344;
  assign new_n347 = ~new_n214 & ~new_n345;
  assign pv198_4_ = ~new_n346 | ~new_n347;
  assign new_n349 = pv96_18_ & new_n207;
  assign new_n350 = ~pv131_18_ & new_n210;
  assign new_n351 = pv131_18_ & new_n212;
  assign new_n352 = ~new_n349 & ~new_n350;
  assign new_n353 = ~new_n214 & ~new_n351;
  assign pv198_22_ = ~new_n352 | ~new_n353;
  assign new_n355 = pv64_8_ & new_n325;
  assign new_n356 = pv32_8_ & new_n327;
  assign new_n357 = ~pv64_8_ & new_n329;
  assign new_n358 = ~new_n355 & ~new_n356;
  assign pv166_8_ = new_n357 | ~new_n358;
  assign new_n360 = pv64_24_ & new_n325;
  assign new_n361 = pv32_24_ & new_n327;
  assign new_n362 = ~pv64_24_ & new_n329;
  assign new_n363 = ~new_n360 & ~new_n361;
  assign pv166_24_ = new_n362 | ~new_n363;
  assign new_n365 = pv32_31_ & new_n207;
  assign new_n366 = ~pv64_31_ & new_n210;
  assign new_n367 = pv64_31_ & new_n212;
  assign new_n368 = ~new_n365 & ~new_n366;
  assign new_n369 = ~new_n214 & ~new_n367;
  assign pv198_3_ = ~new_n368 | ~new_n369;
  assign new_n371 = pv96_19_ & new_n207;
  assign new_n372 = ~pv131_19_ & new_n210;
  assign new_n373 = pv131_19_ & new_n212;
  assign new_n374 = ~new_n371 & ~new_n372;
  assign new_n375 = ~new_n214 & ~new_n373;
  assign pv198_23_ = ~new_n374 | ~new_n375;
  assign new_n377 = pv64_5_ & new_n325;
  assign new_n378 = pv32_5_ & new_n327;
  assign new_n379 = ~pv64_5_ & new_n329;
  assign new_n380 = ~new_n377 & ~new_n378;
  assign pv166_5_ = new_n379 | ~new_n380;
  assign new_n382 = pv64_21_ & new_n325;
  assign new_n383 = pv32_21_ & new_n327;
  assign new_n384 = ~pv64_21_ & new_n329;
  assign new_n385 = ~new_n382 & ~new_n383;
  assign pv166_21_ = new_n384 | ~new_n385;
  assign new_n387 = pv96_2_ & new_n207;
  assign new_n388 = ~pv131_2_ & new_n210;
  assign new_n389 = pv131_2_ & new_n212;
  assign new_n390 = ~new_n387 & ~new_n388;
  assign new_n391 = ~new_n214 & ~new_n389;
  assign pv198_6_ = ~new_n390 | ~new_n391;
  assign new_n393 = pv96_20_ & new_n207;
  assign new_n394 = ~pv131_20_ & new_n210;
  assign new_n395 = pv131_20_ & new_n212;
  assign new_n396 = ~new_n393 & ~new_n394;
  assign new_n397 = ~new_n214 & ~new_n395;
  assign pv198_24_ = ~new_n396 | ~new_n397;
  assign new_n399 = pv64_6_ & new_n325;
  assign new_n400 = pv32_6_ & new_n327;
  assign new_n401 = ~pv64_6_ & new_n329;
  assign new_n402 = ~new_n399 & ~new_n400;
  assign pv166_6_ = new_n401 | ~new_n402;
  assign new_n404 = pv64_22_ & new_n325;
  assign new_n405 = pv32_22_ & new_n327;
  assign new_n406 = ~pv64_22_ & new_n329;
  assign new_n407 = ~new_n404 & ~new_n405;
  assign pv166_22_ = new_n406 | ~new_n407;
  assign new_n409 = pv96_1_ & new_n207;
  assign new_n410 = ~pv131_1_ & new_n210;
  assign new_n411 = pv131_1_ & new_n212;
  assign new_n412 = ~new_n409 & ~new_n410;
  assign new_n413 = ~new_n214 & ~new_n411;
  assign pv198_5_ = ~new_n412 | ~new_n413;
  assign new_n415 = pv96_21_ & new_n207;
  assign new_n416 = ~pv131_21_ & new_n210;
  assign new_n417 = pv131_21_ & new_n212;
  assign new_n418 = ~new_n415 & ~new_n416;
  assign new_n419 = ~new_n214 & ~new_n417;
  assign pv198_25_ = ~new_n418 | ~new_n419;
  assign new_n421 = pv64_14_ & new_n325;
  assign new_n422 = pv32_14_ & new_n327;
  assign new_n423 = ~pv64_14_ & new_n329;
  assign new_n424 = ~new_n421 & ~new_n422;
  assign pv166_14_ = new_n423 | ~new_n424;
  assign new_n426 = pv32_28_ & new_n207;
  assign new_n427 = ~pv64_28_ & new_n210;
  assign new_n428 = pv64_28_ & new_n212;
  assign new_n429 = ~new_n426 & ~new_n427;
  assign new_n430 = ~new_n214 & ~new_n428;
  assign pv198_0_ = ~new_n429 | ~new_n430;
  assign new_n432 = pv96_22_ & new_n207;
  assign new_n433 = ~pv131_22_ & new_n210;
  assign new_n434 = pv131_22_ & new_n212;
  assign new_n435 = ~new_n432 & ~new_n433;
  assign new_n436 = ~new_n214 & ~new_n434;
  assign pv198_26_ = ~new_n435 | ~new_n436;
  assign new_n438 = pv64_13_ & new_n325;
  assign new_n439 = pv32_13_ & new_n327;
  assign new_n440 = ~pv64_13_ & new_n329;
  assign new_n441 = ~new_n438 & ~new_n439;
  assign pv166_13_ = new_n440 | ~new_n441;
  assign new_n443 = pv64_20_ & new_n325;
  assign new_n444 = pv32_20_ & new_n327;
  assign new_n445 = ~pv64_20_ & new_n329;
  assign new_n446 = ~new_n443 & ~new_n444;
  assign pv166_20_ = new_n445 | ~new_n446;
  assign new_n448 = pv96_23_ & new_n207;
  assign new_n449 = ~pv131_23_ & new_n210;
  assign new_n450 = pv131_23_ & new_n212;
  assign new_n451 = ~new_n448 & ~new_n449;
  assign new_n452 = ~new_n214 & ~new_n450;
  assign pv198_27_ = ~new_n451 | ~new_n452;
  assign new_n454 = pv64_9_ & new_n325;
  assign new_n455 = pv32_9_ & new_n327;
  assign new_n456 = ~pv64_9_ & new_n329;
  assign new_n457 = ~new_n454 & ~new_n455;
  assign pv166_9_ = new_n456 | ~new_n457;
  assign new_n459 = pv64_12_ & new_n325;
  assign new_n460 = pv32_12_ & new_n327;
  assign new_n461 = ~pv64_12_ & new_n329;
  assign new_n462 = ~new_n459 & ~new_n460;
  assign pv166_12_ = new_n461 | ~new_n462;
  assign new_n464 = pv32_30_ & new_n207;
  assign new_n465 = ~pv64_30_ & new_n210;
  assign new_n466 = pv64_30_ & new_n212;
  assign new_n467 = ~new_n464 & ~new_n465;
  assign new_n468 = ~new_n214 & ~new_n466;
  assign pv198_2_ = ~new_n467 | ~new_n468;
  assign new_n470 = pv96_24_ & new_n207;
  assign new_n471 = ~pv131_24_ & new_n210;
  assign new_n472 = pv131_24_ & new_n212;
  assign new_n473 = ~new_n470 & ~new_n471;
  assign new_n474 = ~new_n214 & ~new_n472;
  assign pv198_28_ = ~new_n473 | ~new_n474;
  assign new_n476 = pv64_11_ & new_n325;
  assign new_n477 = pv32_11_ & new_n327;
  assign new_n478 = ~pv64_11_ & new_n329;
  assign new_n479 = ~new_n476 & ~new_n477;
  assign pv166_11_ = new_n478 | ~new_n479;
  assign new_n481 = pv32_29_ & new_n207;
  assign new_n482 = ~pv64_29_ & new_n210;
  assign new_n483 = pv64_29_ & new_n212;
  assign new_n484 = ~new_n481 & ~new_n482;
  assign new_n485 = ~new_n214 & ~new_n483;
  assign pv198_1_ = ~new_n484 | ~new_n485;
  assign new_n487 = pv96_25_ & new_n207;
  assign new_n488 = ~pv131_25_ & new_n210;
  assign new_n489 = pv131_25_ & new_n212;
  assign new_n490 = ~new_n487 & ~new_n488;
  assign new_n491 = ~new_n214 & ~new_n489;
  assign pv198_29_ = ~new_n490 | ~new_n491;
  assign new_n493 = pv64_18_ & new_n325;
  assign new_n494 = pv32_18_ & new_n327;
  assign new_n495 = ~pv64_18_ & new_n329;
  assign new_n496 = ~new_n493 & ~new_n494;
  assign pv166_18_ = new_n495 | ~new_n496;
  assign new_n498 = pv64_0_ & new_n325;
  assign new_n499 = pv32_0_ & new_n327;
  assign new_n500 = ~pv64_0_ & new_n329;
  assign new_n501 = ~new_n498 & ~new_n499;
  assign pv166_0_ = new_n500 | ~new_n501;
  assign new_n503 = pv64_17_ & new_n325;
  assign new_n504 = pv32_17_ & new_n327;
  assign new_n505 = ~pv64_17_ & new_n329;
  assign new_n506 = ~new_n503 & ~new_n504;
  assign pv166_17_ = new_n505 | ~new_n506;
  assign new_n508 = pv64_16_ & new_n325;
  assign new_n509 = pv32_16_ & new_n327;
  assign new_n510 = ~pv64_16_ & new_n329;
  assign new_n511 = ~new_n508 & ~new_n509;
  assign pv166_16_ = new_n510 | ~new_n511;
  assign new_n513 = pv64_15_ & new_n325;
  assign new_n514 = pv32_15_ & new_n327;
  assign new_n515 = ~pv64_15_ & new_n329;
  assign new_n516 = ~new_n513 & ~new_n514;
  assign pv166_15_ = new_n515 | ~new_n516;
  assign new_n518 = pv64_3_ & new_n325;
  assign new_n519 = pv32_3_ & new_n327;
  assign new_n520 = ~pv64_3_ & new_n329;
  assign new_n521 = ~new_n518 & ~new_n519;
  assign pv166_3_ = new_n520 | ~new_n521;
  assign new_n523 = pv64_27_ & new_n325;
  assign new_n524 = pv32_27_ & new_n327;
  assign new_n525 = ~pv64_27_ & new_n329;
  assign new_n526 = ~new_n523 & ~new_n524;
  assign pv166_27_ = new_n525 | ~new_n526;
  assign new_n528 = pv96_27_ & new_n207;
  assign new_n529 = ~pv131_27_ & new_n210;
  assign new_n530 = pv131_27_ & new_n212;
  assign new_n531 = ~new_n528 & ~new_n529;
  assign new_n532 = ~new_n214 & ~new_n530;
  assign pv198_31_ = ~new_n531 | ~new_n532;
  assign new_n534 = pv64_4_ & new_n325;
  assign new_n535 = pv32_4_ & new_n327;
  assign new_n536 = ~pv64_4_ & new_n329;
  assign new_n537 = ~new_n534 & ~new_n535;
  assign pv166_4_ = new_n536 | ~new_n537;
  assign new_n539 = pv96_26_ & new_n207;
  assign new_n540 = ~pv131_26_ & new_n210;
  assign new_n541 = pv131_26_ & new_n212;
  assign new_n542 = ~new_n539 & ~new_n540;
  assign new_n543 = ~new_n214 & ~new_n541;
  assign pv198_30_ = ~new_n542 | ~new_n543;
  assign new_n545 = pv64_1_ & new_n325;
  assign new_n546 = pv32_1_ & new_n327;
  assign new_n547 = ~pv64_1_ & new_n329;
  assign new_n548 = ~new_n545 & ~new_n546;
  assign pv166_1_ = new_n547 | ~new_n548;
  assign new_n550 = pv64_25_ & new_n325;
  assign new_n551 = pv32_25_ & new_n327;
  assign new_n552 = ~pv64_25_ & new_n329;
  assign new_n553 = ~new_n550 & ~new_n551;
  assign pv166_25_ = new_n552 | ~new_n553;
  assign new_n555 = pv96_16_ & new_n207;
  assign new_n556 = ~pv131_16_ & new_n210;
  assign new_n557 = pv131_16_ & new_n212;
  assign new_n558 = ~new_n555 & ~new_n556;
  assign new_n559 = ~new_n214 & ~new_n557;
  assign pv198_20_ = ~new_n558 | ~new_n559;
  assign new_n561 = pv64_2_ & new_n325;
  assign new_n562 = pv32_2_ & new_n327;
  assign new_n563 = ~pv64_2_ & new_n329;
  assign new_n564 = ~new_n561 & ~new_n562;
  assign pv166_2_ = new_n563 | ~new_n564;
  assign new_n566 = pv64_19_ & new_n325;
  assign new_n567 = pv32_19_ & new_n327;
  assign new_n568 = ~pv64_19_ & new_n329;
  assign new_n569 = ~new_n566 & ~new_n567;
  assign pv166_19_ = new_n568 | ~new_n569;
  assign new_n571 = pv64_26_ & new_n325;
  assign new_n572 = pv32_26_ & new_n327;
  assign new_n573 = ~pv64_26_ & new_n329;
  assign new_n574 = ~new_n571 & ~new_n572;
  assign pv166_26_ = new_n573 | ~new_n574;
  assign new_n576 = pv96_17_ & new_n207;
  assign new_n577 = ~pv131_17_ & new_n210;
  assign new_n578 = pv131_17_ & new_n212;
  assign new_n579 = ~new_n576 & ~new_n577;
  assign new_n580 = ~new_n214 & ~new_n578;
  assign pv198_21_ = ~new_n579 | ~new_n580;
  assign new_n582 = pv96_7_ & new_n207;
  assign new_n583 = ~pv131_7_ & new_n210;
  assign new_n584 = pv131_7_ & new_n212;
  assign new_n585 = ~new_n582 & ~new_n583;
  assign new_n586 = ~new_n214 & ~new_n584;
  assign pv198_11_ = ~new_n585 | ~new_n586;
  assign new_n588 = pv96_6_ & new_n207;
  assign new_n589 = ~pv131_6_ & new_n210;
  assign new_n590 = pv131_6_ & new_n212;
  assign new_n591 = ~new_n588 & ~new_n589;
  assign new_n592 = ~new_n214 & ~new_n590;
  assign pv198_10_ = ~new_n591 | ~new_n592;
endmodule


