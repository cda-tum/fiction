// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    _1gat_0_, _11gat_3_, _17gat_5_, _95gat_29_, _112gat_34_, _4gat_1_,
    _30gat_9_, _27gat_8_, _8gat_2_, _40gat_12_, _47gat_14_, _69gat_21_,
    _73gat_22_, _89gat_27_, _53gat_16_, _115gat_35_, _37gat_11_,
    _63gat_19_, _99gat_30_, _79gat_24_, _14gat_4_, _102gat_31_, _24gat_7_,
    _82gat_25_, _66gat_20_, _43gat_13_, _92gat_28_, _76gat_23_, _86gat_26_,
    _50gat_15_, _108gat_33_, _21gat_6_, _60gat_18_, _56gat_17_,
    _105gat_32_, _34gat_10_,
    _421gat_188_, _329gat_133_, _223gat_84_, _370gat_163_, _431gat_194_,
    _432gat_195_, _430gat_193_  );
  input  _1gat_0_, _11gat_3_, _17gat_5_, _95gat_29_, _112gat_34_,
    _4gat_1_, _30gat_9_, _27gat_8_, _8gat_2_, _40gat_12_, _47gat_14_,
    _69gat_21_, _73gat_22_, _89gat_27_, _53gat_16_, _115gat_35_,
    _37gat_11_, _63gat_19_, _99gat_30_, _79gat_24_, _14gat_4_, _102gat_31_,
    _24gat_7_, _82gat_25_, _66gat_20_, _43gat_13_, _92gat_28_, _76gat_23_,
    _86gat_26_, _50gat_15_, _108gat_33_, _21gat_6_, _60gat_18_, _56gat_17_,
    _105gat_32_, _34gat_10_;
  output _421gat_188_, _329gat_133_, _223gat_84_, _370gat_163_, _431gat_194_,
    _432gat_195_, _430gat_193_;
  wire new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50,
    new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58,
    new_n59, new_n60, new_n62, new_n63, new_n64, new_n65, new_n66, new_n67,
    new_n68, new_n69, new_n70, new_n71, new_n72, new_n73, new_n74, new_n75,
    new_n76, new_n77, new_n78, new_n79, new_n80, new_n81, new_n82, new_n83,
    new_n84, new_n85, new_n86, new_n87, new_n88, new_n89, new_n90, new_n91,
    new_n92, new_n93, new_n94, new_n95, new_n96, new_n97, new_n98, new_n99,
    new_n100, new_n101, new_n102, new_n103, new_n104, new_n105, new_n106,
    new_n107, new_n108, new_n109, new_n110, new_n111, new_n112, new_n114,
    new_n115, new_n116, new_n117, new_n118, new_n119, new_n120, new_n121,
    new_n122, new_n123, new_n124, new_n125, new_n126, new_n127, new_n128,
    new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n253, new_n254;
  assign new_n44 = ~_47gat_14_ & _43gat_13_;
  assign new_n45 = ~_37gat_11_ & _43gat_13_;
  assign new_n46 = ~_50gat_15_ & _56gat_17_;
  assign new_n47 = ~_11gat_3_ & _17gat_5_;
  assign new_n48 = _30gat_9_ & ~_24gat_7_;
  assign new_n49 = ~_1gat_0_ & _4gat_1_;
  assign new_n50 = _95gat_29_ & ~_89gat_27_;
  assign new_n51 = ~_102gat_31_ & _108gat_33_;
  assign new_n52 = _69gat_21_ & ~_63gat_19_;
  assign new_n53 = _82gat_25_ & ~_76gat_23_;
  assign new_n54 = ~new_n45 & ~new_n46;
  assign new_n55 = ~new_n47 & new_n54;
  assign new_n56 = ~new_n48 & new_n55;
  assign new_n57 = ~new_n49 & new_n56;
  assign new_n58 = ~new_n50 & new_n57;
  assign new_n59 = ~new_n51 & new_n58;
  assign new_n60 = ~new_n52 & new_n59;
  assign _223gat_84_ = new_n53 | ~new_n60;
  assign new_n62 = new_n45 & _223gat_84_;
  assign new_n63 = ~new_n45 & ~_223gat_84_;
  assign new_n64 = ~new_n62 & ~new_n63;
  assign new_n65 = new_n44 & ~new_n64;
  assign new_n66 = ~_60gat_18_ & _56gat_17_;
  assign new_n67 = new_n46 & _223gat_84_;
  assign new_n68 = ~new_n46 & ~_223gat_84_;
  assign new_n69 = ~new_n67 & ~new_n68;
  assign new_n70 = new_n66 & ~new_n69;
  assign new_n71 = _17gat_5_ & ~_21gat_6_;
  assign new_n72 = new_n47 & _223gat_84_;
  assign new_n73 = ~new_n47 & ~_223gat_84_;
  assign new_n74 = ~new_n72 & ~new_n73;
  assign new_n75 = new_n71 & ~new_n74;
  assign new_n76 = _30gat_9_ & ~_34gat_10_;
  assign new_n77 = new_n48 & _223gat_84_;
  assign new_n78 = ~new_n48 & ~_223gat_84_;
  assign new_n79 = ~new_n77 & ~new_n78;
  assign new_n80 = new_n76 & ~new_n79;
  assign new_n81 = _4gat_1_ & ~_8gat_2_;
  assign new_n82 = new_n49 & _223gat_84_;
  assign new_n83 = ~new_n49 & ~_223gat_84_;
  assign new_n84 = ~new_n82 & ~new_n83;
  assign new_n85 = new_n81 & ~new_n84;
  assign new_n86 = _95gat_29_ & ~_99gat_30_;
  assign new_n87 = new_n50 & _223gat_84_;
  assign new_n88 = ~new_n50 & ~_223gat_84_;
  assign new_n89 = ~new_n87 & ~new_n88;
  assign new_n90 = new_n86 & ~new_n89;
  assign new_n91 = ~_112gat_34_ & _108gat_33_;
  assign new_n92 = new_n51 & _223gat_84_;
  assign new_n93 = ~new_n51 & ~_223gat_84_;
  assign new_n94 = ~new_n92 & ~new_n93;
  assign new_n95 = new_n91 & ~new_n94;
  assign new_n96 = _69gat_21_ & ~_73gat_22_;
  assign new_n97 = new_n52 & _223gat_84_;
  assign new_n98 = ~new_n52 & ~_223gat_84_;
  assign new_n99 = ~new_n97 & ~new_n98;
  assign new_n100 = new_n96 & ~new_n99;
  assign new_n101 = _82gat_25_ & ~_86gat_26_;
  assign new_n102 = new_n53 & _223gat_84_;
  assign new_n103 = ~new_n53 & ~_223gat_84_;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = new_n101 & ~new_n104;
  assign new_n106 = ~new_n65 & ~new_n70;
  assign new_n107 = ~new_n75 & new_n106;
  assign new_n108 = ~new_n80 & new_n107;
  assign new_n109 = ~new_n85 & new_n108;
  assign new_n110 = ~new_n90 & new_n109;
  assign new_n111 = ~new_n95 & new_n110;
  assign new_n112 = ~new_n100 & new_n111;
  assign _329gat_133_ = new_n105 | ~new_n112;
  assign new_n114 = _60gat_18_ & _329gat_133_;
  assign new_n115 = ~_53gat_16_ & _43gat_13_;
  assign new_n116 = ~new_n64 & new_n115;
  assign new_n117 = new_n65 & _329gat_133_;
  assign new_n118 = ~new_n65 & ~_329gat_133_;
  assign new_n119 = ~new_n117 & ~new_n118;
  assign new_n120 = new_n116 & ~new_n119;
  assign new_n121 = ~_66gat_20_ & _56gat_17_;
  assign new_n122 = ~new_n69 & new_n121;
  assign new_n123 = new_n70 & _329gat_133_;
  assign new_n124 = ~new_n70 & ~_329gat_133_;
  assign new_n125 = ~new_n123 & ~new_n124;
  assign new_n126 = new_n122 & ~new_n125;
  assign new_n127 = _17gat_5_ & ~_27gat_8_;
  assign new_n128 = ~new_n74 & new_n127;
  assign new_n129 = new_n75 & _329gat_133_;
  assign new_n130 = ~new_n75 & ~_329gat_133_;
  assign new_n131 = ~new_n129 & ~new_n130;
  assign new_n132 = new_n128 & ~new_n131;
  assign new_n133 = _30gat_9_ & ~_40gat_12_;
  assign new_n134 = ~new_n79 & new_n133;
  assign new_n135 = new_n80 & _329gat_133_;
  assign new_n136 = ~new_n80 & ~_329gat_133_;
  assign new_n137 = ~new_n135 & ~new_n136;
  assign new_n138 = new_n134 & ~new_n137;
  assign new_n139 = _4gat_1_ & ~_14gat_4_;
  assign new_n140 = ~new_n84 & new_n139;
  assign new_n141 = new_n85 & _329gat_133_;
  assign new_n142 = ~new_n85 & ~_329gat_133_;
  assign new_n143 = ~new_n141 & ~new_n142;
  assign new_n144 = new_n140 & ~new_n143;
  assign new_n145 = _95gat_29_ & ~_105gat_32_;
  assign new_n146 = ~new_n89 & new_n145;
  assign new_n147 = new_n90 & _329gat_133_;
  assign new_n148 = ~new_n90 & ~_329gat_133_;
  assign new_n149 = ~new_n147 & ~new_n148;
  assign new_n150 = new_n146 & ~new_n149;
  assign new_n151 = ~_115gat_35_ & _108gat_33_;
  assign new_n152 = ~new_n94 & new_n151;
  assign new_n153 = new_n95 & _329gat_133_;
  assign new_n154 = ~new_n95 & ~_329gat_133_;
  assign new_n155 = ~new_n153 & ~new_n154;
  assign new_n156 = new_n152 & ~new_n155;
  assign new_n157 = _69gat_21_ & ~_79gat_24_;
  assign new_n158 = ~new_n99 & new_n157;
  assign new_n159 = new_n100 & _329gat_133_;
  assign new_n160 = ~new_n100 & ~_329gat_133_;
  assign new_n161 = ~new_n159 & ~new_n160;
  assign new_n162 = new_n158 & ~new_n161;
  assign new_n163 = _82gat_25_ & ~_92gat_28_;
  assign new_n164 = ~new_n104 & new_n163;
  assign new_n165 = new_n105 & _329gat_133_;
  assign new_n166 = ~new_n105 & ~_329gat_133_;
  assign new_n167 = ~new_n165 & ~new_n166;
  assign new_n168 = new_n164 & ~new_n167;
  assign new_n169 = ~new_n120 & ~new_n126;
  assign new_n170 = ~new_n132 & new_n169;
  assign new_n171 = ~new_n138 & new_n170;
  assign new_n172 = ~new_n144 & new_n171;
  assign new_n173 = ~new_n150 & new_n172;
  assign new_n174 = ~new_n156 & new_n173;
  assign new_n175 = ~new_n162 & new_n174;
  assign _370gat_163_ = new_n168 | ~new_n175;
  assign new_n177 = _66gat_20_ & _370gat_163_;
  assign new_n178 = _50gat_15_ & _223gat_84_;
  assign new_n179 = _56gat_17_ & ~new_n114;
  assign new_n180 = ~new_n177 & new_n179;
  assign new_n181 = ~new_n178 & new_n180;
  assign new_n182 = _73gat_22_ & _329gat_133_;
  assign new_n183 = _79gat_24_ & _370gat_163_;
  assign new_n184 = _63gat_19_ & _223gat_84_;
  assign new_n185 = _69gat_21_ & ~new_n182;
  assign new_n186 = ~new_n183 & new_n185;
  assign new_n187 = ~new_n184 & new_n186;
  assign new_n188 = _34gat_10_ & _329gat_133_;
  assign new_n189 = _40gat_12_ & _370gat_163_;
  assign new_n190 = _24gat_7_ & _223gat_84_;
  assign new_n191 = _30gat_9_ & ~new_n188;
  assign new_n192 = ~new_n189 & new_n191;
  assign new_n193 = ~new_n190 & new_n192;
  assign new_n194 = _47gat_14_ & _329gat_133_;
  assign new_n195 = _53gat_16_ & _370gat_163_;
  assign new_n196 = _37gat_11_ & _223gat_84_;
  assign new_n197 = _43gat_13_ & ~new_n194;
  assign new_n198 = ~new_n195 & new_n197;
  assign new_n199 = ~new_n196 & new_n198;
  assign new_n200 = _21gat_6_ & _329gat_133_;
  assign new_n201 = _27gat_8_ & _370gat_163_;
  assign new_n202 = _11gat_3_ & _223gat_84_;
  assign new_n203 = _17gat_5_ & ~new_n200;
  assign new_n204 = ~new_n201 & new_n203;
  assign new_n205 = ~new_n202 & new_n204;
  assign new_n206 = _112gat_34_ & _329gat_133_;
  assign new_n207 = _115gat_35_ & _370gat_163_;
  assign new_n208 = _102gat_31_ & _223gat_84_;
  assign new_n209 = _108gat_33_ & ~new_n206;
  assign new_n210 = ~new_n207 & new_n209;
  assign new_n211 = ~new_n208 & new_n210;
  assign new_n212 = _86gat_26_ & _329gat_133_;
  assign new_n213 = _92gat_28_ & _370gat_163_;
  assign new_n214 = _76gat_23_ & _223gat_84_;
  assign new_n215 = _82gat_25_ & ~new_n212;
  assign new_n216 = ~new_n213 & new_n215;
  assign new_n217 = ~new_n214 & new_n216;
  assign new_n218 = _99gat_30_ & _329gat_133_;
  assign new_n219 = _105gat_32_ & _370gat_163_;
  assign new_n220 = _89gat_27_ & _223gat_84_;
  assign new_n221 = _95gat_29_ & ~new_n218;
  assign new_n222 = ~new_n219 & new_n221;
  assign new_n223 = ~new_n220 & new_n222;
  assign new_n224 = ~new_n181 & ~new_n187;
  assign new_n225 = ~new_n193 & new_n224;
  assign new_n226 = ~new_n199 & new_n225;
  assign new_n227 = ~new_n205 & new_n226;
  assign new_n228 = ~new_n211 & new_n227;
  assign new_n229 = ~new_n217 & new_n228;
  assign new_n230 = ~new_n223 & new_n229;
  assign new_n231 = _14gat_4_ & _370gat_163_;
  assign new_n232 = _1gat_0_ & _223gat_84_;
  assign new_n233 = _8gat_2_ & _329gat_133_;
  assign new_n234 = ~new_n231 & ~new_n232;
  assign new_n235 = ~new_n233 & new_n234;
  assign new_n236 = _4gat_1_ & new_n235;
  assign _421gat_188_ = ~new_n230 & ~new_n236;
  assign new_n238 = ~new_n199 & new_n217;
  assign new_n239 = ~new_n181 & new_n238;
  assign new_n240 = ~new_n181 & ~new_n199;
  assign new_n241 = new_n187 & new_n240;
  assign new_n242 = ~new_n193 & new_n241;
  assign new_n243 = ~new_n193 & ~new_n239;
  assign new_n244 = ~new_n242 & new_n243;
  assign _431gat_194_ = new_n205 | ~new_n244;
  assign new_n246 = ~new_n199 & new_n223;
  assign new_n247 = ~new_n217 & new_n246;
  assign new_n248 = ~new_n193 & new_n247;
  assign new_n249 = ~new_n193 & new_n199;
  assign new_n250 = ~new_n248 & ~new_n249;
  assign new_n251 = ~new_n242 & new_n250;
  assign _432gat_195_ = new_n205 | ~new_n251;
  assign new_n253 = ~new_n181 & ~new_n193;
  assign new_n254 = ~new_n249 & new_n253;
  assign _430gat_193_ = new_n205 | ~new_n254;
endmodule


