// Benchmark "b22" written by ABC on Wed Sep  5 10:17:23 2018

module b22 ( clock, 
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28  );
  input  clock;
  input  SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
    SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_,
    SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_,
    SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28;
  reg P1_IR_REG_0_, P1_IR_REG_1_, P1_IR_REG_2_, P1_IR_REG_3_, P1_IR_REG_4_,
    P1_IR_REG_5_, P1_IR_REG_6_, P1_IR_REG_7_, P1_IR_REG_8_, P1_IR_REG_9_,
    P1_IR_REG_10_, P1_IR_REG_11_, P1_IR_REG_12_, P1_IR_REG_13_,
    P1_IR_REG_14_, P1_IR_REG_15_, P1_IR_REG_16_, P1_IR_REG_17_,
    P1_IR_REG_18_, P1_IR_REG_19_, P1_IR_REG_20_, P1_IR_REG_21_,
    P1_IR_REG_22_, P1_IR_REG_23_, P1_IR_REG_24_, P1_IR_REG_25_,
    P1_IR_REG_26_, P1_IR_REG_27_, P1_IR_REG_28_, P1_IR_REG_29_,
    P1_IR_REG_30_, P1_IR_REG_31_, P1_D_REG_0_, P1_D_REG_1_, P1_D_REG_2_,
    P1_D_REG_3_, P1_D_REG_4_, P1_D_REG_5_, P1_D_REG_6_, P1_D_REG_7_,
    P1_D_REG_8_, P1_D_REG_9_, P1_D_REG_10_, P1_D_REG_11_, P1_D_REG_12_,
    P1_D_REG_13_, P1_D_REG_14_, P1_D_REG_15_, P1_D_REG_16_, P1_D_REG_17_,
    P1_D_REG_18_, P1_D_REG_19_, P1_D_REG_20_, P1_D_REG_21_, P1_D_REG_22_,
    P1_D_REG_23_, P1_D_REG_24_, P1_D_REG_25_, P1_D_REG_26_, P1_D_REG_27_,
    P1_D_REG_28_, P1_D_REG_29_, P1_D_REG_30_, P1_D_REG_31_, P1_REG0_REG_0_,
    P1_REG0_REG_1_, P1_REG0_REG_2_, P1_REG0_REG_3_, P1_REG0_REG_4_,
    P1_REG0_REG_5_, P1_REG0_REG_6_, P1_REG0_REG_7_, P1_REG0_REG_8_,
    P1_REG0_REG_9_, P1_REG0_REG_10_, P1_REG0_REG_11_, P1_REG0_REG_12_,
    P1_REG0_REG_13_, P1_REG0_REG_14_, P1_REG0_REG_15_, P1_REG0_REG_16_,
    P1_REG0_REG_17_, P1_REG0_REG_18_, P1_REG0_REG_19_, P1_REG0_REG_20_,
    P1_REG0_REG_21_, P1_REG0_REG_22_, P1_REG0_REG_23_, P1_REG0_REG_24_,
    P1_REG0_REG_25_, P1_REG0_REG_26_, P1_REG0_REG_27_, P1_REG0_REG_28_,
    P1_REG0_REG_29_, P1_REG0_REG_30_, P1_REG0_REG_31_, P1_REG1_REG_0_,
    P1_REG1_REG_1_, P1_REG1_REG_2_, P1_REG1_REG_3_, P1_REG1_REG_4_,
    P1_REG1_REG_5_, P1_REG1_REG_6_, P1_REG1_REG_7_, P1_REG1_REG_8_,
    P1_REG1_REG_9_, P1_REG1_REG_10_, P1_REG1_REG_11_, P1_REG1_REG_12_,
    P1_REG1_REG_13_, P1_REG1_REG_14_, P1_REG1_REG_15_, P1_REG1_REG_16_,
    P1_REG1_REG_17_, P1_REG1_REG_18_, P1_REG1_REG_19_, P1_REG1_REG_20_,
    P1_REG1_REG_21_, P1_REG1_REG_22_, P1_REG1_REG_23_, P1_REG1_REG_24_,
    P1_REG1_REG_25_, P1_REG1_REG_26_, P1_REG1_REG_27_, P1_REG1_REG_28_,
    P1_REG1_REG_29_, P1_REG1_REG_30_, P1_REG1_REG_31_, P1_REG2_REG_0_,
    P1_REG2_REG_1_, P1_REG2_REG_2_, P1_REG2_REG_3_, P1_REG2_REG_4_,
    P1_REG2_REG_5_, P1_REG2_REG_6_, P1_REG2_REG_7_, P1_REG2_REG_8_,
    P1_REG2_REG_9_, P1_REG2_REG_10_, P1_REG2_REG_11_, P1_REG2_REG_12_,
    P1_REG2_REG_13_, P1_REG2_REG_14_, P1_REG2_REG_15_, P1_REG2_REG_16_,
    P1_REG2_REG_17_, P1_REG2_REG_18_, P1_REG2_REG_19_, P1_REG2_REG_20_,
    P1_REG2_REG_21_, P1_REG2_REG_22_, P1_REG2_REG_23_, P1_REG2_REG_24_,
    P1_REG2_REG_25_, P1_REG2_REG_26_, P1_REG2_REG_27_, P1_REG2_REG_28_,
    P1_REG2_REG_29_, P1_REG2_REG_30_, P1_REG2_REG_31_, P1_ADDR_REG_19_,
    P1_ADDR_REG_18_, P1_ADDR_REG_17_, P1_ADDR_REG_16_, P1_ADDR_REG_15_,
    P1_ADDR_REG_14_, P1_ADDR_REG_13_, P1_ADDR_REG_12_, P1_ADDR_REG_11_,
    P1_ADDR_REG_10_, P1_ADDR_REG_9_, P1_ADDR_REG_8_, P1_ADDR_REG_7_,
    P1_ADDR_REG_6_, P1_ADDR_REG_5_, P1_ADDR_REG_4_, P1_ADDR_REG_3_,
    P1_ADDR_REG_2_, P1_ADDR_REG_1_, P1_ADDR_REG_0_, P1_DATAO_REG_0_,
    P1_DATAO_REG_1_, P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_,
    P1_DATAO_REG_5_, P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_,
    P1_DATAO_REG_9_, P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_,
    P1_DATAO_REG_13_, P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_,
    P1_DATAO_REG_17_, P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_,
    P1_DATAO_REG_21_, P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_,
    P1_DATAO_REG_25_, P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_,
    P1_DATAO_REG_29_, P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_B_REG,
    P1_REG3_REG_15_, P1_REG3_REG_26_, P1_REG3_REG_6_, P1_REG3_REG_18_,
    P1_REG3_REG_2_, P1_REG3_REG_11_, P1_REG3_REG_22_, P1_REG3_REG_13_,
    P1_REG3_REG_20_, P1_REG3_REG_0_, P1_REG3_REG_9_, P1_REG3_REG_4_,
    P1_REG3_REG_24_, P1_REG3_REG_17_, P1_REG3_REG_5_, P1_REG3_REG_16_,
    P1_REG3_REG_25_, P1_REG3_REG_12_, P1_REG3_REG_21_, P1_REG3_REG_1_,
    P1_REG3_REG_8_, P1_REG3_REG_28_, P1_REG3_REG_19_, P1_REG3_REG_3_,
    P1_REG3_REG_10_, P1_REG3_REG_23_, P1_REG3_REG_14_, P1_REG3_REG_27_,
    P1_REG3_REG_7_, P1_STATE_REG, P1_RD_REG, P1_WR_REG, P2_IR_REG_0_,
    P2_IR_REG_1_, P2_IR_REG_2_, P2_IR_REG_3_, P2_IR_REG_4_, P2_IR_REG_5_,
    P2_IR_REG_6_, P2_IR_REG_7_, P2_IR_REG_8_, P2_IR_REG_9_, P2_IR_REG_10_,
    P2_IR_REG_11_, P2_IR_REG_12_, P2_IR_REG_13_, P2_IR_REG_14_,
    P2_IR_REG_15_, P2_IR_REG_16_, P2_IR_REG_17_, P2_IR_REG_18_,
    P2_IR_REG_19_, P2_IR_REG_20_, P2_IR_REG_21_, P2_IR_REG_22_,
    P2_IR_REG_23_, P2_IR_REG_24_, P2_IR_REG_25_, P2_IR_REG_26_,
    P2_IR_REG_27_, P2_IR_REG_28_, P2_IR_REG_29_, P2_IR_REG_30_,
    P2_IR_REG_31_, P2_D_REG_0_, P2_D_REG_1_, P2_D_REG_2_, P2_D_REG_3_,
    P2_D_REG_4_, P2_D_REG_5_, P2_D_REG_6_, P2_D_REG_7_, P2_D_REG_8_,
    P2_D_REG_9_, P2_D_REG_10_, P2_D_REG_11_, P2_D_REG_12_, P2_D_REG_13_,
    P2_D_REG_14_, P2_D_REG_15_, P2_D_REG_16_, P2_D_REG_17_, P2_D_REG_18_,
    P2_D_REG_19_, P2_D_REG_20_, P2_D_REG_21_, P2_D_REG_22_, P2_D_REG_23_,
    P2_D_REG_24_, P2_D_REG_25_, P2_D_REG_26_, P2_D_REG_27_, P2_D_REG_28_,
    P2_D_REG_29_, P2_D_REG_30_, P2_D_REG_31_, P2_REG0_REG_0_,
    P2_REG0_REG_1_, P2_REG0_REG_2_, P2_REG0_REG_3_, P2_REG0_REG_4_,
    P2_REG0_REG_5_, P2_REG0_REG_6_, P2_REG0_REG_7_, P2_REG0_REG_8_,
    P2_REG0_REG_9_, P2_REG0_REG_10_, P2_REG0_REG_11_, P2_REG0_REG_12_,
    P2_REG0_REG_13_, P2_REG0_REG_14_, P2_REG0_REG_15_, P2_REG0_REG_16_,
    P2_REG0_REG_17_, P2_REG0_REG_18_, P2_REG0_REG_19_, P2_REG0_REG_20_,
    P2_REG0_REG_21_, P2_REG0_REG_22_, P2_REG0_REG_23_, P2_REG0_REG_24_,
    P2_REG0_REG_25_, P2_REG0_REG_26_, P2_REG0_REG_27_, P2_REG0_REG_28_,
    P2_REG0_REG_29_, P2_REG0_REG_30_, P2_REG0_REG_31_, P2_REG1_REG_0_,
    P2_REG1_REG_1_, P2_REG1_REG_2_, P2_REG1_REG_3_, P2_REG1_REG_4_,
    P2_REG1_REG_5_, P2_REG1_REG_6_, P2_REG1_REG_7_, P2_REG1_REG_8_,
    P2_REG1_REG_9_, P2_REG1_REG_10_, P2_REG1_REG_11_, P2_REG1_REG_12_,
    P2_REG1_REG_13_, P2_REG1_REG_14_, P2_REG1_REG_15_, P2_REG1_REG_16_,
    P2_REG1_REG_17_, P2_REG1_REG_18_, P2_REG1_REG_19_, P2_REG1_REG_20_,
    P2_REG1_REG_21_, P2_REG1_REG_22_, P2_REG1_REG_23_, P2_REG1_REG_24_,
    P2_REG1_REG_25_, P2_REG1_REG_26_, P2_REG1_REG_27_, P2_REG1_REG_28_,
    P2_REG1_REG_29_, P2_REG1_REG_30_, P2_REG1_REG_31_, P2_REG2_REG_0_,
    P2_REG2_REG_1_, P2_REG2_REG_2_, P2_REG2_REG_3_, P2_REG2_REG_4_,
    P2_REG2_REG_5_, P2_REG2_REG_6_, P2_REG2_REG_7_, P2_REG2_REG_8_,
    P2_REG2_REG_9_, P2_REG2_REG_10_, P2_REG2_REG_11_, P2_REG2_REG_12_,
    P2_REG2_REG_13_, P2_REG2_REG_14_, P2_REG2_REG_15_, P2_REG2_REG_16_,
    P2_REG2_REG_17_, P2_REG2_REG_18_, P2_REG2_REG_19_, P2_REG2_REG_20_,
    P2_REG2_REG_21_, P2_REG2_REG_22_, P2_REG2_REG_23_, P2_REG2_REG_24_,
    P2_REG2_REG_25_, P2_REG2_REG_26_, P2_REG2_REG_27_, P2_REG2_REG_28_,
    P2_REG2_REG_29_, P2_REG2_REG_30_, P2_REG2_REG_31_, P2_ADDR_REG_19_,
    P2_ADDR_REG_18_, P2_ADDR_REG_17_, P2_ADDR_REG_16_, P2_ADDR_REG_15_,
    P2_ADDR_REG_14_, P2_ADDR_REG_13_, P2_ADDR_REG_12_, P2_ADDR_REG_11_,
    P2_ADDR_REG_10_, P2_ADDR_REG_9_, P2_ADDR_REG_8_, P2_ADDR_REG_7_,
    P2_ADDR_REG_6_, P2_ADDR_REG_5_, P2_ADDR_REG_4_, P2_ADDR_REG_3_,
    P2_ADDR_REG_2_, P2_ADDR_REG_1_, P2_ADDR_REG_0_, P2_DATAO_REG_0_,
    P2_DATAO_REG_1_, P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_,
    P2_DATAO_REG_5_, P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_,
    P2_DATAO_REG_9_, P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_,
    P2_DATAO_REG_13_, P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_,
    P2_DATAO_REG_17_, P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_,
    P2_DATAO_REG_21_, P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_,
    P2_DATAO_REG_25_, P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_,
    P2_DATAO_REG_29_, P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_B_REG,
    P2_REG3_REG_15_, P2_REG3_REG_26_, P2_REG3_REG_6_, P2_REG3_REG_18_,
    P2_REG3_REG_2_, P2_REG3_REG_11_, P2_REG3_REG_22_, P2_REG3_REG_13_,
    P2_REG3_REG_20_, P2_REG3_REG_0_, P2_REG3_REG_9_, P2_REG3_REG_4_,
    P2_REG3_REG_24_, P2_REG3_REG_17_, P2_REG3_REG_5_, P2_REG3_REG_16_,
    P2_REG3_REG_25_, P2_REG3_REG_12_, P2_REG3_REG_21_, P2_REG3_REG_1_,
    P2_REG3_REG_8_, P2_REG3_REG_28_, P2_REG3_REG_19_, P2_REG3_REG_3_,
    P2_REG3_REG_10_, P2_REG3_REG_23_, P2_REG3_REG_14_, P2_REG3_REG_27_,
    P2_REG3_REG_7_, P2_STATE_REG, P2_RD_REG, P2_WR_REG, P3_IR_REG_0_,
    P3_IR_REG_1_, P3_IR_REG_2_, P3_IR_REG_3_, P3_IR_REG_4_, P3_IR_REG_5_,
    P3_IR_REG_6_, P3_IR_REG_7_, P3_IR_REG_8_, P3_IR_REG_9_, P3_IR_REG_10_,
    P3_IR_REG_11_, P3_IR_REG_12_, P3_IR_REG_13_, P3_IR_REG_14_,
    P3_IR_REG_15_, P3_IR_REG_16_, P3_IR_REG_17_, P3_IR_REG_18_,
    P3_IR_REG_19_, P3_IR_REG_20_, P3_IR_REG_21_, P3_IR_REG_22_,
    P3_IR_REG_23_, P3_IR_REG_24_, P3_IR_REG_25_, P3_IR_REG_26_,
    P3_IR_REG_27_, P3_IR_REG_28_, P3_IR_REG_29_, P3_IR_REG_30_,
    P3_IR_REG_31_, P3_D_REG_0_, P3_D_REG_1_, P3_D_REG_2_, P3_D_REG_3_,
    P3_D_REG_4_, P3_D_REG_5_, P3_D_REG_6_, P3_D_REG_7_, P3_D_REG_8_,
    P3_D_REG_9_, P3_D_REG_10_, P3_D_REG_11_, P3_D_REG_12_, P3_D_REG_13_,
    P3_D_REG_14_, P3_D_REG_15_, P3_D_REG_16_, P3_D_REG_17_, P3_D_REG_18_,
    P3_D_REG_19_, P3_D_REG_20_, P3_D_REG_21_, P3_D_REG_22_, P3_D_REG_23_,
    P3_D_REG_24_, P3_D_REG_25_, P3_D_REG_26_, P3_D_REG_27_, P3_D_REG_28_,
    P3_D_REG_29_, P3_D_REG_30_, P3_D_REG_31_, P3_REG0_REG_0_,
    P3_REG0_REG_1_, P3_REG0_REG_2_, P3_REG0_REG_3_, P3_REG0_REG_4_,
    P3_REG0_REG_5_, P3_REG0_REG_6_, P3_REG0_REG_7_, P3_REG0_REG_8_,
    P3_REG0_REG_9_, P3_REG0_REG_10_, P3_REG0_REG_11_, P3_REG0_REG_12_,
    P3_REG0_REG_13_, P3_REG0_REG_14_, P3_REG0_REG_15_, P3_REG0_REG_16_,
    P3_REG0_REG_17_, P3_REG0_REG_18_, P3_REG0_REG_19_, P3_REG0_REG_20_,
    P3_REG0_REG_21_, P3_REG0_REG_22_, P3_REG0_REG_23_, P3_REG0_REG_24_,
    P3_REG0_REG_25_, P3_REG0_REG_26_, P3_REG0_REG_27_, P3_REG0_REG_28_,
    P3_REG0_REG_29_, P3_REG0_REG_30_, P3_REG0_REG_31_, P3_REG1_REG_0_,
    P3_REG1_REG_1_, P3_REG1_REG_2_, P3_REG1_REG_3_, P3_REG1_REG_4_,
    P3_REG1_REG_5_, P3_REG1_REG_6_, P3_REG1_REG_7_, P3_REG1_REG_8_,
    P3_REG1_REG_9_, P3_REG1_REG_10_, P3_REG1_REG_11_, P3_REG1_REG_12_,
    P3_REG1_REG_13_, P3_REG1_REG_14_, P3_REG1_REG_15_, P3_REG1_REG_16_,
    P3_REG1_REG_17_, P3_REG1_REG_18_, P3_REG1_REG_19_, P3_REG1_REG_20_,
    P3_REG1_REG_21_, P3_REG1_REG_22_, P3_REG1_REG_23_, P3_REG1_REG_24_,
    P3_REG1_REG_25_, P3_REG1_REG_26_, P3_REG1_REG_27_, P3_REG1_REG_28_,
    P3_REG1_REG_29_, P3_REG1_REG_30_, P3_REG1_REG_31_, P3_REG2_REG_0_,
    P3_REG2_REG_1_, P3_REG2_REG_2_, P3_REG2_REG_3_, P3_REG2_REG_4_,
    P3_REG2_REG_5_, P3_REG2_REG_6_, P3_REG2_REG_7_, P3_REG2_REG_8_,
    P3_REG2_REG_9_, P3_REG2_REG_10_, P3_REG2_REG_11_, P3_REG2_REG_12_,
    P3_REG2_REG_13_, P3_REG2_REG_14_, P3_REG2_REG_15_, P3_REG2_REG_16_,
    P3_REG2_REG_17_, P3_REG2_REG_18_, P3_REG2_REG_19_, P3_REG2_REG_20_,
    P3_REG2_REG_21_, P3_REG2_REG_22_, P3_REG2_REG_23_, P3_REG2_REG_24_,
    P3_REG2_REG_25_, P3_REG2_REG_26_, P3_REG2_REG_27_, P3_REG2_REG_28_,
    P3_REG2_REG_29_, P3_REG2_REG_30_, P3_REG2_REG_31_, P3_ADDR_REG_19_,
    P3_ADDR_REG_18_, P3_ADDR_REG_17_, P3_ADDR_REG_16_, P3_ADDR_REG_15_,
    P3_ADDR_REG_14_, P3_ADDR_REG_13_, P3_ADDR_REG_12_, P3_ADDR_REG_11_,
    P3_ADDR_REG_10_, P3_ADDR_REG_9_, P3_ADDR_REG_8_, P3_ADDR_REG_7_,
    P3_ADDR_REG_6_, P3_ADDR_REG_5_, P3_ADDR_REG_4_, P3_ADDR_REG_3_,
    P3_ADDR_REG_2_, P3_ADDR_REG_1_, P3_ADDR_REG_0_, P3_DATAO_REG_0_,
    P3_DATAO_REG_1_, P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_,
    P3_DATAO_REG_5_, P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_,
    P3_DATAO_REG_9_, P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_,
    P3_DATAO_REG_13_, P3_DATAO_REG_14_, P3_DATAO_REG_15_, P3_DATAO_REG_16_,
    P3_DATAO_REG_17_, P3_DATAO_REG_18_, P3_DATAO_REG_19_, P3_DATAO_REG_20_,
    P3_DATAO_REG_21_, P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_,
    P3_DATAO_REG_25_, P3_DATAO_REG_26_, P3_DATAO_REG_27_, P3_DATAO_REG_28_,
    P3_DATAO_REG_29_, P3_DATAO_REG_30_, P3_DATAO_REG_31_, P3_B_REG,
    P3_REG3_REG_15_, P3_REG3_REG_26_, P3_REG3_REG_6_, P3_REG3_REG_18_,
    P3_REG3_REG_2_, P3_REG3_REG_11_, P3_REG3_REG_22_, P3_REG3_REG_13_,
    P3_REG3_REG_20_, P3_REG3_REG_0_, P3_REG3_REG_9_, P3_REG3_REG_4_,
    P3_REG3_REG_24_, P3_REG3_REG_17_, P3_REG3_REG_5_, P3_REG3_REG_16_,
    P3_REG3_REG_25_, P3_REG3_REG_12_, P3_REG3_REG_21_, P3_REG3_REG_1_,
    P3_REG3_REG_8_, P3_REG3_REG_28_, P3_REG3_REG_19_, P3_REG3_REG_3_,
    P3_REG3_REG_10_, P3_REG3_REG_23_, P3_REG3_REG_14_, P3_REG3_REG_27_,
    P3_REG3_REG_7_, P3_STATE_REG, P3_RD_REG, P3_WR_REG;
  wire n2260_1, n2261, n2262, n2263, n2264, n2265_1, n2266, n2267, n2268,
    n2269, n2270_1, n2271, n2272, n2273, n2274, n2275_1, n2276, n2277,
    n2278, n2279, n2280_1, n2281, n2282, n2283, n2284, n2285_1, n2286,
    n2287, n2288, n2289, n2290_1, n2291, n2292, n2293, n2294, n2295_1,
    n2296, n2297, n2298, n2299, n2300_1, n2301, n2302, n2303, n2304,
    n2305_1, n2306, n2307, n2308, n2309, n2310_1, n2311, n2312, n2313,
    n2314, n2315_1, n2316, n2317, n2318, n2319, n2320_1, n2321, n2322,
    n2323, n2324, n2325_1, n2326, n2327, n2328, n2329, n2330_1, n2331,
    n2332, n2333, n2334, n2335_1, n2336, n2337, n2338, n2339, n2340_1,
    n2341, n2342, n2343, n2344, n2345_1, n2346, n2347, n2348, n2349,
    n2350_1, n2351, n2352, n2353, n2354, n2355_1, n2356, n2357, n2358,
    n2359, n2360_1, n2361, n2362, n2363, n2364, n2365_1, n2366, n2367,
    n2368, n2369, n2370_1, n2371, n2372, n2373, n2374, n2375_1, n2376,
    n2377, n2378, n2379, n2380_1, n2381, n2382, n2383, n2384, n2385_1,
    n2386, n2387, n2388, n2389, n2390_1, n2391, n2392, n2393, n2394,
    n2395_1, n2396, n2397, n2398, n2399, n2400_1, n2401, n2402, n2403,
    n2404, n2405_1, n2406, n2407, n2408, n2409, n2410_1, n2411, n2412,
    n2413, n2414, n2415_1, n2416, n2417, n2418, n2419, n2420_1, n2421,
    n2422, n2423, n2424, n2425_1, n2426, n2427, n2428, n2429, n2430_1,
    n2431, n2432, n2433, n2434, n2435_1, n2436, n2437, n2438, n2439,
    n2440_1, n2441, n2442, n2443, n2444, n2445_1, n2446, n2447, n2448,
    n2449, n2450_1, n2451, n2452, n2453, n2454, n2455_1, n2456, n2457,
    n2458, n2459, n2460_1, n2461, n2462, n2463, n2464, n2465_1, n2466,
    n2467, n2468, n2469, n2470_1, n2471, n2472, n2473, n2474, n2475_1,
    n2476, n2477, n2478, n2479, n2480_1, n2481, n2482, n2483, n2484,
    n2485_1, n2486, n2487, n2488, n2489, n2490_1, n2491, n2492, n2493,
    n2494, n2495_1, n2496, n2497, n2499, n2500_1, n2501, n2503, n2504,
    n2505_1, n2506, n2507, n2509, n2510_1, n2511, n2512, n2513, n2515_1,
    n2516, n2517, n2519, n2520_1, n2521, n2523, n2524, n2525_1, n2527,
    n2528, n2529, n2530_1, n2531, n2533, n2534, n2535_1, n2536, n2537,
    n2539, n2540_1, n2541, n2543, n2544, n2545_1, n2546, n2547, n2549,
    n2550_1, n2551, n2553, n2554, n2555_1, n2556, n2557, n2559, n2560_1,
    n2561, n2562, n2563, n2565_1, n2566, n2567, n2569, n2570_1, n2571,
    n2572, n2573, n2575_1, n2576, n2577, n2579, n2580_1, n2581, n2582,
    n2583, n2585_1, n2586, n2587, n2588, n2589, n2590_1, n2591, n2592,
    n2594, n2595_1, n2597, n2598, n2599, n2601, n2602, n2603, n2605_1,
    n2606, n2607, n2608, n2609, n2610_1, n2611, n2612, n2613, n2614,
    n2615_1, n2616, n2617, n2618, n2619, n2620_1, n2621, n2622, n2623,
    n2624, n2625_1, n2626, n2628, n2629, n2630_1, n2631, n2632, n2633,
    n2634, n2635_1, n2636, n2637, n2638, n2639, n2640_1, n2641, n2642,
    n2643, n2644, n2645_1, n2646, n2647, n2648, n2649, n2650_1, n2651,
    n2652, n2654, n2655_1, n2656, n2657, n2658, n2659, n2660_1, n2661,
    n2662, n2663, n2664, n2665_1, n2666, n2667, n2668, n2669, n2670_1,
    n2671, n2672, n2673, n2674, n2675_1, n2676, n2677, n2679, n2680_1,
    n2681, n2682, n2683, n2684, n2685_1, n2686, n2687, n2688, n2689,
    n2690_1, n2691, n2692, n2693, n2694, n2695_1, n2696, n2697, n2698,
    n2699, n2700_1, n2701, n2702, n2703, n2704, n2705_1, n2706, n2707,
    n2708, n2710_1, n2711, n2712, n2713, n2714, n2715_1, n2716, n2717,
    n2718, n2719, n2720_1, n2721, n2722, n2723, n2724, n2725_1, n2726,
    n2727, n2728, n2729, n2730_1, n2731, n2732, n2733, n2734, n2735_1,
    n2736, n2738, n2739, n2740_1, n2741, n2742, n2743, n2744, n2745_1,
    n2746, n2747, n2748, n2749, n2750_1, n2751, n2752, n2753, n2754,
    n2755_1, n2756, n2757, n2758, n2759, n2760_1, n2762, n2763, n2764,
    n2765_1, n2766, n2767, n2768, n2769, n2770_1, n2771, n2772, n2773,
    n2774, n2775_1, n2776, n2777, n2778, n2779, n2780_1, n2781, n2782,
    n2783, n2784, n2785_1, n2786, n2787, n2788, n2790_1, n2791, n2792,
    n2793, n2794, n2795_1, n2796, n2797, n2798, n2799, n2800_1, n2801,
    n2802, n2803, n2804, n2805_1, n2806, n2807, n2808, n2809, n2810_1,
    n2811, n2812, n2813, n2814, n2815_1, n2817, n2818, n2819, n2820_1,
    n2821, n2822, n2823, n2824, n2825_1, n2826, n2827, n2828, n2829,
    n2830_1, n2831, n2832, n2833, n2834, n2835_1, n2836, n2837, n2838,
    n2839, n2840_1, n2841, n2842, n2843, n2845_1, n2846, n2847, n2848,
    n2849, n2850_1, n2851, n2852, n2853, n2854, n2855_1, n2856, n2857,
    n2858, n2859, n2860_1, n2861, n2862, n2863, n2864, n2865_1, n2866,
    n2867, n2868, n2869, n2870_1, n2872, n2873, n2874, n2875_1, n2876,
    n2877, n2878, n2879, n2880_1, n2881, n2882, n2883, n2884, n2885_1,
    n2886, n2887, n2888, n2889, n2890_1, n2891, n2892, n2893, n2894,
    n2895_1, n2896, n2897, n2898, n2900_1, n2901, n2902, n2903, n2904,
    n2905_1, n2906, n2907, n2908, n2909, n2910_1, n2911, n2912, n2913,
    n2914, n2915_1, n2916, n2917, n2918, n2919, n2920_1, n2921, n2922,
    n2923, n2924, n2925_1, n2927, n2928, n2929, n2930_1, n2931, n2932,
    n2933, n2934, n2935_1, n2936, n2937, n2938, n2939, n2940_1, n2941,
    n2942, n2943, n2944, n2945_1, n2946, n2947, n2948, n2949, n2950_1,
    n2951, n2952, n2954, n2955_1, n2956, n2957, n2958, n2959, n2960_1,
    n2961, n2962, n2963, n2964, n2965_1, n2966, n2967, n2968, n2969,
    n2970_1, n2971, n2972, n2973, n2974, n2975_1, n2976, n2977, n2978,
    n2979, n2981, n2982, n2983, n2984, n2985_1, n2986, n2987, n2988, n2989,
    n2990_1, n2991, n2992, n2993, n2994, n2995_1, n2996, n2997, n2998,
    n2999, n3000_1, n3001, n3002, n3003, n3004, n3005_1, n3006, n3007,
    n3009, n3010_1, n3011, n3012, n3013, n3014, n3015_1, n3016, n3017,
    n3018, n3019, n3020_1, n3021, n3022, n3023, n3024, n3025_1, n3026,
    n3027, n3028, n3029, n3030_1, n3031, n3032, n3033, n3034, n3036, n3037,
    n3038, n3039, n3040_1, n3041, n3042, n3043, n3044, n3045_1, n3046,
    n3047, n3048, n3049, n3050_1, n3051, n3052, n3053, n3054, n3055_1,
    n3056, n3057, n3058, n3059, n3060_1, n3061, n3062, n3063, n3064,
    n3065_1, n3066, n3067, n3068, n3069, n3070_1, n3071, n3072, n3073,
    n3074, n3075_1, n3077, n3078, n3079, n3080_1, n3081, n3082, n3083,
    n3084, n3085_1, n3086, n3087, n3088, n3089, n3090_1, n3091, n3092,
    n3093, n3094, n3095_1, n3096, n3097, n3098, n3099, n3101, n3102, n3103,
    n3104, n3105_1, n3106, n3107, n3108, n3109, n3110_1, n3111, n3112,
    n3113, n3114, n3115_1, n3116, n3117, n3118, n3119, n3120_1, n3121,
    n3122, n3123, n3124, n3125_1, n3126, n3127, n3128, n3129, n3130_1,
    n3131, n3132, n3133, n3135_1, n3136, n3137, n3138, n3139, n3140_1,
    n3141, n3142, n3143, n3144, n3145_1, n3146, n3147, n3148, n3149,
    n3150_1, n3151, n3152, n3153, n3154, n3155_1, n3156, n3157, n3158,
    n3159, n3160_1, n3161, n3162, n3163, n3164, n3165_1, n3166, n3167,
    n3168, n3169, n3170_1, n3172, n3173, n3174, n3175_1, n3176, n3177,
    n3178, n3179, n3180_1, n3181, n3182, n3183, n3184, n3185_1, n3186,
    n3187, n3188, n3189, n3190_1, n3191, n3192, n3193, n3194, n3195_1,
    n3196, n3197, n3198, n3199, n3200_1, n3201, n3202, n3203, n3204,
    n3205_1, n3206, n3207, n3209, n3210_1, n3211, n3212, n3213, n3214,
    n3215_1, n3216, n3217, n3218, n3219, n3220_1, n3221, n3222, n3223,
    n3224, n3225_1, n3226, n3227, n3228, n3229, n3230_1, n3231, n3233,
    n3234, n3235_1, n3236, n3237, n3238, n3239, n3240_1, n3241, n3242,
    n3243, n3244, n3245_1, n3246, n3247, n3248, n3249, n3250_1, n3251,
    n3252, n3253, n3254, n3255_1, n3256, n3257, n3258, n3259, n3260_1,
    n3261, n3262, n3263, n3264, n3265_1, n3266, n3267, n3268, n3270_1,
    n3271, n3272, n3273, n3274, n3275_1, n3276, n3277, n3278, n3279,
    n3280_1, n3281, n3282, n3283, n3284, n3285_1, n3286, n3287, n3288,
    n3289, n3290_1, n3291, n3292, n3293, n3294, n3295_1, n3296, n3297,
    n3298, n3299, n3300_1, n3301, n3302, n3303, n3304, n3305_1, n3306,
    n3307, n3308, n3309, n3310_1, n3312, n3313, n3314, n3315_1, n3316,
    n3317, n3318, n3319, n3320_1, n3321, n3322, n3323, n3324, n3325_1,
    n3326, n3327, n3328, n3329, n3330_1, n3331, n3332, n3333, n3334,
    n3335_1, n3336, n3337, n3338, n3339, n3340_1, n3341, n3342, n3343,
    n3344, n3345_1, n3346, n3347, n3348, n3349, n3350_1, n3352, n3353,
    n3354, n3355_1, n3356, n3357, n3358, n3359, n3360_1, n3361, n3362,
    n3363, n3364, n3365_1, n3366, n3367, n3368, n3369, n3370_1, n3371,
    n3372, n3373, n3374, n3376, n3377, n3378, n3379, n3380_1, n3381, n3382,
    n3383, n3384, n3385_1, n3386, n3387, n3388, n3389, n3390_1, n3391,
    n3392, n3393, n3394, n3395_1, n3396, n3397, n3398, n3399, n3400_1,
    n3401, n3402, n3403, n3404, n3405_1, n3406, n3407, n3408, n3409,
    n3410_1, n3411, n3412, n3413, n3414, n3415_1, n3416, n3417, n3419,
    n3420_1, n3421, n3422, n3423, n3424, n3425_1, n3426, n3427, n3428,
    n3429, n3430_1, n3431, n3432, n3433, n3434, n3435_1, n3436, n3437,
    n3438, n3439, n3440_1, n3441, n3443, n3444, n3445_1, n3446, n3447,
    n3448, n3449, n3450_1, n3451, n3452, n3453, n3454, n3455_1, n3456,
    n3457, n3458, n3459, n3460_1, n3461, n3462, n3463, n3464, n3465_1,
    n3466, n3467, n3468, n3469, n3470_1, n3471, n3472, n3473, n3474,
    n3475_1, n3476, n3477, n3478, n3479, n3480_1, n3481, n3482, n3483,
    n3484, n3485_1, n3486, n3488, n3489, n3490_1, n3491, n3492, n3493,
    n3494, n3495_1, n3496, n3497, n3498, n3499, n3500_1, n3501, n3502,
    n3503, n3504, n3505_1, n3506, n3507, n3508, n3509, n3510_1, n3511,
    n3512, n3513, n3514, n3515_1, n3517, n3518, n3519, n3520_1, n3521,
    n3522, n3523, n3524, n3525_1, n3526, n3527, n3528, n3529, n3530_1,
    n3531, n3532, n3533, n3534, n3535_1, n3536, n3537, n3538, n3539, n3541,
    n3542, n3543, n3544, n3545_1, n3546, n3547, n3548, n3549, n3550_1,
    n3551, n3552, n3553, n3554, n3555_1, n3556, n3557, n3558, n3559,
    n3560_1, n3561, n3562, n3563, n3564, n3565_1, n3566, n3567, n3568,
    n3569, n3570_1, n3572, n3573, n3574, n3575_1, n3576, n3577, n3578,
    n3579, n3580_1, n3581, n3582, n3583, n3584, n3585_1, n3586, n3587,
    n3588, n3589, n3590_1, n3591, n3592, n3593, n3594, n3595_1, n3596,
    n3597, n3599, n3600_1, n3601, n3633, n3634, n3635_1, n3636, n3637,
    n3638, n3639, n3640_1, n3641, n3642, n3643, n3644, n3645_1, n3646,
    n3647, n3648, n3649, n3650_1, n3651, n3652, n3653, n3654, n3655_1,
    n3656, n3657, n3658, n3659, n3660_1, n3661, n3662, n3663, n3664,
    n3665_1, n3666, n3667, n3668, n3669, n3670_1, n3671, n3672, n3673,
    n3674, n3675_1, n3676, n3677, n3678, n3679, n3680_1, n3681, n3682,
    n3683, n3684, n3685_1, n3686, n3687, n3688, n3689, n3690_1, n3691,
    n3692, n3693, n3694, n3695_1, n3696, n3697, n3698, n3699, n3700_1,
    n3701, n3702, n3703, n3704, n3705_1, n3706, n3707, n3708, n3709,
    n3710_1, n3711, n3712, n3713, n3714, n3715_1, n3716, n3717, n3718,
    n3719, n3720_1, n3721, n3722, n3723, n3724, n3725_1, n3726, n3727,
    n3728, n3729, n3730_1, n3731, n3732, n3733, n3734, n3735_1, n3736,
    n3737, n3738, n3739, n3740_1, n3741, n3742, n3743, n3744, n3745_1,
    n3746, n3747, n3748, n3749, n3750_1, n3751, n3752, n3753, n3754,
    n3755_1, n3756, n3757, n3758, n3759, n3760_1, n3761, n3762, n3763,
    n3764, n3765_1, n3766, n3767, n3768, n3769, n3770_1, n3771, n3772,
    n3773, n3774, n3775_1, n3776, n3777, n3778, n3779, n3780_1, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4125, n4126, n4127,
    n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
    n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
    n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
    n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
    n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
    n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
    n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5117, n5118, n5119, n5120, n5121, n5122,
    n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
    n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5690, n5691, n5692, n5693,
    n5695, n5696, n5698, n5699, n5701, n5702, n5704, n5705, n5707, n5708,
    n5710, n5711, n5713, n5714, n5716, n5717, n5719, n5720, n5722, n5723,
    n5725, n5726, n5728, n5729, n5731, n5732, n5734, n5735, n5737, n5738,
    n5740, n5741, n5743, n5744, n5746, n5747, n5749, n5750, n5752, n5753,
    n5755, n5756, n5758, n5759, n5761, n5762, n5764, n5765, n5767, n5768,
    n5770, n5771, n5773, n5774, n5776, n5777, n5779, n5780, n5782, n5783,
    n5785, n5786, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
    n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
    n6011, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6130,
    n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6193, n6194, n6195,
    n6196, n6197, n6198, n6200, n6201, n6202, n6203, n6204, n6206, n6207,
    n6208, n6209, n6210, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
    n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
    n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
    n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
    n6522, n6523, n6524, n6525, n6526, n6527, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
    n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
    n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7090, n7091, n7093, n7094, n7096, n7097, n7099, n7100, n7102, n7103,
    n7105, n7106, n7108, n7109, n7111, n7112, n7114, n7115, n7117, n7118,
    n7120, n7121, n7123, n7124, n7126, n7127, n7129, n7130, n7132, n7133,
    n7135, n7136, n7138, n7139, n7141, n7142, n7144, n7145, n7147, n7148,
    n7150, n7151, n7153, n7154, n7156, n7157, n7159, n7160, n7162, n7163,
    n7165, n7166, n7168, n7169, n7171, n7172, n7174, n7175, n7177, n7178,
    n7180, n7181, n7183, n7184, n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
    n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
    n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
    n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
    n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
    n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
    n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
    n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
    n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
    n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
    n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
    n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
    n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
    n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
    n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
    n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
    n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
    n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
    n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
    n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
    n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
    n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
    n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
    n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
    n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
    n7842, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
    n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
    n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
    n8506, n8507, n8508, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
    n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
    n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
    n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
    n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
    n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
    n8704, n8705, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
    n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
    n8746, n8747, n8748, n8749, n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
    n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
    n8928, n8929, n8930, n8931, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
    n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
    n9315, n9316, n9317, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
    n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
    n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9773, n9774, n9775, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
    n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
    n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
    n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
    n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
    n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
    n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
    n10212, n10213, n10214, n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10364, n10365, n10366, n10367,
    n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
    n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
    n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
    n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
    n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
    n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10641,
    n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
    n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
    n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
    n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
    n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
    n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
    n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
    n10979, n10980, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
    n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
    n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11115, n11116,
    n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
    n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
    n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
    n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11184, n11185, n11186, n11187, n11188, n11189,
    n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
    n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
    n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
    n11308, n11309, n11310, n11311, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11378, n11379, n11380, n11381,
    n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
    n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
    n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11449, n11450, n11451, n11452, n11453, n11454,
    n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
    n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
    n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
    n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
    n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
    n11509, n11510, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
    n11538, n11540, n11541, n11542, n11543, n11545, n11546, n11548, n11549,
    n11551, n11552, n11554, n11555, n11557, n11558, n11560, n11561, n11563,
    n11564, n11566, n11567, n11569, n11570, n11572, n11573, n11575, n11576,
    n11578, n11579, n11581, n11582, n11584, n11585, n11587, n11588, n11590,
    n11591, n11593, n11594, n11596, n11597, n11599, n11600, n11602, n11603,
    n11605, n11606, n11608, n11609, n11611, n11612, n11614, n11615, n11617,
    n11618, n11620, n11621, n11623, n11624, n11626, n11627, n11629, n11630,
    n11632, n11633, n11635, n11636, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
    n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11694, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
    n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822, n11824, n11825, n11826,
    n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11857, n11858, n11859, n11860, n11861, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
    n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11902, n11903, n11904,
    n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
    n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11928, n11929, n11930, n11931, n11932, n11933,
    n11934, n11935, n11936, n11937, n11938, n11939, n11941, n11942, n11943,
    n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
    n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978, n11980, n11981, n11982,
    n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
    n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12043, n12044, n12045, n12046, n12047, n12048, n12050, n12051,
    n12052, n12053, n12054, n12056, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
    n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12292, n12293, n12294, n12295, n12296, n12297,
    n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
    n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
    n12325, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
    n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
    n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
    n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
    n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524, n12526, n12527, n12528,
    n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
    n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
    n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12647, n12648,
    n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
    n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
    n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
    n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764, n12766, n12767, n12768,
    n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
    n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
    n12796, n12797, n12798, n12799, n12800, n12801, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12897,
    n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
    n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
    n12934, n12935, n12936, n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13008,
    n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
    n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
    n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
    n13037, n13038, n13040, n13041, n13043, n13044, n13046, n13047, n13049,
    n13050, n13052, n13053, n13055, n13056, n13058, n13059, n13061, n13062,
    n13064, n13065, n13067, n13068, n13070, n13071, n13073, n13074, n13076,
    n13077, n13079, n13080, n13082, n13083, n13085, n13086, n13088, n13089,
    n13091, n13092, n13094, n13095, n13097, n13098, n13100, n13101, n13103,
    n13104, n13106, n13107, n13109, n13110, n13112, n13113, n13115, n13116,
    n13118, n13119, n13121, n13122, n13124, n13125, n13127, n13128, n13130,
    n13131, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
    n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
    n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
    n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
    n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
    n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
    n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
    n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
    n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
    n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
    n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
    n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
    n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
    n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
    n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
    n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
    n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
    n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
    n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
    n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
    n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
    n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
    n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
    n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
    n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
    n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
    n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
    n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
    n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
    n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
    n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
    n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
    n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
    n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
    n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
    n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
    n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
    n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
    n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
    n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
    n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
    n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
    n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
    n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
    n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
    n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
    n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
    n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
    n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
    n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
    n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
    n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
    n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
    n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
    n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
    n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
    n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14275, n14276, n14277, n14278, n14279, n14280,
    n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
    n14290, n14291, n14292, n14293, n14294, n14295, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
    n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
    n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
    n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14421, n14422,
    n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
    n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
    n14460, n14461, n14462, n14463, n14464, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14485, n14486, n14487, n14488,
    n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
    n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
    n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14570, n14571, n14572, n14573,
    n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
    n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
    n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
    n14657, n14658, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
    n14676, n14677, n14678, n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
    n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
    n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
    n14761, n14762, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14786, n14787, n14788, n14789,
    n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
    n14808, n14810, n14811, n14813, n14814, n14815, n14816, n14817, n14818,
    n14819, n14820, n14821, n14822, n14823, n14824, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14843, n14844, n14845, n14846, n14847,
    n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
    n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14909, n14910, n14911, n14912, n14913,
    n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
    n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
    n14970, n14971, n14972, n14974, n14975, n14976, n14977, n14978, n14979,
    n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
    n14998, n14999, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
    n15017, n15018, n15019, n15020, n15021, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
    n15036, n15037, n15038, n15039, n15040, n15041, n15043, n15044, n15045,
    n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
    n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
    n15083, n15084, n15085, n15086, n15087, n15088, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
    n15149, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
    n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
    n15196, n15197, n15198, n15199, n15200, n15201, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
    n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15242, n15243,
    n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
    n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
    n15262, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
    n15281, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
    n15319, n15320, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15345, n15346, n15347,
    n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362, n15364, n15365, n15366,
    n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
    n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
    n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
    n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
    n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
    n15461, n15462, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
    n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
    n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15517,
    n15518, n15519, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
    n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
    n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
    n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
    n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
    n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
    n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
    n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
    n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15733, n15734, n15735, n15736, n15737, n15738,
    n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
    n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
    n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
    n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
    n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
    n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
    n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
    n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
    n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
    n15839, n15840, n15841, n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15903,
    n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
    n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
    n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
    n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
    n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
    n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
    n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
    n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
    n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
    n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
    n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
    n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
    n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16158, n16159,
    n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
    n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
    n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
    n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
    n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
    n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
    n16214, n16215, n16216, n16217, n16218, n16219, n16221, n16222, n16223,
    n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
    n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
    n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
    n16278, n16279, n16280, n16281, n16282, n16283, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
    n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
    n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
    n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
    n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
    n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
    n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
    n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
    n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
    n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
    n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
    n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
    n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
    n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
    n16543, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
    n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
    n16662, n16663, n16664, n16665, n16666, n16667, n16669, n16670, n16671,
    n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
    n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
    n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
    n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
    n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
    n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
    n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
    n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868, n16870, n16871, n16872,
    n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
    n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
    n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
    n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
    n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
    n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
    n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
    n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
    n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
    n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17109, n17110,
    n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
    n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
    n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
    n17165, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
    n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
    n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
    n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
    n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
    n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
    n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
    n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
    n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
    n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
    n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17408, n17409, n17410, n17411, n17412,
    n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
    n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
    n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
    n17467, n17468, n17469, n17470, n17471, n17473, n17474, n17475, n17476,
    n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
    n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
    n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
    n17531, n17532, n17533, n17534, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17549, n17550,
    n17551, n17552, n17553, n17555, n17556, n17557, n17558, n17559, n17560,
    n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17572, n17573, n17575, n17576, n17578, n17579, n17581, n17582,
    n17584, n17585, n17587, n17588, n17590, n17591, n17593, n17594, n17596,
    n17597, n17599, n17600, n17602, n17603, n17605, n17606, n17608, n17609,
    n17611, n17612, n17614, n17615, n17617, n17618, n17620, n17621, n17623,
    n17624, n17626, n17627, n17629, n17630, n17632, n17633, n17635, n17636,
    n17638, n17639, n17641, n17642, n17644, n17645, n17647, n17648, n17650,
    n17651, n17653, n17654, n17656, n17657, n17659, n17660, n17662, n17663,
    n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
    n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
    n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
    n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
    n17722, n17723, n17724, n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17737, n17738, n17739, n17740, n17741,
    n17742, n17743, n17744, n17745, n17746, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17770, n17771,
    n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17781,
    n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
    n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
    n17801, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
    n17821, n17822, n17823, n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17847, n17848, n17849, n17850,
    n17851, n17852, n17853, n17854, n17855, n17856, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
    n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17935, n17936, n17937, n17938, n17939,
    n17940, n17941, n17942, n17943, n17944, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17968, n17969,
    n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
    n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
    n18010, n18011, n18012, n18013, n18014, n18016, n18017, n18018, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
    n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
    n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
    n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
    n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
    n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
    n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
    n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
    n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
    n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
    n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206, n18208, n18209, n18210,
    n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
    n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
    n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
    n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
    n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
    n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
    n18373, n18374, n18375, n18376, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
    n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
    n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
    n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
    n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
    n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18540,
    n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
    n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
    n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
    n18568, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
    n18633, n18634, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
    n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
    n18661, n18662, n18663, n18664, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18731, n18732, n18733, n18734, n18735,
    n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
    n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
    n18754, n18755, n18756, n18757, n18758, n18759, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18827, n18828,
    n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
    n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
    n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18892, n18893,
    n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
    n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
    n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
    n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18982, n18983, n18985, n18986, n18988,
    n18989, n18991, n18992, n18994, n18995, n18997, n18998, n19000, n19001,
    n19003, n19004, n19006, n19007, n19009, n19010, n19012, n19013, n19015,
    n19016, n19018, n19019, n19021, n19022, n19024, n19025, n19027, n19028,
    n19030, n19031, n19033, n19034, n19036, n19037, n19039, n19040, n19042,
    n19043, n19045, n19046, n19048, n19049, n19051, n19052, n19054, n19055,
    n19057, n19058, n19060, n19061, n19063, n19064, n19066, n19067, n19069,
    n19070, n19072, n19073, n19075, n19076, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
    n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
    n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
    n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
    n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
    n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
    n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
    n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
    n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
    n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
    n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
    n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
    n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
    n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
    n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
    n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
    n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
    n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
    n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
    n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
    n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
    n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
    n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
    n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
    n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
    n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19863, n19864, n19865,
    n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
    n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
    n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
    n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
    n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
    n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
    n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
    n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
    n20028, n20029, n20030, n20031, n20032, n20034, n20035, n20036, n20037,
    n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
    n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
    n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
    n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
    n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
    n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
    n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
    n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
    n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
    n20146, n20147, n20148, n20149, n20150, n20151, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
    n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
    n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
    n20212, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
    n20231, n20232, n20233, n20234, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
    n20250, n20251, n20252, n20253, n20254, n20256, n20257, n20258, n20259,
    n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
    n20278, n20279, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
    n20297, n20298, n20299, n20300, n20301, n20302, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
    n20316, n20317, n20318, n20319, n20321, n20322, n20323, n20324, n20325,
    n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
    n20335, n20336, n20337, n20338, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20359, n20360, n20361, n20362, n20363,
    n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378, n20380, n20381, n20382,
    n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
    n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
    n20401, n20402, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
    n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20443, n20444, n20445, n20446, n20447, n20448,
    n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
    n20458, n20459, n20460, n20461, n20462, n20463, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
    n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20509, n20510, n20511, n20512, n20513, n20514,
    n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
    n20524, n20525, n20526, n20527, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
    n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
    n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594, n20596, n20597, n20598,
    n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
    n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
    n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20640, n20641, n20642, n20643, n20644, n20645,
    n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20659, n20660, n20661, n20662, n20663, n20664,
    n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
    n20674, n20675, n20676, n20677, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
    n20693, n20694, n20695, n20696, n20697, n20698, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
    n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20721,
    n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
    n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
    n20740, n20741, n20742, n20743, n20745, n20746, n110, n115, n120, n125,
    n130, n135, n140, n145, n150, n155, n160, n165, n170, n175, n180, n185,
    n190, n195, n200, n205, n210, n215, n220, n225, n230, n235, n240, n245,
    n250, n255, n260, n265, n270, n275, n280, n285, n290, n295, n300, n305,
    n310, n315, n320, n325, n330, n335, n340, n345, n350, n355, n360, n365,
    n370, n375, n380, n385, n390, n395, n400, n405, n410, n415, n420, n425,
    n430, n435, n440, n445, n450, n455, n460, n465, n470, n475, n480, n485,
    n490, n495, n500, n505, n510, n515, n520, n525, n530, n535, n540, n545,
    n550, n555, n560, n565, n570, n575, n580, n585, n590, n595, n600, n605,
    n610, n615, n620, n625, n630, n635, n640, n645, n650, n655, n660, n665,
    n670, n675, n680, n685, n690, n695, n700, n705, n710, n715, n720, n725,
    n730, n735, n740, n745, n750, n755, n760, n765, n770, n775, n780, n785,
    n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840, n845,
    n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900, n905,
    n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960, n965,
    n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015, n1020,
    n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070,
    n1075, n1080, n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1120,
    n1125, n1130, n1135, n1140, n1145, n1150, n1155, n1160, n1165, n1170,
    n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220,
    n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270,
    n1275, n1280, n1285, n1290, n1295, n1300, n1305, n1310, n1315, n1320,
    n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365, n1370,
    n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415, n1420,
    n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465, n1470,
    n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515, n1520,
    n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570,
    n1575, n1580, n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620,
    n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670,
    n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720,
    n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770,
    n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820,
    n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870,
    n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920,
    n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970,
    n1975, n1980, n1985, n1990, n1995, n2000, n2005, n2010, n2015, n2020,
    n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070,
    n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120,
    n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165, n2170,
    n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210, n2215, n2220,
    n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260, n2265, n2270,
    n2275, n2280, n2285, n2290, n2295, n2300, n2305, n2310, n2315, n2320,
    n2325, n2330, n2335, n2340, n2345, n2350, n2355, n2360, n2365, n2370,
    n2375, n2380, n2385, n2390, n2395, n2400, n2405, n2410, n2415, n2420,
    n2425, n2430, n2435, n2440, n2445, n2450, n2455, n2460, n2465, n2470,
    n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520,
    n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570,
    n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620,
    n2625, n2630, n2635, n2640, n2645, n2650, n2655, n2660, n2665, n2670,
    n2675, n2680, n2685, n2690, n2695, n2700, n2705, n2710, n2715, n2720,
    n2725, n2730, n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770,
    n2775, n2780, n2785, n2790, n2795, n2800, n2805, n2810, n2815, n2820,
    n2825, n2830, n2835, n2840, n2845, n2850, n2855, n2860, n2865, n2870,
    n2875, n2880, n2885, n2890, n2895, n2900, n2905, n2910, n2915, n2920,
    n2925, n2930, n2935, n2940, n2945, n2950, n2955, n2960, n2965, n2970,
    n2975, n2980, n2985, n2990, n2995, n3000, n3005, n3010, n3015, n3020,
    n3025, n3030, n3035, n3040, n3045, n3050, n3055, n3060, n3065, n3070,
    n3075, n3080, n3085, n3090, n3095, n3100, n3105, n3110, n3115, n3120,
    n3125, n3130, n3135, n3140, n3145, n3150, n3155, n3160, n3165, n3170,
    n3175, n3180, n3185, n3190, n3195, n3200, n3205, n3210, n3215, n3220,
    n3225, n3230, n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270,
    n3275, n3280, n3285, n3290, n3295, n3300, n3305, n3310, n3315, n3320,
    n3325, n3330, n3335, n3340, n3345, n3350, n3355, n3360, n3365, n3370,
    n3375, n3380, n3385, n3390, n3395, n3400, n3405, n3410, n3415, n3420,
    n3425, n3430, n3435, n3440, n3445, n3450, n3455, n3460, n3465, n3470,
    n3475, n3480, n3485, n3490, n3495, n3500, n3505, n3510, n3515, n3520,
    n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570,
    n3575, n3580, n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620,
    n3625, n3630, n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670,
    n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720,
    n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770,
    n3775, n3780;
  assign n2260_1 = P1_ADDR_REG_17_ & ~P3_ADDR_REG_17_;
  assign n2261 = ~P1_ADDR_REG_17_ & P3_ADDR_REG_17_;
  assign n2262 = ~n2260_1 & ~n2261;
  assign n2263 = P1_ADDR_REG_16_ & ~P3_ADDR_REG_16_;
  assign n2264 = ~P1_ADDR_REG_16_ & P3_ADDR_REG_16_;
  assign n2265_1 = P1_ADDR_REG_15_ & ~P3_ADDR_REG_15_;
  assign n2266 = ~P1_ADDR_REG_15_ & P3_ADDR_REG_15_;
  assign n2267 = P1_ADDR_REG_14_ & ~P3_ADDR_REG_14_;
  assign n2268 = ~P1_ADDR_REG_14_ & P3_ADDR_REG_14_;
  assign n2269 = P1_ADDR_REG_13_ & ~P3_ADDR_REG_13_;
  assign n2270_1 = ~P1_ADDR_REG_13_ & P3_ADDR_REG_13_;
  assign n2271 = P1_ADDR_REG_12_ & ~P3_ADDR_REG_12_;
  assign n2272 = ~P1_ADDR_REG_12_ & P3_ADDR_REG_12_;
  assign n2273 = P1_ADDR_REG_11_ & ~P3_ADDR_REG_11_;
  assign n2274 = ~P1_ADDR_REG_11_ & P3_ADDR_REG_11_;
  assign n2275_1 = P1_ADDR_REG_10_ & ~P3_ADDR_REG_10_;
  assign n2276 = ~P1_ADDR_REG_10_ & P3_ADDR_REG_10_;
  assign n2277 = P1_ADDR_REG_9_ & ~P3_ADDR_REG_9_;
  assign n2278 = ~P1_ADDR_REG_9_ & P3_ADDR_REG_9_;
  assign n2279 = P1_ADDR_REG_8_ & ~P3_ADDR_REG_8_;
  assign n2280_1 = ~P1_ADDR_REG_8_ & P3_ADDR_REG_8_;
  assign n2281 = P1_ADDR_REG_7_ & ~P3_ADDR_REG_7_;
  assign n2282 = ~P1_ADDR_REG_7_ & P3_ADDR_REG_7_;
  assign n2283 = P1_ADDR_REG_6_ & ~P3_ADDR_REG_6_;
  assign n2284 = ~P1_ADDR_REG_6_ & P3_ADDR_REG_6_;
  assign n2285_1 = P1_ADDR_REG_5_ & ~P3_ADDR_REG_5_;
  assign n2286 = ~P1_ADDR_REG_5_ & P3_ADDR_REG_5_;
  assign n2287 = P1_ADDR_REG_4_ & ~P3_ADDR_REG_4_;
  assign n2288 = ~P1_ADDR_REG_4_ & P3_ADDR_REG_4_;
  assign n2289 = P1_ADDR_REG_3_ & ~P3_ADDR_REG_3_;
  assign n2290_1 = ~P1_ADDR_REG_3_ & P3_ADDR_REG_3_;
  assign n2291 = P1_ADDR_REG_2_ & ~P3_ADDR_REG_2_;
  assign n2292 = ~P1_ADDR_REG_2_ & P3_ADDR_REG_2_;
  assign n2293 = ~P1_ADDR_REG_0_ & P3_ADDR_REG_0_;
  assign n2294 = P1_ADDR_REG_1_ & ~n2293;
  assign n2295_1 = ~P1_ADDR_REG_1_ & n2293;
  assign n2296 = ~P3_ADDR_REG_1_ & ~n2295_1;
  assign n2297 = ~n2294 & ~n2296;
  assign n2298 = ~n2292 & ~n2297;
  assign n2299 = ~n2291 & ~n2298;
  assign n2300_1 = ~n2290_1 & ~n2299;
  assign n2301 = ~n2289 & ~n2300_1;
  assign n2302 = ~n2288 & ~n2301;
  assign n2303 = ~n2287 & ~n2302;
  assign n2304 = ~n2286 & ~n2303;
  assign n2305_1 = ~n2285_1 & ~n2304;
  assign n2306 = ~n2284 & ~n2305_1;
  assign n2307 = ~n2283 & ~n2306;
  assign n2308 = ~n2282 & ~n2307;
  assign n2309 = ~n2281 & ~n2308;
  assign n2310_1 = ~n2280_1 & ~n2309;
  assign n2311 = ~n2279 & ~n2310_1;
  assign n2312 = ~n2278 & ~n2311;
  assign n2313 = ~n2277 & ~n2312;
  assign n2314 = ~n2276 & ~n2313;
  assign n2315_1 = ~n2275_1 & ~n2314;
  assign n2316 = ~n2274 & ~n2315_1;
  assign n2317 = ~n2273 & ~n2316;
  assign n2318 = ~n2272 & ~n2317;
  assign n2319 = ~n2271 & ~n2318;
  assign n2320_1 = ~n2270_1 & ~n2319;
  assign n2321 = ~n2269 & ~n2320_1;
  assign n2322 = ~n2268 & ~n2321;
  assign n2323 = ~n2267 & ~n2322;
  assign n2324 = ~n2266 & ~n2323;
  assign n2325_1 = ~n2265_1 & ~n2324;
  assign n2326 = ~n2264 & ~n2325_1;
  assign n2327 = ~n2263 & ~n2326;
  assign n2328 = ~n2262 & ~n2327;
  assign n2329 = n2262 & n2327;
  assign n2330_1 = ~n2328 & ~n2329;
  assign n2331 = P2_ADDR_REG_17_ & ~n2330_1;
  assign n2332 = ~P2_ADDR_REG_17_ & n2330_1;
  assign n2333 = ~n2263 & ~n2264;
  assign n2334 = ~n2325_1 & ~n2333;
  assign n2335_1 = n2325_1 & n2333;
  assign n2336 = ~n2334 & ~n2335_1;
  assign n2337 = P2_ADDR_REG_16_ & ~n2336;
  assign n2338 = ~P2_ADDR_REG_16_ & n2336;
  assign n2339 = ~n2271 & ~n2272;
  assign n2340_1 = ~n2317 & ~n2339;
  assign n2341 = n2317 & n2339;
  assign n2342 = ~n2340_1 & ~n2341;
  assign n2343 = P2_ADDR_REG_12_ & ~n2342;
  assign n2344 = ~P2_ADDR_REG_12_ & n2342;
  assign n2345_1 = ~n2273 & ~n2274;
  assign n2346 = ~n2315_1 & ~n2345_1;
  assign n2347 = n2315_1 & n2345_1;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = P2_ADDR_REG_11_ & ~n2348;
  assign n2350_1 = ~P2_ADDR_REG_11_ & n2348;
  assign n2351 = ~n2277 & ~n2278;
  assign n2352 = ~n2311 & ~n2351;
  assign n2353 = n2311 & n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355_1 = P2_ADDR_REG_9_ & ~n2354;
  assign n2356 = ~P2_ADDR_REG_9_ & n2354;
  assign n2357 = ~n2281 & ~n2282;
  assign n2358 = ~n2307 & ~n2357;
  assign n2359 = n2307 & n2357;
  assign n2360_1 = ~n2358 & ~n2359;
  assign n2361 = P2_ADDR_REG_7_ & ~n2360_1;
  assign n2362 = ~P2_ADDR_REG_7_ & n2360_1;
  assign n2363 = ~n2283 & ~n2284;
  assign n2364 = ~n2305_1 & ~n2363;
  assign n2365_1 = n2305_1 & n2363;
  assign n2366 = ~n2364 & ~n2365_1;
  assign n2367 = P2_ADDR_REG_6_ & ~n2366;
  assign n2368 = ~P2_ADDR_REG_6_ & n2366;
  assign n2369 = ~n2287 & ~n2288;
  assign n2370_1 = ~n2301 & ~n2369;
  assign n2371 = n2301 & n2369;
  assign n2372 = ~n2370_1 & ~n2371;
  assign n2373 = P2_ADDR_REG_4_ & ~n2372;
  assign n2374 = ~P2_ADDR_REG_4_ & n2372;
  assign n2375_1 = ~n2291 & ~n2292;
  assign n2376 = ~n2297 & ~n2375_1;
  assign n2377 = n2297 & n2375_1;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = P2_ADDR_REG_2_ & ~n2378;
  assign n2380_1 = ~P2_ADDR_REG_2_ & n2378;
  assign n2381 = P1_ADDR_REG_1_ & ~P3_ADDR_REG_1_;
  assign n2382 = ~P1_ADDR_REG_1_ & P3_ADDR_REG_1_;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2293 & ~n2383;
  assign n2385_1 = n2293 & n2383;
  assign n2386 = ~n2384 & ~n2385_1;
  assign n2387 = P1_ADDR_REG_0_ & ~P3_ADDR_REG_0_;
  assign n2388 = ~n2293 & ~n2387;
  assign n2389 = P2_ADDR_REG_0_ & ~n2388;
  assign n2390_1 = ~n2386 & n2389;
  assign n2391 = n2386 & ~n2389;
  assign n2392 = P2_ADDR_REG_1_ & ~n2391;
  assign n2393 = ~n2390_1 & ~n2392;
  assign n2394 = ~n2380_1 & ~n2393;
  assign n2395_1 = ~n2379 & ~n2394;
  assign n2396 = P2_ADDR_REG_3_ & ~n2395_1;
  assign n2397 = ~n2289 & ~n2290_1;
  assign n2398 = ~n2299 & ~n2397;
  assign n2399 = n2299 & n2397;
  assign n2400_1 = ~n2398 & ~n2399;
  assign n2401 = ~P2_ADDR_REG_3_ & n2395_1;
  assign n2402 = ~n2400_1 & ~n2401;
  assign n2403 = ~n2396 & ~n2402;
  assign n2404 = ~n2374 & ~n2403;
  assign n2405_1 = ~n2373 & ~n2404;
  assign n2406 = P2_ADDR_REG_5_ & ~n2405_1;
  assign n2407 = ~n2285_1 & ~n2286;
  assign n2408 = ~n2303 & ~n2407;
  assign n2409 = n2303 & n2407;
  assign n2410_1 = ~n2408 & ~n2409;
  assign n2411 = ~P2_ADDR_REG_5_ & n2405_1;
  assign n2412 = ~n2410_1 & ~n2411;
  assign n2413 = ~n2406 & ~n2412;
  assign n2414 = ~n2368 & ~n2413;
  assign n2415_1 = ~n2367 & ~n2414;
  assign n2416 = ~n2362 & ~n2415_1;
  assign n2417 = ~n2361 & ~n2416;
  assign n2418 = P2_ADDR_REG_8_ & ~n2417;
  assign n2419 = ~n2279 & ~n2280_1;
  assign n2420_1 = ~n2309 & ~n2419;
  assign n2421 = n2309 & n2419;
  assign n2422 = ~n2420_1 & ~n2421;
  assign n2423 = ~P2_ADDR_REG_8_ & n2417;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425_1 = ~n2418 & ~n2424;
  assign n2426 = ~n2356 & ~n2425_1;
  assign n2427 = ~n2355_1 & ~n2426;
  assign n2428 = P2_ADDR_REG_10_ & ~n2427;
  assign n2429 = ~n2275_1 & ~n2276;
  assign n2430_1 = ~n2313 & ~n2429;
  assign n2431 = n2313 & n2429;
  assign n2432 = ~n2430_1 & ~n2431;
  assign n2433 = ~P2_ADDR_REG_10_ & n2427;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435_1 = ~n2428 & ~n2434;
  assign n2436 = ~n2350_1 & ~n2435_1;
  assign n2437 = ~n2349 & ~n2436;
  assign n2438 = ~n2344 & ~n2437;
  assign n2439 = ~n2343 & ~n2438;
  assign n2440_1 = P2_ADDR_REG_13_ & ~n2439;
  assign n2441 = ~n2269 & ~n2270_1;
  assign n2442 = ~n2319 & ~n2441;
  assign n2443 = n2319 & n2441;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445_1 = ~P2_ADDR_REG_13_ & n2439;
  assign n2446 = ~n2444 & ~n2445_1;
  assign n2447 = ~n2440_1 & ~n2446;
  assign n2448 = P2_ADDR_REG_14_ & ~n2447;
  assign n2449 = ~n2267 & ~n2268;
  assign n2450_1 = ~n2321 & ~n2449;
  assign n2451 = n2321 & n2449;
  assign n2452 = ~n2450_1 & ~n2451;
  assign n2453 = ~P2_ADDR_REG_14_ & n2447;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455_1 = ~n2448 & ~n2454;
  assign n2456 = P2_ADDR_REG_15_ & ~n2455_1;
  assign n2457 = ~n2265_1 & ~n2266;
  assign n2458 = ~n2323 & ~n2457;
  assign n2459 = n2323 & n2457;
  assign n2460_1 = ~n2458 & ~n2459;
  assign n2461 = ~P2_ADDR_REG_15_ & n2455_1;
  assign n2462 = ~n2460_1 & ~n2461;
  assign n2463 = ~n2456 & ~n2462;
  assign n2464 = ~n2338 & ~n2463;
  assign n2465_1 = ~n2337 & ~n2464;
  assign n2466 = ~n2332 & ~n2465_1;
  assign n2467 = ~n2331 & ~n2466;
  assign n2468 = ~P2_ADDR_REG_18_ & n2467;
  assign n2469 = P2_ADDR_REG_18_ & ~n2467;
  assign n2470_1 = P1_ADDR_REG_18_ & ~P3_ADDR_REG_18_;
  assign n2471 = ~P1_ADDR_REG_18_ & P3_ADDR_REG_18_;
  assign n2472 = ~n2470_1 & ~n2471;
  assign n2473 = ~n2261 & ~n2327;
  assign n2474 = ~n2260_1 & ~n2473;
  assign n2475_1 = ~n2472 & ~n2474;
  assign n2476 = n2472 & n2474;
  assign n2477 = ~n2475_1 & ~n2476;
  assign n2478 = ~n2469 & n2477;
  assign n2479 = P1_ADDR_REG_19_ & ~P3_ADDR_REG_19_;
  assign n2480_1 = ~P1_ADDR_REG_19_ & P3_ADDR_REG_19_;
  assign n2481 = ~n2479 & ~n2480_1;
  assign n2482 = ~n2470_1 & n2474;
  assign n2483 = ~n2471 & ~n2481;
  assign n2484 = ~n2482 & n2483;
  assign n2485_1 = ~n2471 & ~n2474;
  assign n2486 = ~n2470_1 & n2481;
  assign n2487 = ~n2485_1 & n2486;
  assign n2488 = ~n2484 & ~n2487;
  assign n2489 = ~P2_ADDR_REG_19_ & ~n2488;
  assign n2490_1 = P2_ADDR_REG_19_ & n2488;
  assign n2491 = ~n2489 & ~n2490_1;
  assign n2492 = ~n2468 & ~n2478;
  assign n2493 = ~n2491 & n2492;
  assign n2494 = ~n2468 & ~n2477;
  assign n2495_1 = ~n2469 & ~n2494;
  assign n2496 = ~n2489 & n2495_1;
  assign n2497 = ~n2490_1 & n2496;
  assign SUB_1596_U4 = ~n2493 & ~n2497;
  assign n2499 = ~n2468 & ~n2469;
  assign n2500_1 = ~n2477 & ~n2499;
  assign n2501 = n2477 & n2499;
  assign SUB_1596_U62 = n2500_1 | n2501;
  assign n2503 = ~P2_ADDR_REG_17_ & ~n2330_1;
  assign n2504 = P2_ADDR_REG_17_ & n2330_1;
  assign n2505_1 = ~n2503 & ~n2504;
  assign n2506 = n2465_1 & ~n2505_1;
  assign n2507 = ~n2465_1 & n2505_1;
  assign SUB_1596_U63 = n2506 | n2507;
  assign n2509 = ~P2_ADDR_REG_16_ & ~n2336;
  assign n2510_1 = P2_ADDR_REG_16_ & n2336;
  assign n2511 = ~n2509 & ~n2510_1;
  assign n2512 = n2463 & ~n2511;
  assign n2513 = ~n2463 & n2511;
  assign SUB_1596_U64 = n2512 | n2513;
  assign n2515_1 = ~n2456 & ~n2461;
  assign n2516 = ~n2460_1 & ~n2515_1;
  assign n2517 = n2460_1 & n2515_1;
  assign SUB_1596_U65 = n2516 | n2517;
  assign n2519 = ~n2448 & ~n2453;
  assign n2520_1 = ~n2452 & ~n2519;
  assign n2521 = n2452 & n2519;
  assign SUB_1596_U66 = n2520_1 | n2521;
  assign n2523 = ~n2440_1 & ~n2445_1;
  assign n2524 = ~n2444 & ~n2523;
  assign n2525_1 = n2444 & n2523;
  assign SUB_1596_U67 = n2524 | n2525_1;
  assign n2527 = ~P2_ADDR_REG_12_ & ~n2342;
  assign n2528 = P2_ADDR_REG_12_ & n2342;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530_1 = n2437 & ~n2529;
  assign n2531 = ~n2437 & n2529;
  assign SUB_1596_U68 = n2530_1 | n2531;
  assign n2533 = ~P2_ADDR_REG_11_ & ~n2348;
  assign n2534 = P2_ADDR_REG_11_ & n2348;
  assign n2535_1 = ~n2533 & ~n2534;
  assign n2536 = n2435_1 & ~n2535_1;
  assign n2537 = ~n2435_1 & n2535_1;
  assign SUB_1596_U69 = n2536 | n2537;
  assign n2539 = ~n2428 & ~n2433;
  assign n2540_1 = ~n2432 & ~n2539;
  assign n2541 = n2432 & n2539;
  assign SUB_1596_U70 = n2540_1 | n2541;
  assign n2543 = ~P2_ADDR_REG_9_ & ~n2354;
  assign n2544 = P2_ADDR_REG_9_ & n2354;
  assign n2545_1 = ~n2543 & ~n2544;
  assign n2546 = n2425_1 & ~n2545_1;
  assign n2547 = ~n2425_1 & n2545_1;
  assign SUB_1596_U54 = n2546 | n2547;
  assign n2549 = ~n2418 & ~n2423;
  assign n2550_1 = ~n2422 & ~n2549;
  assign n2551 = n2422 & n2549;
  assign SUB_1596_U55 = n2550_1 | n2551;
  assign n2553 = ~P2_ADDR_REG_7_ & ~n2360_1;
  assign n2554 = P2_ADDR_REG_7_ & n2360_1;
  assign n2555_1 = ~n2553 & ~n2554;
  assign n2556 = n2415_1 & ~n2555_1;
  assign n2557 = ~n2415_1 & n2555_1;
  assign SUB_1596_U56 = n2556 | n2557;
  assign n2559 = ~P2_ADDR_REG_6_ & ~n2366;
  assign n2560_1 = P2_ADDR_REG_6_ & n2366;
  assign n2561 = ~n2559 & ~n2560_1;
  assign n2562 = n2413 & ~n2561;
  assign n2563 = ~n2413 & n2561;
  assign SUB_1596_U57 = n2562 | n2563;
  assign n2565_1 = ~n2406 & ~n2411;
  assign n2566 = ~n2410_1 & ~n2565_1;
  assign n2567 = n2410_1 & n2565_1;
  assign SUB_1596_U58 = n2566 | n2567;
  assign n2569 = ~P2_ADDR_REG_4_ & ~n2372;
  assign n2570_1 = P2_ADDR_REG_4_ & n2372;
  assign n2571 = ~n2569 & ~n2570_1;
  assign n2572 = n2403 & ~n2571;
  assign n2573 = ~n2403 & n2571;
  assign SUB_1596_U59 = n2572 | n2573;
  assign n2575_1 = ~n2396 & ~n2401;
  assign n2576 = ~n2400_1 & ~n2575_1;
  assign n2577 = n2400_1 & n2575_1;
  assign SUB_1596_U60 = n2576 | n2577;
  assign n2579 = ~P2_ADDR_REG_2_ & ~n2378;
  assign n2580_1 = P2_ADDR_REG_2_ & n2378;
  assign n2581 = ~n2579 & ~n2580_1;
  assign n2582 = n2393 & ~n2581;
  assign n2583 = ~n2393 & n2581;
  assign SUB_1596_U61 = n2582 | n2583;
  assign n2585_1 = P2_ADDR_REG_1_ & n2390_1;
  assign n2586 = ~n2386 & ~n2389;
  assign n2587 = ~P2_ADDR_REG_1_ & n2586;
  assign n2588 = ~P2_ADDR_REG_1_ & n2389;
  assign n2589 = P2_ADDR_REG_1_ & ~n2389;
  assign n2590_1 = ~n2588 & ~n2589;
  assign n2591 = n2386 & ~n2590_1;
  assign n2592 = ~n2585_1 & ~n2587;
  assign SUB_1596_U5 = n2591 | ~n2592;
  assign n2594 = ~P2_ADDR_REG_0_ & ~n2388;
  assign n2595_1 = P2_ADDR_REG_0_ & n2388;
  assign SUB_1596_U53 = n2594 | n2595_1;
  assign n2597 = P1_RD_REG & ~P2_RD_REG;
  assign n2598 = ~P1_RD_REG & P2_RD_REG;
  assign n2599 = ~n2597 & ~n2598;
  assign U29 = P3_RD_REG | n2599;
  assign n2601 = P1_WR_REG & ~P2_WR_REG;
  assign n2602 = ~P1_WR_REG & P2_WR_REG;
  assign n2603 = ~n2601 & ~n2602;
  assign U28 = P3_WR_REG | n2603;
  assign n2605_1 = ~P1_IR_REG_31_ & P1_STATE_REG;
  assign n2606 = P1_STATE_REG & ~n2605_1;
  assign n2607 = P1_IR_REG_0_ & n2606;
  assign n2608 = P1_IR_REG_0_ & n2605_1;
  assign n2609 = ~P1_ADDR_REG_19_ & ~P2_ADDR_REG_19_;
  assign n2610_1 = P3_ADDR_REG_19_ & n2609;
  assign n2611 = ~P1_RD_REG & n2610_1;
  assign n2612 = P1_ADDR_REG_19_ & P2_ADDR_REG_19_;
  assign n2613 = ~P3_ADDR_REG_19_ & n2612;
  assign n2614 = ~P2_RD_REG & n2613;
  assign n2615_1 = ~n2611 & ~n2614;
  assign n2616 = P2_DATAO_REG_0_ & n2615_1;
  assign n2617 = P1_DATAO_REG_0_ & n2615_1;
  assign n2618 = P2_DATAO_REG_0_ & ~n2615_1;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620_1 = SI_0_ & n2619;
  assign n2621 = ~SI_0_ & ~n2619;
  assign n2622 = ~n2620_1 & ~n2621;
  assign n2623 = ~n2615_1 & ~n2622;
  assign n2624 = ~n2616 & ~n2623;
  assign n2625_1 = ~P1_STATE_REG & ~n2624;
  assign n2626 = ~n2607 & ~n2608;
  assign n110 = n2625_1 | ~n2626;
  assign n2628 = P1_IR_REG_0_ & ~P1_IR_REG_1_;
  assign n2629 = ~P1_IR_REG_0_ & P1_IR_REG_1_;
  assign n2630_1 = ~n2628 & ~n2629;
  assign n2631 = n2606 & ~n2630_1;
  assign n2632 = P1_IR_REG_1_ & n2605_1;
  assign n2633 = P2_DATAO_REG_1_ & n2615_1;
  assign n2634 = SI_1_ & SI_0_;
  assign n2635_1 = ~n2619 & n2634;
  assign n2636 = P1_DATAO_REG_1_ & n2615_1;
  assign n2637 = P2_DATAO_REG_1_ & ~n2615_1;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = n2635_1 & ~n2638;
  assign n2640_1 = SI_0_ & ~n2619;
  assign n2641 = SI_1_ & ~n2640_1;
  assign n2642 = n2638 & n2641;
  assign n2643 = ~n2639 & ~n2642;
  assign n2644 = n2638 & n2640_1;
  assign n2645_1 = ~n2638 & ~n2640_1;
  assign n2646 = ~n2644 & ~n2645_1;
  assign n2647 = ~SI_1_ & ~n2646;
  assign n2648 = n2643 & ~n2647;
  assign n2649 = ~n2615_1 & ~n2648;
  assign n2650_1 = ~n2633 & ~n2649;
  assign n2651 = ~P1_STATE_REG & ~n2650_1;
  assign n2652 = ~n2631 & ~n2632;
  assign n115 = n2651 | ~n2652;
  assign n2654 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_;
  assign n2655_1 = P1_IR_REG_2_ & ~n2654;
  assign n2656 = ~P1_IR_REG_2_ & n2654;
  assign n2657 = ~n2655_1 & ~n2656;
  assign n2658 = n2606 & n2657;
  assign n2659 = P1_IR_REG_2_ & n2605_1;
  assign n2660_1 = P2_DATAO_REG_2_ & n2615_1;
  assign n2661 = SI_1_ & ~n2638;
  assign n2662 = ~n2638 & n2640_1;
  assign n2663 = ~n2635_1 & ~n2661;
  assign n2664 = ~n2662 & n2663;
  assign n2665_1 = P1_DATAO_REG_2_ & n2615_1;
  assign n2666 = P2_DATAO_REG_2_ & ~n2615_1;
  assign n2667 = ~n2665_1 & ~n2666;
  assign n2668 = SI_2_ & n2667;
  assign n2669 = ~SI_2_ & ~n2667;
  assign n2670_1 = ~n2668 & ~n2669;
  assign n2671 = n2664 & ~n2670_1;
  assign n2672 = ~n2664 & n2670_1;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~n2615_1 & ~n2673;
  assign n2675_1 = ~n2660_1 & ~n2674;
  assign n2676 = ~P1_STATE_REG & ~n2675_1;
  assign n2677 = ~n2658 & ~n2659;
  assign n120 = n2676 | ~n2677;
  assign n2679 = P1_IR_REG_3_ & ~n2656;
  assign n2680_1 = ~P1_IR_REG_3_ & n2656;
  assign n2681 = ~n2679 & ~n2680_1;
  assign n2682 = n2606 & n2681;
  assign n2683 = P1_IR_REG_3_ & n2605_1;
  assign n2684 = P2_DATAO_REG_3_ & n2615_1;
  assign n2685_1 = ~SI_2_ & n2667;
  assign n2686 = n2661 & ~n2685_1;
  assign n2687 = SI_1_ & ~n2685_1;
  assign n2688 = n2640_1 & n2687;
  assign n2689 = ~n2619 & ~n2638;
  assign n2690_1 = SI_0_ & ~n2685_1;
  assign n2691 = n2689 & n2690_1;
  assign n2692 = SI_2_ & ~n2667;
  assign n2693 = ~n2686 & ~n2688;
  assign n2694 = ~n2691 & n2693;
  assign n2695_1 = ~n2692 & n2694;
  assign n2696 = P1_DATAO_REG_3_ & n2615_1;
  assign n2697 = P2_DATAO_REG_3_ & ~n2615_1;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = SI_3_ & n2698;
  assign n2700_1 = ~SI_3_ & ~n2698;
  assign n2701 = ~n2699 & ~n2700_1;
  assign n2702 = n2695_1 & ~n2701;
  assign n2703 = ~n2695_1 & n2701;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705_1 = ~n2615_1 & ~n2704;
  assign n2706 = ~n2684 & ~n2705_1;
  assign n2707 = ~P1_STATE_REG & ~n2706;
  assign n2708 = ~n2682 & ~n2683;
  assign n125 = n2707 | ~n2708;
  assign n2710_1 = P1_IR_REG_4_ & ~n2680_1;
  assign n2711 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign n2712 = n2656 & n2711;
  assign n2713 = ~n2710_1 & ~n2712;
  assign n2714 = n2606 & n2713;
  assign n2715_1 = P1_IR_REG_4_ & n2605_1;
  assign n2716 = P2_DATAO_REG_4_ & n2615_1;
  assign n2717 = ~SI_3_ & n2698;
  assign n2718 = n2692 & ~n2717;
  assign n2719 = SI_3_ & ~n2698;
  assign n2720_1 = ~n2718 & ~n2719;
  assign n2721 = ~n2685_1 & ~n2717;
  assign n2722 = ~n2664 & n2721;
  assign n2723 = n2720_1 & ~n2722;
  assign n2724 = P1_DATAO_REG_4_ & n2615_1;
  assign n2725_1 = P2_DATAO_REG_4_ & ~n2615_1;
  assign n2726 = ~n2724 & ~n2725_1;
  assign n2727 = SI_4_ & n2726;
  assign n2728 = ~SI_4_ & ~n2726;
  assign n2729 = ~n2727 & ~n2728;
  assign n2730_1 = n2723 & ~n2729;
  assign n2731 = ~n2723 & n2729;
  assign n2732 = ~n2730_1 & ~n2731;
  assign n2733 = ~n2615_1 & ~n2732;
  assign n2734 = ~n2716 & ~n2733;
  assign n2735_1 = ~P1_STATE_REG & ~n2734;
  assign n2736 = ~n2714 & ~n2715_1;
  assign n130 = n2735_1 | ~n2736;
  assign n2738 = ~P1_IR_REG_5_ & n2712;
  assign n2739 = P1_IR_REG_5_ & ~n2712;
  assign n2740_1 = ~n2738 & ~n2739;
  assign n2741 = n2606 & n2740_1;
  assign n2742 = P1_IR_REG_5_ & n2605_1;
  assign n2743 = P2_DATAO_REG_5_ & n2615_1;
  assign n2744 = SI_4_ & ~n2726;
  assign n2745_1 = ~SI_4_ & n2726;
  assign n2746 = ~n2723 & ~n2745_1;
  assign n2747 = ~n2744 & ~n2746;
  assign n2748 = P1_DATAO_REG_5_ & n2615_1;
  assign n2749 = P2_DATAO_REG_5_ & ~n2615_1;
  assign n2750_1 = ~n2748 & ~n2749;
  assign n2751 = SI_5_ & n2750_1;
  assign n2752 = ~SI_5_ & ~n2750_1;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = n2747 & ~n2753;
  assign n2755_1 = ~n2747 & n2753;
  assign n2756 = ~n2754 & ~n2755_1;
  assign n2757 = ~n2615_1 & ~n2756;
  assign n2758 = ~n2743 & ~n2757;
  assign n2759 = ~P1_STATE_REG & ~n2758;
  assign n2760_1 = ~n2741 & ~n2742;
  assign n135 = n2759 | ~n2760_1;
  assign n2762 = P1_IR_REG_6_ & ~n2738;
  assign n2763 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_;
  assign n2764 = n2712 & n2763;
  assign n2765_1 = ~n2762 & ~n2764;
  assign n2766 = n2606 & n2765_1;
  assign n2767 = P1_IR_REG_6_ & n2605_1;
  assign n2768 = P2_DATAO_REG_6_ & n2615_1;
  assign n2769 = ~SI_5_ & n2750_1;
  assign n2770_1 = n2744 & ~n2769;
  assign n2771 = SI_5_ & ~n2750_1;
  assign n2772 = ~n2770_1 & ~n2771;
  assign n2773 = ~n2745_1 & ~n2769;
  assign n2774 = ~n2723 & n2773;
  assign n2775_1 = n2772 & ~n2774;
  assign n2776 = P1_DATAO_REG_6_ & n2615_1;
  assign n2777 = P2_DATAO_REG_6_ & ~n2615_1;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = SI_6_ & n2778;
  assign n2780_1 = ~SI_6_ & ~n2778;
  assign n2781 = ~n2779 & ~n2780_1;
  assign n2782 = n2775_1 & ~n2781;
  assign n2783 = ~n2775_1 & n2781;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785_1 = ~n2615_1 & ~n2784;
  assign n2786 = ~n2768 & ~n2785_1;
  assign n2787 = ~P1_STATE_REG & ~n2786;
  assign n2788 = ~n2766 & ~n2767;
  assign n140 = n2787 | ~n2788;
  assign n2790_1 = P1_IR_REG_7_ & ~n2764;
  assign n2791 = ~P1_IR_REG_7_ & n2764;
  assign n2792 = ~n2790_1 & ~n2791;
  assign n2793 = n2606 & n2792;
  assign n2794 = P1_IR_REG_7_ & n2605_1;
  assign n2795_1 = P2_DATAO_REG_7_ & n2615_1;
  assign n2796 = ~SI_6_ & n2778;
  assign n2797 = ~n2772 & ~n2796;
  assign n2798 = SI_6_ & ~n2778;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800_1 = n2773 & ~n2796;
  assign n2801 = ~n2723 & n2800_1;
  assign n2802 = n2799 & ~n2801;
  assign n2803 = P1_DATAO_REG_7_ & n2615_1;
  assign n2804 = P2_DATAO_REG_7_ & ~n2615_1;
  assign n2805_1 = ~n2803 & ~n2804;
  assign n2806 = SI_7_ & n2805_1;
  assign n2807 = ~SI_7_ & ~n2805_1;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n2802 & ~n2808;
  assign n2810_1 = ~n2802 & n2808;
  assign n2811 = ~n2809 & ~n2810_1;
  assign n2812 = ~n2615_1 & ~n2811;
  assign n2813 = ~n2795_1 & ~n2812;
  assign n2814 = ~P1_STATE_REG & ~n2813;
  assign n2815_1 = ~n2793 & ~n2794;
  assign n145 = n2814 | ~n2815_1;
  assign n2817 = P1_IR_REG_8_ & ~n2791;
  assign n2818 = ~P1_IR_REG_7_ & ~P1_IR_REG_8_;
  assign n2819 = ~P1_IR_REG_5_ & n2711;
  assign n2820_1 = ~P1_IR_REG_6_ & n2819;
  assign n2821 = n2656 & n2818;
  assign n2822 = n2820_1 & n2821;
  assign n2823 = ~n2817 & ~n2822;
  assign n2824 = n2606 & n2823;
  assign n2825_1 = P1_IR_REG_8_ & n2605_1;
  assign n2826 = P2_DATAO_REG_8_ & n2615_1;
  assign n2827 = ~SI_7_ & n2805_1;
  assign n2828 = ~n2802 & ~n2827;
  assign n2829 = SI_7_ & ~n2805_1;
  assign n2830_1 = ~n2828 & ~n2829;
  assign n2831 = P1_DATAO_REG_8_ & n2615_1;
  assign n2832 = P2_DATAO_REG_8_ & ~n2615_1;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = SI_8_ & n2833;
  assign n2835_1 = ~SI_8_ & ~n2833;
  assign n2836 = ~n2834 & ~n2835_1;
  assign n2837 = n2830_1 & ~n2836;
  assign n2838 = ~n2830_1 & n2836;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840_1 = ~n2615_1 & ~n2839;
  assign n2841 = ~n2826 & ~n2840_1;
  assign n2842 = ~P1_STATE_REG & ~n2841;
  assign n2843 = ~n2824 & ~n2825_1;
  assign n150 = n2842 | ~n2843;
  assign n2845_1 = ~P1_IR_REG_9_ & n2822;
  assign n2846 = P1_IR_REG_9_ & ~n2822;
  assign n2847 = ~n2845_1 & ~n2846;
  assign n2848 = n2606 & n2847;
  assign n2849 = P1_IR_REG_9_ & n2605_1;
  assign n2850_1 = P2_DATAO_REG_9_ & n2615_1;
  assign n2851 = ~SI_8_ & n2833;
  assign n2852 = n2829 & ~n2851;
  assign n2853 = SI_8_ & ~n2833;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855_1 = ~n2827 & ~n2851;
  assign n2856 = ~n2802 & n2855_1;
  assign n2857 = n2854 & ~n2856;
  assign n2858 = P1_DATAO_REG_9_ & n2615_1;
  assign n2859 = P2_DATAO_REG_9_ & ~n2615_1;
  assign n2860_1 = ~n2858 & ~n2859;
  assign n2861 = SI_9_ & n2860_1;
  assign n2862 = ~SI_9_ & ~n2860_1;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = n2857 & ~n2863;
  assign n2865_1 = ~n2857 & n2863;
  assign n2866 = ~n2864 & ~n2865_1;
  assign n2867 = ~n2615_1 & ~n2866;
  assign n2868 = ~n2850_1 & ~n2867;
  assign n2869 = ~P1_STATE_REG & ~n2868;
  assign n2870_1 = ~n2848 & ~n2849;
  assign n155 = n2869 | ~n2870_1;
  assign n2872 = P1_IR_REG_10_ & ~n2845_1;
  assign n2873 = ~P1_IR_REG_9_ & ~P1_IR_REG_10_;
  assign n2874 = n2822 & n2873;
  assign n2875_1 = ~n2872 & ~n2874;
  assign n2876 = n2606 & n2875_1;
  assign n2877 = P1_IR_REG_10_ & n2605_1;
  assign n2878 = P2_DATAO_REG_10_ & n2615_1;
  assign n2879 = ~SI_9_ & n2860_1;
  assign n2880_1 = ~n2854 & ~n2879;
  assign n2881 = SI_9_ & ~n2860_1;
  assign n2882 = ~n2880_1 & ~n2881;
  assign n2883 = n2855_1 & ~n2879;
  assign n2884 = ~n2802 & n2883;
  assign n2885_1 = n2882 & ~n2884;
  assign n2886 = P1_DATAO_REG_10_ & n2615_1;
  assign n2887 = P2_DATAO_REG_10_ & ~n2615_1;
  assign n2888 = ~n2886 & ~n2887;
  assign n2889 = SI_10_ & n2888;
  assign n2890_1 = ~SI_10_ & ~n2888;
  assign n2891 = ~n2889 & ~n2890_1;
  assign n2892 = n2885_1 & ~n2891;
  assign n2893 = ~n2885_1 & n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895_1 = ~n2615_1 & ~n2894;
  assign n2896 = ~n2878 & ~n2895_1;
  assign n2897 = ~P1_STATE_REG & ~n2896;
  assign n2898 = ~n2876 & ~n2877;
  assign n160 = n2897 | ~n2898;
  assign n2900_1 = P1_IR_REG_11_ & ~n2874;
  assign n2901 = ~P1_IR_REG_11_ & n2874;
  assign n2902 = ~n2900_1 & ~n2901;
  assign n2903 = n2606 & n2902;
  assign n2904 = P1_IR_REG_11_ & n2605_1;
  assign n2905_1 = P2_DATAO_REG_11_ & n2615_1;
  assign n2906 = ~SI_10_ & n2888;
  assign n2907 = ~n2882 & ~n2906;
  assign n2908 = SI_10_ & ~n2888;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910_1 = n2883 & ~n2906;
  assign n2911 = ~n2802 & n2910_1;
  assign n2912 = n2909 & ~n2911;
  assign n2913 = P1_DATAO_REG_11_ & n2615_1;
  assign n2914 = P2_DATAO_REG_11_ & ~n2615_1;
  assign n2915_1 = ~n2913 & ~n2914;
  assign n2916 = SI_11_ & n2915_1;
  assign n2917 = ~SI_11_ & ~n2915_1;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = n2912 & ~n2918;
  assign n2920_1 = ~n2912 & n2918;
  assign n2921 = ~n2919 & ~n2920_1;
  assign n2922 = ~n2615_1 & ~n2921;
  assign n2923 = ~n2905_1 & ~n2922;
  assign n2924 = ~P1_STATE_REG & ~n2923;
  assign n2925_1 = ~n2903 & ~n2904;
  assign n165 = n2924 | ~n2925_1;
  assign n2927 = P1_IR_REG_12_ & ~n2901;
  assign n2928 = ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign n2929 = ~P1_IR_REG_12_ & n2928;
  assign n2930_1 = ~P1_IR_REG_9_ & n2929;
  assign n2931 = n2822 & n2930_1;
  assign n2932 = ~n2927 & ~n2931;
  assign n2933 = n2606 & n2932;
  assign n2934 = P1_IR_REG_12_ & n2605_1;
  assign n2935_1 = P2_DATAO_REG_12_ & n2615_1;
  assign n2936 = ~SI_11_ & n2915_1;
  assign n2937 = ~n2912 & ~n2936;
  assign n2938 = SI_11_ & ~n2915_1;
  assign n2939 = ~n2937 & ~n2938;
  assign n2940_1 = P1_DATAO_REG_12_ & n2615_1;
  assign n2941 = P2_DATAO_REG_12_ & ~n2615_1;
  assign n2942 = ~n2940_1 & ~n2941;
  assign n2943 = SI_12_ & n2942;
  assign n2944 = ~SI_12_ & ~n2942;
  assign n2945_1 = ~n2943 & ~n2944;
  assign n2946 = n2939 & ~n2945_1;
  assign n2947 = ~n2939 & n2945_1;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n2615_1 & ~n2948;
  assign n2950_1 = ~n2935_1 & ~n2949;
  assign n2951 = ~P1_STATE_REG & ~n2950_1;
  assign n2952 = ~n2933 & ~n2934;
  assign n170 = n2951 | ~n2952;
  assign n2954 = ~P1_IR_REG_13_ & n2931;
  assign n2955_1 = P1_IR_REG_13_ & ~n2931;
  assign n2956 = ~n2954 & ~n2955_1;
  assign n2957 = n2606 & n2956;
  assign n2958 = P1_IR_REG_13_ & n2605_1;
  assign n2959 = P2_DATAO_REG_13_ & n2615_1;
  assign n2960_1 = ~SI_12_ & n2942;
  assign n2961 = n2938 & ~n2960_1;
  assign n2962 = SI_12_ & ~n2942;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = ~n2936 & ~n2960_1;
  assign n2965_1 = ~n2912 & n2964;
  assign n2966 = n2963 & ~n2965_1;
  assign n2967 = P1_DATAO_REG_13_ & n2615_1;
  assign n2968 = P2_DATAO_REG_13_ & ~n2615_1;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970_1 = SI_13_ & n2969;
  assign n2971 = ~SI_13_ & ~n2969;
  assign n2972 = ~n2970_1 & ~n2971;
  assign n2973 = n2966 & ~n2972;
  assign n2974 = ~n2966 & n2972;
  assign n2975_1 = ~n2973 & ~n2974;
  assign n2976 = ~n2615_1 & ~n2975_1;
  assign n2977 = ~n2959 & ~n2976;
  assign n2978 = ~P1_STATE_REG & ~n2977;
  assign n2979 = ~n2957 & ~n2958;
  assign n175 = n2978 | ~n2979;
  assign n2981 = P1_IR_REG_14_ & ~n2954;
  assign n2982 = ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign n2983 = n2931 & n2982;
  assign n2984 = ~n2981 & ~n2983;
  assign n2985_1 = n2606 & n2984;
  assign n2986 = P1_IR_REG_14_ & n2605_1;
  assign n2987 = P2_DATAO_REG_14_ & n2615_1;
  assign n2988 = ~SI_13_ & n2969;
  assign n2989 = ~n2963 & ~n2988;
  assign n2990_1 = SI_13_ & ~n2969;
  assign n2991 = ~n2989 & ~n2990_1;
  assign n2992 = n2964 & ~n2988;
  assign n2993 = ~n2912 & n2992;
  assign n2994 = n2991 & ~n2993;
  assign n2995_1 = P1_DATAO_REG_14_ & n2615_1;
  assign n2996 = P2_DATAO_REG_14_ & ~n2615_1;
  assign n2997 = ~n2995_1 & ~n2996;
  assign n2998 = SI_14_ & n2997;
  assign n2999 = ~SI_14_ & ~n2997;
  assign n3000_1 = ~n2998 & ~n2999;
  assign n3001 = n2994 & ~n3000_1;
  assign n3002 = ~n2994 & n3000_1;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = ~n2615_1 & ~n3003;
  assign n3005_1 = ~n2987 & ~n3004;
  assign n3006 = ~P1_STATE_REG & ~n3005_1;
  assign n3007 = ~n2985_1 & ~n2986;
  assign n180 = n3006 | ~n3007;
  assign n3009 = P1_IR_REG_15_ & ~n2983;
  assign n3010_1 = ~P1_IR_REG_15_ & n2983;
  assign n3011 = ~n3009 & ~n3010_1;
  assign n3012 = n2606 & n3011;
  assign n3013 = P1_IR_REG_15_ & n2605_1;
  assign n3014 = P2_DATAO_REG_15_ & n2615_1;
  assign n3015_1 = ~SI_14_ & n2997;
  assign n3016 = ~n2991 & ~n3015_1;
  assign n3017 = SI_14_ & ~n2997;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = n2992 & ~n3015_1;
  assign n3020_1 = ~n2912 & n3019;
  assign n3021 = n3018 & ~n3020_1;
  assign n3022 = P1_DATAO_REG_15_ & n2615_1;
  assign n3023 = P2_DATAO_REG_15_ & ~n2615_1;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025_1 = SI_15_ & n3024;
  assign n3026 = ~SI_15_ & ~n3024;
  assign n3027 = ~n3025_1 & ~n3026;
  assign n3028 = n3021 & ~n3027;
  assign n3029 = ~n3021 & n3027;
  assign n3030_1 = ~n3028 & ~n3029;
  assign n3031 = ~n2615_1 & ~n3030_1;
  assign n3032 = ~n3014 & ~n3031;
  assign n3033 = ~P1_STATE_REG & ~n3032;
  assign n3034 = ~n3012 & ~n3013;
  assign n185 = n3033 | ~n3034;
  assign n3036 = P1_IR_REG_16_ & ~n3010_1;
  assign n3037 = ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign n3038 = ~P1_IR_REG_8_ & n3037;
  assign n3039 = ~P1_IR_REG_9_ & n3038;
  assign n3040_1 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_;
  assign n3041 = ~P1_IR_REG_4_ & n3040_1;
  assign n3042 = ~P1_IR_REG_5_ & n3041;
  assign n3043 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_;
  assign n3044 = ~P1_IR_REG_1_ & n3043;
  assign n3045_1 = ~P1_IR_REG_0_ & n3044;
  assign n3046 = ~P1_IR_REG_12_ & n2982;
  assign n3047 = ~P1_IR_REG_10_ & n3046;
  assign n3048 = ~P1_IR_REG_11_ & n3047;
  assign n3049 = n3039 & n3042;
  assign n3050_1 = n3045_1 & n3049;
  assign n3051 = n3048 & n3050_1;
  assign n3052 = ~n3036 & ~n3051;
  assign n3053 = n2606 & n3052;
  assign n3054 = P1_IR_REG_16_ & n2605_1;
  assign n3055_1 = P2_DATAO_REG_16_ & n2615_1;
  assign n3056 = ~SI_15_ & n3024;
  assign n3057 = ~n3018 & ~n3056;
  assign n3058 = SI_15_ & ~n3024;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060_1 = n3019 & ~n3056;
  assign n3061 = ~n2912 & n3060_1;
  assign n3062 = n3059 & ~n3061;
  assign n3063 = P1_DATAO_REG_16_ & n2615_1;
  assign n3064 = P2_DATAO_REG_16_ & ~n2615_1;
  assign n3065_1 = ~n3063 & ~n3064;
  assign n3066 = SI_16_ & n3065_1;
  assign n3067 = ~SI_16_ & ~n3065_1;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = n3062 & ~n3068;
  assign n3070_1 = ~n3062 & n3068;
  assign n3071 = ~n3069 & ~n3070_1;
  assign n3072 = ~n2615_1 & ~n3071;
  assign n3073 = ~n3055_1 & ~n3072;
  assign n3074 = ~P1_STATE_REG & ~n3073;
  assign n3075_1 = ~n3053 & ~n3054;
  assign n190 = n3074 | ~n3075_1;
  assign n3077 = ~P1_IR_REG_17_ & n3051;
  assign n3078 = P1_IR_REG_17_ & ~n3051;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080_1 = n2606 & n3079;
  assign n3081 = P1_IR_REG_17_ & n2605_1;
  assign n3082 = P2_DATAO_REG_17_ & n2615_1;
  assign n3083 = SI_16_ & ~n3065_1;
  assign n3084 = ~SI_16_ & n3065_1;
  assign n3085_1 = ~n3062 & ~n3084;
  assign n3086 = ~n3083 & ~n3085_1;
  assign n3087 = P1_DATAO_REG_17_ & n2615_1;
  assign n3088 = P2_DATAO_REG_17_ & ~n2615_1;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090_1 = SI_17_ & n3089;
  assign n3091 = ~SI_17_ & ~n3089;
  assign n3092 = ~n3090_1 & ~n3091;
  assign n3093 = n3086 & ~n3092;
  assign n3094 = ~n3086 & n3092;
  assign n3095_1 = ~n3093 & ~n3094;
  assign n3096 = ~n2615_1 & ~n3095_1;
  assign n3097 = ~n3082 & ~n3096;
  assign n3098 = ~P1_STATE_REG & ~n3097;
  assign n3099 = ~n3080_1 & ~n3081;
  assign n195 = n3098 | ~n3099;
  assign n3101 = P1_IR_REG_18_ & ~n3077;
  assign n3102 = ~P1_IR_REG_4_ & ~P1_IR_REG_5_;
  assign n3103 = ~P1_IR_REG_3_ & n3102;
  assign n3104 = ~P1_IR_REG_0_ & n3103;
  assign n3105_1 = ~P1_IR_REG_2_ & n3104;
  assign n3106 = ~P1_IR_REG_1_ & ~P1_IR_REG_18_;
  assign n3107 = ~P1_IR_REG_17_ & n3106;
  assign n3108 = ~P1_IR_REG_15_ & n3107;
  assign n3109 = ~P1_IR_REG_16_ & n3108;
  assign n3110_1 = n3039 & n3105_1;
  assign n3111 = n3109 & n3110_1;
  assign n3112 = n3048 & n3111;
  assign n3113 = ~n3101 & ~n3112;
  assign n3114 = n2606 & n3113;
  assign n3115_1 = P1_IR_REG_18_ & n2605_1;
  assign n3116 = P2_DATAO_REG_18_ & n2615_1;
  assign n3117 = SI_17_ & ~n3089;
  assign n3118 = ~SI_17_ & n3089;
  assign n3119 = ~n3086 & ~n3118;
  assign n3120_1 = ~n3117 & ~n3119;
  assign n3121 = P1_DATAO_REG_18_ & n2615_1;
  assign n3122 = P2_DATAO_REG_18_ & ~n2615_1;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = SI_18_ & n3123;
  assign n3125_1 = ~SI_18_ & ~n3123;
  assign n3126 = ~n3124 & ~n3125_1;
  assign n3127 = n3120_1 & ~n3126;
  assign n3128 = ~n3120_1 & n3126;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130_1 = ~n2615_1 & ~n3129;
  assign n3131 = ~n3116 & ~n3130_1;
  assign n3132 = ~P1_STATE_REG & ~n3131;
  assign n3133 = ~n3114 & ~n3115_1;
  assign n200 = n3132 | ~n3133;
  assign n3135_1 = P1_IR_REG_19_ & ~n3112;
  assign n3136 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign n3137 = ~P1_IR_REG_7_ & n3136;
  assign n3138 = ~P1_IR_REG_5_ & n3137;
  assign n3139 = ~P1_IR_REG_6_ & n3138;
  assign n3140_1 = ~P1_IR_REG_2_ & n2711;
  assign n3141 = ~P1_IR_REG_1_ & n3140_1;
  assign n3142 = ~P1_IR_REG_0_ & n3141;
  assign n3143 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign n3144 = ~P1_IR_REG_17_ & n3143;
  assign n3145_1 = ~P1_IR_REG_15_ & n3144;
  assign n3146 = ~P1_IR_REG_16_ & n3145_1;
  assign n3147 = n3139 & n3142;
  assign n3148 = n3146 & n3147;
  assign n3149 = n3048 & n3148;
  assign n3150_1 = ~n3135_1 & ~n3149;
  assign n3151 = n2606 & n3150_1;
  assign n3152 = P1_IR_REG_19_ & n2605_1;
  assign n3153 = P2_DATAO_REG_19_ & n2615_1;
  assign n3154 = SI_18_ & ~n3123;
  assign n3155_1 = ~SI_18_ & n3123;
  assign n3156 = ~n3120_1 & ~n3155_1;
  assign n3157 = ~n3154 & ~n3156;
  assign n3158 = P1_DATAO_REG_19_ & n2615_1;
  assign n3159 = P2_DATAO_REG_19_ & ~n2615_1;
  assign n3160_1 = ~n3158 & ~n3159;
  assign n3161 = SI_19_ & n3160_1;
  assign n3162 = ~SI_19_ & ~n3160_1;
  assign n3163 = ~n3161 & ~n3162;
  assign n3164 = n3157 & ~n3163;
  assign n3165_1 = ~n3157 & n3163;
  assign n3166 = ~n3164 & ~n3165_1;
  assign n3167 = ~n2615_1 & ~n3166;
  assign n3168 = ~n3153 & ~n3167;
  assign n3169 = ~P1_STATE_REG & ~n3168;
  assign n3170_1 = ~n3151 & ~n3152;
  assign n205 = n3169 | ~n3170_1;
  assign n3172 = P1_IR_REG_20_ & ~n3149;
  assign n3173 = ~P1_IR_REG_13_ & ~P1_IR_REG_15_;
  assign n3174 = ~P1_IR_REG_14_ & n3173;
  assign n3175_1 = ~P1_IR_REG_10_ & ~P1_IR_REG_12_;
  assign n3176 = ~P1_IR_REG_11_ & n3175_1;
  assign n3177 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_;
  assign n3178 = ~P1_IR_REG_18_ & n3177;
  assign n3179 = ~P1_IR_REG_16_ & n3178;
  assign n3180_1 = ~P1_IR_REG_17_ & n3179;
  assign n3181 = ~P1_IR_REG_0_ & n3140_1;
  assign n3182 = ~P1_IR_REG_20_ & n3181;
  assign n3183 = n3174 & n3176;
  assign n3184 = n3180_1 & n3183;
  assign n3185_1 = n3139 & n3184;
  assign n3186 = n3182 & n3185_1;
  assign n3187 = ~n3172 & ~n3186;
  assign n3188 = n2606 & n3187;
  assign n3189 = P1_IR_REG_20_ & n2605_1;
  assign n3190_1 = P2_DATAO_REG_20_ & n2615_1;
  assign n3191 = SI_19_ & ~n3160_1;
  assign n3192 = ~SI_19_ & n3160_1;
  assign n3193 = ~n3157 & ~n3192;
  assign n3194 = ~n3191 & ~n3193;
  assign n3195_1 = P1_DATAO_REG_20_ & n2615_1;
  assign n3196 = P2_DATAO_REG_20_ & ~n2615_1;
  assign n3197 = ~n3195_1 & ~n3196;
  assign n3198 = SI_20_ & n3197;
  assign n3199 = ~SI_20_ & ~n3197;
  assign n3200_1 = ~n3198 & ~n3199;
  assign n3201 = n3194 & ~n3200_1;
  assign n3202 = ~n3194 & n3200_1;
  assign n3203 = ~n3201 & ~n3202;
  assign n3204 = ~n2615_1 & ~n3203;
  assign n3205_1 = ~n3190_1 & ~n3204;
  assign n3206 = ~P1_STATE_REG & ~n3205_1;
  assign n3207 = ~n3188 & ~n3189;
  assign n210 = n3206 | ~n3207;
  assign n3209 = ~P1_IR_REG_21_ & n3186;
  assign n3210_1 = P1_IR_REG_21_ & ~n3186;
  assign n3211 = ~n3209 & ~n3210_1;
  assign n3212 = n2606 & n3211;
  assign n3213 = P1_IR_REG_21_ & n2605_1;
  assign n3214 = P2_DATAO_REG_21_ & n2615_1;
  assign n3215_1 = SI_20_ & ~n3197;
  assign n3216 = ~SI_20_ & n3197;
  assign n3217 = ~n3194 & ~n3216;
  assign n3218 = ~n3215_1 & ~n3217;
  assign n3219 = P1_DATAO_REG_21_ & n2615_1;
  assign n3220_1 = P2_DATAO_REG_21_ & ~n2615_1;
  assign n3221 = ~n3219 & ~n3220_1;
  assign n3222 = SI_21_ & n3221;
  assign n3223 = ~SI_21_ & ~n3221;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225_1 = n3218 & ~n3224;
  assign n3226 = ~n3218 & n3224;
  assign n3227 = ~n3225_1 & ~n3226;
  assign n3228 = ~n2615_1 & ~n3227;
  assign n3229 = ~n3214 & ~n3228;
  assign n3230_1 = ~P1_STATE_REG & ~n3229;
  assign n3231 = ~n3212 & ~n3213;
  assign n215 = n3230_1 | ~n3231;
  assign n3233 = ~P1_IR_REG_2_ & ~P1_IR_REG_4_;
  assign n3234 = ~P1_IR_REG_3_ & n3233;
  assign n3235_1 = ~P1_IR_REG_0_ & ~P1_IR_REG_21_;
  assign n3236 = ~P1_IR_REG_20_ & n3235_1;
  assign n3237 = n3234 & n3236;
  assign n3238 = n3139 & n3237;
  assign n3239 = n3180_1 & n3238;
  assign n3240_1 = n3183 & n3239;
  assign n3241 = P1_IR_REG_22_ & ~n3240_1;
  assign n3242 = ~P1_IR_REG_19_ & ~P1_IR_REG_20_;
  assign n3243 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign n3244 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign n3245_1 = n3242 & n3243;
  assign n3246 = n3244 & n3245_1;
  assign n3247 = n3051 & n3246;
  assign n3248 = ~n3241 & ~n3247;
  assign n3249 = n2606 & n3248;
  assign n3250_1 = P1_IR_REG_22_ & n2605_1;
  assign n3251 = P2_DATAO_REG_22_ & n2615_1;
  assign n3252 = SI_21_ & ~n3221;
  assign n3253 = ~SI_21_ & n3221;
  assign n3254 = ~n3218 & ~n3253;
  assign n3255_1 = ~n3252 & ~n3254;
  assign n3256 = P1_DATAO_REG_22_ & n2615_1;
  assign n3257 = P2_DATAO_REG_22_ & ~n2615_1;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = SI_22_ & n3258;
  assign n3260_1 = ~SI_22_ & ~n3258;
  assign n3261 = ~n3259 & ~n3260_1;
  assign n3262 = n3255_1 & ~n3261;
  assign n3263 = ~n3255_1 & n3261;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265_1 = ~n2615_1 & ~n3264;
  assign n3266 = ~n3251 & ~n3265_1;
  assign n3267 = ~P1_STATE_REG & ~n3266;
  assign n3268 = ~n3249 & ~n3250_1;
  assign n220 = n3267 | ~n3268;
  assign n3270_1 = P1_IR_REG_23_ & ~n3247;
  assign n3271 = ~P1_IR_REG_7_ & ~P1_IR_REG_9_;
  assign n3272 = ~P1_IR_REG_8_ & n3271;
  assign n3273 = ~P1_IR_REG_4_ & ~P1_IR_REG_6_;
  assign n3274 = ~P1_IR_REG_5_ & n3273;
  assign n3275_1 = ~P1_IR_REG_3_ & ~P1_IR_REG_23_;
  assign n3276 = ~P1_IR_REG_2_ & n3275_1;
  assign n3277 = ~P1_IR_REG_20_ & ~P1_IR_REG_22_;
  assign n3278 = ~P1_IR_REG_21_ & n3277;
  assign n3279 = n3272 & n3274;
  assign n3280_1 = n3276 & n3279;
  assign n3281 = n3278 & n3280_1;
  assign n3282 = ~P1_IR_REG_0_ & ~P1_IR_REG_19_;
  assign n3283 = ~P1_IR_REG_1_ & n3282;
  assign n3284 = ~P1_IR_REG_16_ & ~P1_IR_REG_18_;
  assign n3285_1 = ~P1_IR_REG_17_ & n3284;
  assign n3286 = n3283 & n3285_1;
  assign n3287 = n3174 & n3286;
  assign n3288 = n3176 & n3287;
  assign n3289 = n3281 & n3288;
  assign n3290_1 = ~n3270_1 & ~n3289;
  assign n3291 = n2606 & n3290_1;
  assign n3292 = P1_IR_REG_23_ & n2605_1;
  assign n3293 = P2_DATAO_REG_23_ & n2615_1;
  assign n3294 = SI_22_ & ~n3258;
  assign n3295_1 = ~SI_22_ & n3258;
  assign n3296 = ~n3255_1 & ~n3295_1;
  assign n3297 = ~n3294 & ~n3296;
  assign n3298 = P1_DATAO_REG_23_ & n2615_1;
  assign n3299 = P2_DATAO_REG_23_ & ~n2615_1;
  assign n3300_1 = ~n3298 & ~n3299;
  assign n3301 = SI_23_ & n3300_1;
  assign n3302 = ~SI_23_ & ~n3300_1;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = n3297 & ~n3303;
  assign n3305_1 = ~n3297 & n3303;
  assign n3306 = ~n3304 & ~n3305_1;
  assign n3307 = ~n2615_1 & ~n3306;
  assign n3308 = ~n3293 & ~n3307;
  assign n3309 = ~P1_STATE_REG & ~n3308;
  assign n3310_1 = ~n3291 & ~n3292;
  assign n225 = n3309 | ~n3310_1;
  assign n3312 = P1_IR_REG_24_ & ~n3289;
  assign n3313 = ~P1_IR_REG_3_ & ~P1_IR_REG_24_;
  assign n3314 = ~P1_IR_REG_2_ & n3313;
  assign n3315_1 = ~P1_IR_REG_21_ & ~P1_IR_REG_23_;
  assign n3316 = ~P1_IR_REG_22_ & n3315_1;
  assign n3317 = n3279 & n3314;
  assign n3318 = n3316 & n3317;
  assign n3319 = ~P1_IR_REG_1_ & ~P1_IR_REG_20_;
  assign n3320_1 = ~P1_IR_REG_0_ & n3319;
  assign n3321 = ~P1_IR_REG_17_ & ~P1_IR_REG_19_;
  assign n3322 = ~P1_IR_REG_18_ & n3321;
  assign n3323 = ~P1_IR_REG_14_ & ~P1_IR_REG_16_;
  assign n3324 = ~P1_IR_REG_15_ & n3323;
  assign n3325_1 = ~P1_IR_REG_13_ & n2929;
  assign n3326 = n3320_1 & n3322;
  assign n3327 = n3324 & n3326;
  assign n3328 = n3325_1 & n3327;
  assign n3329 = n3318 & n3328;
  assign n3330_1 = ~n3312 & ~n3329;
  assign n3331 = n2606 & n3330_1;
  assign n3332 = P1_IR_REG_24_ & n2605_1;
  assign n3333 = P2_DATAO_REG_24_ & n2615_1;
  assign n3334 = SI_23_ & ~n3300_1;
  assign n3335_1 = ~SI_23_ & n3300_1;
  assign n3336 = ~n3297 & ~n3335_1;
  assign n3337 = ~n3334 & ~n3336;
  assign n3338 = P1_DATAO_REG_24_ & n2615_1;
  assign n3339 = P2_DATAO_REG_24_ & ~n2615_1;
  assign n3340_1 = ~n3338 & ~n3339;
  assign n3341 = SI_24_ & n3340_1;
  assign n3342 = ~SI_24_ & ~n3340_1;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = n3337 & ~n3343;
  assign n3345_1 = ~n3337 & n3343;
  assign n3346 = ~n3344 & ~n3345_1;
  assign n3347 = ~n2615_1 & ~n3346;
  assign n3348 = ~n3333 & ~n3347;
  assign n3349 = ~P1_STATE_REG & ~n3348;
  assign n3350_1 = ~n3331 & ~n3332;
  assign n230 = n3349 | ~n3350_1;
  assign n3352 = ~P1_IR_REG_25_ & n3329;
  assign n3353 = P1_IR_REG_25_ & ~n3329;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355_1 = n2606 & n3354;
  assign n3356 = P1_IR_REG_25_ & n2605_1;
  assign n3357 = P2_DATAO_REG_25_ & n2615_1;
  assign n3358 = SI_24_ & ~n3340_1;
  assign n3359 = ~SI_24_ & n3340_1;
  assign n3360_1 = ~n3337 & ~n3359;
  assign n3361 = ~n3358 & ~n3360_1;
  assign n3362 = P1_DATAO_REG_25_ & n2615_1;
  assign n3363 = P2_DATAO_REG_25_ & ~n2615_1;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365_1 = SI_25_ & n3364;
  assign n3366 = ~SI_25_ & ~n3364;
  assign n3367 = ~n3365_1 & ~n3366;
  assign n3368 = n3361 & ~n3367;
  assign n3369 = ~n3361 & n3367;
  assign n3370_1 = ~n3368 & ~n3369;
  assign n3371 = ~n2615_1 & ~n3370_1;
  assign n3372 = ~n3357 & ~n3371;
  assign n3373 = ~P1_STATE_REG & ~n3372;
  assign n3374 = ~n3355_1 & ~n3356;
  assign n235 = n3373 | ~n3374;
  assign n3376 = ~P1_IR_REG_3_ & ~P1_IR_REG_25_;
  assign n3377 = ~P1_IR_REG_2_ & n3376;
  assign n3378 = ~P1_IR_REG_23_ & n3244;
  assign n3379 = ~P1_IR_REG_24_ & n3378;
  assign n3380_1 = n3279 & n3377;
  assign n3381 = n3379 & n3380_1;
  assign n3382 = n3328 & n3381;
  assign n3383 = P1_IR_REG_26_ & ~n3382;
  assign n3384 = ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign n3385_1 = ~P1_IR_REG_2_ & n3384;
  assign n3386 = ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign n3387 = ~P1_IR_REG_24_ & n3386;
  assign n3388 = ~P1_IR_REG_25_ & n3387;
  assign n3389 = n3279 & n3385_1;
  assign n3390_1 = n3388 & n3389;
  assign n3391 = ~P1_IR_REG_19_ & n3243;
  assign n3392 = ~P1_IR_REG_1_ & n3391;
  assign n3393 = n3236 & n3392;
  assign n3394 = n3324 & n3393;
  assign n3395_1 = n3325_1 & n3394;
  assign n3396 = n3390_1 & n3395_1;
  assign n3397 = ~n3383 & ~n3396;
  assign n3398 = n2606 & n3397;
  assign n3399 = P1_IR_REG_26_ & n2605_1;
  assign n3400_1 = P2_DATAO_REG_26_ & n2615_1;
  assign n3401 = SI_25_ & ~n3364;
  assign n3402 = ~SI_25_ & n3364;
  assign n3403 = ~n3361 & ~n3402;
  assign n3404 = ~n3401 & ~n3403;
  assign n3405_1 = P1_DATAO_REG_26_ & n2615_1;
  assign n3406 = P2_DATAO_REG_26_ & ~n2615_1;
  assign n3407 = ~n3405_1 & ~n3406;
  assign n3408 = SI_26_ & n3407;
  assign n3409 = ~SI_26_ & ~n3407;
  assign n3410_1 = ~n3408 & ~n3409;
  assign n3411 = n3404 & ~n3410_1;
  assign n3412 = ~n3404 & n3410_1;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n2615_1 & ~n3413;
  assign n3415_1 = ~n3400_1 & ~n3414;
  assign n3416 = ~P1_STATE_REG & ~n3415_1;
  assign n3417 = ~n3398 & ~n3399;
  assign n240 = n3416 | ~n3417;
  assign n3419 = ~P1_IR_REG_27_ & ~n3396;
  assign n3420_1 = P1_IR_REG_27_ & n3396;
  assign n3421 = ~n3419 & ~n3420_1;
  assign n3422 = n2606 & ~n3421;
  assign n3423 = P1_IR_REG_27_ & n2605_1;
  assign n3424 = P2_DATAO_REG_27_ & n2615_1;
  assign n3425_1 = SI_26_ & ~n3407;
  assign n3426 = ~SI_26_ & n3407;
  assign n3427 = ~n3404 & ~n3426;
  assign n3428 = ~n3425_1 & ~n3427;
  assign n3429 = P1_DATAO_REG_27_ & n2615_1;
  assign n3430_1 = P2_DATAO_REG_27_ & ~n2615_1;
  assign n3431 = ~n3429 & ~n3430_1;
  assign n3432 = SI_27_ & n3431;
  assign n3433 = ~SI_27_ & ~n3431;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435_1 = n3428 & ~n3434;
  assign n3436 = ~n3428 & n3434;
  assign n3437 = ~n3435_1 & ~n3436;
  assign n3438 = ~n2615_1 & ~n3437;
  assign n3439 = ~n3424 & ~n3438;
  assign n3440_1 = ~P1_STATE_REG & ~n3439;
  assign n3441 = ~n3422 & ~n3423;
  assign n245 = n3440_1 | ~n3441;
  assign n3443 = ~P1_IR_REG_2_ & ~P1_IR_REG_26_;
  assign n3444 = ~P1_IR_REG_27_ & n3443;
  assign n3445_1 = n2820_1 & n3272;
  assign n3446 = n3444 & n3445_1;
  assign n3447 = n3388 & n3446;
  assign n3448 = n3395_1 & n3447;
  assign n3449 = P1_IR_REG_28_ & ~n3448;
  assign n3450_1 = ~P1_IR_REG_2_ & ~P1_IR_REG_27_;
  assign n3451 = ~P1_IR_REG_28_ & n3450_1;
  assign n3452 = ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign n3453 = ~P1_IR_REG_25_ & n3452;
  assign n3454 = ~P1_IR_REG_26_ & n3453;
  assign n3455_1 = n3445_1 & n3451;
  assign n3456 = n3454 & n3455_1;
  assign n3457 = ~P1_IR_REG_1_ & n3143;
  assign n3458 = ~P1_IR_REG_0_ & n3457;
  assign n3459 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign n3460_1 = ~P1_IR_REG_16_ & n3459;
  assign n3461 = ~P1_IR_REG_17_ & n3460_1;
  assign n3462 = n3278 & n3458;
  assign n3463 = n3461 & n3462;
  assign n3464 = n3325_1 & n3463;
  assign n3465_1 = n3456 & n3464;
  assign n3466 = ~n3449 & ~n3465_1;
  assign n3467 = n2606 & n3466;
  assign n3468 = P1_IR_REG_28_ & n2605_1;
  assign n3469 = P2_DATAO_REG_28_ & n2615_1;
  assign n3470_1 = SI_27_ & ~n3431;
  assign n3471 = ~SI_27_ & n3431;
  assign n3472 = ~n3428 & ~n3471;
  assign n3473 = ~n3470_1 & ~n3472;
  assign n3474 = P1_DATAO_REG_28_ & n2615_1;
  assign n3475_1 = P2_DATAO_REG_28_ & ~n2615_1;
  assign n3476 = ~n3474 & ~n3475_1;
  assign n3477 = SI_28_ & n3476;
  assign n3478 = ~SI_28_ & ~n3476;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480_1 = n3473 & ~n3479;
  assign n3481 = ~n3473 & n3479;
  assign n3482 = ~n3480_1 & ~n3481;
  assign n3483 = ~n2615_1 & ~n3482;
  assign n3484 = ~n3469 & ~n3483;
  assign n3485_1 = ~P1_STATE_REG & ~n3484;
  assign n3486 = ~n3467 & ~n3468;
  assign n250 = n3485_1 | ~n3486;
  assign n3488 = P1_IR_REG_29_ & ~n3465_1;
  assign n3489 = ~P1_IR_REG_27_ & ~P1_IR_REG_28_;
  assign n3490_1 = ~P1_IR_REG_29_ & n3489;
  assign n3491 = ~P1_IR_REG_2_ & n3490_1;
  assign n3492 = n3445_1 & n3491;
  assign n3493 = n3454 & n3492;
  assign n3494 = n3464 & n3493;
  assign n3495_1 = ~n3488 & ~n3494;
  assign n3496 = n2606 & n3495_1;
  assign n3497 = P1_IR_REG_29_ & n2605_1;
  assign n3498 = P2_DATAO_REG_29_ & n2615_1;
  assign n3499 = SI_28_ & ~n3476;
  assign n3500_1 = ~SI_28_ & n3476;
  assign n3501 = ~n3473 & ~n3500_1;
  assign n3502 = ~n3499 & ~n3501;
  assign n3503 = P1_DATAO_REG_29_ & n2615_1;
  assign n3504 = P2_DATAO_REG_29_ & ~n2615_1;
  assign n3505_1 = ~n3503 & ~n3504;
  assign n3506 = SI_29_ & n3505_1;
  assign n3507 = ~SI_29_ & ~n3505_1;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = n3502 & ~n3508;
  assign n3510_1 = ~n3502 & n3508;
  assign n3511 = ~n3509 & ~n3510_1;
  assign n3512 = ~n2615_1 & ~n3511;
  assign n3513 = ~n3498 & ~n3512;
  assign n3514 = ~P1_STATE_REG & ~n3513;
  assign n3515_1 = ~n3496 & ~n3497;
  assign n255 = n3514 | ~n3515_1;
  assign n3517 = ~P1_IR_REG_30_ & n3494;
  assign n3518 = P1_IR_REG_30_ & ~n3494;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520_1 = n2606 & n3519;
  assign n3521 = P1_IR_REG_30_ & n2605_1;
  assign n3522 = P2_DATAO_REG_30_ & n2615_1;
  assign n3523 = SI_29_ & ~n3505_1;
  assign n3524 = ~SI_29_ & n3505_1;
  assign n3525_1 = ~n3502 & ~n3524;
  assign n3526 = ~n3523 & ~n3525_1;
  assign n3527 = P1_DATAO_REG_30_ & n2615_1;
  assign n3528 = P2_DATAO_REG_30_ & ~n2615_1;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530_1 = SI_30_ & n3529;
  assign n3531 = ~SI_30_ & ~n3529;
  assign n3532 = ~n3530_1 & ~n3531;
  assign n3533 = n3526 & ~n3532;
  assign n3534 = ~n3526 & n3532;
  assign n3535_1 = ~n3533 & ~n3534;
  assign n3536 = ~n2615_1 & ~n3535_1;
  assign n3537 = ~n3522 & ~n3536;
  assign n3538 = ~P1_STATE_REG & ~n3537;
  assign n3539 = ~n3520_1 & ~n3521;
  assign n260 = n3538 | ~n3539;
  assign n3541 = P1_IR_REG_31_ & n3517;
  assign n3542 = ~P1_IR_REG_31_ & ~n3517;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = n2606 & ~n3543;
  assign n3545_1 = P1_IR_REG_31_ & n2605_1;
  assign n3546 = P2_DATAO_REG_31_ & n2615_1;
  assign n3547 = P1_DATAO_REG_31_ & n2615_1;
  assign n3548 = P2_DATAO_REG_31_ & ~n2615_1;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550_1 = SI_31_ & n3549;
  assign n3551 = ~SI_31_ & ~n3549;
  assign n3552 = ~n3550_1 & ~n3551;
  assign n3553 = SI_30_ & ~n3529;
  assign n3554 = n3552 & ~n3553;
  assign n3555_1 = ~n3523 & n3554;
  assign n3556 = ~n3525_1 & n3555_1;
  assign n3557 = SI_30_ & ~n3552;
  assign n3558 = ~n3529 & n3557;
  assign n3559 = ~SI_30_ & n3552;
  assign n3560_1 = n3529 & n3559;
  assign n3561 = ~n3558 & ~n3560_1;
  assign n3562 = ~n3556 & n3561;
  assign n3563 = ~SI_30_ & n3529;
  assign n3564 = ~n3552 & ~n3563;
  assign n3565_1 = ~n3526 & n3564;
  assign n3566 = n3562 & ~n3565_1;
  assign n3567 = ~n2615_1 & n3566;
  assign n3568 = ~n3546 & ~n3567;
  assign n3569 = ~P1_STATE_REG & ~n3568;
  assign n3570_1 = ~n3544 & ~n3545_1;
  assign n265 = n3569 | ~n3570_1;
  assign n3572 = P1_IR_REG_31_ & n3290_1;
  assign n3573 = P1_IR_REG_23_ & ~P1_IR_REG_31_;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575_1 = P1_STATE_REG & n3574;
  assign n3576 = P1_IR_REG_31_ & n3330_1;
  assign n3577 = P1_IR_REG_24_ & ~P1_IR_REG_31_;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = P1_IR_REG_31_ & n3397;
  assign n3580_1 = P1_IR_REG_26_ & ~P1_IR_REG_31_;
  assign n3581 = ~n3579 & ~n3580_1;
  assign n3582 = P1_IR_REG_31_ & n3354;
  assign n3583 = P1_IR_REG_25_ & ~P1_IR_REG_31_;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585_1 = ~n3578 & ~n3581;
  assign n3586 = ~n3584 & n3585_1;
  assign n3587 = n3575_1 & ~n3586;
  assign n3588 = ~n3581 & n3584;
  assign n3589 = n3578 & n3588;
  assign n3590_1 = P1_B_REG & n3589;
  assign n3591 = ~P1_B_REG & ~n3578;
  assign n3592 = ~n3590_1 & ~n3591;
  assign n3593 = ~n3581 & n3592;
  assign n3594 = n3587 & ~n3593;
  assign n3595_1 = n3578 & ~n3588;
  assign n3596 = n3594 & ~n3595_1;
  assign n3597 = P1_D_REG_0_ & ~n3594;
  assign n270 = n3596 | n3597;
  assign n3599 = n3584 & ~n3588;
  assign n3600_1 = n3594 & ~n3599;
  assign n3601 = P1_D_REG_1_ & ~n3594;
  assign n275 = n3600_1 | n3601;
  assign n280 = P1_D_REG_2_ & ~n3594;
  assign n285 = P1_D_REG_3_ & ~n3594;
  assign n290 = P1_D_REG_4_ & ~n3594;
  assign n295 = P1_D_REG_5_ & ~n3594;
  assign n300 = P1_D_REG_6_ & ~n3594;
  assign n305 = P1_D_REG_7_ & ~n3594;
  assign n310 = P1_D_REG_8_ & ~n3594;
  assign n315 = P1_D_REG_9_ & ~n3594;
  assign n320 = P1_D_REG_10_ & ~n3594;
  assign n325 = P1_D_REG_11_ & ~n3594;
  assign n330 = P1_D_REG_12_ & ~n3594;
  assign n335 = P1_D_REG_13_ & ~n3594;
  assign n340 = P1_D_REG_14_ & ~n3594;
  assign n345 = P1_D_REG_15_ & ~n3594;
  assign n350 = P1_D_REG_16_ & ~n3594;
  assign n355 = P1_D_REG_17_ & ~n3594;
  assign n360 = P1_D_REG_18_ & ~n3594;
  assign n365 = P1_D_REG_19_ & ~n3594;
  assign n370 = P1_D_REG_20_ & ~n3594;
  assign n375 = P1_D_REG_21_ & ~n3594;
  assign n380 = P1_D_REG_22_ & ~n3594;
  assign n385 = P1_D_REG_23_ & ~n3594;
  assign n390 = P1_D_REG_24_ & ~n3594;
  assign n395 = P1_D_REG_25_ & ~n3594;
  assign n400 = P1_D_REG_26_ & ~n3594;
  assign n405 = P1_D_REG_27_ & ~n3594;
  assign n410 = P1_D_REG_28_ & ~n3594;
  assign n415 = P1_D_REG_29_ & ~n3594;
  assign n420 = P1_D_REG_30_ & ~n3594;
  assign n425 = P1_D_REG_31_ & ~n3594;
  assign n3633 = P1_D_REG_0_ & n3593;
  assign n3634 = n3578 & n3581;
  assign n3635_1 = ~n3593 & ~n3634;
  assign n3636 = ~n3633 & ~n3635_1;
  assign n3637 = n3587 & n3636;
  assign n3638 = ~n3593 & ~n3599;
  assign n3639 = P1_D_REG_1_ & n3593;
  assign n3640_1 = ~n3638 & ~n3639;
  assign n3641 = P1_IR_REG_31_ & n3248;
  assign n3642 = P1_IR_REG_22_ & ~P1_IR_REG_31_;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = P1_IR_REG_31_ & n3211;
  assign n3645_1 = P1_IR_REG_21_ & ~P1_IR_REG_31_;
  assign n3646 = ~n3644 & ~n3645_1;
  assign n3647 = P1_IR_REG_31_ & n3187;
  assign n3648 = P1_IR_REG_20_ & ~P1_IR_REG_31_;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650_1 = n3646 & n3649;
  assign n3651 = n3643 & ~n3650_1;
  assign n3652 = ~n3643 & n3646;
  assign n3653 = P1_IR_REG_31_ & n3150_1;
  assign n3654 = P1_IR_REG_19_ & ~P1_IR_REG_31_;
  assign n3655_1 = ~n3653 & ~n3654;
  assign n3656 = n3649 & n3655_1;
  assign n3657 = ~n3651 & ~n3652;
  assign n3658 = ~n3656 & n3657;
  assign n3659 = n3640_1 & ~n3658;
  assign n3660_1 = P1_D_REG_8_ & n3593;
  assign n3661 = P1_D_REG_7_ & n3593;
  assign n3662 = P1_D_REG_9_ & n3593;
  assign n3663 = ~n3660_1 & ~n3661;
  assign n3664 = ~n3662 & n3663;
  assign n3665_1 = P1_D_REG_6_ & n3593;
  assign n3666 = P1_D_REG_5_ & n3593;
  assign n3667 = P1_D_REG_4_ & n3593;
  assign n3668 = P1_D_REG_3_ & n3593;
  assign n3669 = ~n3665_1 & ~n3666;
  assign n3670_1 = ~n3667 & n3669;
  assign n3671 = ~n3668 & n3670_1;
  assign n3672 = P1_D_REG_31_ & n3593;
  assign n3673 = P1_D_REG_30_ & n3593;
  assign n3674 = P1_D_REG_2_ & n3593;
  assign n3675_1 = P1_D_REG_29_ & n3593;
  assign n3676 = ~n3672 & ~n3673;
  assign n3677 = ~n3674 & n3676;
  assign n3678 = ~n3675_1 & n3677;
  assign n3679 = P1_D_REG_28_ & n3593;
  assign n3680_1 = P1_D_REG_27_ & n3593;
  assign n3681 = P1_D_REG_26_ & n3593;
  assign n3682 = P1_D_REG_25_ & n3593;
  assign n3683 = ~n3679 & ~n3680_1;
  assign n3684 = ~n3681 & n3683;
  assign n3685_1 = ~n3682 & n3684;
  assign n3686 = n3664 & n3671;
  assign n3687 = n3678 & n3686;
  assign n3688 = n3685_1 & n3687;
  assign n3689 = P1_D_REG_23_ & n3593;
  assign n3690_1 = P1_D_REG_22_ & n3593;
  assign n3691 = P1_D_REG_24_ & n3593;
  assign n3692 = ~n3689 & ~n3690_1;
  assign n3693 = ~n3691 & n3692;
  assign n3694 = P1_D_REG_21_ & n3593;
  assign n3695_1 = P1_D_REG_20_ & n3593;
  assign n3696 = P1_D_REG_19_ & n3593;
  assign n3697 = P1_D_REG_18_ & n3593;
  assign n3698 = ~n3694 & ~n3695_1;
  assign n3699 = ~n3696 & n3698;
  assign n3700_1 = ~n3697 & n3699;
  assign n3701 = P1_D_REG_17_ & n3593;
  assign n3702 = P1_D_REG_16_ & n3593;
  assign n3703 = P1_D_REG_15_ & n3593;
  assign n3704 = P1_D_REG_14_ & n3593;
  assign n3705_1 = ~n3701 & ~n3702;
  assign n3706 = ~n3703 & n3705_1;
  assign n3707 = ~n3704 & n3706;
  assign n3708 = P1_D_REG_13_ & n3593;
  assign n3709 = P1_D_REG_12_ & n3593;
  assign n3710_1 = P1_D_REG_11_ & n3593;
  assign n3711 = P1_D_REG_10_ & n3593;
  assign n3712 = ~n3708 & ~n3709;
  assign n3713 = ~n3710_1 & n3712;
  assign n3714 = ~n3711 & n3713;
  assign n3715_1 = n3693 & n3700_1;
  assign n3716 = n3707 & n3715_1;
  assign n3717 = n3714 & n3716;
  assign n3718 = n3688 & n3717;
  assign n3719 = n3659 & n3718;
  assign n3720_1 = n3637 & n3719;
  assign n3721 = P1_IR_REG_31_ & ~n3421;
  assign n3722 = P1_IR_REG_27_ & ~P1_IR_REG_31_;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = P1_IR_REG_31_ & n3466;
  assign n3725_1 = P1_IR_REG_28_ & ~P1_IR_REG_31_;
  assign n3726 = ~n3724 & ~n3725_1;
  assign n3727 = n3723 & n3726;
  assign n3728 = P1_IR_REG_0_ & P1_IR_REG_31_;
  assign n3729 = P1_IR_REG_0_ & ~P1_IR_REG_31_;
  assign n3730_1 = ~n3728 & ~n3729;
  assign n3731 = n3727 & ~n3730_1;
  assign n3732 = ~n2624 & ~n3727;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = n3646 & ~n3655_1;
  assign n3735_1 = n3643 & n3734;
  assign n3736 = n3646 & n3655_1;
  assign n3737 = n3643 & n3736;
  assign n3738 = ~n3649 & n3737;
  assign n3739 = ~n3735_1 & ~n3738;
  assign n3740_1 = ~n3733 & ~n3739;
  assign n3741 = ~n3643 & ~n3646;
  assign n3742 = n3726 & n3741;
  assign n3743 = P1_IR_REG_31_ & n3519;
  assign n3744 = P1_IR_REG_30_ & ~P1_IR_REG_31_;
  assign n3745_1 = ~n3743 & ~n3744;
  assign n3746 = P1_IR_REG_31_ & n3495_1;
  assign n3747 = P1_IR_REG_29_ & ~P1_IR_REG_31_;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = ~n3745_1 & ~n3748;
  assign n3750_1 = P1_REG3_REG_1_ & n3749;
  assign n3751 = n3745_1 & n3748;
  assign n3752 = P1_REG0_REG_1_ & n3751;
  assign n3753 = n3745_1 & ~n3748;
  assign n3754 = P1_REG1_REG_1_ & n3753;
  assign n3755_1 = ~n3745_1 & n3748;
  assign n3756 = P1_REG2_REG_1_ & n3755_1;
  assign n3757 = ~n3750_1 & ~n3752;
  assign n3758 = ~n3754 & n3757;
  assign n3759 = ~n3756 & n3758;
  assign n3760_1 = n3742 & ~n3759;
  assign n3761 = P1_REG3_REG_0_ & n3749;
  assign n3762 = P1_REG2_REG_0_ & n3755_1;
  assign n3763 = P1_REG1_REG_0_ & n3753;
  assign n3764 = P1_REG0_REG_0_ & n3751;
  assign n3765_1 = ~n3761 & ~n3762;
  assign n3766 = ~n3763 & n3765_1;
  assign n3767 = ~n3764 & n3766;
  assign n3768 = ~n3733 & n3767;
  assign n3769 = n3733 & ~n3767;
  assign n3770_1 = ~n3768 & ~n3769;
  assign n3771 = n3649 & ~n3655_1;
  assign n3772 = n3643 & n3771;
  assign n3773 = ~n3770_1 & n3772;
  assign n3774 = n3643 & n3649;
  assign n3775_1 = n3646 & n3774;
  assign n3776 = ~n3733 & n3775_1;
  assign n3777 = ~n3773 & ~n3776;
  assign n3778 = ~n3643 & n3736;
  assign n3779 = n3649 & n3778;
  assign n3780_1 = ~n3770_1 & n3779;
  assign n3781 = ~n3649 & n3655_1;
  assign n3782 = ~n3646 & n3781;
  assign n3783 = ~n3770_1 & n3782;
  assign n3784 = ~n3646 & n3656;
  assign n3785 = n3643 & n3784;
  assign n3786 = ~n3770_1 & n3785;
  assign n3787 = ~n3649 & ~n3655_1;
  assign n3788 = ~n3646 & n3787;
  assign n3789 = ~n3770_1 & n3788;
  assign n3790 = ~n3643 & n3781;
  assign n3791 = ~n3770_1 & n3790;
  assign n3792 = ~n3789 & ~n3791;
  assign n3793 = ~n3643 & n3787;
  assign n3794 = ~n3770_1 & n3793;
  assign n3795 = ~n3643 & n3771;
  assign n3796 = ~n3770_1 & n3795;
  assign n3797 = ~n3794 & ~n3796;
  assign n3798 = ~n3780_1 & ~n3783;
  assign n3799 = ~n3786 & n3798;
  assign n3800 = n3792 & n3799;
  assign n3801 = n3797 & n3800;
  assign n3802 = ~n3740_1 & ~n3760_1;
  assign n3803 = n3777 & n3802;
  assign n3804 = n3801 & n3803;
  assign n3805 = n3720_1 & ~n3804;
  assign n3806 = P1_REG0_REG_0_ & ~n3720_1;
  assign n430 = n3805 | n3806;
  assign n3808 = P1_IR_REG_31_ & ~n2630_1;
  assign n3809 = P1_IR_REG_1_ & ~P1_IR_REG_31_;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = n3727 & ~n3810;
  assign n3812 = ~n2650_1 & ~n3727;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = ~n3733 & n3813;
  assign n3815 = n3733 & ~n3813;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = n3775_1 & ~n3816;
  assign n3818 = P1_REG3_REG_2_ & n3749;
  assign n3819 = P1_REG0_REG_2_ & n3751;
  assign n3820 = P1_REG1_REG_2_ & n3753;
  assign n3821 = P1_REG2_REG_2_ & n3755_1;
  assign n3822 = ~n3818 & ~n3819;
  assign n3823 = ~n3820 & n3822;
  assign n3824 = ~n3821 & n3823;
  assign n3825 = n3742 & ~n3824;
  assign n3826 = ~n3739 & ~n3813;
  assign n3827 = ~n3759 & ~n3813;
  assign n3828 = n3759 & n3813;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~n3733 & ~n3767;
  assign n3831 = n3829 & ~n3830;
  assign n3832 = ~n3829 & n3830;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = n3772 & ~n3833;
  assign n3835 = ~n3817 & ~n3825;
  assign n3836 = ~n3826 & n3835;
  assign n3837 = ~n3834 & n3836;
  assign n3838 = ~n3759 & n3813;
  assign n3839 = n3759 & ~n3813;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = ~n3768 & ~n3840;
  assign n3842 = n3768 & n3840;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = n3795 & ~n3843;
  assign n3845 = ~n3726 & n3741;
  assign n3846 = ~n3767 & n3845;
  assign n3847 = n3790 & ~n3833;
  assign n3848 = n3793 & ~n3843;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n3785 & ~n3833;
  assign n3851 = n3779 & ~n3833;
  assign n3852 = n3782 & ~n3843;
  assign n3853 = n3788 & ~n3843;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~n3850 & ~n3851;
  assign n3856 = n3854 & n3855;
  assign n3857 = ~n3844 & ~n3846;
  assign n3858 = n3849 & n3857;
  assign n3859 = n3856 & n3858;
  assign n3860 = n3837 & n3859;
  assign n3861 = n3720_1 & ~n3860;
  assign n3862 = P1_REG0_REG_1_ & ~n3720_1;
  assign n435 = n3861 | n3862;
  assign n3864 = P1_IR_REG_31_ & n2657;
  assign n3865 = P1_IR_REG_2_ & ~P1_IR_REG_31_;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n3727 & ~n3866;
  assign n3868 = ~n2675_1 & ~n3727;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = n3733 & n3813;
  assign n3871 = ~n3869 & ~n3870;
  assign n3872 = n3869 & n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = n3775_1 & n3873;
  assign n3875 = ~P1_REG3_REG_3_ & n3749;
  assign n3876 = P1_REG0_REG_3_ & n3751;
  assign n3877 = P1_REG1_REG_3_ & n3753;
  assign n3878 = P1_REG2_REG_3_ & n3755_1;
  assign n3879 = ~n3875 & ~n3876;
  assign n3880 = ~n3877 & n3879;
  assign n3881 = ~n3878 & n3880;
  assign n3882 = n3742 & ~n3881;
  assign n3883 = ~n3739 & ~n3869;
  assign n3884 = ~n3824 & ~n3869;
  assign n3885 = n3824 & n3869;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~n3828 & n3830;
  assign n3888 = ~n3827 & ~n3887;
  assign n3889 = n3886 & ~n3888;
  assign n3890 = n3824 & ~n3869;
  assign n3891 = ~n3824 & n3869;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = ~n3827 & n3892;
  assign n3894 = ~n3887 & n3893;
  assign n3895 = ~n3889 & ~n3894;
  assign n3896 = n3772 & n3895;
  assign n3897 = ~n3874 & ~n3882;
  assign n3898 = ~n3883 & n3897;
  assign n3899 = ~n3896 & n3898;
  assign n3900 = ~n3759 & ~n3768;
  assign n3901 = n3759 & n3768;
  assign n3902 = n3813 & ~n3901;
  assign n3903 = ~n3900 & ~n3902;
  assign n3904 = n3892 & n3903;
  assign n3905 = ~n3892 & ~n3903;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = n3795 & ~n3906;
  assign n3908 = ~n3759 & n3845;
  assign n3909 = n3790 & n3895;
  assign n3910 = n3793 & ~n3906;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = n3785 & n3895;
  assign n3913 = n3779 & n3895;
  assign n3914 = n3782 & ~n3906;
  assign n3915 = n3788 & ~n3906;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = ~n3912 & ~n3913;
  assign n3918 = n3916 & n3917;
  assign n3919 = ~n3907 & ~n3908;
  assign n3920 = n3911 & n3919;
  assign n3921 = n3918 & n3920;
  assign n3922 = n3899 & n3921;
  assign n3923 = n3720_1 & ~n3922;
  assign n3924 = P1_REG0_REG_2_ & ~n3720_1;
  assign n440 = n3923 | n3924;
  assign n3926 = P1_IR_REG_31_ & n2681;
  assign n3927 = P1_IR_REG_3_ & ~P1_IR_REG_31_;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = n3727 & ~n3928;
  assign n3930 = ~n2706 & ~n3727;
  assign n3931 = ~n3929 & ~n3930;
  assign n3932 = ~n3872 & ~n3931;
  assign n3933 = n3872 & n3931;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = n3775_1 & n3934;
  assign n3936 = ~P1_REG3_REG_4_ & P1_REG3_REG_3_;
  assign n3937 = P1_REG3_REG_4_ & ~P1_REG3_REG_3_;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = n3749 & ~n3938;
  assign n3940 = P1_REG0_REG_4_ & n3751;
  assign n3941 = P1_REG1_REG_4_ & n3753;
  assign n3942 = P1_REG2_REG_4_ & n3755_1;
  assign n3943 = ~n3939 & ~n3940;
  assign n3944 = ~n3941 & n3943;
  assign n3945 = ~n3942 & n3944;
  assign n3946 = n3742 & ~n3945;
  assign n3947 = ~n3739 & ~n3931;
  assign n3948 = n3827 & ~n3885;
  assign n3949 = ~n3884 & ~n3948;
  assign n3950 = ~n3885 & n3887;
  assign n3951 = n3949 & ~n3950;
  assign n3952 = n3881 & ~n3931;
  assign n3953 = ~n3881 & n3931;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = n3951 & ~n3954;
  assign n3956 = ~n3881 & ~n3931;
  assign n3957 = n3881 & n3931;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = ~n3951 & ~n3958;
  assign n3960 = ~n3955 & ~n3959;
  assign n3961 = n3772 & ~n3960;
  assign n3962 = ~n3935 & ~n3946;
  assign n3963 = ~n3947 & n3962;
  assign n3964 = ~n3961 & n3963;
  assign n3965 = ~n3890 & ~n3954;
  assign n3966 = ~n3891 & n3903;
  assign n3967 = n3965 & ~n3966;
  assign n3968 = ~n3891 & n3954;
  assign n3969 = ~n3890 & ~n3903;
  assign n3970 = n3968 & ~n3969;
  assign n3971 = ~n3967 & ~n3970;
  assign n3972 = n3795 & ~n3971;
  assign n3973 = ~n3824 & n3845;
  assign n3974 = n3790 & ~n3960;
  assign n3975 = n3793 & ~n3971;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = n3785 & ~n3960;
  assign n3978 = n3779 & ~n3960;
  assign n3979 = n3782 & ~n3971;
  assign n3980 = n3788 & ~n3971;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = ~n3977 & ~n3978;
  assign n3983 = n3981 & n3982;
  assign n3984 = ~n3972 & ~n3973;
  assign n3985 = n3976 & n3984;
  assign n3986 = n3983 & n3985;
  assign n3987 = n3964 & n3986;
  assign n3988 = n3720_1 & ~n3987;
  assign n3989 = P1_REG0_REG_3_ & ~n3720_1;
  assign n445 = n3988 | n3989;
  assign n3991 = P1_IR_REG_31_ & n2713;
  assign n3992 = P1_IR_REG_4_ & ~P1_IR_REG_31_;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = n3727 & ~n3993;
  assign n3995 = ~n2734 & ~n3727;
  assign n3996 = ~n3994 & ~n3995;
  assign n3997 = ~n3933 & ~n3996;
  assign n3998 = n3933 & n3996;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = n3775_1 & n3999;
  assign n4001 = P1_REG3_REG_4_ & P1_REG3_REG_3_;
  assign n4002 = ~P1_REG3_REG_5_ & n4001;
  assign n4003 = P1_REG3_REG_5_ & ~n4001;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = n3749 & ~n4004;
  assign n4006 = P1_REG0_REG_5_ & n3751;
  assign n4007 = P1_REG1_REG_5_ & n3753;
  assign n4008 = P1_REG2_REG_5_ & n3755_1;
  assign n4009 = ~n4005 & ~n4006;
  assign n4010 = ~n4007 & n4009;
  assign n4011 = ~n4008 & n4010;
  assign n4012 = n3742 & ~n4011;
  assign n4013 = ~n3739 & ~n3996;
  assign n4014 = n3945 & ~n3996;
  assign n4015 = ~n3945 & n3996;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n3885 & ~n3957;
  assign n4018 = n3887 & n4017;
  assign n4019 = ~n3956 & ~n4018;
  assign n4020 = ~n3949 & ~n3957;
  assign n4021 = n4019 & ~n4020;
  assign n4022 = ~n4016 & n4021;
  assign n4023 = n3945 & n3996;
  assign n4024 = ~n3945 & ~n3996;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~n4021 & ~n4025;
  assign n4027 = ~n4022 & ~n4026;
  assign n4028 = n3772 & ~n4027;
  assign n4029 = ~n4000 & ~n4012;
  assign n4030 = ~n4013 & n4029;
  assign n4031 = ~n4028 & n4030;
  assign n4032 = n3881 & ~n3891;
  assign n4033 = n3931 & ~n4032;
  assign n4034 = ~n3881 & n3891;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = ~n3890 & ~n3952;
  assign n4037 = ~n3903 & n4036;
  assign n4038 = n4035 & ~n4037;
  assign n4039 = n4016 & n4038;
  assign n4040 = ~n4016 & ~n4038;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = n3795 & ~n4041;
  assign n4043 = n3845 & ~n3881;
  assign n4044 = n3790 & ~n4027;
  assign n4045 = n3793 & ~n4041;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = n3785 & ~n4027;
  assign n4048 = n3779 & ~n4027;
  assign n4049 = n3782 & ~n4041;
  assign n4050 = n3788 & ~n4041;
  assign n4051 = ~n4049 & ~n4050;
  assign n4052 = ~n4047 & ~n4048;
  assign n4053 = n4051 & n4052;
  assign n4054 = ~n4042 & ~n4043;
  assign n4055 = n4046 & n4054;
  assign n4056 = n4053 & n4055;
  assign n4057 = n4031 & n4056;
  assign n4058 = n3720_1 & ~n4057;
  assign n4059 = P1_REG0_REG_4_ & ~n3720_1;
  assign n450 = n4058 | n4059;
  assign n4061 = P1_IR_REG_31_ & n2740_1;
  assign n4062 = P1_IR_REG_5_ & ~P1_IR_REG_31_;
  assign n4063 = ~n4061 & ~n4062;
  assign n4064 = n3727 & ~n4063;
  assign n4065 = ~n2758 & ~n3727;
  assign n4066 = ~n4064 & ~n4065;
  assign n4067 = n3998 & n4066;
  assign n4068 = ~n3998 & ~n4066;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = n3775_1 & n4069;
  assign n4071 = P1_REG3_REG_5_ & n4001;
  assign n4072 = ~P1_REG3_REG_6_ & n4071;
  assign n4073 = P1_REG3_REG_6_ & ~n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n3749 & ~n4074;
  assign n4076 = P1_REG0_REG_6_ & n3751;
  assign n4077 = P1_REG1_REG_6_ & n3753;
  assign n4078 = P1_REG2_REG_6_ & n3755_1;
  assign n4079 = ~n4075 & ~n4076;
  assign n4080 = ~n4077 & n4079;
  assign n4081 = ~n4078 & n4080;
  assign n4082 = n3742 & ~n4081;
  assign n4083 = ~n3739 & ~n4066;
  assign n4084 = ~n4011 & ~n4066;
  assign n4085 = n4011 & n4066;
  assign n4086 = ~n4023 & ~n4085;
  assign n4087 = ~n4084 & n4086;
  assign n4088 = n4021 & ~n4024;
  assign n4089 = n4087 & ~n4088;
  assign n4090 = n4011 & ~n4066;
  assign n4091 = ~n4011 & n4066;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = ~n4024 & n4092;
  assign n4094 = ~n4021 & ~n4023;
  assign n4095 = n4093 & ~n4094;
  assign n4096 = ~n4089 & ~n4095;
  assign n4097 = n3772 & n4096;
  assign n4098 = ~n4070 & ~n4082;
  assign n4099 = ~n4083 & n4098;
  assign n4100 = ~n4097 & n4099;
  assign n4101 = ~n4014 & ~n4038;
  assign n4102 = ~n4015 & ~n4101;
  assign n4103 = n4092 & n4102;
  assign n4104 = ~n4092 & ~n4102;
  assign n4105 = ~n4103 & ~n4104;
  assign n4106 = n3795 & ~n4105;
  assign n4107 = n3845 & ~n3945;
  assign n4108 = n3790 & n4096;
  assign n4109 = n3793 & ~n4105;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = n3785 & n4096;
  assign n4112 = n3779 & n4096;
  assign n4113 = n3782 & ~n4105;
  assign n4114 = n3788 & ~n4105;
  assign n4115 = ~n4113 & ~n4114;
  assign n4116 = ~n4111 & ~n4112;
  assign n4117 = n4115 & n4116;
  assign n4118 = ~n4106 & ~n4107;
  assign n4119 = n4110 & n4118;
  assign n4120 = n4117 & n4119;
  assign n4121 = n4100 & n4120;
  assign n4122 = n3720_1 & ~n4121;
  assign n4123 = P1_REG0_REG_5_ & ~n3720_1;
  assign n455 = n4122 | n4123;
  assign n4125 = P1_IR_REG_31_ & n2765_1;
  assign n4126 = P1_IR_REG_6_ & ~P1_IR_REG_31_;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = n3727 & ~n4127;
  assign n4129 = ~n2786 & ~n3727;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = ~n4067 & ~n4130;
  assign n4132 = n4066 & n4130;
  assign n4133 = n3998 & n4132;
  assign n4134 = ~n4131 & ~n4133;
  assign n4135 = n3775_1 & n4134;
  assign n4136 = P1_REG3_REG_6_ & n4071;
  assign n4137 = ~P1_REG3_REG_7_ & n4136;
  assign n4138 = P1_REG3_REG_7_ & ~n4136;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = n3749 & ~n4139;
  assign n4141 = P1_REG0_REG_7_ & n3751;
  assign n4142 = P1_REG1_REG_7_ & n3753;
  assign n4143 = P1_REG2_REG_7_ & n3755_1;
  assign n4144 = ~n4140 & ~n4141;
  assign n4145 = ~n4142 & n4144;
  assign n4146 = ~n4143 & n4145;
  assign n4147 = n3742 & ~n4146;
  assign n4148 = ~n3739 & ~n4130;
  assign n4149 = n4081 & ~n4130;
  assign n4150 = ~n4081 & n4130;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = n4024 & ~n4066;
  assign n4153 = ~n4024 & n4066;
  assign n4154 = ~n4011 & ~n4153;
  assign n4155 = ~n4152 & ~n4154;
  assign n4156 = n3884 & ~n3957;
  assign n4157 = ~n3956 & ~n4156;
  assign n4158 = ~n3888 & n4017;
  assign n4159 = n4157 & ~n4158;
  assign n4160 = n4086 & ~n4159;
  assign n4161 = n4155 & ~n4160;
  assign n4162 = ~n4151 & n4161;
  assign n4163 = n4081 & n4130;
  assign n4164 = ~n4081 & ~n4130;
  assign n4165 = ~n4163 & ~n4164;
  assign n4166 = ~n4161 & ~n4165;
  assign n4167 = ~n4162 & ~n4166;
  assign n4168 = n3772 & ~n4167;
  assign n4169 = ~n4135 & ~n4147;
  assign n4170 = ~n4148 & n4169;
  assign n4171 = ~n4168 & n4170;
  assign n4172 = ~n4090 & ~n4151;
  assign n4173 = ~n4091 & n4102;
  assign n4174 = n4172 & ~n4173;
  assign n4175 = ~n4091 & ~n4150;
  assign n4176 = ~n4149 & n4175;
  assign n4177 = ~n4090 & ~n4102;
  assign n4178 = n4176 & ~n4177;
  assign n4179 = ~n4174 & ~n4178;
  assign n4180 = n3795 & ~n4179;
  assign n4181 = n3845 & ~n4011;
  assign n4182 = n3790 & ~n4167;
  assign n4183 = n3793 & ~n4179;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = n3785 & ~n4167;
  assign n4186 = n3779 & ~n4167;
  assign n4187 = n3782 & ~n4179;
  assign n4188 = n3788 & ~n4179;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~n4185 & ~n4186;
  assign n4191 = n4189 & n4190;
  assign n4192 = ~n4180 & ~n4181;
  assign n4193 = n4184 & n4192;
  assign n4194 = n4191 & n4193;
  assign n4195 = n4171 & n4194;
  assign n4196 = n3720_1 & ~n4195;
  assign n4197 = P1_REG0_REG_6_ & ~n3720_1;
  assign n460 = n4196 | n4197;
  assign n4199 = P1_IR_REG_31_ & n2792;
  assign n4200 = P1_IR_REG_7_ & ~P1_IR_REG_31_;
  assign n4201 = ~n4199 & ~n4200;
  assign n4202 = n3727 & ~n4201;
  assign n4203 = ~n2813 & ~n3727;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = ~n4133 & ~n4204;
  assign n4206 = n4133 & n4204;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = n3775_1 & n4207;
  assign n4209 = P1_REG3_REG_7_ & n4136;
  assign n4210 = ~P1_REG3_REG_8_ & n4209;
  assign n4211 = P1_REG3_REG_8_ & ~n4209;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = n3749 & ~n4212;
  assign n4214 = P1_REG0_REG_8_ & n3751;
  assign n4215 = P1_REG1_REG_8_ & n3753;
  assign n4216 = P1_REG2_REG_8_ & n3755_1;
  assign n4217 = ~n4213 & ~n4214;
  assign n4218 = ~n4215 & n4217;
  assign n4219 = ~n4216 & n4218;
  assign n4220 = n3742 & ~n4219;
  assign n4221 = ~n3739 & ~n4204;
  assign n4222 = ~n4146 & ~n4204;
  assign n4223 = n4146 & n4204;
  assign n4224 = ~n4163 & ~n4223;
  assign n4225 = ~n4222 & n4224;
  assign n4226 = n4161 & ~n4164;
  assign n4227 = n4225 & ~n4226;
  assign n4228 = n4146 & ~n4204;
  assign n4229 = ~n4146 & n4204;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = ~n4164 & n4230;
  assign n4232 = ~n4161 & ~n4163;
  assign n4233 = n4231 & ~n4232;
  assign n4234 = ~n4227 & ~n4233;
  assign n4235 = n3772 & n4234;
  assign n4236 = ~n4208 & ~n4220;
  assign n4237 = ~n4221 & n4236;
  assign n4238 = ~n4235 & n4237;
  assign n4239 = ~n4090 & ~n4149;
  assign n4240 = n4015 & n4239;
  assign n4241 = n4175 & ~n4240;
  assign n4242 = ~n4149 & ~n4241;
  assign n4243 = n4101 & n4239;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = n4230 & n4244;
  assign n4246 = ~n4230 & ~n4244;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = n3795 & ~n4247;
  assign n4249 = n3845 & ~n4081;
  assign n4250 = n3790 & n4234;
  assign n4251 = n3793 & ~n4247;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = n3785 & n4234;
  assign n4254 = n3779 & n4234;
  assign n4255 = n3782 & ~n4247;
  assign n4256 = n3788 & ~n4247;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n4253 & ~n4254;
  assign n4259 = n4257 & n4258;
  assign n4260 = ~n4248 & ~n4249;
  assign n4261 = n4252 & n4260;
  assign n4262 = n4259 & n4261;
  assign n4263 = n4238 & n4262;
  assign n4264 = n3720_1 & ~n4263;
  assign n4265 = P1_REG0_REG_7_ & ~n3720_1;
  assign n465 = n4264 | n4265;
  assign n4267 = P1_IR_REG_31_ & n2823;
  assign n4268 = P1_IR_REG_8_ & ~P1_IR_REG_31_;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = n3727 & ~n4269;
  assign n4271 = ~n2841 & ~n3727;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = ~n4206 & ~n4272;
  assign n4274 = n4206 & n4272;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = n3775_1 & n4275;
  assign n4277 = P1_REG1_REG_9_ & n3753;
  assign n4278 = P1_REG0_REG_9_ & n3751;
  assign n4279 = P1_REG2_REG_9_ & n3755_1;
  assign n4280 = P1_REG3_REG_8_ & n4209;
  assign n4281 = ~P1_REG3_REG_9_ & n4280;
  assign n4282 = P1_REG3_REG_9_ & ~n4280;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = n3749 & ~n4283;
  assign n4285 = ~n4277 & ~n4278;
  assign n4286 = ~n4279 & n4285;
  assign n4287 = ~n4284 & n4286;
  assign n4288 = n3742 & ~n4287;
  assign n4289 = ~n3739 & ~n4272;
  assign n4290 = n4164 & ~n4204;
  assign n4291 = ~n4164 & n4204;
  assign n4292 = ~n4146 & ~n4291;
  assign n4293 = ~n4290 & ~n4292;
  assign n4294 = ~n4161 & n4224;
  assign n4295 = n4293 & ~n4294;
  assign n4296 = n4219 & ~n4272;
  assign n4297 = ~n4219 & n4272;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = n4295 & ~n4298;
  assign n4300 = n4219 & n4272;
  assign n4301 = ~n4219 & ~n4272;
  assign n4302 = ~n4300 & ~n4301;
  assign n4303 = ~n4295 & ~n4302;
  assign n4304 = ~n4299 & ~n4303;
  assign n4305 = n3772 & ~n4304;
  assign n4306 = ~n4276 & ~n4288;
  assign n4307 = ~n4289 & n4306;
  assign n4308 = ~n4305 & n4307;
  assign n4309 = ~n4228 & ~n4298;
  assign n4310 = ~n4229 & n4244;
  assign n4311 = n4309 & ~n4310;
  assign n4312 = ~n4229 & n4298;
  assign n4313 = ~n4228 & ~n4244;
  assign n4314 = n4312 & ~n4313;
  assign n4315 = ~n4311 & ~n4314;
  assign n4316 = n3795 & ~n4315;
  assign n4317 = n3845 & ~n4146;
  assign n4318 = n3790 & ~n4304;
  assign n4319 = n3793 & ~n4315;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = n3785 & ~n4304;
  assign n4322 = n3779 & ~n4304;
  assign n4323 = n3782 & ~n4315;
  assign n4324 = n3788 & ~n4315;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4321 & ~n4322;
  assign n4327 = n4325 & n4326;
  assign n4328 = ~n4316 & ~n4317;
  assign n4329 = n4320 & n4328;
  assign n4330 = n4327 & n4329;
  assign n4331 = n4308 & n4330;
  assign n4332 = n3720_1 & ~n4331;
  assign n4333 = P1_REG0_REG_8_ & ~n3720_1;
  assign n470 = n4332 | n4333;
  assign n4335 = P1_IR_REG_31_ & n2847;
  assign n4336 = P1_IR_REG_9_ & ~P1_IR_REG_31_;
  assign n4337 = ~n4335 & ~n4336;
  assign n4338 = n3727 & ~n4337;
  assign n4339 = ~n2868 & ~n3727;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = n4274 & n4340;
  assign n4342 = ~n4274 & ~n4340;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = n3775_1 & n4343;
  assign n4345 = P1_REG1_REG_10_ & n3753;
  assign n4346 = P1_REG0_REG_10_ & n3751;
  assign n4347 = P1_REG2_REG_10_ & n3755_1;
  assign n4348 = P1_REG3_REG_9_ & n4280;
  assign n4349 = ~P1_REG3_REG_10_ & n4348;
  assign n4350 = P1_REG3_REG_10_ & ~n4348;
  assign n4351 = ~n4349 & ~n4350;
  assign n4352 = n3749 & ~n4351;
  assign n4353 = ~n4345 & ~n4346;
  assign n4354 = ~n4347 & n4353;
  assign n4355 = ~n4352 & n4354;
  assign n4356 = n3742 & ~n4355;
  assign n4357 = ~n3739 & ~n4340;
  assign n4358 = n4287 & ~n4340;
  assign n4359 = ~n4287 & n4340;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~n4295 & ~n4300;
  assign n4362 = ~n4301 & ~n4361;
  assign n4363 = ~n4360 & n4362;
  assign n4364 = n4287 & n4340;
  assign n4365 = ~n4287 & ~n4340;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4362 & ~n4366;
  assign n4368 = ~n4363 & ~n4367;
  assign n4369 = n3772 & ~n4368;
  assign n4370 = ~n4344 & ~n4356;
  assign n4371 = ~n4357 & n4370;
  assign n4372 = ~n4369 & n4371;
  assign n4373 = n4219 & ~n4229;
  assign n4374 = n4272 & ~n4373;
  assign n4375 = ~n4219 & n4229;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = ~n4228 & ~n4296;
  assign n4378 = ~n4244 & n4377;
  assign n4379 = n4376 & ~n4378;
  assign n4380 = n4360 & n4379;
  assign n4381 = ~n4360 & ~n4379;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = n3795 & ~n4382;
  assign n4384 = n3845 & ~n4219;
  assign n4385 = n3790 & ~n4368;
  assign n4386 = n3793 & ~n4382;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = n3785 & ~n4368;
  assign n4389 = n3779 & ~n4368;
  assign n4390 = n3782 & ~n4382;
  assign n4391 = n3788 & ~n4382;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = ~n4388 & ~n4389;
  assign n4394 = n4392 & n4393;
  assign n4395 = ~n4383 & ~n4384;
  assign n4396 = n4387 & n4395;
  assign n4397 = n4394 & n4396;
  assign n4398 = n4372 & n4397;
  assign n4399 = n3720_1 & ~n4398;
  assign n4400 = P1_REG0_REG_9_ & ~n3720_1;
  assign n475 = n4399 | n4400;
  assign n4402 = P1_IR_REG_31_ & n2875_1;
  assign n4403 = P1_IR_REG_10_ & ~P1_IR_REG_31_;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = n3727 & ~n4404;
  assign n4406 = ~n2896 & ~n3727;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = ~n4341 & ~n4407;
  assign n4409 = n4340 & n4407;
  assign n4410 = n4274 & n4409;
  assign n4411 = ~n4408 & ~n4410;
  assign n4412 = n3775_1 & n4411;
  assign n4413 = P1_REG1_REG_11_ & n3753;
  assign n4414 = P1_REG0_REG_11_ & n3751;
  assign n4415 = P1_REG2_REG_11_ & n3755_1;
  assign n4416 = P1_REG3_REG_10_ & n4348;
  assign n4417 = ~P1_REG3_REG_11_ & n4416;
  assign n4418 = P1_REG3_REG_11_ & ~n4416;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = n3749 & ~n4419;
  assign n4421 = ~n4413 & ~n4414;
  assign n4422 = ~n4415 & n4421;
  assign n4423 = ~n4420 & n4422;
  assign n4424 = n3742 & ~n4423;
  assign n4425 = ~n3739 & ~n4407;
  assign n4426 = ~n4355 & ~n4407;
  assign n4427 = n4355 & n4407;
  assign n4428 = ~n4364 & ~n4427;
  assign n4429 = ~n4426 & n4428;
  assign n4430 = n4362 & ~n4365;
  assign n4431 = n4429 & ~n4430;
  assign n4432 = n4355 & ~n4407;
  assign n4433 = ~n4355 & n4407;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4365 & n4434;
  assign n4436 = ~n4362 & ~n4364;
  assign n4437 = n4435 & ~n4436;
  assign n4438 = ~n4431 & ~n4437;
  assign n4439 = n3772 & n4438;
  assign n4440 = ~n4412 & ~n4424;
  assign n4441 = ~n4425 & n4440;
  assign n4442 = ~n4439 & n4441;
  assign n4443 = ~n4358 & ~n4379;
  assign n4444 = ~n4359 & ~n4443;
  assign n4445 = n4434 & n4444;
  assign n4446 = ~n4434 & ~n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n3795 & ~n4447;
  assign n4449 = n3845 & ~n4287;
  assign n4450 = n3790 & n4438;
  assign n4451 = n3793 & ~n4447;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = n3785 & n4438;
  assign n4454 = n3779 & n4438;
  assign n4455 = n3782 & ~n4447;
  assign n4456 = n3788 & ~n4447;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n4453 & ~n4454;
  assign n4459 = n4457 & n4458;
  assign n4460 = ~n4448 & ~n4449;
  assign n4461 = n4452 & n4460;
  assign n4462 = n4459 & n4461;
  assign n4463 = n4442 & n4462;
  assign n4464 = n3720_1 & ~n4463;
  assign n4465 = P1_REG0_REG_10_ & ~n3720_1;
  assign n480 = n4464 | n4465;
  assign n4467 = P1_IR_REG_31_ & n2902;
  assign n4468 = P1_IR_REG_11_ & ~P1_IR_REG_31_;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n3727 & ~n4469;
  assign n4471 = ~n2923 & ~n3727;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = ~n3739 & ~n4472;
  assign n4474 = ~n4410 & ~n4472;
  assign n4475 = n4410 & n4472;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = n3775_1 & n4476;
  assign n4478 = ~n4365 & ~n4426;
  assign n4479 = n4301 & n4428;
  assign n4480 = n4478 & ~n4479;
  assign n4481 = ~n4427 & ~n4480;
  assign n4482 = ~n4300 & n4428;
  assign n4483 = ~n4295 & n4482;
  assign n4484 = ~n4481 & ~n4483;
  assign n4485 = n4423 & ~n4472;
  assign n4486 = ~n4423 & n4472;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = n4484 & ~n4487;
  assign n4489 = n4423 & n4472;
  assign n4490 = ~n4423 & ~n4472;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = ~n4484 & ~n4491;
  assign n4493 = ~n4488 & ~n4492;
  assign n4494 = n3772 & ~n4493;
  assign n4495 = P1_REG1_REG_12_ & n3753;
  assign n4496 = P1_REG0_REG_12_ & n3751;
  assign n4497 = P1_REG2_REG_12_ & n3755_1;
  assign n4498 = P1_REG3_REG_11_ & n4416;
  assign n4499 = ~P1_REG3_REG_12_ & n4498;
  assign n4500 = P1_REG3_REG_12_ & ~n4498;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = n3749 & ~n4501;
  assign n4503 = ~n4495 & ~n4496;
  assign n4504 = ~n4497 & n4503;
  assign n4505 = ~n4502 & n4504;
  assign n4506 = n3742 & ~n4505;
  assign n4507 = ~n4473 & ~n4477;
  assign n4508 = ~n4494 & n4507;
  assign n4509 = ~n4506 & n4508;
  assign n4510 = ~n4432 & ~n4487;
  assign n4511 = ~n4433 & n4444;
  assign n4512 = n4510 & ~n4511;
  assign n4513 = ~n4433 & ~n4486;
  assign n4514 = ~n4485 & n4513;
  assign n4515 = ~n4432 & ~n4444;
  assign n4516 = n4514 & ~n4515;
  assign n4517 = ~n4512 & ~n4516;
  assign n4518 = n3795 & ~n4517;
  assign n4519 = n3845 & ~n4355;
  assign n4520 = n3790 & ~n4493;
  assign n4521 = n3793 & ~n4517;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = n3785 & ~n4493;
  assign n4524 = n3779 & ~n4493;
  assign n4525 = n3782 & ~n4517;
  assign n4526 = n3788 & ~n4517;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = ~n4523 & ~n4524;
  assign n4529 = n4527 & n4528;
  assign n4530 = ~n4518 & ~n4519;
  assign n4531 = n4522 & n4530;
  assign n4532 = n4529 & n4531;
  assign n4533 = n4509 & n4532;
  assign n4534 = n3720_1 & ~n4533;
  assign n4535 = P1_REG0_REG_11_ & ~n3720_1;
  assign n485 = n4534 | n4535;
  assign n4537 = P1_IR_REG_31_ & n2932;
  assign n4538 = P1_IR_REG_12_ & ~P1_IR_REG_31_;
  assign n4539 = ~n4537 & ~n4538;
  assign n4540 = n3727 & ~n4539;
  assign n4541 = ~n2950_1 & ~n3727;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n3739 & ~n4542;
  assign n4544 = n4505 & ~n4542;
  assign n4545 = ~n4505 & n4542;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~n4484 & ~n4489;
  assign n4548 = ~n4490 & ~n4547;
  assign n4549 = ~n4546 & n4548;
  assign n4550 = n4505 & n4542;
  assign n4551 = ~n4505 & ~n4542;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4548 & ~n4552;
  assign n4554 = ~n4549 & ~n4553;
  assign n4555 = n3772 & ~n4554;
  assign n4556 = ~n4475 & ~n4542;
  assign n4557 = n4475 & n4542;
  assign n4558 = ~n4556 & ~n4557;
  assign n4559 = n3775_1 & n4558;
  assign n4560 = P1_REG1_REG_13_ & n3753;
  assign n4561 = P1_REG0_REG_13_ & n3751;
  assign n4562 = P1_REG2_REG_13_ & n3755_1;
  assign n4563 = P1_REG3_REG_12_ & n4498;
  assign n4564 = ~P1_REG3_REG_13_ & n4563;
  assign n4565 = P1_REG3_REG_13_ & ~n4563;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n3749 & ~n4566;
  assign n4568 = ~n4560 & ~n4561;
  assign n4569 = ~n4562 & n4568;
  assign n4570 = ~n4567 & n4569;
  assign n4571 = n3742 & ~n4570;
  assign n4572 = ~n4543 & ~n4555;
  assign n4573 = ~n4559 & n4572;
  assign n4574 = ~n4571 & n4573;
  assign n4575 = ~n4432 & ~n4485;
  assign n4576 = n4359 & n4575;
  assign n4577 = n4513 & ~n4576;
  assign n4578 = ~n4485 & ~n4577;
  assign n4579 = ~n4358 & n4575;
  assign n4580 = ~n4379 & n4579;
  assign n4581 = ~n4578 & ~n4580;
  assign n4582 = ~n4546 & ~n4581;
  assign n4583 = n4546 & n4581;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = n3795 & ~n4584;
  assign n4586 = n3845 & ~n4423;
  assign n4587 = n3790 & ~n4554;
  assign n4588 = n3793 & ~n4584;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = n3785 & ~n4554;
  assign n4591 = n3779 & ~n4554;
  assign n4592 = n3782 & ~n4584;
  assign n4593 = n3788 & ~n4584;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = ~n4590 & ~n4591;
  assign n4596 = n4594 & n4595;
  assign n4597 = ~n4585 & ~n4586;
  assign n4598 = n4589 & n4597;
  assign n4599 = n4596 & n4598;
  assign n4600 = n4574 & n4599;
  assign n4601 = n3720_1 & ~n4600;
  assign n4602 = P1_REG0_REG_12_ & ~n3720_1;
  assign n490 = n4601 | n4602;
  assign n4604 = P1_IR_REG_31_ & n2956;
  assign n4605 = P1_IR_REG_13_ & ~P1_IR_REG_31_;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = n3727 & ~n4606;
  assign n4608 = ~n2977 & ~n3727;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = ~n3739 & ~n4609;
  assign n4611 = n4557 & n4609;
  assign n4612 = ~n4557 & ~n4609;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = n3775_1 & n4613;
  assign n4615 = ~n4570 & ~n4609;
  assign n4616 = n4570 & n4609;
  assign n4617 = ~n4550 & ~n4616;
  assign n4618 = ~n4615 & n4617;
  assign n4619 = n4548 & ~n4551;
  assign n4620 = n4618 & ~n4619;
  assign n4621 = n4570 & ~n4609;
  assign n4622 = ~n4570 & n4609;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = ~n4551 & n4623;
  assign n4625 = ~n4548 & ~n4550;
  assign n4626 = n4624 & ~n4625;
  assign n4627 = ~n4620 & ~n4626;
  assign n4628 = n3772 & n4627;
  assign n4629 = P1_REG1_REG_14_ & n3753;
  assign n4630 = P1_REG0_REG_14_ & n3751;
  assign n4631 = P1_REG2_REG_14_ & n3755_1;
  assign n4632 = P1_REG3_REG_13_ & n4563;
  assign n4633 = ~P1_REG3_REG_14_ & n4632;
  assign n4634 = P1_REG3_REG_14_ & ~n4632;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = n3749 & ~n4635;
  assign n4637 = ~n4629 & ~n4630;
  assign n4638 = ~n4631 & n4637;
  assign n4639 = ~n4636 & n4638;
  assign n4640 = n3742 & ~n4639;
  assign n4641 = ~n4610 & ~n4614;
  assign n4642 = ~n4628 & n4641;
  assign n4643 = ~n4640 & n4642;
  assign n4644 = ~n4544 & ~n4581;
  assign n4645 = ~n4545 & ~n4644;
  assign n4646 = ~n4623 & ~n4645;
  assign n4647 = n4623 & n4645;
  assign n4648 = ~n4646 & ~n4647;
  assign n4649 = n3795 & ~n4648;
  assign n4650 = n3845 & ~n4505;
  assign n4651 = n3790 & n4627;
  assign n4652 = n3793 & ~n4648;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = n3785 & n4627;
  assign n4655 = n3779 & n4627;
  assign n4656 = n3782 & ~n4648;
  assign n4657 = n3788 & ~n4648;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n4654 & ~n4655;
  assign n4660 = n4658 & n4659;
  assign n4661 = ~n4649 & ~n4650;
  assign n4662 = n4653 & n4661;
  assign n4663 = n4660 & n4662;
  assign n4664 = n4643 & n4663;
  assign n4665 = n3720_1 & ~n4664;
  assign n4666 = P1_REG0_REG_13_ & ~n3720_1;
  assign n495 = n4665 | n4666;
  assign n4668 = P1_IR_REG_31_ & n2984;
  assign n4669 = P1_IR_REG_14_ & ~P1_IR_REG_31_;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = n3727 & ~n4670;
  assign n4672 = ~n3005_1 & ~n3727;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = ~n3739 & ~n4673;
  assign n4675 = ~n4551 & ~n4615;
  assign n4676 = n4490 & n4617;
  assign n4677 = n4675 & ~n4676;
  assign n4678 = ~n4616 & ~n4677;
  assign n4679 = n4547 & n4617;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = n4639 & ~n4673;
  assign n4682 = ~n4639 & n4673;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = n4680 & ~n4683;
  assign n4685 = ~n4680 & n4683;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = n3772 & ~n4686;
  assign n4688 = ~n4611 & ~n4673;
  assign n4689 = n4609 & n4673;
  assign n4690 = n4557 & n4689;
  assign n4691 = ~n4688 & ~n4690;
  assign n4692 = n3775_1 & n4691;
  assign n4693 = P1_REG1_REG_15_ & n3753;
  assign n4694 = P1_REG0_REG_15_ & n3751;
  assign n4695 = P1_REG2_REG_15_ & n3755_1;
  assign n4696 = P1_REG3_REG_14_ & n4632;
  assign n4697 = ~P1_REG3_REG_15_ & n4696;
  assign n4698 = P1_REG3_REG_15_ & ~n4696;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = n3749 & ~n4699;
  assign n4701 = ~n4693 & ~n4694;
  assign n4702 = ~n4695 & n4701;
  assign n4703 = ~n4700 & n4702;
  assign n4704 = n3742 & ~n4703;
  assign n4705 = ~n4674 & ~n4687;
  assign n4706 = ~n4692 & n4705;
  assign n4707 = ~n4704 & n4706;
  assign n4708 = ~n4621 & ~n4645;
  assign n4709 = ~n4622 & ~n4708;
  assign n4710 = n4683 & n4709;
  assign n4711 = ~n4683 & ~n4709;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = n3795 & ~n4712;
  assign n4714 = n3845 & ~n4570;
  assign n4715 = n3790 & ~n4686;
  assign n4716 = n3793 & ~n4712;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = n3785 & ~n4686;
  assign n4719 = n3779 & ~n4686;
  assign n4720 = n3782 & ~n4712;
  assign n4721 = n3788 & ~n4712;
  assign n4722 = ~n4720 & ~n4721;
  assign n4723 = ~n4718 & ~n4719;
  assign n4724 = n4722 & n4723;
  assign n4725 = ~n4713 & ~n4714;
  assign n4726 = n4717 & n4725;
  assign n4727 = n4724 & n4726;
  assign n4728 = n4707 & n4727;
  assign n4729 = n3720_1 & ~n4728;
  assign n4730 = P1_REG0_REG_14_ & ~n3720_1;
  assign n500 = n4729 | n4730;
  assign n4732 = P1_IR_REG_31_ & n3011;
  assign n4733 = P1_IR_REG_15_ & ~P1_IR_REG_31_;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = n3727 & ~n4734;
  assign n4736 = ~n3032 & ~n3727;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = ~n4690 & ~n4737;
  assign n4739 = n4690 & n4737;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = n3775_1 & n4740;
  assign n4742 = P1_REG1_REG_16_ & n3753;
  assign n4743 = P1_REG0_REG_16_ & n3751;
  assign n4744 = P1_REG2_REG_16_ & n3755_1;
  assign n4745 = P1_REG3_REG_15_ & n4696;
  assign n4746 = ~P1_REG3_REG_16_ & n4745;
  assign n4747 = P1_REG3_REG_16_ & ~n4745;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = n3749 & ~n4748;
  assign n4750 = ~n4742 & ~n4743;
  assign n4751 = ~n4744 & n4750;
  assign n4752 = ~n4749 & n4751;
  assign n4753 = n3742 & ~n4752;
  assign n4754 = ~n3739 & ~n4737;
  assign n4755 = ~n4639 & ~n4673;
  assign n4756 = n4639 & n4673;
  assign n4757 = ~n4680 & ~n4756;
  assign n4758 = ~n4755 & ~n4757;
  assign n4759 = n4703 & ~n4737;
  assign n4760 = ~n4703 & n4737;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = n4758 & ~n4761;
  assign n4763 = ~n4758 & n4761;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = n3772 & ~n4764;
  assign n4766 = ~n4741 & ~n4753;
  assign n4767 = ~n4754 & n4766;
  assign n4768 = ~n4765 & n4767;
  assign n4769 = ~n4681 & ~n4709;
  assign n4770 = ~n4682 & ~n4769;
  assign n4771 = n4761 & n4770;
  assign n4772 = ~n4761 & ~n4770;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = n3795 & ~n4773;
  assign n4775 = n3845 & ~n4639;
  assign n4776 = n3790 & ~n4764;
  assign n4777 = n3793 & ~n4773;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = n3785 & ~n4764;
  assign n4780 = n3779 & ~n4764;
  assign n4781 = n3782 & ~n4773;
  assign n4782 = n3788 & ~n4773;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = ~n4779 & ~n4780;
  assign n4785 = n4783 & n4784;
  assign n4786 = ~n4774 & ~n4775;
  assign n4787 = n4778 & n4786;
  assign n4788 = n4785 & n4787;
  assign n4789 = n4768 & n4788;
  assign n4790 = n3720_1 & ~n4789;
  assign n4791 = P1_REG0_REG_15_ & ~n3720_1;
  assign n505 = n4790 | n4791;
  assign n4793 = P1_IR_REG_31_ & n3052;
  assign n4794 = P1_IR_REG_16_ & ~P1_IR_REG_31_;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = n3727 & ~n4795;
  assign n4797 = ~n3073 & ~n3727;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n4739 & ~n4798;
  assign n4800 = n4739 & n4798;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = n3775_1 & n4801;
  assign n4803 = P1_REG1_REG_17_ & n3753;
  assign n4804 = P1_REG0_REG_17_ & n3751;
  assign n4805 = P1_REG2_REG_17_ & n3755_1;
  assign n4806 = P1_REG3_REG_16_ & n4745;
  assign n4807 = ~P1_REG3_REG_17_ & n4806;
  assign n4808 = P1_REG3_REG_17_ & ~n4806;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = n3749 & ~n4809;
  assign n4811 = ~n4803 & ~n4804;
  assign n4812 = ~n4805 & n4811;
  assign n4813 = ~n4810 & n4812;
  assign n4814 = n3742 & ~n4813;
  assign n4815 = ~n3739 & ~n4798;
  assign n4816 = n4752 & ~n4798;
  assign n4817 = ~n4752 & n4798;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = ~n4703 & ~n4737;
  assign n4820 = n4703 & n4737;
  assign n4821 = ~n4758 & ~n4820;
  assign n4822 = ~n4819 & ~n4821;
  assign n4823 = ~n4818 & n4822;
  assign n4824 = n4752 & n4798;
  assign n4825 = ~n4752 & ~n4798;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = ~n4822 & ~n4826;
  assign n4828 = ~n4823 & ~n4827;
  assign n4829 = n3772 & ~n4828;
  assign n4830 = ~n4802 & ~n4814;
  assign n4831 = ~n4815 & n4830;
  assign n4832 = ~n4829 & n4831;
  assign n4833 = ~n4759 & ~n4818;
  assign n4834 = ~n4760 & n4770;
  assign n4835 = n4833 & ~n4834;
  assign n4836 = ~n4759 & ~n4770;
  assign n4837 = ~n4760 & ~n4817;
  assign n4838 = ~n4816 & ~n4836;
  assign n4839 = n4837 & n4838;
  assign n4840 = ~n4835 & ~n4839;
  assign n4841 = n3795 & ~n4840;
  assign n4842 = n3845 & ~n4703;
  assign n4843 = n3790 & ~n4828;
  assign n4844 = n3793 & ~n4840;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = n3785 & ~n4828;
  assign n4847 = n3779 & ~n4828;
  assign n4848 = n3782 & ~n4840;
  assign n4849 = n3788 & ~n4840;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4846 & ~n4847;
  assign n4852 = n4850 & n4851;
  assign n4853 = ~n4841 & ~n4842;
  assign n4854 = n4845 & n4853;
  assign n4855 = n4852 & n4854;
  assign n4856 = n4832 & n4855;
  assign n4857 = n3720_1 & ~n4856;
  assign n4858 = P1_REG0_REG_16_ & ~n3720_1;
  assign n510 = n4857 | n4858;
  assign n4860 = P1_IR_REG_31_ & n3079;
  assign n4861 = P1_IR_REG_17_ & ~P1_IR_REG_31_;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = n3727 & ~n4862;
  assign n4864 = ~n3097 & ~n3727;
  assign n4865 = ~n4863 & ~n4864;
  assign n4866 = ~n3739 & ~n4865;
  assign n4867 = ~n4813 & ~n4865;
  assign n4868 = n4822 & ~n4825;
  assign n4869 = n4813 & n4865;
  assign n4870 = ~n4824 & ~n4869;
  assign n4871 = ~n4867 & ~n4868;
  assign n4872 = n4870 & n4871;
  assign n4873 = n4813 & ~n4865;
  assign n4874 = ~n4813 & n4865;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n4825 & n4875;
  assign n4877 = ~n4822 & ~n4824;
  assign n4878 = n4876 & ~n4877;
  assign n4879 = ~n4872 & ~n4878;
  assign n4880 = n3772 & n4879;
  assign n4881 = n4800 & n4865;
  assign n4882 = ~n4800 & ~n4865;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = n3775_1 & n4883;
  assign n4885 = P1_REG1_REG_18_ & n3753;
  assign n4886 = P1_REG0_REG_18_ & n3751;
  assign n4887 = P1_REG2_REG_18_ & n3755_1;
  assign n4888 = P1_REG3_REG_17_ & n4806;
  assign n4889 = ~P1_REG3_REG_18_ & n4888;
  assign n4890 = P1_REG3_REG_18_ & ~n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = n3749 & ~n4891;
  assign n4893 = ~n4885 & ~n4886;
  assign n4894 = ~n4887 & n4893;
  assign n4895 = ~n4892 & n4894;
  assign n4896 = n3742 & ~n4895;
  assign n4897 = ~n4866 & ~n4880;
  assign n4898 = ~n4884 & n4897;
  assign n4899 = ~n4896 & n4898;
  assign n4900 = n4682 & ~n4759;
  assign n4901 = n4837 & ~n4900;
  assign n4902 = ~n4816 & ~n4901;
  assign n4903 = ~n4681 & ~n4759;
  assign n4904 = ~n4709 & n4903;
  assign n4905 = ~n4816 & n4904;
  assign n4906 = ~n4902 & ~n4905;
  assign n4907 = ~n4875 & ~n4906;
  assign n4908 = n4875 & n4906;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = n3795 & ~n4909;
  assign n4911 = n3845 & ~n4752;
  assign n4912 = n3790 & n4879;
  assign n4913 = n3793 & ~n4909;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = n3785 & n4879;
  assign n4916 = n3779 & n4879;
  assign n4917 = n3782 & ~n4909;
  assign n4918 = n3788 & ~n4909;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = ~n4915 & ~n4916;
  assign n4921 = n4919 & n4920;
  assign n4922 = ~n4910 & ~n4911;
  assign n4923 = n4914 & n4922;
  assign n4924 = n4921 & n4923;
  assign n4925 = n4899 & n4924;
  assign n4926 = n3720_1 & ~n4925;
  assign n4927 = P1_REG0_REG_17_ & ~n3720_1;
  assign n515 = n4926 | n4927;
  assign n4929 = P1_IR_REG_31_ & n3113;
  assign n4930 = P1_IR_REG_18_ & ~P1_IR_REG_31_;
  assign n4931 = ~n4929 & ~n4930;
  assign n4932 = n3727 & ~n4931;
  assign n4933 = ~n3131 & ~n3727;
  assign n4934 = ~n4932 & ~n4933;
  assign n4935 = ~n3739 & ~n4934;
  assign n4936 = n4825 & ~n4865;
  assign n4937 = ~n4825 & n4865;
  assign n4938 = ~n4813 & ~n4937;
  assign n4939 = ~n4936 & ~n4938;
  assign n4940 = ~n4822 & n4870;
  assign n4941 = n4939 & ~n4940;
  assign n4942 = n4895 & ~n4934;
  assign n4943 = ~n4895 & n4934;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = n4941 & ~n4944;
  assign n4946 = n4895 & n4934;
  assign n4947 = ~n4895 & ~n4934;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = ~n4941 & ~n4948;
  assign n4950 = ~n4945 & ~n4949;
  assign n4951 = n3772 & ~n4950;
  assign n4952 = ~n4881 & ~n4934;
  assign n4953 = n4865 & n4934;
  assign n4954 = n4800 & n4953;
  assign n4955 = ~n4952 & ~n4954;
  assign n4956 = n3775_1 & n4955;
  assign n4957 = P1_REG1_REG_19_ & n3753;
  assign n4958 = P1_REG0_REG_19_ & n3751;
  assign n4959 = P1_REG2_REG_19_ & n3755_1;
  assign n4960 = P1_REG3_REG_18_ & n4888;
  assign n4961 = ~P1_REG3_REG_19_ & n4960;
  assign n4962 = P1_REG3_REG_19_ & ~n4960;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = n3749 & ~n4963;
  assign n4965 = ~n4957 & ~n4958;
  assign n4966 = ~n4959 & n4965;
  assign n4967 = ~n4964 & n4966;
  assign n4968 = n3742 & ~n4967;
  assign n4969 = ~n4935 & ~n4951;
  assign n4970 = ~n4956 & n4969;
  assign n4971 = ~n4968 & n4970;
  assign n4972 = ~n4873 & ~n4906;
  assign n4973 = ~n4874 & ~n4972;
  assign n4974 = ~n4944 & ~n4973;
  assign n4975 = n4944 & n4973;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = n3795 & ~n4976;
  assign n4978 = n3845 & ~n4813;
  assign n4979 = n3790 & ~n4950;
  assign n4980 = n3793 & ~n4976;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n3785 & ~n4950;
  assign n4983 = n3779 & ~n4950;
  assign n4984 = n3782 & ~n4976;
  assign n4985 = n3788 & ~n4976;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = ~n4982 & ~n4983;
  assign n4988 = n4986 & n4987;
  assign n4989 = ~n4977 & ~n4978;
  assign n4990 = n4981 & n4989;
  assign n4991 = n4988 & n4990;
  assign n4992 = n4971 & n4991;
  assign n4993 = n3720_1 & ~n4992;
  assign n4994 = P1_REG0_REG_18_ & ~n3720_1;
  assign n520 = n4993 | n4994;
  assign n4996 = ~n3655_1 & n3727;
  assign n4997 = ~n3168 & ~n3727;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n4954 & n4998;
  assign n5000 = ~n4954 & ~n4998;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = n3775_1 & n5001;
  assign n5003 = P1_REG1_REG_20_ & n3753;
  assign n5004 = P1_REG0_REG_20_ & n3751;
  assign n5005 = P1_REG2_REG_20_ & n3755_1;
  assign n5006 = P1_REG3_REG_19_ & n4960;
  assign n5007 = ~P1_REG3_REG_20_ & n5006;
  assign n5008 = P1_REG3_REG_20_ & ~n5006;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = n3749 & ~n5009;
  assign n5011 = ~n5003 & ~n5004;
  assign n5012 = ~n5005 & n5011;
  assign n5013 = ~n5010 & n5012;
  assign n5014 = n3742 & ~n5013;
  assign n5015 = ~n3739 & ~n4998;
  assign n5016 = n4967 & ~n4998;
  assign n5017 = ~n4967 & n4998;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = ~n4941 & ~n4946;
  assign n5020 = ~n4947 & ~n5019;
  assign n5021 = ~n5018 & n5020;
  assign n5022 = n4967 & n4998;
  assign n5023 = ~n4967 & ~n4998;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = ~n5020 & ~n5024;
  assign n5026 = ~n5021 & ~n5025;
  assign n5027 = n3772 & ~n5026;
  assign n5028 = ~n5002 & ~n5014;
  assign n5029 = ~n5015 & n5028;
  assign n5030 = ~n5027 & n5029;
  assign n5031 = ~n4895 & ~n4973;
  assign n5032 = n4895 & n4973;
  assign n5033 = n4934 & ~n5032;
  assign n5034 = ~n5031 & ~n5033;
  assign n5035 = ~n5018 & ~n5034;
  assign n5036 = n5018 & n5034;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = n3795 & ~n5037;
  assign n5039 = n3845 & ~n4895;
  assign n5040 = n3790 & ~n5026;
  assign n5041 = n3793 & ~n5037;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = n3785 & ~n5026;
  assign n5044 = n3779 & ~n5026;
  assign n5045 = n3782 & ~n5037;
  assign n5046 = n3788 & ~n5037;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = ~n5043 & ~n5044;
  assign n5049 = n5047 & n5048;
  assign n5050 = ~n5038 & ~n5039;
  assign n5051 = n5042 & n5050;
  assign n5052 = n5049 & n5051;
  assign n5053 = n5030 & n5052;
  assign n5054 = n3720_1 & ~n5053;
  assign n5055 = P1_REG0_REG_19_ & ~n3720_1;
  assign n525 = n5054 | n5055;
  assign n5057 = ~n3205_1 & ~n3727;
  assign n5058 = ~n4999 & n5057;
  assign n5059 = n4998 & ~n5057;
  assign n5060 = n4954 & n5059;
  assign n5061 = ~n5058 & ~n5060;
  assign n5062 = n3775_1 & n5061;
  assign n5063 = P1_REG1_REG_21_ & n3753;
  assign n5064 = P1_REG0_REG_21_ & n3751;
  assign n5065 = P1_REG2_REG_21_ & n3755_1;
  assign n5066 = P1_REG3_REG_20_ & n5006;
  assign n5067 = ~P1_REG3_REG_21_ & n5066;
  assign n5068 = P1_REG3_REG_21_ & ~n5066;
  assign n5069 = ~n5067 & ~n5068;
  assign n5070 = n3749 & ~n5069;
  assign n5071 = ~n5063 & ~n5064;
  assign n5072 = ~n5065 & n5071;
  assign n5073 = ~n5070 & n5072;
  assign n5074 = n3742 & ~n5073;
  assign n5075 = ~n3739 & n5057;
  assign n5076 = ~n5013 & n5057;
  assign n5077 = n5020 & ~n5023;
  assign n5078 = n5013 & ~n5057;
  assign n5079 = ~n5022 & ~n5078;
  assign n5080 = ~n5076 & ~n5077;
  assign n5081 = n5079 & n5080;
  assign n5082 = ~n5020 & ~n5022;
  assign n5083 = n5013 & n5057;
  assign n5084 = ~n5013 & ~n5057;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = ~n5023 & ~n5082;
  assign n5087 = n5085 & n5086;
  assign n5088 = ~n5081 & ~n5087;
  assign n5089 = n3772 & n5088;
  assign n5090 = ~n5062 & ~n5074;
  assign n5091 = ~n5075 & n5090;
  assign n5092 = ~n5089 & n5091;
  assign n5093 = ~n5016 & ~n5034;
  assign n5094 = ~n5017 & ~n5093;
  assign n5095 = ~n5085 & ~n5094;
  assign n5096 = n5085 & n5094;
  assign n5097 = ~n5095 & ~n5096;
  assign n5098 = n3795 & ~n5097;
  assign n5099 = n3845 & ~n4967;
  assign n5100 = n3790 & n5088;
  assign n5101 = n3793 & ~n5097;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = n3785 & n5088;
  assign n5104 = n3779 & n5088;
  assign n5105 = n3782 & ~n5097;
  assign n5106 = n3788 & ~n5097;
  assign n5107 = ~n5105 & ~n5106;
  assign n5108 = ~n5103 & ~n5104;
  assign n5109 = n5107 & n5108;
  assign n5110 = ~n5098 & ~n5099;
  assign n5111 = n5102 & n5110;
  assign n5112 = n5109 & n5111;
  assign n5113 = n5092 & n5112;
  assign n5114 = n3720_1 & ~n5113;
  assign n5115 = P1_REG0_REG_20_ & ~n3720_1;
  assign n530 = n5114 | n5115;
  assign n5117 = ~n3229 & ~n3727;
  assign n5118 = n5060 & ~n5117;
  assign n5119 = ~n5060 & n5117;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = n3775_1 & n5120;
  assign n5122 = P1_REG1_REG_22_ & n3753;
  assign n5123 = P1_REG0_REG_22_ & n3751;
  assign n5124 = P1_REG2_REG_22_ & n3755_1;
  assign n5125 = P1_REG3_REG_21_ & n5066;
  assign n5126 = ~P1_REG3_REG_22_ & n5125;
  assign n5127 = P1_REG3_REG_22_ & ~n5125;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = n3749 & ~n5128;
  assign n5130 = ~n5122 & ~n5123;
  assign n5131 = ~n5124 & n5130;
  assign n5132 = ~n5129 & n5131;
  assign n5133 = n3742 & ~n5132;
  assign n5134 = ~n3739 & n5117;
  assign n5135 = n5073 & n5117;
  assign n5136 = ~n5073 & ~n5117;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = ~n5020 & n5079;
  assign n5139 = ~n5023 & ~n5057;
  assign n5140 = n5023 & n5057;
  assign n5141 = n5013 & ~n5140;
  assign n5142 = ~n5139 & ~n5141;
  assign n5143 = ~n5138 & ~n5142;
  assign n5144 = ~n5137 & ~n5143;
  assign n5145 = n5137 & ~n5142;
  assign n5146 = ~n5138 & n5145;
  assign n5147 = ~n5144 & ~n5146;
  assign n5148 = n3772 & n5147;
  assign n5149 = ~n5121 & ~n5133;
  assign n5150 = ~n5134 & n5149;
  assign n5151 = ~n5148 & n5150;
  assign n5152 = ~n5083 & ~n5094;
  assign n5153 = ~n5084 & ~n5152;
  assign n5154 = n5137 & n5153;
  assign n5155 = ~n5137 & ~n5153;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = n3795 & ~n5156;
  assign n5158 = n3845 & ~n5013;
  assign n5159 = n3790 & n5147;
  assign n5160 = n3793 & ~n5156;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = n3785 & n5147;
  assign n5163 = n3779 & n5147;
  assign n5164 = n3782 & ~n5156;
  assign n5165 = n3788 & ~n5156;
  assign n5166 = ~n5164 & ~n5165;
  assign n5167 = ~n5162 & ~n5163;
  assign n5168 = n5166 & n5167;
  assign n5169 = ~n5157 & ~n5158;
  assign n5170 = n5161 & n5169;
  assign n5171 = n5168 & n5170;
  assign n5172 = n5151 & n5171;
  assign n5173 = n3720_1 & ~n5172;
  assign n5174 = P1_REG0_REG_21_ & ~n3720_1;
  assign n535 = n5173 | n5174;
  assign n5176 = ~n3266 & ~n3727;
  assign n5177 = ~n5118 & n5176;
  assign n5178 = n5118 & ~n5176;
  assign n5179 = ~n5177 & ~n5178;
  assign n5180 = n3775_1 & n5179;
  assign n5181 = P1_REG1_REG_23_ & n3753;
  assign n5182 = P1_REG0_REG_23_ & n3751;
  assign n5183 = P1_REG2_REG_23_ & n3755_1;
  assign n5184 = P1_REG3_REG_22_ & n5125;
  assign n5185 = ~P1_REG3_REG_23_ & n5184;
  assign n5186 = P1_REG3_REG_23_ & ~n5184;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = n3749 & ~n5187;
  assign n5189 = ~n5181 & ~n5182;
  assign n5190 = ~n5183 & n5189;
  assign n5191 = ~n5188 & n5190;
  assign n5192 = n3742 & ~n5191;
  assign n5193 = ~n3739 & n5176;
  assign n5194 = n5073 & ~n5117;
  assign n5195 = n4947 & n5079;
  assign n5196 = ~n5142 & ~n5195;
  assign n5197 = ~n5194 & ~n5196;
  assign n5198 = ~n5073 & n5117;
  assign n5199 = ~n5197 & ~n5198;
  assign n5200 = ~n4946 & n5079;
  assign n5201 = ~n4941 & ~n5194;
  assign n5202 = n5200 & n5201;
  assign n5203 = n5199 & ~n5202;
  assign n5204 = n5132 & n5176;
  assign n5205 = ~n5132 & ~n5176;
  assign n5206 = ~n5204 & ~n5205;
  assign n5207 = n5203 & ~n5206;
  assign n5208 = ~n5203 & n5206;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n3772 & ~n5209;
  assign n5211 = ~n5180 & ~n5192;
  assign n5212 = ~n5193 & n5211;
  assign n5213 = ~n5210 & n5212;
  assign n5214 = ~n5135 & ~n5153;
  assign n5215 = ~n5136 & ~n5214;
  assign n5216 = n5206 & n5215;
  assign n5217 = ~n5206 & ~n5215;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = n3795 & ~n5218;
  assign n5220 = n3845 & ~n5073;
  assign n5221 = n3790 & ~n5209;
  assign n5222 = n3793 & ~n5218;
  assign n5223 = ~n5221 & ~n5222;
  assign n5224 = n3785 & ~n5209;
  assign n5225 = n3779 & ~n5209;
  assign n5226 = n3782 & ~n5218;
  assign n5227 = n3788 & ~n5218;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = ~n5224 & ~n5225;
  assign n5230 = n5228 & n5229;
  assign n5231 = ~n5219 & ~n5220;
  assign n5232 = n5223 & n5231;
  assign n5233 = n5230 & n5232;
  assign n5234 = n5213 & n5233;
  assign n5235 = n3720_1 & ~n5234;
  assign n5236 = P1_REG0_REG_22_ & ~n3720_1;
  assign n540 = n5235 | n5236;
  assign n5238 = ~n3308 & ~n3727;
  assign n5239 = n5178 & ~n5238;
  assign n5240 = ~n5178 & n5238;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = n3775_1 & n5241;
  assign n5243 = P1_REG1_REG_24_ & n3753;
  assign n5244 = P1_REG0_REG_24_ & n3751;
  assign n5245 = P1_REG2_REG_24_ & n3755_1;
  assign n5246 = P1_REG3_REG_23_ & n5184;
  assign n5247 = ~P1_REG3_REG_24_ & n5246;
  assign n5248 = P1_REG3_REG_24_ & ~n5246;
  assign n5249 = ~n5247 & ~n5248;
  assign n5250 = n3749 & ~n5249;
  assign n5251 = ~n5243 & ~n5244;
  assign n5252 = ~n5245 & n5251;
  assign n5253 = ~n5250 & n5252;
  assign n5254 = n3742 & ~n5253;
  assign n5255 = ~n3739 & n5238;
  assign n5256 = ~n5132 & n5176;
  assign n5257 = n5132 & ~n5176;
  assign n5258 = ~n5203 & ~n5257;
  assign n5259 = ~n5256 & ~n5258;
  assign n5260 = n5191 & n5238;
  assign n5261 = ~n5191 & ~n5238;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = n5259 & ~n5262;
  assign n5264 = ~n5259 & n5262;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = n3772 & ~n5265;
  assign n5267 = ~n5242 & ~n5254;
  assign n5268 = ~n5255 & n5267;
  assign n5269 = ~n5266 & n5268;
  assign n5270 = ~n5204 & ~n5262;
  assign n5271 = ~n5205 & n5215;
  assign n5272 = n5270 & ~n5271;
  assign n5273 = ~n5204 & ~n5215;
  assign n5274 = ~n5205 & ~n5261;
  assign n5275 = ~n5260 & ~n5273;
  assign n5276 = n5274 & n5275;
  assign n5277 = ~n5272 & ~n5276;
  assign n5278 = n3795 & ~n5277;
  assign n5279 = n3845 & ~n5132;
  assign n5280 = n3790 & ~n5265;
  assign n5281 = n3793 & ~n5277;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = n3785 & ~n5265;
  assign n5284 = n3779 & ~n5265;
  assign n5285 = n3782 & ~n5277;
  assign n5286 = n3788 & ~n5277;
  assign n5287 = ~n5285 & ~n5286;
  assign n5288 = ~n5283 & ~n5284;
  assign n5289 = n5287 & n5288;
  assign n5290 = ~n5278 & ~n5279;
  assign n5291 = n5282 & n5290;
  assign n5292 = n5289 & n5291;
  assign n5293 = n5269 & n5292;
  assign n5294 = n3720_1 & ~n5293;
  assign n5295 = P1_REG0_REG_23_ & ~n3720_1;
  assign n545 = n5294 | n5295;
  assign n5297 = ~n3348 & ~n3727;
  assign n5298 = ~n5239 & n5297;
  assign n5299 = n5239 & ~n5297;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = n3775_1 & n5300;
  assign n5302 = P1_REG1_REG_25_ & n3753;
  assign n5303 = P1_REG0_REG_25_ & n3751;
  assign n5304 = P1_REG2_REG_25_ & n3755_1;
  assign n5305 = P1_REG3_REG_24_ & n5246;
  assign n5306 = ~P1_REG3_REG_25_ & n5305;
  assign n5307 = P1_REG3_REG_25_ & ~n5305;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = n3749 & ~n5308;
  assign n5310 = ~n5302 & ~n5303;
  assign n5311 = ~n5304 & n5310;
  assign n5312 = ~n5309 & n5311;
  assign n5313 = n3742 & ~n5312;
  assign n5314 = ~n3739 & n5297;
  assign n5315 = ~n5191 & n5238;
  assign n5316 = n5191 & ~n5238;
  assign n5317 = ~n5259 & ~n5316;
  assign n5318 = ~n5315 & ~n5317;
  assign n5319 = n5253 & n5297;
  assign n5320 = ~n5253 & ~n5297;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = n5318 & ~n5321;
  assign n5323 = n5253 & ~n5297;
  assign n5324 = ~n5253 & n5297;
  assign n5325 = ~n5323 & ~n5324;
  assign n5326 = ~n5318 & ~n5325;
  assign n5327 = ~n5322 & ~n5326;
  assign n5328 = n3772 & ~n5327;
  assign n5329 = ~n5301 & ~n5313;
  assign n5330 = ~n5314 & n5329;
  assign n5331 = ~n5328 & n5330;
  assign n5332 = n5136 & ~n5204;
  assign n5333 = n5274 & ~n5332;
  assign n5334 = ~n5260 & ~n5333;
  assign n5335 = ~n5135 & ~n5204;
  assign n5336 = ~n5153 & n5335;
  assign n5337 = ~n5260 & n5336;
  assign n5338 = ~n5334 & ~n5337;
  assign n5339 = ~n5321 & ~n5338;
  assign n5340 = n5321 & n5338;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = n3795 & ~n5341;
  assign n5343 = n3845 & ~n5191;
  assign n5344 = n3790 & ~n5327;
  assign n5345 = n3793 & ~n5341;
  assign n5346 = ~n5344 & ~n5345;
  assign n5347 = n3785 & ~n5327;
  assign n5348 = n3779 & ~n5327;
  assign n5349 = n3782 & ~n5341;
  assign n5350 = n3788 & ~n5341;
  assign n5351 = ~n5349 & ~n5350;
  assign n5352 = ~n5347 & ~n5348;
  assign n5353 = n5351 & n5352;
  assign n5354 = ~n5342 & ~n5343;
  assign n5355 = n5346 & n5354;
  assign n5356 = n5353 & n5355;
  assign n5357 = n5331 & n5356;
  assign n5358 = n3720_1 & ~n5357;
  assign n5359 = P1_REG0_REG_24_ & ~n3720_1;
  assign n550 = n5358 | n5359;
  assign n5361 = ~n3372 & ~n3727;
  assign n5362 = n5299 & ~n5361;
  assign n5363 = ~n5299 & n5361;
  assign n5364 = ~n5362 & ~n5363;
  assign n5365 = n3775_1 & n5364;
  assign n5366 = P1_REG1_REG_26_ & n3753;
  assign n5367 = P1_REG0_REG_26_ & n3751;
  assign n5368 = P1_REG2_REG_26_ & n3755_1;
  assign n5369 = P1_REG3_REG_25_ & n5305;
  assign n5370 = ~P1_REG3_REG_26_ & n5369;
  assign n5371 = P1_REG3_REG_26_ & ~n5369;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = n3749 & ~n5372;
  assign n5374 = ~n5366 & ~n5367;
  assign n5375 = ~n5368 & n5374;
  assign n5376 = ~n5373 & n5375;
  assign n5377 = n3742 & ~n5376;
  assign n5378 = ~n3739 & n5361;
  assign n5379 = n5312 & n5361;
  assign n5380 = ~n5312 & ~n5361;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = ~n5318 & ~n5323;
  assign n5383 = ~n5324 & ~n5382;
  assign n5384 = ~n5381 & n5383;
  assign n5385 = n5312 & ~n5361;
  assign n5386 = ~n5312 & n5361;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = ~n5383 & ~n5387;
  assign n5389 = ~n5384 & ~n5388;
  assign n5390 = n3772 & ~n5389;
  assign n5391 = ~n5365 & ~n5377;
  assign n5392 = ~n5378 & n5391;
  assign n5393 = ~n5390 & n5392;
  assign n5394 = ~n5319 & ~n5338;
  assign n5395 = ~n5320 & ~n5394;
  assign n5396 = ~n5381 & ~n5395;
  assign n5397 = n5381 & n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = n3795 & ~n5398;
  assign n5400 = n3845 & ~n5253;
  assign n5401 = n3790 & ~n5389;
  assign n5402 = n3793 & ~n5398;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = n3785 & ~n5389;
  assign n5405 = n3779 & ~n5389;
  assign n5406 = n3782 & ~n5398;
  assign n5407 = n3788 & ~n5398;
  assign n5408 = ~n5406 & ~n5407;
  assign n5409 = ~n5404 & ~n5405;
  assign n5410 = n5408 & n5409;
  assign n5411 = ~n5399 & ~n5400;
  assign n5412 = n5403 & n5411;
  assign n5413 = n5410 & n5412;
  assign n5414 = n5393 & n5413;
  assign n5415 = n3720_1 & ~n5414;
  assign n5416 = P1_REG0_REG_25_ & ~n3720_1;
  assign n555 = n5415 | n5416;
  assign n5418 = ~n3415_1 & ~n3727;
  assign n5419 = ~n5362 & n5418;
  assign n5420 = n5362 & ~n5418;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = n3775_1 & n5421;
  assign n5423 = P1_REG1_REG_27_ & n3753;
  assign n5424 = P1_REG0_REG_27_ & n3751;
  assign n5425 = P1_REG2_REG_27_ & n3755_1;
  assign n5426 = P1_REG3_REG_26_ & n5369;
  assign n5427 = ~P1_REG3_REG_27_ & n5426;
  assign n5428 = P1_REG3_REG_27_ & ~n5426;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = n3749 & ~n5429;
  assign n5431 = ~n5423 & ~n5424;
  assign n5432 = ~n5425 & n5431;
  assign n5433 = ~n5430 & n5432;
  assign n5434 = n3742 & ~n5433;
  assign n5435 = ~n3739 & n5418;
  assign n5436 = n5383 & ~n5386;
  assign n5437 = ~n5376 & n5418;
  assign n5438 = ~n5385 & n5418;
  assign n5439 = ~n5376 & ~n5385;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = ~n5436 & ~n5437;
  assign n5442 = ~n5440 & n5441;
  assign n5443 = ~n5383 & ~n5385;
  assign n5444 = n5376 & n5418;
  assign n5445 = ~n5376 & ~n5418;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = ~n5386 & ~n5443;
  assign n5448 = n5446 & n5447;
  assign n5449 = ~n5442 & ~n5448;
  assign n5450 = n3772 & n5449;
  assign n5451 = ~n5422 & ~n5434;
  assign n5452 = ~n5435 & n5451;
  assign n5453 = ~n5450 & n5452;
  assign n5454 = ~n5379 & ~n5395;
  assign n5455 = ~n5380 & ~n5454;
  assign n5456 = n5446 & n5455;
  assign n5457 = ~n5446 & ~n5455;
  assign n5458 = ~n5456 & ~n5457;
  assign n5459 = n3795 & ~n5458;
  assign n5460 = n3845 & ~n5312;
  assign n5461 = n3790 & n5449;
  assign n5462 = n3793 & ~n5458;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = n3785 & n5449;
  assign n5465 = n3779 & n5449;
  assign n5466 = n3782 & ~n5458;
  assign n5467 = n3788 & ~n5458;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = ~n5464 & ~n5465;
  assign n5470 = n5468 & n5469;
  assign n5471 = ~n5459 & ~n5460;
  assign n5472 = n5463 & n5471;
  assign n5473 = n5470 & n5472;
  assign n5474 = n5453 & n5473;
  assign n5475 = n3720_1 & ~n5474;
  assign n5476 = P1_REG0_REG_26_ & ~n3720_1;
  assign n560 = n5475 | n5476;
  assign n5478 = ~n3439 & ~n3727;
  assign n5479 = n5420 & ~n5478;
  assign n5480 = ~n5420 & n5478;
  assign n5481 = ~n5479 & ~n5480;
  assign n5482 = n3775_1 & n5481;
  assign n5483 = P1_REG1_REG_28_ & n3753;
  assign n5484 = P1_REG0_REG_28_ & n3751;
  assign n5485 = P1_REG2_REG_28_ & n3755_1;
  assign n5486 = P1_REG3_REG_27_ & n5426;
  assign n5487 = ~P1_REG3_REG_28_ & n5486;
  assign n5488 = P1_REG3_REG_28_ & ~n5486;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = n3749 & ~n5489;
  assign n5491 = ~n5483 & ~n5484;
  assign n5492 = ~n5485 & n5491;
  assign n5493 = ~n5490 & n5492;
  assign n5494 = n3742 & ~n5493;
  assign n5495 = ~n3739 & n5478;
  assign n5496 = ~n5324 & ~n5386;
  assign n5497 = ~n5440 & ~n5496;
  assign n5498 = n5382 & ~n5440;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = ~n5437 & n5499;
  assign n5501 = n5433 & n5478;
  assign n5502 = ~n5433 & ~n5478;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = n5500 & ~n5503;
  assign n5505 = ~n5500 & n5503;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = n3772 & ~n5506;
  assign n5508 = ~n5482 & ~n5494;
  assign n5509 = ~n5495 & n5508;
  assign n5510 = ~n5507 & n5509;
  assign n5511 = ~n5444 & ~n5503;
  assign n5512 = ~n5445 & n5455;
  assign n5513 = n5511 & ~n5512;
  assign n5514 = ~n5445 & n5503;
  assign n5515 = ~n5444 & ~n5455;
  assign n5516 = n5514 & ~n5515;
  assign n5517 = ~n5513 & ~n5516;
  assign n5518 = n3795 & ~n5517;
  assign n5519 = n3845 & ~n5376;
  assign n5520 = n3790 & ~n5506;
  assign n5521 = n3793 & ~n5517;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = n3785 & ~n5506;
  assign n5524 = n3779 & ~n5506;
  assign n5525 = n3782 & ~n5517;
  assign n5526 = n3788 & ~n5517;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = ~n5523 & ~n5524;
  assign n5529 = n5527 & n5528;
  assign n5530 = ~n5518 & ~n5519;
  assign n5531 = n5522 & n5530;
  assign n5532 = n5529 & n5531;
  assign n5533 = n5510 & n5532;
  assign n5534 = n3720_1 & ~n5533;
  assign n5535 = P1_REG0_REG_27_ & ~n3720_1;
  assign n565 = n5534 | n5535;
  assign n5537 = ~n3484 & ~n3727;
  assign n5538 = ~n5479 & n5537;
  assign n5539 = n5479 & ~n5537;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = n3775_1 & n5540;
  assign n5542 = P1_REG0_REG_29_ & n3751;
  assign n5543 = P1_REG1_REG_29_ & n3753;
  assign n5544 = P1_REG2_REG_29_ & n3755_1;
  assign n5545 = P1_REG3_REG_28_ & P1_REG3_REG_27_;
  assign n5546 = n5426 & n5545;
  assign n5547 = n3749 & n5546;
  assign n5548 = ~n5542 & ~n5543;
  assign n5549 = ~n5544 & n5548;
  assign n5550 = ~n5547 & n5549;
  assign n5551 = n3742 & ~n5550;
  assign n5552 = ~n3739 & n5537;
  assign n5553 = n5433 & ~n5478;
  assign n5554 = n5437 & ~n5553;
  assign n5555 = ~n5323 & ~n5553;
  assign n5556 = ~n5318 & ~n5440;
  assign n5557 = n5555 & n5556;
  assign n5558 = n5497 & ~n5553;
  assign n5559 = ~n5433 & n5478;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = ~n5554 & ~n5557;
  assign n5562 = n5560 & n5561;
  assign n5563 = n5493 & n5537;
  assign n5564 = ~n5493 & ~n5537;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = n5562 & ~n5565;
  assign n5567 = ~n5562 & n5565;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = n3772 & ~n5568;
  assign n5570 = ~n5541 & ~n5551;
  assign n5571 = ~n5552 & n5570;
  assign n5572 = ~n5569 & n5571;
  assign n5573 = n5433 & ~n5445;
  assign n5574 = ~n5478 & ~n5573;
  assign n5575 = ~n5433 & n5445;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = ~n5501 & n5515;
  assign n5578 = n5576 & ~n5577;
  assign n5579 = ~n5565 & ~n5578;
  assign n5580 = n5565 & n5578;
  assign n5581 = ~n5579 & ~n5580;
  assign n5582 = n3795 & ~n5581;
  assign n5583 = n3845 & ~n5433;
  assign n5584 = n3790 & ~n5568;
  assign n5585 = n3793 & ~n5581;
  assign n5586 = ~n5584 & ~n5585;
  assign n5587 = n3785 & ~n5568;
  assign n5588 = n3779 & ~n5568;
  assign n5589 = n3782 & ~n5581;
  assign n5590 = n3788 & ~n5581;
  assign n5591 = ~n5589 & ~n5590;
  assign n5592 = ~n5587 & ~n5588;
  assign n5593 = n5591 & n5592;
  assign n5594 = ~n5582 & ~n5583;
  assign n5595 = n5586 & n5594;
  assign n5596 = n5593 & n5595;
  assign n5597 = n5572 & n5596;
  assign n5598 = n3720_1 & ~n5597;
  assign n5599 = P1_REG0_REG_28_ & ~n3720_1;
  assign n570 = n5598 | n5599;
  assign n5601 = ~n3513 & ~n3727;
  assign n5602 = n5539 & ~n5601;
  assign n5603 = ~n5539 & n5601;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = n3775_1 & n5604;
  assign n5606 = ~n3739 & n5601;
  assign n5607 = n5537 & ~n5562;
  assign n5608 = ~n5493 & ~n5562;
  assign n5609 = ~n5493 & n5537;
  assign n5610 = ~n5607 & ~n5608;
  assign n5611 = ~n5609 & n5610;
  assign n5612 = n5550 & n5601;
  assign n5613 = ~n5550 & ~n5601;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = n5611 & ~n5614;
  assign n5616 = ~n5611 & n5614;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = n3772 & ~n5617;
  assign n5619 = ~n5605 & ~n5606;
  assign n5620 = ~n5618 & n5619;
  assign n5621 = n3785 & ~n5617;
  assign n5622 = n3779 & ~n5617;
  assign n5623 = n5493 & n5614;
  assign n5624 = n5537 & n5623;
  assign n5625 = ~n5493 & ~n5614;
  assign n5626 = ~n5537 & n5625;
  assign n5627 = ~n5624 & ~n5626;
  assign n5628 = ~n5563 & ~n5614;
  assign n5629 = ~n5578 & n5628;
  assign n5630 = ~n5564 & n5576;
  assign n5631 = ~n5577 & n5614;
  assign n5632 = n5630 & n5631;
  assign n5633 = n5627 & ~n5629;
  assign n5634 = ~n5632 & n5633;
  assign n5635 = n3782 & ~n5634;
  assign n5636 = n3788 & ~n5634;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = ~n5621 & ~n5622;
  assign n5639 = n5637 & n5638;
  assign n5640 = n3845 & ~n5493;
  assign n5641 = ~P1_B_REG & n3726;
  assign n5642 = ~n3727 & ~n5641;
  assign n5643 = n3741 & ~n5642;
  assign n5644 = P1_REG1_REG_30_ & n3753;
  assign n5645 = P1_REG0_REG_30_ & n3751;
  assign n5646 = P1_REG2_REG_30_ & n3755_1;
  assign n5647 = ~n5644 & ~n5645;
  assign n5648 = ~n5646 & n5647;
  assign n5649 = n5643 & ~n5648;
  assign n5650 = n3795 & ~n5634;
  assign n5651 = n3793 & ~n5634;
  assign n5652 = n3790 & ~n5617;
  assign n5653 = ~n5640 & ~n5649;
  assign n5654 = ~n5650 & n5653;
  assign n5655 = ~n5651 & n5654;
  assign n5656 = ~n5652 & n5655;
  assign n5657 = n5639 & n5656;
  assign n5658 = n5620 & n5657;
  assign n5659 = n3720_1 & ~n5658;
  assign n5660 = P1_REG0_REG_29_ & ~n3720_1;
  assign n575 = n5659 | n5660;
  assign n5662 = ~n3537 & ~n3727;
  assign n5663 = ~n3739 & n5662;
  assign n5664 = P1_REG1_REG_31_ & n3753;
  assign n5665 = P1_REG0_REG_31_ & n3751;
  assign n5666 = P1_REG2_REG_31_ & n3755_1;
  assign n5667 = ~n5664 & ~n5665;
  assign n5668 = ~n5666 & n5667;
  assign n5669 = n5643 & ~n5668;
  assign n5670 = ~n5602 & n5662;
  assign n5671 = n5602 & ~n5662;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = n3775_1 & n5672;
  assign n5674 = ~n5663 & ~n5669;
  assign n5675 = ~n5673 & n5674;
  assign n5676 = n3720_1 & ~n5675;
  assign n5677 = P1_REG0_REG_30_ & ~n3720_1;
  assign n580 = n5676 | n5677;
  assign n5679 = ~n3568 & ~n3727;
  assign n5680 = ~n3739 & n5679;
  assign n5681 = n5671 & ~n5679;
  assign n5682 = ~n5671 & n5679;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = n3775_1 & n5683;
  assign n5685 = ~n5669 & ~n5680;
  assign n5686 = ~n5684 & n5685;
  assign n5687 = n3720_1 & ~n5686;
  assign n5688 = P1_REG0_REG_31_ & ~n3720_1;
  assign n585 = n5687 | n5688;
  assign n5690 = n3587 & ~n3636;
  assign n5691 = n3719 & n5690;
  assign n5692 = ~n3804 & n5691;
  assign n5693 = P1_REG1_REG_0_ & ~n5691;
  assign n590 = n5692 | n5693;
  assign n5695 = ~n3860 & n5691;
  assign n5696 = P1_REG1_REG_1_ & ~n5691;
  assign n595 = n5695 | n5696;
  assign n5698 = ~n3922 & n5691;
  assign n5699 = P1_REG1_REG_2_ & ~n5691;
  assign n600 = n5698 | n5699;
  assign n5701 = ~n3987 & n5691;
  assign n5702 = P1_REG1_REG_3_ & ~n5691;
  assign n605 = n5701 | n5702;
  assign n5704 = ~n4057 & n5691;
  assign n5705 = P1_REG1_REG_4_ & ~n5691;
  assign n610 = n5704 | n5705;
  assign n5707 = ~n4121 & n5691;
  assign n5708 = P1_REG1_REG_5_ & ~n5691;
  assign n615 = n5707 | n5708;
  assign n5710 = ~n4195 & n5691;
  assign n5711 = P1_REG1_REG_6_ & ~n5691;
  assign n620 = n5710 | n5711;
  assign n5713 = ~n4263 & n5691;
  assign n5714 = P1_REG1_REG_7_ & ~n5691;
  assign n625 = n5713 | n5714;
  assign n5716 = ~n4331 & n5691;
  assign n5717 = P1_REG1_REG_8_ & ~n5691;
  assign n630 = n5716 | n5717;
  assign n5719 = ~n4398 & n5691;
  assign n5720 = P1_REG1_REG_9_ & ~n5691;
  assign n635 = n5719 | n5720;
  assign n5722 = ~n4463 & n5691;
  assign n5723 = P1_REG1_REG_10_ & ~n5691;
  assign n640 = n5722 | n5723;
  assign n5725 = ~n4533 & n5691;
  assign n5726 = P1_REG1_REG_11_ & ~n5691;
  assign n645 = n5725 | n5726;
  assign n5728 = ~n4600 & n5691;
  assign n5729 = P1_REG1_REG_12_ & ~n5691;
  assign n650 = n5728 | n5729;
  assign n5731 = ~n4664 & n5691;
  assign n5732 = P1_REG1_REG_13_ & ~n5691;
  assign n655 = n5731 | n5732;
  assign n5734 = ~n4728 & n5691;
  assign n5735 = P1_REG1_REG_14_ & ~n5691;
  assign n660 = n5734 | n5735;
  assign n5737 = ~n4789 & n5691;
  assign n5738 = P1_REG1_REG_15_ & ~n5691;
  assign n665 = n5737 | n5738;
  assign n5740 = ~n4856 & n5691;
  assign n5741 = P1_REG1_REG_16_ & ~n5691;
  assign n670 = n5740 | n5741;
  assign n5743 = ~n4925 & n5691;
  assign n5744 = P1_REG1_REG_17_ & ~n5691;
  assign n675 = n5743 | n5744;
  assign n5746 = ~n4992 & n5691;
  assign n5747 = P1_REG1_REG_18_ & ~n5691;
  assign n680 = n5746 | n5747;
  assign n5749 = ~n5053 & n5691;
  assign n5750 = P1_REG1_REG_19_ & ~n5691;
  assign n685 = n5749 | n5750;
  assign n5752 = ~n5113 & n5691;
  assign n5753 = P1_REG1_REG_20_ & ~n5691;
  assign n690 = n5752 | n5753;
  assign n5755 = ~n5172 & n5691;
  assign n5756 = P1_REG1_REG_21_ & ~n5691;
  assign n695 = n5755 | n5756;
  assign n5758 = ~n5234 & n5691;
  assign n5759 = P1_REG1_REG_22_ & ~n5691;
  assign n700 = n5758 | n5759;
  assign n5761 = ~n5293 & n5691;
  assign n5762 = P1_REG1_REG_23_ & ~n5691;
  assign n705 = n5761 | n5762;
  assign n5764 = ~n5357 & n5691;
  assign n5765 = P1_REG1_REG_24_ & ~n5691;
  assign n710 = n5764 | n5765;
  assign n5767 = ~n5414 & n5691;
  assign n5768 = P1_REG1_REG_25_ & ~n5691;
  assign n715 = n5767 | n5768;
  assign n5770 = ~n5474 & n5691;
  assign n5771 = P1_REG1_REG_26_ & ~n5691;
  assign n720 = n5770 | n5771;
  assign n5773 = ~n5533 & n5691;
  assign n5774 = P1_REG1_REG_27_ & ~n5691;
  assign n725 = n5773 | n5774;
  assign n5776 = ~n5597 & n5691;
  assign n5777 = P1_REG1_REG_28_ & ~n5691;
  assign n730 = n5776 | n5777;
  assign n5779 = ~n5658 & n5691;
  assign n5780 = P1_REG1_REG_29_ & ~n5691;
  assign n735 = n5779 | n5780;
  assign n5782 = ~n5675 & n5691;
  assign n5783 = P1_REG1_REG_30_ & ~n5691;
  assign n740 = n5782 | n5783;
  assign n5785 = ~n5686 & n5691;
  assign n5786 = P1_REG1_REG_31_ & ~n5691;
  assign n745 = n5785 | n5786;
  assign n5788 = n3649 & n3737;
  assign n5789 = n3649 & n3735_1;
  assign n5790 = ~n3656 & n3741;
  assign n5791 = n3636 & ~n5790;
  assign n5792 = ~n3640_1 & n5791;
  assign n5793 = n3718 & n5792;
  assign n5794 = ~n5789 & ~n5793;
  assign n5795 = n3587 & ~n5794;
  assign n5796 = n5788 & n5795;
  assign n5797 = ~n3733 & n5796;
  assign n5798 = n3643 & n3787;
  assign n5799 = n3646 & n5798;
  assign n5800 = ~n3738 & ~n5799;
  assign n5801 = n5795 & ~n5800;
  assign n5802 = ~n3733 & n5801;
  assign n5803 = ~n3801 & n5795;
  assign n5804 = P1_REG2_REG_0_ & ~n5795;
  assign n5805 = ~n5803 & ~n5804;
  assign n5806 = ~n5797 & ~n5802;
  assign n5807 = n5805 & n5806;
  assign n5808 = n5789 & n5795;
  assign n5809 = P1_REG3_REG_0_ & n5808;
  assign n5810 = n3742 & n5795;
  assign n5811 = ~n3759 & n5810;
  assign n5812 = ~n3646 & n3771;
  assign n5813 = n5795 & n5812;
  assign n5814 = ~n3770_1 & n5813;
  assign n5815 = ~n5809 & ~n5811;
  assign n5816 = ~n5814 & n5815;
  assign n750 = ~n5807 | ~n5816;
  assign n5818 = ~n3816 & n5796;
  assign n5819 = ~n3813 & n5801;
  assign n5820 = ~n3859 & n5795;
  assign n5821 = P1_REG2_REG_1_ & ~n5795;
  assign n5822 = ~n5820 & ~n5821;
  assign n5823 = ~n5818 & ~n5819;
  assign n5824 = n5822 & n5823;
  assign n5825 = P1_REG3_REG_1_ & n5808;
  assign n5826 = ~n3824 & n5810;
  assign n5827 = ~n3833 & n5813;
  assign n5828 = ~n5825 & ~n5826;
  assign n5829 = ~n5827 & n5828;
  assign n755 = ~n5824 | ~n5829;
  assign n5831 = n3873 & n5796;
  assign n5832 = ~n3869 & n5801;
  assign n5833 = ~n3921 & n5795;
  assign n5834 = P1_REG2_REG_2_ & ~n5795;
  assign n5835 = ~n5833 & ~n5834;
  assign n5836 = ~n5831 & ~n5832;
  assign n5837 = n5835 & n5836;
  assign n5838 = P1_REG3_REG_2_ & n5808;
  assign n5839 = ~n3881 & n5810;
  assign n5840 = n3895 & n5813;
  assign n5841 = ~n5838 & ~n5839;
  assign n5842 = ~n5840 & n5841;
  assign n760 = ~n5837 | ~n5842;
  assign n5844 = n3934 & n5796;
  assign n5845 = ~n3931 & n5801;
  assign n5846 = ~n3986 & n5795;
  assign n5847 = P1_REG2_REG_3_ & ~n5795;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = ~n5844 & ~n5845;
  assign n5850 = n5848 & n5849;
  assign n5851 = ~P1_REG3_REG_3_ & n5808;
  assign n5852 = ~n3945 & n5810;
  assign n5853 = ~n3960 & n5813;
  assign n5854 = ~n5851 & ~n5852;
  assign n5855 = ~n5853 & n5854;
  assign n765 = ~n5850 | ~n5855;
  assign n5857 = n3999 & n5796;
  assign n5858 = ~n3996 & n5801;
  assign n5859 = ~n4056 & n5795;
  assign n5860 = P1_REG2_REG_4_ & ~n5795;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = ~n5857 & ~n5858;
  assign n5863 = n5861 & n5862;
  assign n5864 = ~n3938 & n5808;
  assign n5865 = ~n4011 & n5810;
  assign n5866 = ~n4027 & n5813;
  assign n5867 = ~n5864 & ~n5865;
  assign n5868 = ~n5866 & n5867;
  assign n770 = ~n5863 | ~n5868;
  assign n5870 = n4069 & n5796;
  assign n5871 = ~n4066 & n5801;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = ~n4004 & n5808;
  assign n5874 = ~n4081 & n5810;
  assign n5875 = n4096 & n5813;
  assign n5876 = ~n5873 & ~n5874;
  assign n5877 = ~n5875 & n5876;
  assign n5878 = ~n4120 & n5795;
  assign n5879 = P1_REG2_REG_5_ & ~n5795;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = n5872 & n5877;
  assign n775 = ~n5880 | ~n5881;
  assign n5883 = n4134 & n5796;
  assign n5884 = ~n4130 & n5801;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = ~n4074 & n5808;
  assign n5887 = ~n4146 & n5810;
  assign n5888 = ~n4167 & n5813;
  assign n5889 = ~n5886 & ~n5887;
  assign n5890 = ~n5888 & n5889;
  assign n5891 = ~n4194 & n5795;
  assign n5892 = P1_REG2_REG_6_ & ~n5795;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = n5885 & n5890;
  assign n780 = ~n5893 | ~n5894;
  assign n5896 = n4207 & n5796;
  assign n5897 = ~n4204 & n5801;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = ~n4139 & n5808;
  assign n5900 = ~n4219 & n5810;
  assign n5901 = n4234 & n5813;
  assign n5902 = ~n5899 & ~n5900;
  assign n5903 = ~n5901 & n5902;
  assign n5904 = ~n4262 & n5795;
  assign n5905 = P1_REG2_REG_7_ & ~n5795;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = n5898 & n5903;
  assign n785 = ~n5906 | ~n5907;
  assign n5909 = n4275 & n5796;
  assign n5910 = ~n4272 & n5801;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = ~n4212 & n5808;
  assign n5913 = ~n4287 & n5810;
  assign n5914 = ~n4304 & n5813;
  assign n5915 = ~n5912 & ~n5913;
  assign n5916 = ~n5914 & n5915;
  assign n5917 = ~n4330 & n5795;
  assign n5918 = P1_REG2_REG_8_ & ~n5795;
  assign n5919 = ~n5917 & ~n5918;
  assign n5920 = n5911 & n5916;
  assign n790 = ~n5919 | ~n5920;
  assign n5922 = ~n4283 & n5808;
  assign n5923 = ~n4355 & n5810;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = n4343 & n5796;
  assign n5926 = ~n4340 & n5801;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n4368 & n5813;
  assign n5929 = ~n4397 & n5795;
  assign n5930 = P1_REG2_REG_9_ & ~n5795;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = n5924 & n5927;
  assign n5933 = ~n5928 & n5932;
  assign n795 = ~n5931 | ~n5933;
  assign n5935 = ~n4351 & n5808;
  assign n5936 = ~n4423 & n5810;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = n4411 & n5796;
  assign n5939 = ~n4407 & n5801;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = n4438 & n5813;
  assign n5942 = ~n4462 & n5795;
  assign n5943 = P1_REG2_REG_10_ & ~n5795;
  assign n5944 = ~n5942 & ~n5943;
  assign n5945 = n5937 & n5940;
  assign n5946 = ~n5941 & n5945;
  assign n800 = ~n5944 | ~n5946;
  assign n5948 = n4476 & n5796;
  assign n5949 = ~n4472 & n5801;
  assign n5950 = ~n5948 & ~n5949;
  assign n5951 = ~n4419 & n5808;
  assign n5952 = ~n4505 & n5810;
  assign n5953 = ~n4493 & n5813;
  assign n5954 = ~n5951 & ~n5952;
  assign n5955 = ~n5953 & n5954;
  assign n5956 = ~n4532 & n5795;
  assign n5957 = P1_REG2_REG_11_ & ~n5795;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = n5950 & n5955;
  assign n805 = ~n5958 | ~n5959;
  assign n5961 = n4558 & n5796;
  assign n5962 = ~n4542 & n5801;
  assign n5963 = ~n5961 & ~n5962;
  assign n5964 = ~n4501 & n5808;
  assign n5965 = ~n4570 & n5810;
  assign n5966 = ~n4554 & n5813;
  assign n5967 = ~n5964 & ~n5965;
  assign n5968 = ~n5966 & n5967;
  assign n5969 = ~n4599 & n5795;
  assign n5970 = P1_REG2_REG_12_ & ~n5795;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = n5963 & n5968;
  assign n810 = ~n5971 | ~n5972;
  assign n5974 = n4613 & n5796;
  assign n5975 = ~n4609 & n5801;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~n4566 & n5808;
  assign n5978 = ~n4639 & n5810;
  assign n5979 = n4627 & n5813;
  assign n5980 = ~n5977 & ~n5978;
  assign n5981 = ~n5979 & n5980;
  assign n5982 = ~n4663 & n5795;
  assign n5983 = P1_REG2_REG_13_ & ~n5795;
  assign n5984 = ~n5982 & ~n5983;
  assign n5985 = n5976 & n5981;
  assign n815 = ~n5984 | ~n5985;
  assign n5987 = n4691 & n5796;
  assign n5988 = ~n4673 & n5801;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = ~n4635 & n5808;
  assign n5991 = ~n4703 & n5810;
  assign n5992 = ~n4686 & n5813;
  assign n5993 = ~n5990 & ~n5991;
  assign n5994 = ~n5992 & n5993;
  assign n5995 = ~n4727 & n5795;
  assign n5996 = P1_REG2_REG_14_ & ~n5795;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = n5989 & n5994;
  assign n820 = ~n5997 | ~n5998;
  assign n6000 = ~n4699 & n5808;
  assign n6001 = ~n4752 & n5810;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = n4740 & n5796;
  assign n6004 = ~n4737 & n5801;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = ~n4764 & n5813;
  assign n6007 = ~n4788 & n5795;
  assign n6008 = P1_REG2_REG_15_ & ~n5795;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = n6002 & n6005;
  assign n6011 = ~n6006 & n6010;
  assign n825 = ~n6009 | ~n6011;
  assign n6013 = ~n4748 & n5808;
  assign n6014 = ~n4813 & n5810;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = n4801 & n5796;
  assign n6017 = ~n4798 & n5801;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019 = ~n4828 & n5813;
  assign n6020 = ~n4855 & n5795;
  assign n6021 = P1_REG2_REG_16_ & ~n5795;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = n6015 & n6018;
  assign n6024 = ~n6019 & n6023;
  assign n830 = ~n6022 | ~n6024;
  assign n6026 = n4883 & n5796;
  assign n6027 = ~n4865 & n5801;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = ~n4809 & n5808;
  assign n6030 = ~n4895 & n5810;
  assign n6031 = n4879 & n5813;
  assign n6032 = ~n6029 & ~n6030;
  assign n6033 = ~n6031 & n6032;
  assign n6034 = ~n4924 & n5795;
  assign n6035 = P1_REG2_REG_17_ & ~n5795;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = n6028 & n6033;
  assign n835 = ~n6036 | ~n6037;
  assign n6039 = n4955 & n5796;
  assign n6040 = ~n4934 & n5801;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = ~n4891 & n5808;
  assign n6043 = ~n4967 & n5810;
  assign n6044 = ~n4950 & n5813;
  assign n6045 = ~n6042 & ~n6043;
  assign n6046 = ~n6044 & n6045;
  assign n6047 = ~n4991 & n5795;
  assign n6048 = P1_REG2_REG_18_ & ~n5795;
  assign n6049 = ~n6047 & ~n6048;
  assign n6050 = n6041 & n6046;
  assign n840 = ~n6049 | ~n6050;
  assign n6052 = ~n4963 & n5808;
  assign n6053 = ~n5013 & n5810;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = n5001 & n5796;
  assign n6056 = ~n4998 & n5801;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n5026 & n5813;
  assign n6059 = ~n5052 & n5795;
  assign n6060 = P1_REG2_REG_19_ & ~n5795;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = n6054 & n6057;
  assign n6063 = ~n6058 & n6062;
  assign n845 = ~n6061 | ~n6063;
  assign n6065 = ~n5009 & n5808;
  assign n6066 = ~n5073 & n5810;
  assign n6067 = ~n6065 & ~n6066;
  assign n6068 = n5061 & n5796;
  assign n6069 = n5057 & n5801;
  assign n6070 = ~n6068 & ~n6069;
  assign n6071 = n5088 & n5813;
  assign n6072 = ~n5112 & n5795;
  assign n6073 = P1_REG2_REG_20_ & ~n5795;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = n6067 & n6070;
  assign n6076 = ~n6071 & n6075;
  assign n850 = ~n6074 | ~n6076;
  assign n6078 = ~n5069 & n5808;
  assign n6079 = ~n5132 & n5810;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = n5120 & n5796;
  assign n6082 = n5117 & n5801;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = n5147 & n5813;
  assign n6085 = ~n5171 & n5795;
  assign n6086 = P1_REG2_REG_21_ & ~n5795;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = n6080 & n6083;
  assign n6089 = ~n6084 & n6088;
  assign n855 = ~n6087 | ~n6089;
  assign n6091 = ~n5128 & n5808;
  assign n6092 = ~n5191 & n5810;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = n5179 & n5796;
  assign n6095 = n5176 & n5801;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n5209 & n5813;
  assign n6098 = ~n5233 & n5795;
  assign n6099 = P1_REG2_REG_22_ & ~n5795;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = n6093 & n6096;
  assign n6102 = ~n6097 & n6101;
  assign n860 = ~n6100 | ~n6102;
  assign n6104 = ~n5187 & n5808;
  assign n6105 = ~n5253 & n5810;
  assign n6106 = ~n6104 & ~n6105;
  assign n6107 = n5241 & n5796;
  assign n6108 = n5238 & n5801;
  assign n6109 = ~n6107 & ~n6108;
  assign n6110 = ~n5265 & n5813;
  assign n6111 = ~n5292 & n5795;
  assign n6112 = P1_REG2_REG_23_ & ~n5795;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = n6106 & n6109;
  assign n6115 = ~n6110 & n6114;
  assign n865 = ~n6113 | ~n6115;
  assign n6117 = ~n5249 & n5808;
  assign n6118 = ~n5312 & n5810;
  assign n6119 = ~n6117 & ~n6118;
  assign n6120 = n5300 & n5796;
  assign n6121 = n5297 & n5801;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = ~n5327 & n5813;
  assign n6124 = ~n5356 & n5795;
  assign n6125 = P1_REG2_REG_24_ & ~n5795;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = n6119 & n6122;
  assign n6128 = ~n6123 & n6127;
  assign n870 = ~n6126 | ~n6128;
  assign n6130 = ~n5308 & n5808;
  assign n6131 = ~n5376 & n5810;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = n5364 & n5796;
  assign n6134 = n5361 & n5801;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = ~n5389 & n5813;
  assign n6137 = ~n5413 & n5795;
  assign n6138 = P1_REG2_REG_25_ & ~n5795;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = n6132 & n6135;
  assign n6141 = ~n6136 & n6140;
  assign n875 = ~n6139 | ~n6141;
  assign n6143 = ~n5372 & n5808;
  assign n6144 = ~n5433 & n5810;
  assign n6145 = ~n6143 & ~n6144;
  assign n6146 = n5421 & n5796;
  assign n6147 = n5418 & n5801;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = n5449 & n5813;
  assign n6150 = ~n5473 & n5795;
  assign n6151 = P1_REG2_REG_26_ & ~n5795;
  assign n6152 = ~n6150 & ~n6151;
  assign n6153 = n6145 & n6148;
  assign n6154 = ~n6149 & n6153;
  assign n880 = ~n6152 | ~n6154;
  assign n6156 = ~n5429 & n5808;
  assign n6157 = ~n5493 & n5810;
  assign n6158 = ~n6156 & ~n6157;
  assign n6159 = n5481 & n5796;
  assign n6160 = n5478 & n5801;
  assign n6161 = ~n6159 & ~n6160;
  assign n6162 = ~n5506 & n5813;
  assign n6163 = ~n5532 & n5795;
  assign n6164 = P1_REG2_REG_27_ & ~n5795;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = n6158 & n6161;
  assign n6167 = ~n6162 & n6166;
  assign n885 = ~n6165 | ~n6167;
  assign n6169 = ~n5489 & n5808;
  assign n6170 = ~n5550 & n5810;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = n5540 & n5796;
  assign n6173 = n5537 & n5801;
  assign n6174 = ~n6172 & ~n6173;
  assign n6175 = ~n5568 & n5813;
  assign n6176 = ~n5596 & n5795;
  assign n6177 = P1_REG2_REG_28_ & ~n5795;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = n6171 & n6174;
  assign n6180 = ~n6175 & n6179;
  assign n890 = ~n6178 | ~n6180;
  assign n6182 = n5601 & n5801;
  assign n6183 = n5546 & n5808;
  assign n6184 = n5604 & n5796;
  assign n6185 = ~n5617 & n5813;
  assign n6186 = ~n5657 & n5795;
  assign n6187 = P1_REG2_REG_29_ & ~n5795;
  assign n6188 = ~n6186 & ~n6187;
  assign n6189 = ~n6182 & ~n6183;
  assign n6190 = ~n6184 & n6189;
  assign n6191 = ~n6185 & n6190;
  assign n895 = ~n6188 | ~n6191;
  assign n6193 = n5669 & n5795;
  assign n6194 = P1_REG2_REG_30_ & ~n5795;
  assign n6195 = ~n6193 & ~n6194;
  assign n6196 = n5662 & n5801;
  assign n6197 = n5672 & n5796;
  assign n6198 = n6195 & ~n6196;
  assign n900 = n6197 | ~n6198;
  assign n6200 = P1_REG2_REG_31_ & ~n5795;
  assign n6201 = ~n6193 & ~n6200;
  assign n6202 = n5679 & n5801;
  assign n6203 = n5683 & n5796;
  assign n6204 = n6201 & ~n6202;
  assign n905 = n6203 | ~n6204;
  assign n6206 = P1_STATE_REG & ~n3574;
  assign n6207 = n3574 & n3586;
  assign n6208 = ~n3586 & ~n3741;
  assign n6209 = n3574 & ~n6208;
  assign n6210 = ~n3727 & ~n6209;
  assign n1325 = ~P1_STATE_REG | n6210;
  assign n6212 = ~n6207 & ~n1325;
  assign n6213 = n6206 & ~n6212;
  assign n6214 = ~n3723 & ~n3726;
  assign n6215 = n6213 & n6214;
  assign n6216 = ~P1_REG2_REG_18_ & n4931;
  assign n6217 = P1_REG2_REG_19_ & n3655_1;
  assign n6218 = ~P1_REG2_REG_19_ & ~n3655_1;
  assign n6219 = ~n6217 & ~n6218;
  assign n6220 = P1_REG2_REG_16_ & ~n4795;
  assign n6221 = P1_REG2_REG_17_ & n6220;
  assign n6222 = ~P1_REG2_REG_17_ & ~n6220;
  assign n6223 = ~n4862 & ~n6222;
  assign n6224 = ~P1_REG2_REG_16_ & n4795;
  assign n6225 = ~P1_REG2_REG_17_ & n4862;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = P1_REG2_REG_15_ & ~n4734;
  assign n6228 = ~P1_REG2_REG_15_ & n4734;
  assign n6229 = P1_REG2_REG_14_ & ~n4670;
  assign n6230 = ~P1_REG2_REG_14_ & n4670;
  assign n6231 = ~P1_REG2_REG_13_ & n4606;
  assign n6232 = P1_REG2_REG_13_ & ~n4606;
  assign n6233 = P1_REG2_REG_12_ & ~n4539;
  assign n6234 = P1_REG2_REG_11_ & ~n4469;
  assign n6235 = ~P1_REG2_REG_12_ & n4539;
  assign n6236 = ~n6231 & ~n6235;
  assign n6237 = n6234 & n6236;
  assign n6238 = ~n6232 & ~n6233;
  assign n6239 = ~n6237 & n6238;
  assign n6240 = ~n6231 & ~n6239;
  assign n6241 = ~P1_REG2_REG_11_ & n4469;
  assign n6242 = ~P1_REG2_REG_10_ & n4404;
  assign n6243 = P1_REG2_REG_10_ & ~n4404;
  assign n6244 = P1_REG2_REG_9_ & ~n4337;
  assign n6245 = P1_REG2_REG_8_ & ~n4269;
  assign n6246 = ~P1_REG2_REG_9_ & n4337;
  assign n6247 = ~n6242 & ~n6246;
  assign n6248 = n6245 & n6247;
  assign n6249 = ~n6243 & ~n6244;
  assign n6250 = ~n6248 & n6249;
  assign n6251 = ~n6242 & ~n6250;
  assign n6252 = ~P1_REG2_REG_8_ & n4269;
  assign n6253 = P1_REG2_REG_6_ & ~n4127;
  assign n6254 = P1_REG2_REG_7_ & n6253;
  assign n6255 = ~P1_REG2_REG_7_ & ~n6253;
  assign n6256 = ~n4201 & ~n6255;
  assign n6257 = ~P1_REG2_REG_6_ & n4127;
  assign n6258 = ~P1_REG2_REG_7_ & n4201;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = P1_REG2_REG_4_ & ~n3993;
  assign n6261 = P1_REG2_REG_5_ & n6260;
  assign n6262 = ~P1_REG2_REG_5_ & ~n6260;
  assign n6263 = ~n4063 & ~n6262;
  assign n6264 = ~P1_REG2_REG_4_ & n3993;
  assign n6265 = ~P1_REG2_REG_5_ & n4063;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = P1_REG2_REG_3_ & ~n3928;
  assign n6268 = ~P1_REG2_REG_3_ & n3928;
  assign n6269 = P1_REG2_REG_2_ & ~n3866;
  assign n6270 = ~n6268 & n6269;
  assign n6271 = ~P1_REG2_REG_2_ & n3866;
  assign n6272 = ~n6268 & ~n6271;
  assign n6273 = P1_REG2_REG_0_ & ~n3730_1;
  assign n6274 = ~P1_REG2_REG_1_ & n3810;
  assign n6275 = n6273 & ~n6274;
  assign n6276 = P1_REG2_REG_1_ & ~n3810;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = n6272 & ~n6277;
  assign n6279 = ~n6267 & ~n6270;
  assign n6280 = ~n6278 & n6279;
  assign n6281 = n6266 & ~n6280;
  assign n6282 = ~n6261 & ~n6263;
  assign n6283 = ~n6281 & n6282;
  assign n6284 = n6259 & ~n6283;
  assign n6285 = ~n6254 & ~n6256;
  assign n6286 = ~n6284 & n6285;
  assign n6287 = n6247 & ~n6252;
  assign n6288 = ~n6286 & n6287;
  assign n6289 = ~n6251 & ~n6288;
  assign n6290 = n6236 & ~n6241;
  assign n6291 = ~n6289 & n6290;
  assign n6292 = ~n6240 & ~n6291;
  assign n6293 = ~n6230 & ~n6292;
  assign n6294 = ~n6229 & ~n6293;
  assign n6295 = ~n6228 & ~n6294;
  assign n6296 = ~n6227 & ~n6295;
  assign n6297 = n6226 & ~n6296;
  assign n6298 = ~n6221 & ~n6223;
  assign n6299 = ~n6297 & n6298;
  assign n6300 = P1_REG2_REG_18_ & ~n4931;
  assign n6301 = n6299 & ~n6300;
  assign n6302 = ~n6216 & ~n6219;
  assign n6303 = ~n6301 & n6302;
  assign n6304 = ~n6216 & ~n6299;
  assign n6305 = n6219 & ~n6300;
  assign n6306 = ~n6304 & n6305;
  assign n6307 = ~n6303 & ~n6306;
  assign n6308 = n6215 & n6307;
  assign n6309 = P1_REG3_REG_19_ & ~P1_STATE_REG;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = P1_ADDR_REG_19_ & n6212;
  assign n6312 = n3726 & n6213;
  assign n6313 = ~n3655_1 & n6312;
  assign n6314 = n3723 & n6213;
  assign n6315 = ~P1_REG1_REG_18_ & n4931;
  assign n6316 = P1_REG1_REG_19_ & n3655_1;
  assign n6317 = ~P1_REG1_REG_19_ & ~n3655_1;
  assign n6318 = ~n6316 & ~n6317;
  assign n6319 = P1_REG1_REG_16_ & ~n4795;
  assign n6320 = P1_REG1_REG_17_ & n6319;
  assign n6321 = ~P1_REG1_REG_17_ & ~n6319;
  assign n6322 = ~n4862 & ~n6321;
  assign n6323 = ~P1_REG1_REG_16_ & n4795;
  assign n6324 = ~P1_REG1_REG_17_ & n4862;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = P1_REG1_REG_15_ & ~n4734;
  assign n6327 = ~P1_REG1_REG_15_ & n4734;
  assign n6328 = P1_REG1_REG_14_ & ~n4670;
  assign n6329 = ~P1_REG1_REG_14_ & n4670;
  assign n6330 = ~P1_REG1_REG_13_ & n4606;
  assign n6331 = P1_REG1_REG_13_ & ~n4606;
  assign n6332 = P1_REG1_REG_12_ & ~n4539;
  assign n6333 = P1_REG1_REG_11_ & ~n4469;
  assign n6334 = ~P1_REG1_REG_12_ & n4539;
  assign n6335 = ~n6330 & ~n6334;
  assign n6336 = n6333 & n6335;
  assign n6337 = ~n6331 & ~n6332;
  assign n6338 = ~n6336 & n6337;
  assign n6339 = ~n6330 & ~n6338;
  assign n6340 = ~P1_REG1_REG_11_ & n4469;
  assign n6341 = ~P1_REG1_REG_10_ & n4404;
  assign n6342 = P1_REG1_REG_10_ & ~n4404;
  assign n6343 = P1_REG1_REG_9_ & ~n4337;
  assign n6344 = P1_REG1_REG_8_ & ~n4269;
  assign n6345 = ~P1_REG1_REG_9_ & n4337;
  assign n6346 = ~n6341 & ~n6345;
  assign n6347 = n6344 & n6346;
  assign n6348 = ~n6342 & ~n6343;
  assign n6349 = ~n6347 & n6348;
  assign n6350 = ~n6341 & ~n6349;
  assign n6351 = ~P1_REG1_REG_8_ & n4269;
  assign n6352 = P1_REG1_REG_6_ & ~n4127;
  assign n6353 = P1_REG1_REG_7_ & n6352;
  assign n6354 = ~P1_REG1_REG_7_ & ~n6352;
  assign n6355 = ~n4201 & ~n6354;
  assign n6356 = ~P1_REG1_REG_6_ & n4127;
  assign n6357 = ~P1_REG1_REG_7_ & n4201;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = P1_REG1_REG_4_ & ~n3993;
  assign n6360 = P1_REG1_REG_5_ & n6359;
  assign n6361 = ~P1_REG1_REG_5_ & ~n6359;
  assign n6362 = ~n4063 & ~n6361;
  assign n6363 = ~P1_REG1_REG_4_ & n3993;
  assign n6364 = ~P1_REG1_REG_5_ & n4063;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = P1_REG1_REG_3_ & ~n3928;
  assign n6367 = ~P1_REG1_REG_3_ & n3928;
  assign n6368 = P1_REG1_REG_2_ & ~n3866;
  assign n6369 = ~n6367 & n6368;
  assign n6370 = ~P1_REG1_REG_2_ & n3866;
  assign n6371 = ~n6367 & ~n6370;
  assign n6372 = P1_REG1_REG_0_ & ~n3730_1;
  assign n6373 = ~P1_REG1_REG_1_ & n3810;
  assign n6374 = n6372 & ~n6373;
  assign n6375 = P1_REG1_REG_1_ & ~n3810;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = n6371 & ~n6376;
  assign n6378 = ~n6366 & ~n6369;
  assign n6379 = ~n6377 & n6378;
  assign n6380 = n6365 & ~n6379;
  assign n6381 = ~n6360 & ~n6362;
  assign n6382 = ~n6380 & n6381;
  assign n6383 = n6358 & ~n6382;
  assign n6384 = ~n6353 & ~n6355;
  assign n6385 = ~n6383 & n6384;
  assign n6386 = n6346 & ~n6351;
  assign n6387 = ~n6385 & n6386;
  assign n6388 = ~n6350 & ~n6387;
  assign n6389 = n6335 & ~n6340;
  assign n6390 = ~n6388 & n6389;
  assign n6391 = ~n6339 & ~n6390;
  assign n6392 = ~n6329 & ~n6391;
  assign n6393 = ~n6328 & ~n6392;
  assign n6394 = ~n6327 & ~n6393;
  assign n6395 = ~n6326 & ~n6394;
  assign n6396 = n6325 & ~n6395;
  assign n6397 = ~n6320 & ~n6322;
  assign n6398 = ~n6396 & n6397;
  assign n6399 = P1_REG1_REG_18_ & ~n4931;
  assign n6400 = n6398 & ~n6399;
  assign n6401 = ~n6315 & ~n6318;
  assign n6402 = ~n6400 & n6401;
  assign n6403 = ~n6315 & ~n6398;
  assign n6404 = n6318 & ~n6399;
  assign n6405 = ~n6403 & n6404;
  assign n6406 = ~n6402 & ~n6405;
  assign n6407 = n6314 & n6406;
  assign n6408 = ~n6311 & ~n6313;
  assign n6409 = ~n6407 & n6408;
  assign n6410 = n3587 & ~n6212;
  assign n6411 = ~n3782 & ~n5812;
  assign n6412 = ~n3788 & n6411;
  assign n6413 = ~n3790 & ~n3793;
  assign n6414 = ~n3784 & n6413;
  assign n6415 = ~n3643 & n3656;
  assign n6416 = ~n3795 & ~n6415;
  assign n6417 = ~n5788 & n6416;
  assign n6418 = n6412 & n6414;
  assign n6419 = n6417 & n6418;
  assign n6420 = n5800 & n6419;
  assign n6421 = ~n5789 & n6420;
  assign n6422 = n3726 & ~n6421;
  assign n6423 = ~n3655_1 & n6422;
  assign n6424 = n6214 & ~n6421;
  assign n6425 = n6307 & n6424;
  assign n6426 = n3723 & ~n6421;
  assign n6427 = n6406 & n6426;
  assign n6428 = ~n6423 & ~n6425;
  assign n6429 = ~n6427 & n6428;
  assign n6430 = n6410 & ~n6429;
  assign n6431 = n6310 & n6409;
  assign n910 = n6430 | ~n6431;
  assign n6433 = P1_REG2_REG_18_ & n4931;
  assign n6434 = ~P1_REG2_REG_18_ & ~n4931;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = n6299 & ~n6435;
  assign n6437 = ~n6299 & n6435;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = n6215 & ~n6438;
  assign n6440 = P1_REG3_REG_18_ & ~P1_STATE_REG;
  assign n6441 = ~n6439 & ~n6440;
  assign n6442 = P1_ADDR_REG_18_ & n6212;
  assign n6443 = ~n4931 & n6312;
  assign n6444 = P1_REG1_REG_18_ & n4931;
  assign n6445 = ~P1_REG1_REG_18_ & ~n4931;
  assign n6446 = ~n6444 & ~n6445;
  assign n6447 = n6398 & ~n6446;
  assign n6448 = ~n6398 & n6446;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = n6314 & ~n6449;
  assign n6451 = ~n6442 & ~n6443;
  assign n6452 = ~n6450 & n6451;
  assign n6453 = ~n4931 & n6422;
  assign n6454 = n6424 & ~n6438;
  assign n6455 = n6426 & ~n6449;
  assign n6456 = ~n6453 & ~n6454;
  assign n6457 = ~n6455 & n6456;
  assign n6458 = n6410 & ~n6457;
  assign n6459 = n6441 & n6452;
  assign n915 = n6458 | ~n6459;
  assign n6461 = P1_REG2_REG_17_ & ~n4862;
  assign n6462 = ~n6220 & n6296;
  assign n6463 = n6226 & ~n6461;
  assign n6464 = ~n6462 & n6463;
  assign n6465 = P1_REG2_REG_17_ & n4862;
  assign n6466 = ~P1_REG2_REG_17_ & ~n4862;
  assign n6467 = ~n6224 & ~n6296;
  assign n6468 = ~n6465 & ~n6466;
  assign n6469 = ~n6220 & n6468;
  assign n6470 = ~n6467 & n6469;
  assign n6471 = ~n6464 & ~n6470;
  assign n6472 = n6215 & n6471;
  assign n6473 = P1_REG3_REG_17_ & ~P1_STATE_REG;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = P1_ADDR_REG_17_ & n6212;
  assign n6476 = ~n4862 & n6312;
  assign n6477 = P1_REG1_REG_17_ & ~n4862;
  assign n6478 = ~n6319 & n6395;
  assign n6479 = n6325 & ~n6477;
  assign n6480 = ~n6478 & n6479;
  assign n6481 = P1_REG1_REG_17_ & n4862;
  assign n6482 = ~P1_REG1_REG_17_ & ~n4862;
  assign n6483 = ~n6323 & ~n6395;
  assign n6484 = ~n6481 & ~n6482;
  assign n6485 = ~n6319 & n6484;
  assign n6486 = ~n6483 & n6485;
  assign n6487 = ~n6480 & ~n6486;
  assign n6488 = n6314 & n6487;
  assign n6489 = ~n6475 & ~n6476;
  assign n6490 = ~n6488 & n6489;
  assign n6491 = ~n4862 & n6422;
  assign n6492 = n6424 & n6471;
  assign n6493 = n6426 & n6487;
  assign n6494 = ~n6491 & ~n6492;
  assign n6495 = ~n6493 & n6494;
  assign n6496 = n6410 & ~n6495;
  assign n6497 = n6474 & n6490;
  assign n920 = n6496 | ~n6497;
  assign n6499 = P1_REG2_REG_16_ & n4795;
  assign n6500 = ~P1_REG2_REG_16_ & ~n4795;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = n6296 & ~n6501;
  assign n6503 = ~n6220 & ~n6224;
  assign n6504 = ~n6296 & ~n6503;
  assign n6505 = ~n6502 & ~n6504;
  assign n6506 = n6215 & ~n6505;
  assign n6507 = P1_REG3_REG_16_ & ~P1_STATE_REG;
  assign n6508 = ~n6506 & ~n6507;
  assign n6509 = P1_ADDR_REG_16_ & n6212;
  assign n6510 = ~n4795 & n6312;
  assign n6511 = P1_REG1_REG_16_ & n4795;
  assign n6512 = ~P1_REG1_REG_16_ & ~n4795;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = n6395 & ~n6513;
  assign n6515 = ~n6319 & ~n6323;
  assign n6516 = ~n6395 & ~n6515;
  assign n6517 = ~n6514 & ~n6516;
  assign n6518 = n6314 & ~n6517;
  assign n6519 = ~n6509 & ~n6510;
  assign n6520 = ~n6518 & n6519;
  assign n6521 = ~n4795 & n6422;
  assign n6522 = n6424 & ~n6505;
  assign n6523 = n6426 & ~n6517;
  assign n6524 = ~n6521 & ~n6522;
  assign n6525 = ~n6523 & n6524;
  assign n6526 = n6410 & ~n6525;
  assign n6527 = n6508 & n6520;
  assign n925 = n6526 | ~n6527;
  assign n6529 = P1_REG2_REG_15_ & n4734;
  assign n6530 = ~P1_REG2_REG_15_ & ~n4734;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = n6294 & ~n6531;
  assign n6533 = ~n6294 & n6531;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = n6215 & ~n6534;
  assign n6536 = P1_REG3_REG_15_ & ~P1_STATE_REG;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = P1_ADDR_REG_15_ & n6212;
  assign n6539 = ~n4734 & n6312;
  assign n6540 = P1_REG1_REG_15_ & n4734;
  assign n6541 = ~P1_REG1_REG_15_ & ~n4734;
  assign n6542 = ~n6540 & ~n6541;
  assign n6543 = n6393 & ~n6542;
  assign n6544 = ~n6393 & n6542;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = n6314 & ~n6545;
  assign n6547 = ~n6538 & ~n6539;
  assign n6548 = ~n6546 & n6547;
  assign n6549 = ~n4734 & n6422;
  assign n6550 = n6424 & ~n6534;
  assign n6551 = n6426 & ~n6545;
  assign n6552 = ~n6549 & ~n6550;
  assign n6553 = ~n6551 & n6552;
  assign n6554 = n6410 & ~n6553;
  assign n6555 = n6537 & n6548;
  assign n930 = n6554 | ~n6555;
  assign n6557 = P1_REG2_REG_14_ & n4670;
  assign n6558 = ~P1_REG2_REG_14_ & ~n4670;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = n6292 & ~n6559;
  assign n6561 = ~n6292 & n6559;
  assign n6562 = ~n6560 & ~n6561;
  assign n6563 = n6215 & ~n6562;
  assign n6564 = P1_REG3_REG_14_ & ~P1_STATE_REG;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = P1_ADDR_REG_14_ & n6212;
  assign n6567 = ~n4670 & n6312;
  assign n6568 = P1_REG1_REG_14_ & n4670;
  assign n6569 = ~P1_REG1_REG_14_ & ~n4670;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = n6391 & ~n6570;
  assign n6572 = ~n6391 & n6570;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = n6314 & ~n6573;
  assign n6575 = ~n6566 & ~n6567;
  assign n6576 = ~n6574 & n6575;
  assign n6577 = ~n4670 & n6422;
  assign n6578 = n6424 & ~n6562;
  assign n6579 = n6426 & ~n6573;
  assign n6580 = ~n6577 & ~n6578;
  assign n6581 = ~n6579 & n6580;
  assign n6582 = n6410 & ~n6581;
  assign n6583 = n6565 & n6576;
  assign n935 = n6582 | ~n6583;
  assign n6585 = ~n6241 & ~n6289;
  assign n6586 = ~n6234 & ~n6585;
  assign n6587 = ~n6233 & n6586;
  assign n6588 = ~n6232 & n6236;
  assign n6589 = ~n6587 & n6588;
  assign n6590 = P1_REG2_REG_13_ & n4606;
  assign n6591 = ~P1_REG2_REG_13_ & ~n4606;
  assign n6592 = ~n6235 & ~n6586;
  assign n6593 = ~n6590 & ~n6591;
  assign n6594 = ~n6233 & n6593;
  assign n6595 = ~n6592 & n6594;
  assign n6596 = ~n6589 & ~n6595;
  assign n6597 = n6215 & n6596;
  assign n6598 = P1_REG3_REG_13_ & ~P1_STATE_REG;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = P1_ADDR_REG_13_ & n6212;
  assign n6601 = ~n4606 & n6312;
  assign n6602 = ~n6340 & ~n6388;
  assign n6603 = ~n6333 & ~n6602;
  assign n6604 = ~n6332 & n6603;
  assign n6605 = ~n6331 & n6335;
  assign n6606 = ~n6604 & n6605;
  assign n6607 = P1_REG1_REG_13_ & n4606;
  assign n6608 = ~P1_REG1_REG_13_ & ~n4606;
  assign n6609 = ~n6334 & ~n6603;
  assign n6610 = ~n6607 & ~n6608;
  assign n6611 = ~n6332 & n6610;
  assign n6612 = ~n6609 & n6611;
  assign n6613 = ~n6606 & ~n6612;
  assign n6614 = n6314 & n6613;
  assign n6615 = ~n6600 & ~n6601;
  assign n6616 = ~n6614 & n6615;
  assign n6617 = ~n4606 & n6422;
  assign n6618 = n6424 & n6596;
  assign n6619 = n6426 & n6613;
  assign n6620 = ~n6617 & ~n6618;
  assign n6621 = ~n6619 & n6620;
  assign n6622 = n6410 & ~n6621;
  assign n6623 = n6599 & n6616;
  assign n940 = n6622 | ~n6623;
  assign n6625 = P1_REG2_REG_12_ & n4539;
  assign n6626 = ~P1_REG2_REG_12_ & ~n4539;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = n6586 & ~n6627;
  assign n6629 = ~n6233 & ~n6235;
  assign n6630 = ~n6586 & ~n6629;
  assign n6631 = ~n6628 & ~n6630;
  assign n6632 = n6215 & ~n6631;
  assign n6633 = P1_REG3_REG_12_ & ~P1_STATE_REG;
  assign n6634 = ~n6632 & ~n6633;
  assign n6635 = P1_ADDR_REG_12_ & n6212;
  assign n6636 = ~n4539 & n6312;
  assign n6637 = P1_REG1_REG_12_ & n4539;
  assign n6638 = ~P1_REG1_REG_12_ & ~n4539;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = n6603 & ~n6639;
  assign n6641 = ~n6332 & ~n6334;
  assign n6642 = ~n6603 & ~n6641;
  assign n6643 = ~n6640 & ~n6642;
  assign n6644 = n6314 & ~n6643;
  assign n6645 = ~n6635 & ~n6636;
  assign n6646 = ~n6644 & n6645;
  assign n6647 = ~n4539 & n6422;
  assign n6648 = n6424 & ~n6631;
  assign n6649 = n6426 & ~n6643;
  assign n6650 = ~n6647 & ~n6648;
  assign n6651 = ~n6649 & n6650;
  assign n6652 = n6410 & ~n6651;
  assign n6653 = n6634 & n6646;
  assign n945 = n6652 | ~n6653;
  assign n6655 = P1_REG2_REG_11_ & n4469;
  assign n6656 = ~P1_REG2_REG_11_ & ~n4469;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = n6289 & ~n6657;
  assign n6659 = ~n6234 & ~n6241;
  assign n6660 = ~n6289 & ~n6659;
  assign n6661 = ~n6658 & ~n6660;
  assign n6662 = n6215 & ~n6661;
  assign n6663 = P1_REG3_REG_11_ & ~P1_STATE_REG;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = P1_ADDR_REG_11_ & n6212;
  assign n6666 = ~n4469 & n6312;
  assign n6667 = P1_REG1_REG_11_ & n4469;
  assign n6668 = ~P1_REG1_REG_11_ & ~n4469;
  assign n6669 = ~n6667 & ~n6668;
  assign n6670 = n6388 & ~n6669;
  assign n6671 = ~n6333 & ~n6340;
  assign n6672 = ~n6388 & ~n6671;
  assign n6673 = ~n6670 & ~n6672;
  assign n6674 = n6314 & ~n6673;
  assign n6675 = ~n6665 & ~n6666;
  assign n6676 = ~n6674 & n6675;
  assign n6677 = ~n4469 & n6422;
  assign n6678 = n6424 & ~n6661;
  assign n6679 = n6426 & ~n6673;
  assign n6680 = ~n6677 & ~n6678;
  assign n6681 = ~n6679 & n6680;
  assign n6682 = n6410 & ~n6681;
  assign n6683 = n6664 & n6676;
  assign n950 = n6682 | ~n6683;
  assign n6685 = ~n6252 & ~n6286;
  assign n6686 = ~n6245 & ~n6685;
  assign n6687 = ~n6244 & n6686;
  assign n6688 = ~n6243 & n6247;
  assign n6689 = ~n6687 & n6688;
  assign n6690 = P1_REG2_REG_10_ & n4404;
  assign n6691 = ~P1_REG2_REG_10_ & ~n4404;
  assign n6692 = ~n6246 & ~n6686;
  assign n6693 = ~n6690 & ~n6691;
  assign n6694 = ~n6244 & n6693;
  assign n6695 = ~n6692 & n6694;
  assign n6696 = ~n6689 & ~n6695;
  assign n6697 = n6215 & n6696;
  assign n6698 = P1_REG3_REG_10_ & ~P1_STATE_REG;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = P1_ADDR_REG_10_ & n6212;
  assign n6701 = ~n4404 & n6312;
  assign n6702 = ~n6351 & ~n6385;
  assign n6703 = ~n6344 & ~n6702;
  assign n6704 = ~n6343 & n6703;
  assign n6705 = ~n6342 & n6346;
  assign n6706 = ~n6704 & n6705;
  assign n6707 = P1_REG1_REG_10_ & n4404;
  assign n6708 = ~P1_REG1_REG_10_ & ~n4404;
  assign n6709 = ~n6345 & ~n6703;
  assign n6710 = ~n6707 & ~n6708;
  assign n6711 = ~n6343 & n6710;
  assign n6712 = ~n6709 & n6711;
  assign n6713 = ~n6706 & ~n6712;
  assign n6714 = n6314 & n6713;
  assign n6715 = ~n6700 & ~n6701;
  assign n6716 = ~n6714 & n6715;
  assign n6717 = ~n4404 & n6422;
  assign n6718 = n6424 & n6696;
  assign n6719 = n6426 & n6713;
  assign n6720 = ~n6717 & ~n6718;
  assign n6721 = ~n6719 & n6720;
  assign n6722 = n6410 & ~n6721;
  assign n6723 = n6699 & n6716;
  assign n955 = n6722 | ~n6723;
  assign n6725 = P1_REG2_REG_9_ & n4337;
  assign n6726 = ~P1_REG2_REG_9_ & ~n4337;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = n6686 & ~n6727;
  assign n6729 = ~n6244 & ~n6246;
  assign n6730 = ~n6686 & ~n6729;
  assign n6731 = ~n6728 & ~n6730;
  assign n6732 = n6215 & ~n6731;
  assign n6733 = P1_REG3_REG_9_ & ~P1_STATE_REG;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = P1_ADDR_REG_9_ & n6212;
  assign n6736 = ~n4337 & n6312;
  assign n6737 = P1_REG1_REG_9_ & n4337;
  assign n6738 = ~P1_REG1_REG_9_ & ~n4337;
  assign n6739 = ~n6737 & ~n6738;
  assign n6740 = n6703 & ~n6739;
  assign n6741 = ~n6343 & ~n6345;
  assign n6742 = ~n6703 & ~n6741;
  assign n6743 = ~n6740 & ~n6742;
  assign n6744 = n6314 & ~n6743;
  assign n6745 = ~n6735 & ~n6736;
  assign n6746 = ~n6744 & n6745;
  assign n6747 = ~n4337 & n6422;
  assign n6748 = n6424 & ~n6731;
  assign n6749 = n6426 & ~n6743;
  assign n6750 = ~n6747 & ~n6748;
  assign n6751 = ~n6749 & n6750;
  assign n6752 = n6410 & ~n6751;
  assign n6753 = n6734 & n6746;
  assign n960 = n6752 | ~n6753;
  assign n6755 = P1_REG2_REG_8_ & n4269;
  assign n6756 = ~P1_REG2_REG_8_ & ~n4269;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = n6286 & ~n6757;
  assign n6759 = ~n6245 & ~n6252;
  assign n6760 = ~n6286 & ~n6759;
  assign n6761 = ~n6758 & ~n6760;
  assign n6762 = n6215 & ~n6761;
  assign n6763 = P1_REG3_REG_8_ & ~P1_STATE_REG;
  assign n6764 = ~n6762 & ~n6763;
  assign n6765 = P1_ADDR_REG_8_ & n6212;
  assign n6766 = ~n4269 & n6312;
  assign n6767 = P1_REG1_REG_8_ & n4269;
  assign n6768 = ~P1_REG1_REG_8_ & ~n4269;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = n6385 & ~n6769;
  assign n6771 = ~n6344 & ~n6351;
  assign n6772 = ~n6385 & ~n6771;
  assign n6773 = ~n6770 & ~n6772;
  assign n6774 = n6314 & ~n6773;
  assign n6775 = ~n6765 & ~n6766;
  assign n6776 = ~n6774 & n6775;
  assign n6777 = ~n4269 & n6422;
  assign n6778 = n6424 & ~n6761;
  assign n6779 = n6426 & ~n6773;
  assign n6780 = ~n6777 & ~n6778;
  assign n6781 = ~n6779 & n6780;
  assign n6782 = n6410 & ~n6781;
  assign n6783 = n6764 & n6776;
  assign n965 = n6782 | ~n6783;
  assign n6785 = P1_REG2_REG_7_ & ~n4201;
  assign n6786 = ~n6253 & n6283;
  assign n6787 = n6259 & ~n6785;
  assign n6788 = ~n6786 & n6787;
  assign n6789 = P1_REG2_REG_7_ & n4201;
  assign n6790 = ~P1_REG2_REG_7_ & ~n4201;
  assign n6791 = ~n6257 & ~n6283;
  assign n6792 = ~n6789 & ~n6790;
  assign n6793 = ~n6253 & n6792;
  assign n6794 = ~n6791 & n6793;
  assign n6795 = ~n6788 & ~n6794;
  assign n6796 = n6215 & n6795;
  assign n6797 = P1_REG3_REG_7_ & ~P1_STATE_REG;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = P1_ADDR_REG_7_ & n6212;
  assign n6800 = ~n4201 & n6312;
  assign n6801 = P1_REG1_REG_7_ & ~n4201;
  assign n6802 = ~n6352 & n6382;
  assign n6803 = n6358 & ~n6801;
  assign n6804 = ~n6802 & n6803;
  assign n6805 = P1_REG1_REG_7_ & n4201;
  assign n6806 = ~P1_REG1_REG_7_ & ~n4201;
  assign n6807 = ~n6356 & ~n6382;
  assign n6808 = ~n6805 & ~n6806;
  assign n6809 = ~n6352 & n6808;
  assign n6810 = ~n6807 & n6809;
  assign n6811 = ~n6804 & ~n6810;
  assign n6812 = n6314 & n6811;
  assign n6813 = ~n6799 & ~n6800;
  assign n6814 = ~n6812 & n6813;
  assign n6815 = ~n4201 & n6422;
  assign n6816 = n6424 & n6795;
  assign n6817 = n6426 & n6811;
  assign n6818 = ~n6815 & ~n6816;
  assign n6819 = ~n6817 & n6818;
  assign n6820 = n6410 & ~n6819;
  assign n6821 = n6798 & n6814;
  assign n970 = n6820 | ~n6821;
  assign n6823 = P1_REG2_REG_6_ & n4127;
  assign n6824 = ~P1_REG2_REG_6_ & ~n4127;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = n6283 & ~n6825;
  assign n6827 = ~n6253 & ~n6257;
  assign n6828 = ~n6283 & ~n6827;
  assign n6829 = ~n6826 & ~n6828;
  assign n6830 = n6215 & ~n6829;
  assign n6831 = P1_REG3_REG_6_ & ~P1_STATE_REG;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = P1_REG1_REG_6_ & n4127;
  assign n6834 = ~P1_REG1_REG_6_ & ~n4127;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = n6382 & ~n6835;
  assign n6837 = ~n6352 & ~n6356;
  assign n6838 = ~n6382 & ~n6837;
  assign n6839 = ~n6836 & ~n6838;
  assign n6840 = n6314 & ~n6839;
  assign n6841 = ~n4127 & n6312;
  assign n6842 = P1_ADDR_REG_6_ & n6212;
  assign n6843 = ~n6840 & ~n6841;
  assign n6844 = ~n6842 & n6843;
  assign n6845 = ~n4127 & n6422;
  assign n6846 = n6424 & ~n6829;
  assign n6847 = n6426 & ~n6839;
  assign n6848 = ~n6845 & ~n6846;
  assign n6849 = ~n6847 & n6848;
  assign n6850 = n6410 & ~n6849;
  assign n6851 = n6832 & n6844;
  assign n975 = n6850 | ~n6851;
  assign n6853 = P1_REG2_REG_5_ & ~n4063;
  assign n6854 = n6272 & n6275;
  assign n6855 = ~n6271 & n6276;
  assign n6856 = ~n6269 & ~n6855;
  assign n6857 = ~n6268 & ~n6856;
  assign n6858 = ~n6267 & ~n6854;
  assign n6859 = ~n6857 & n6858;
  assign n6860 = ~n6260 & n6859;
  assign n6861 = n6266 & ~n6853;
  assign n6862 = ~n6860 & n6861;
  assign n6863 = P1_REG2_REG_5_ & n4063;
  assign n6864 = ~P1_REG2_REG_5_ & ~n4063;
  assign n6865 = ~n6264 & ~n6859;
  assign n6866 = ~n6863 & ~n6864;
  assign n6867 = ~n6260 & n6866;
  assign n6868 = ~n6865 & n6867;
  assign n6869 = ~n6862 & ~n6868;
  assign n6870 = n6215 & n6869;
  assign n6871 = P1_REG3_REG_5_ & ~P1_STATE_REG;
  assign n6872 = ~n6870 & ~n6871;
  assign n6873 = ~n4063 & n6422;
  assign n6874 = n6424 & n6869;
  assign n6875 = P1_REG1_REG_5_ & ~n4063;
  assign n6876 = n6371 & n6374;
  assign n6877 = ~n6370 & n6375;
  assign n6878 = ~n6368 & ~n6877;
  assign n6879 = ~n6367 & ~n6878;
  assign n6880 = ~n6366 & ~n6876;
  assign n6881 = ~n6879 & n6880;
  assign n6882 = ~n6359 & n6881;
  assign n6883 = n6365 & ~n6875;
  assign n6884 = ~n6882 & n6883;
  assign n6885 = P1_REG1_REG_5_ & n4063;
  assign n6886 = ~P1_REG1_REG_5_ & ~n4063;
  assign n6887 = ~n6363 & ~n6881;
  assign n6888 = ~n6885 & ~n6886;
  assign n6889 = ~n6359 & n6888;
  assign n6890 = ~n6887 & n6889;
  assign n6891 = ~n6884 & ~n6890;
  assign n6892 = n6426 & n6891;
  assign n6893 = ~n6873 & ~n6874;
  assign n6894 = ~n6892 & n6893;
  assign n6895 = n6410 & ~n6894;
  assign n6896 = n6314 & n6891;
  assign n6897 = ~n4063 & n6312;
  assign n6898 = P1_ADDR_REG_5_ & n6212;
  assign n6899 = ~n6896 & ~n6897;
  assign n6900 = ~n6898 & n6899;
  assign n6901 = n6872 & ~n6895;
  assign n980 = ~n6900 | ~n6901;
  assign n6903 = ~n3993 & n6422;
  assign n6904 = P1_REG2_REG_4_ & n3993;
  assign n6905 = ~P1_REG2_REG_4_ & ~n3993;
  assign n6906 = ~n6904 & ~n6905;
  assign n6907 = n6859 & ~n6906;
  assign n6908 = ~n6260 & ~n6264;
  assign n6909 = ~n6859 & ~n6908;
  assign n6910 = ~n6907 & ~n6909;
  assign n6911 = n6424 & ~n6910;
  assign n6912 = P1_REG1_REG_4_ & n3993;
  assign n6913 = ~P1_REG1_REG_4_ & ~n3993;
  assign n6914 = ~n6912 & ~n6913;
  assign n6915 = n6881 & ~n6914;
  assign n6916 = ~n6359 & ~n6363;
  assign n6917 = ~n6881 & ~n6916;
  assign n6918 = ~n6915 & ~n6917;
  assign n6919 = n6426 & ~n6918;
  assign n6920 = ~n6903 & ~n6911;
  assign n6921 = ~n6919 & n6920;
  assign n6922 = n6410 & ~n6921;
  assign n6923 = P1_REG3_REG_4_ & ~P1_STATE_REG;
  assign n1330 = P1_STATE_REG & n6207;
  assign n6925 = P1_REG2_REG_0_ & n6214;
  assign n6926 = n3730_1 & n6925;
  assign n6927 = ~P1_REG2_REG_0_ & ~n3723;
  assign n6928 = ~n3726 & ~n6927;
  assign n6929 = ~n3730_1 & ~n6928;
  assign n6930 = ~n3646 & ~n3649;
  assign n6931 = ~n3734 & ~n6930;
  assign n6932 = n3643 & n3646;
  assign n6933 = ~n3586 & n6932;
  assign n6934 = n6931 & ~n6933;
  assign n6935 = ~n3586 & ~n6934;
  assign n6936 = n3586 & ~n3730_1;
  assign n6937 = ~n3784 & ~n5812;
  assign n6938 = ~n3586 & ~n6937;
  assign n6939 = ~n3733 & n6938;
  assign n6940 = ~n6936 & ~n6939;
  assign n6941 = ~n3781 & ~n6415;
  assign n6942 = ~n3788 & n6941;
  assign n6943 = ~n3586 & ~n6942;
  assign n6944 = ~n3586 & n3734;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = ~n3767 & ~n6945;
  assign n6947 = n6940 & ~n6946;
  assign n6948 = n6935 & n6947;
  assign n6949 = ~n6935 & ~n6947;
  assign n6950 = ~n6948 & ~n6949;
  assign n6951 = ~n3767 & n6938;
  assign n6952 = P1_REG1_REG_0_ & n3586;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = ~n6933 & n6945;
  assign n6955 = ~n3733 & ~n6954;
  assign n6956 = n6953 & ~n6955;
  assign n6957 = ~n6935 & ~n6956;
  assign n6958 = n6935 & n6956;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6950 & n6959;
  assign n6961 = n6950 & ~n6959;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = n3723 & ~n3726;
  assign n6964 = ~n6962 & n6963;
  assign n6965 = ~n6926 & ~n6929;
  assign n6966 = ~n6964 & n6965;
  assign n6967 = n1330 & ~n6966;
  assign n6968 = ~n6923 & ~n6967;
  assign n6969 = n6215 & ~n6910;
  assign n6970 = n6968 & ~n6969;
  assign n6971 = n6314 & ~n6918;
  assign n6972 = ~n3993 & n6312;
  assign n6973 = P1_ADDR_REG_4_ & n6212;
  assign n6974 = ~n6971 & ~n6972;
  assign n6975 = ~n6973 & n6974;
  assign n6976 = ~n6922 & n6970;
  assign n985 = ~n6975 | ~n6976;
  assign n6978 = ~n6271 & n6275;
  assign n6979 = n6856 & ~n6978;
  assign n6980 = P1_REG2_REG_3_ & n3928;
  assign n6981 = ~P1_REG2_REG_3_ & ~n3928;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = n6979 & ~n6982;
  assign n6984 = ~n6267 & ~n6268;
  assign n6985 = ~n6979 & ~n6984;
  assign n6986 = ~n6983 & ~n6985;
  assign n6987 = n6215 & ~n6986;
  assign n6988 = P1_REG3_REG_3_ & ~P1_STATE_REG;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = ~n3928 & n6422;
  assign n6991 = n6424 & ~n6986;
  assign n6992 = ~n6370 & n6374;
  assign n6993 = n6878 & ~n6992;
  assign n6994 = P1_REG1_REG_3_ & n3928;
  assign n6995 = ~P1_REG1_REG_3_ & ~n3928;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = n6993 & ~n6996;
  assign n6998 = ~n6366 & ~n6367;
  assign n6999 = ~n6993 & ~n6998;
  assign n7000 = ~n6997 & ~n6999;
  assign n7001 = n6426 & ~n7000;
  assign n7002 = ~n6990 & ~n6991;
  assign n7003 = ~n7001 & n7002;
  assign n7004 = n6410 & ~n7003;
  assign n7005 = n6314 & ~n7000;
  assign n7006 = ~n3928 & n6312;
  assign n7007 = P1_ADDR_REG_3_ & n6212;
  assign n7008 = ~n7005 & ~n7006;
  assign n7009 = ~n7007 & n7008;
  assign n7010 = n6989 & ~n7004;
  assign n990 = ~n7009 | ~n7010;
  assign n7012 = ~n3866 & n6422;
  assign n7013 = ~n6269 & ~n6271;
  assign n7014 = ~n6277 & n7013;
  assign n7015 = P1_REG2_REG_2_ & n3866;
  assign n7016 = ~P1_REG2_REG_2_ & ~n3866;
  assign n7017 = n6277 & ~n7015;
  assign n7018 = ~n7016 & n7017;
  assign n7019 = ~n7014 & ~n7018;
  assign n7020 = n6424 & n7019;
  assign n7021 = ~n6368 & ~n6370;
  assign n7022 = ~n6376 & n7021;
  assign n7023 = P1_REG1_REG_2_ & n3866;
  assign n7024 = ~P1_REG1_REG_2_ & ~n3866;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = ~n6375 & n7025;
  assign n7027 = ~n6374 & n7026;
  assign n7028 = ~n7022 & ~n7027;
  assign n7029 = n6426 & n7028;
  assign n7030 = ~n7012 & ~n7020;
  assign n7031 = ~n7029 & n7030;
  assign n7032 = n6410 & ~n7031;
  assign n7033 = P1_REG3_REG_2_ & ~P1_STATE_REG;
  assign n7034 = ~n6967 & ~n7033;
  assign n7035 = n6215 & n7019;
  assign n7036 = n7034 & ~n7035;
  assign n7037 = n6314 & n7028;
  assign n7038 = ~n3866 & n6312;
  assign n7039 = P1_ADDR_REG_2_ & n6212;
  assign n7040 = ~n7037 & ~n7038;
  assign n7041 = ~n7039 & n7040;
  assign n7042 = ~n7032 & n7036;
  assign n995 = ~n7041 | ~n7042;
  assign n7044 = ~n6274 & ~n6276;
  assign n7045 = ~n6273 & n7044;
  assign n7046 = n6273 & ~n7044;
  assign n7047 = ~n7045 & ~n7046;
  assign n7048 = n6215 & ~n7047;
  assign n7049 = P1_REG3_REG_1_ & ~P1_STATE_REG;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = ~n3810 & n6422;
  assign n7052 = n6424 & ~n7047;
  assign n7053 = ~n6373 & ~n6375;
  assign n7054 = ~n6372 & n7053;
  assign n7055 = n6372 & ~n7053;
  assign n7056 = ~n7054 & ~n7055;
  assign n7057 = n6426 & ~n7056;
  assign n7058 = ~n7051 & ~n7052;
  assign n7059 = ~n7057 & n7058;
  assign n7060 = n6410 & ~n7059;
  assign n7061 = n6314 & ~n7056;
  assign n7062 = ~n3810 & n6312;
  assign n7063 = P1_ADDR_REG_1_ & n6212;
  assign n7064 = ~n7061 & ~n7062;
  assign n7065 = ~n7063 & n7064;
  assign n7066 = n7050 & ~n7060;
  assign n1000 = ~n7065 | ~n7066;
  assign n7068 = P1_REG2_REG_0_ & n3730_1;
  assign n7069 = ~P1_REG2_REG_0_ & ~n3730_1;
  assign n7070 = ~n7068 & ~n7069;
  assign n7071 = n6215 & ~n7070;
  assign n7072 = P1_REG3_REG_0_ & ~P1_STATE_REG;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = ~n3730_1 & n6422;
  assign n7075 = n6424 & ~n7070;
  assign n7076 = P1_REG1_REG_0_ & n3730_1;
  assign n7077 = ~P1_REG1_REG_0_ & ~n3730_1;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = n6426 & ~n7078;
  assign n7080 = ~n7074 & ~n7075;
  assign n7081 = ~n7079 & n7080;
  assign n7082 = n6410 & ~n7081;
  assign n7083 = n6314 & ~n7078;
  assign n7084 = ~n3730_1 & n6312;
  assign n7085 = P1_ADDR_REG_0_ & n6212;
  assign n7086 = ~n7083 & ~n7084;
  assign n7087 = ~n7085 & n7086;
  assign n7088 = n7073 & ~n7082;
  assign n1005 = ~n7087 | ~n7088;
  assign n7090 = ~n3767 & n1330;
  assign n7091 = P1_DATAO_REG_0_ & ~n1330;
  assign n1010 = n7090 | n7091;
  assign n7093 = ~n3759 & n1330;
  assign n7094 = P1_DATAO_REG_1_ & ~n1330;
  assign n1015 = n7093 | n7094;
  assign n7096 = ~n3824 & n1330;
  assign n7097 = P1_DATAO_REG_2_ & ~n1330;
  assign n1020 = n7096 | n7097;
  assign n7099 = ~n3881 & n1330;
  assign n7100 = P1_DATAO_REG_3_ & ~n1330;
  assign n1025 = n7099 | n7100;
  assign n7102 = ~n3945 & n1330;
  assign n7103 = P1_DATAO_REG_4_ & ~n1330;
  assign n1030 = n7102 | n7103;
  assign n7105 = ~n4011 & n1330;
  assign n7106 = P1_DATAO_REG_5_ & ~n1330;
  assign n1035 = n7105 | n7106;
  assign n7108 = ~n4081 & n1330;
  assign n7109 = P1_DATAO_REG_6_ & ~n1330;
  assign n1040 = n7108 | n7109;
  assign n7111 = ~n4146 & n1330;
  assign n7112 = P1_DATAO_REG_7_ & ~n1330;
  assign n1045 = n7111 | n7112;
  assign n7114 = ~n4219 & n1330;
  assign n7115 = P1_DATAO_REG_8_ & ~n1330;
  assign n1050 = n7114 | n7115;
  assign n7117 = ~n4287 & n1330;
  assign n7118 = P1_DATAO_REG_9_ & ~n1330;
  assign n1055 = n7117 | n7118;
  assign n7120 = ~n4355 & n1330;
  assign n7121 = P1_DATAO_REG_10_ & ~n1330;
  assign n1060 = n7120 | n7121;
  assign n7123 = ~n4423 & n1330;
  assign n7124 = P1_DATAO_REG_11_ & ~n1330;
  assign n1065 = n7123 | n7124;
  assign n7126 = ~n4505 & n1330;
  assign n7127 = P1_DATAO_REG_12_ & ~n1330;
  assign n1070 = n7126 | n7127;
  assign n7129 = ~n4570 & n1330;
  assign n7130 = P1_DATAO_REG_13_ & ~n1330;
  assign n1075 = n7129 | n7130;
  assign n7132 = ~n4639 & n1330;
  assign n7133 = P1_DATAO_REG_14_ & ~n1330;
  assign n1080 = n7132 | n7133;
  assign n7135 = ~n4703 & n1330;
  assign n7136 = P1_DATAO_REG_15_ & ~n1330;
  assign n1085 = n7135 | n7136;
  assign n7138 = ~n4752 & n1330;
  assign n7139 = P1_DATAO_REG_16_ & ~n1330;
  assign n1090 = n7138 | n7139;
  assign n7141 = ~n4813 & n1330;
  assign n7142 = P1_DATAO_REG_17_ & ~n1330;
  assign n1095 = n7141 | n7142;
  assign n7144 = ~n4895 & n1330;
  assign n7145 = P1_DATAO_REG_18_ & ~n1330;
  assign n1100 = n7144 | n7145;
  assign n7147 = ~n4967 & n1330;
  assign n7148 = P1_DATAO_REG_19_ & ~n1330;
  assign n1105 = n7147 | n7148;
  assign n7150 = ~n5013 & n1330;
  assign n7151 = P1_DATAO_REG_20_ & ~n1330;
  assign n1110 = n7150 | n7151;
  assign n7153 = ~n5073 & n1330;
  assign n7154 = P1_DATAO_REG_21_ & ~n1330;
  assign n1115 = n7153 | n7154;
  assign n7156 = ~n5132 & n1330;
  assign n7157 = P1_DATAO_REG_22_ & ~n1330;
  assign n1120 = n7156 | n7157;
  assign n7159 = ~n5191 & n1330;
  assign n7160 = P1_DATAO_REG_23_ & ~n1330;
  assign n1125 = n7159 | n7160;
  assign n7162 = ~n5253 & n1330;
  assign n7163 = P1_DATAO_REG_24_ & ~n1330;
  assign n1130 = n7162 | n7163;
  assign n7165 = ~n5312 & n1330;
  assign n7166 = P1_DATAO_REG_25_ & ~n1330;
  assign n1135 = n7165 | n7166;
  assign n7168 = ~n5376 & n1330;
  assign n7169 = P1_DATAO_REG_26_ & ~n1330;
  assign n1140 = n7168 | n7169;
  assign n7171 = ~n5433 & n1330;
  assign n7172 = P1_DATAO_REG_27_ & ~n1330;
  assign n1145 = n7171 | n7172;
  assign n7174 = ~n5493 & n1330;
  assign n7175 = P1_DATAO_REG_28_ & ~n1330;
  assign n1150 = n7174 | n7175;
  assign n7177 = ~n5550 & n1330;
  assign n7178 = P1_DATAO_REG_29_ & ~n1330;
  assign n1155 = n7177 | n7178;
  assign n7180 = ~n5648 & n1330;
  assign n7181 = P1_DATAO_REG_30_ & ~n1330;
  assign n1160 = n7180 | n7181;
  assign n7183 = ~n5668 & n1330;
  assign n7184 = P1_DATAO_REG_31_ & ~n1330;
  assign n1165 = n7183 | n7184;
  assign n7186 = ~n3574 & ~n3643;
  assign n7187 = ~n3643 & n3784;
  assign n7188 = n6214 & n7187;
  assign n7189 = n3574 & ~n7188;
  assign n7190 = P1_STATE_REG & ~n6207;
  assign n7191 = ~n7186 & ~n7189;
  assign n7192 = n7190 & n7191;
  assign n7193 = P1_B_REG & ~n7192;
  assign n7194 = ~n3735_1 & ~n3778;
  assign n7195 = n3643 & n3781;
  assign n7196 = ~n3793 & ~n7195;
  assign n7197 = ~n5648 & n5668;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = n7194 & ~n7198;
  assign n7200 = ~n5668 & ~n7199;
  assign n7201 = n5648 & ~n5668;
  assign n7202 = ~n7197 & ~n7201;
  assign n7203 = ~n7196 & n7197;
  assign n7204 = n7202 & n7203;
  assign n7205 = ~n7200 & ~n7204;
  assign n7206 = ~n3574 & n7187;
  assign n7207 = ~n3643 & n3734;
  assign n7208 = ~n3737 & ~n7207;
  assign n7209 = ~n3785 & n7208;
  assign n7210 = ~n5812 & ~n7206;
  assign n7211 = n7209 & n7210;
  assign n7212 = ~n3790 & ~n5798;
  assign n7213 = n7211 & n7212;
  assign n7214 = n5679 & ~n7213;
  assign n7215 = n7205 & ~n7214;
  assign n7216 = ~n7197 & ~n7212;
  assign n7217 = n7211 & ~n7216;
  assign n7218 = ~n5668 & ~n7217;
  assign n7219 = n7197 & ~n7212;
  assign n7220 = n7202 & n7219;
  assign n7221 = n7194 & n7196;
  assign n7222 = n5679 & ~n7221;
  assign n7223 = ~n7218 & ~n7220;
  assign n7224 = ~n7222 & n7223;
  assign n7225 = ~n7215 & n7224;
  assign n7226 = n7215 & ~n7224;
  assign n7227 = ~n7225 & ~n7226;
  assign n7228 = ~n5648 & ~n7217;
  assign n7229 = n5648 & n7219;
  assign n7230 = n5662 & ~n7221;
  assign n7231 = ~n7228 & ~n7229;
  assign n7232 = ~n7230 & n7231;
  assign n7233 = ~n5648 & ~n7199;
  assign n7234 = n5648 & n7203;
  assign n7235 = ~n7233 & ~n7234;
  assign n7236 = n5662 & ~n7213;
  assign n7237 = n7235 & ~n7236;
  assign n7238 = n7227 & n7232;
  assign n7239 = ~n7237 & n7238;
  assign n7240 = n3574 & n7187;
  assign n7241 = n7224 & n7240;
  assign n7242 = ~n7215 & n7241;
  assign n7243 = ~n7224 & ~n7240;
  assign n7244 = n7215 & n7243;
  assign n7245 = ~n7242 & ~n7244;
  assign n7246 = ~n7232 & n7237;
  assign n7247 = n5601 & ~n7213;
  assign n7248 = ~n5550 & n7203;
  assign n7249 = ~n5550 & ~n7199;
  assign n7250 = ~n3574 & ~n7249;
  assign n7251 = ~n7247 & ~n7248;
  assign n7252 = n7250 & n7251;
  assign n7253 = n5601 & ~n7221;
  assign n7254 = ~n5550 & n7219;
  assign n7255 = ~n7253 & ~n7254;
  assign n7256 = ~n5550 & ~n7217;
  assign n7257 = n3574 & ~n5493;
  assign n7258 = n7255 & ~n7256;
  assign n7259 = ~n7257 & n7258;
  assign n7260 = n7227 & ~n7246;
  assign n7261 = ~n7252 & n7260;
  assign n7262 = n7259 & n7261;
  assign n7263 = ~n7239 & n7245;
  assign n7264 = ~n7262 & n7263;
  assign n7265 = n5478 & ~n7213;
  assign n7266 = ~n5433 & n7203;
  assign n7267 = ~n5433 & ~n7199;
  assign n7268 = ~n3574 & ~n7267;
  assign n7269 = ~n7265 & ~n7266;
  assign n7270 = n7268 & n7269;
  assign n7271 = n3574 & ~n5376;
  assign n7272 = ~n5433 & ~n7217;
  assign n7273 = n5478 & ~n7221;
  assign n7274 = ~n5433 & n7219;
  assign n7275 = ~n7273 & ~n7274;
  assign n7276 = ~n7271 & ~n7272;
  assign n7277 = n7275 & n7276;
  assign n7278 = ~n7270 & n7277;
  assign n7279 = n3574 & ~n5433;
  assign n7280 = ~n5493 & ~n7217;
  assign n7281 = n5537 & ~n7221;
  assign n7282 = ~n5493 & n7219;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 = ~n7279 & ~n7280;
  assign n7285 = n7283 & n7284;
  assign n7286 = ~n7278 & ~n7285;
  assign n7287 = n3574 & ~n5312;
  assign n7288 = ~n5376 & ~n7217;
  assign n7289 = n5418 & ~n7221;
  assign n7290 = ~n5376 & n7219;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n7287 & ~n7288;
  assign n7293 = n7291 & n7292;
  assign n7294 = n5418 & ~n7213;
  assign n7295 = ~n5376 & n7203;
  assign n7296 = ~n5376 & ~n7199;
  assign n7297 = ~n3574 & ~n7296;
  assign n7298 = ~n7294 & ~n7295;
  assign n7299 = n7297 & n7298;
  assign n7300 = ~n7293 & n7299;
  assign n7301 = n7270 & ~n7277;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = n5361 & ~n7213;
  assign n7304 = ~n5312 & n7203;
  assign n7305 = ~n5312 & ~n7199;
  assign n7306 = ~n3574 & ~n7305;
  assign n7307 = ~n7303 & ~n7304;
  assign n7308 = n7306 & n7307;
  assign n7309 = n3574 & ~n5253;
  assign n7310 = ~n5312 & ~n7217;
  assign n7311 = n5361 & ~n7221;
  assign n7312 = ~n5312 & n7219;
  assign n7313 = ~n7311 & ~n7312;
  assign n7314 = ~n7309 & ~n7310;
  assign n7315 = n7313 & n7314;
  assign n7316 = ~n7308 & n7315;
  assign n7317 = n7293 & ~n7299;
  assign n7318 = ~n7316 & ~n7317;
  assign n7319 = n3574 & ~n5191;
  assign n7320 = ~n5253 & ~n7217;
  assign n7321 = n5297 & ~n7221;
  assign n7322 = ~n5253 & n7219;
  assign n7323 = ~n7321 & ~n7322;
  assign n7324 = ~n7319 & ~n7320;
  assign n7325 = n7323 & n7324;
  assign n7326 = n5297 & ~n7213;
  assign n7327 = ~n5253 & n7203;
  assign n7328 = ~n5253 & ~n7199;
  assign n7329 = ~n3574 & ~n7328;
  assign n7330 = ~n7326 & ~n7327;
  assign n7331 = n7329 & n7330;
  assign n7332 = ~n7325 & n7331;
  assign n7333 = n7308 & ~n7315;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = n5238 & ~n7213;
  assign n7336 = ~n5191 & n7203;
  assign n7337 = ~n5191 & ~n7199;
  assign n7338 = ~n3574 & ~n7337;
  assign n7339 = ~n7335 & ~n7336;
  assign n7340 = n7338 & n7339;
  assign n7341 = n3574 & ~n5132;
  assign n7342 = ~n5191 & ~n7217;
  assign n7343 = n5238 & ~n7221;
  assign n7344 = ~n5191 & n7219;
  assign n7345 = ~n7343 & ~n7344;
  assign n7346 = ~n7341 & ~n7342;
  assign n7347 = n7345 & n7346;
  assign n7348 = ~n7340 & n7347;
  assign n7349 = n7325 & ~n7331;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = n3574 & ~n5073;
  assign n7352 = ~n5132 & ~n7217;
  assign n7353 = n5176 & ~n7221;
  assign n7354 = ~n5132 & n7219;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = ~n7351 & ~n7352;
  assign n7357 = n7355 & n7356;
  assign n7358 = n5176 & ~n7213;
  assign n7359 = ~n5132 & n7203;
  assign n7360 = ~n5132 & ~n7199;
  assign n7361 = ~n3574 & ~n7360;
  assign n7362 = ~n7358 & ~n7359;
  assign n7363 = n7361 & n7362;
  assign n7364 = ~n7357 & n7363;
  assign n7365 = n7340 & ~n7347;
  assign n7366 = ~n7364 & ~n7365;
  assign n7367 = n5117 & ~n7213;
  assign n7368 = ~n5073 & n7203;
  assign n7369 = ~n5073 & ~n7199;
  assign n7370 = ~n3574 & ~n7369;
  assign n7371 = ~n7367 & ~n7368;
  assign n7372 = n7370 & n7371;
  assign n7373 = n3574 & ~n5013;
  assign n7374 = ~n5073 & ~n7217;
  assign n7375 = n5117 & ~n7221;
  assign n7376 = ~n5073 & n7219;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = ~n7373 & ~n7374;
  assign n7379 = n7377 & n7378;
  assign n7380 = ~n7372 & n7379;
  assign n7381 = n7357 & ~n7363;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = n3574 & ~n4967;
  assign n7384 = ~n5013 & ~n7217;
  assign n7385 = n5057 & ~n7221;
  assign n7386 = ~n5013 & n7219;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = ~n7383 & ~n7384;
  assign n7389 = n7387 & n7388;
  assign n7390 = n5057 & ~n7213;
  assign n7391 = ~n5013 & n7203;
  assign n7392 = ~n5013 & ~n7199;
  assign n7393 = ~n3574 & ~n7392;
  assign n7394 = ~n7390 & ~n7391;
  assign n7395 = n7393 & n7394;
  assign n7396 = ~n7389 & n7395;
  assign n7397 = n7372 & ~n7379;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = ~n4998 & ~n7213;
  assign n7400 = ~n4967 & n7203;
  assign n7401 = ~n4967 & ~n7199;
  assign n7402 = ~n3574 & ~n7401;
  assign n7403 = ~n7399 & ~n7400;
  assign n7404 = n7402 & n7403;
  assign n7405 = n3574 & ~n4895;
  assign n7406 = ~n4967 & ~n7217;
  assign n7407 = ~n4998 & ~n7221;
  assign n7408 = ~n4967 & n7219;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = ~n7405 & ~n7406;
  assign n7411 = n7409 & n7410;
  assign n7412 = ~n7404 & n7411;
  assign n7413 = n7389 & ~n7395;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = n3574 & ~n4813;
  assign n7416 = ~n4895 & ~n7217;
  assign n7417 = ~n4934 & ~n7221;
  assign n7418 = ~n4895 & n7219;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = ~n7415 & ~n7416;
  assign n7421 = n7419 & n7420;
  assign n7422 = ~n4934 & ~n7213;
  assign n7423 = ~n4895 & n7203;
  assign n7424 = ~n4895 & ~n7199;
  assign n7425 = ~n3574 & ~n7424;
  assign n7426 = ~n7422 & ~n7423;
  assign n7427 = n7425 & n7426;
  assign n7428 = ~n7421 & n7427;
  assign n7429 = n7404 & ~n7411;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~n4865 & ~n7213;
  assign n7432 = ~n4813 & n7203;
  assign n7433 = ~n4813 & ~n7199;
  assign n7434 = ~n3574 & ~n7433;
  assign n7435 = ~n7431 & ~n7432;
  assign n7436 = n7434 & n7435;
  assign n7437 = n3574 & ~n4752;
  assign n7438 = ~n4813 & ~n7217;
  assign n7439 = ~n4865 & ~n7221;
  assign n7440 = ~n4813 & n7219;
  assign n7441 = ~n7439 & ~n7440;
  assign n7442 = ~n7437 & ~n7438;
  assign n7443 = n7441 & n7442;
  assign n7444 = ~n7436 & n7443;
  assign n7445 = n7421 & ~n7427;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = n3574 & ~n4703;
  assign n7448 = ~n4752 & ~n7217;
  assign n7449 = ~n4798 & ~n7221;
  assign n7450 = ~n4752 & n7219;
  assign n7451 = ~n7449 & ~n7450;
  assign n7452 = ~n7447 & ~n7448;
  assign n7453 = n7451 & n7452;
  assign n7454 = ~n4798 & ~n7213;
  assign n7455 = ~n4752 & n7203;
  assign n7456 = ~n4752 & ~n7199;
  assign n7457 = ~n3574 & ~n7456;
  assign n7458 = ~n7454 & ~n7455;
  assign n7459 = n7457 & n7458;
  assign n7460 = ~n7453 & n7459;
  assign n7461 = n7436 & ~n7443;
  assign n7462 = ~n7460 & ~n7461;
  assign n7463 = ~n4737 & ~n7213;
  assign n7464 = ~n4703 & n7203;
  assign n7465 = ~n4703 & ~n7199;
  assign n7466 = ~n3574 & ~n7465;
  assign n7467 = ~n7463 & ~n7464;
  assign n7468 = n7466 & n7467;
  assign n7469 = n3574 & ~n4639;
  assign n7470 = ~n4703 & ~n7217;
  assign n7471 = ~n4737 & ~n7221;
  assign n7472 = ~n4703 & n7219;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = ~n7469 & ~n7470;
  assign n7475 = n7473 & n7474;
  assign n7476 = ~n7468 & n7475;
  assign n7477 = n7453 & ~n7459;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = n3574 & ~n4570;
  assign n7480 = ~n4639 & ~n7217;
  assign n7481 = ~n4673 & ~n7221;
  assign n7482 = ~n4639 & n7219;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n7479 & ~n7480;
  assign n7485 = n7483 & n7484;
  assign n7486 = ~n4673 & ~n7213;
  assign n7487 = ~n4639 & n7203;
  assign n7488 = ~n4639 & ~n7199;
  assign n7489 = ~n3574 & ~n7488;
  assign n7490 = ~n7486 & ~n7487;
  assign n7491 = n7489 & n7490;
  assign n7492 = ~n7485 & n7491;
  assign n7493 = n7468 & ~n7475;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~n4609 & ~n7213;
  assign n7496 = ~n4570 & n7203;
  assign n7497 = ~n4570 & ~n7199;
  assign n7498 = ~n3574 & ~n7497;
  assign n7499 = ~n7495 & ~n7496;
  assign n7500 = n7498 & n7499;
  assign n7501 = n3574 & ~n4505;
  assign n7502 = ~n4570 & ~n7217;
  assign n7503 = ~n4609 & ~n7221;
  assign n7504 = ~n4570 & n7219;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n7501 & ~n7502;
  assign n7507 = n7505 & n7506;
  assign n7508 = ~n7500 & n7507;
  assign n7509 = n7485 & ~n7491;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = n3574 & ~n4423;
  assign n7512 = ~n4505 & ~n7217;
  assign n7513 = ~n4542 & ~n7221;
  assign n7514 = ~n4505 & n7219;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7511 & ~n7512;
  assign n7517 = n7515 & n7516;
  assign n7518 = ~n4542 & ~n7213;
  assign n7519 = ~n4505 & n7203;
  assign n7520 = ~n4505 & ~n7199;
  assign n7521 = ~n3574 & ~n7520;
  assign n7522 = ~n7518 & ~n7519;
  assign n7523 = n7521 & n7522;
  assign n7524 = ~n7517 & n7523;
  assign n7525 = n7500 & ~n7507;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = ~n4472 & ~n7213;
  assign n7528 = ~n4423 & n7203;
  assign n7529 = ~n4423 & ~n7199;
  assign n7530 = ~n3574 & ~n7529;
  assign n7531 = ~n7527 & ~n7528;
  assign n7532 = n7530 & n7531;
  assign n7533 = n3574 & ~n4355;
  assign n7534 = ~n4423 & ~n7217;
  assign n7535 = ~n4472 & ~n7221;
  assign n7536 = ~n4423 & n7219;
  assign n7537 = ~n7535 & ~n7536;
  assign n7538 = ~n7533 & ~n7534;
  assign n7539 = n7537 & n7538;
  assign n7540 = ~n7532 & n7539;
  assign n7541 = n7517 & ~n7523;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = n3574 & ~n4287;
  assign n7544 = ~n4355 & ~n7217;
  assign n7545 = ~n4407 & ~n7221;
  assign n7546 = ~n4355 & n7219;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = ~n7543 & ~n7544;
  assign n7549 = n7547 & n7548;
  assign n7550 = ~n4407 & ~n7213;
  assign n7551 = ~n4355 & n7203;
  assign n7552 = ~n4355 & ~n7199;
  assign n7553 = ~n3574 & ~n7552;
  assign n7554 = ~n7550 & ~n7551;
  assign n7555 = n7553 & n7554;
  assign n7556 = ~n7549 & n7555;
  assign n7557 = n7532 & ~n7539;
  assign n7558 = ~n7556 & ~n7557;
  assign n7559 = ~n4340 & ~n7213;
  assign n7560 = ~n4287 & n7203;
  assign n7561 = ~n3574 & ~n7560;
  assign n7562 = ~n4287 & ~n7199;
  assign n7563 = n7561 & ~n7562;
  assign n7564 = ~n7559 & n7563;
  assign n7565 = n3574 & ~n4219;
  assign n7566 = ~n4287 & n7219;
  assign n7567 = ~n7565 & ~n7566;
  assign n7568 = ~n4287 & ~n7217;
  assign n7569 = ~n4340 & ~n7221;
  assign n7570 = n7567 & ~n7568;
  assign n7571 = ~n7569 & n7570;
  assign n7572 = ~n7564 & n7571;
  assign n7573 = n7549 & ~n7555;
  assign n7574 = ~n7572 & ~n7573;
  assign n7575 = n3574 & ~n4146;
  assign n7576 = ~n4219 & n7219;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = ~n4219 & ~n7217;
  assign n7579 = ~n4272 & ~n7221;
  assign n7580 = n7577 & ~n7578;
  assign n7581 = ~n7579 & n7580;
  assign n7582 = ~n4272 & ~n7213;
  assign n7583 = ~n4219 & n7203;
  assign n7584 = ~n3574 & ~n7583;
  assign n7585 = ~n4219 & ~n7199;
  assign n7586 = n7584 & ~n7585;
  assign n7587 = ~n7582 & n7586;
  assign n7588 = ~n7581 & n7587;
  assign n7589 = n7564 & ~n7571;
  assign n7590 = ~n7588 & ~n7589;
  assign n7591 = ~n4204 & ~n7213;
  assign n7592 = ~n4146 & n7203;
  assign n7593 = ~n3574 & ~n7592;
  assign n7594 = ~n4146 & ~n7199;
  assign n7595 = n7593 & ~n7594;
  assign n7596 = ~n7591 & n7595;
  assign n7597 = n3574 & ~n4081;
  assign n7598 = ~n4146 & ~n7217;
  assign n7599 = ~n4204 & ~n7221;
  assign n7600 = ~n4146 & n7219;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = ~n7597 & ~n7598;
  assign n7603 = n7601 & n7602;
  assign n7604 = ~n7596 & n7603;
  assign n7605 = n7581 & ~n7587;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = n3574 & ~n4011;
  assign n7608 = ~n4081 & ~n7217;
  assign n7609 = ~n4130 & ~n7221;
  assign n7610 = ~n4081 & n7219;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = ~n7607 & ~n7608;
  assign n7613 = n7611 & n7612;
  assign n7614 = ~n4130 & ~n7213;
  assign n7615 = ~n4081 & n7203;
  assign n7616 = ~n3574 & ~n7615;
  assign n7617 = ~n4081 & ~n7199;
  assign n7618 = n7616 & ~n7617;
  assign n7619 = ~n7614 & n7618;
  assign n7620 = ~n7613 & n7619;
  assign n7621 = n7596 & ~n7603;
  assign n7622 = ~n7620 & ~n7621;
  assign n7623 = ~n4066 & ~n7213;
  assign n7624 = ~n4011 & n7203;
  assign n7625 = ~n3574 & ~n7624;
  assign n7626 = ~n4011 & ~n7199;
  assign n7627 = n7625 & ~n7626;
  assign n7628 = ~n7623 & n7627;
  assign n7629 = n3574 & ~n3945;
  assign n7630 = ~n4011 & ~n7217;
  assign n7631 = ~n4066 & ~n7221;
  assign n7632 = ~n4011 & n7219;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = ~n7629 & ~n7630;
  assign n7635 = n7633 & n7634;
  assign n7636 = ~n7628 & n7635;
  assign n7637 = n7613 & ~n7619;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = n3574 & ~n3881;
  assign n7640 = ~n3945 & ~n7217;
  assign n7641 = ~n3996 & ~n7221;
  assign n7642 = ~n3945 & n7219;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7639 & ~n7640;
  assign n7645 = n7643 & n7644;
  assign n7646 = ~n3996 & ~n7213;
  assign n7647 = ~n3945 & n7203;
  assign n7648 = ~n3574 & ~n7647;
  assign n7649 = ~n3945 & ~n7199;
  assign n7650 = n7648 & ~n7649;
  assign n7651 = ~n7646 & n7650;
  assign n7652 = ~n7645 & n7651;
  assign n7653 = n7628 & ~n7635;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~n3931 & ~n7213;
  assign n7656 = ~n3881 & n7203;
  assign n7657 = ~n3574 & ~n7656;
  assign n7658 = ~n3881 & ~n7199;
  assign n7659 = n7657 & ~n7658;
  assign n7660 = ~n7655 & n7659;
  assign n7661 = ~n3931 & ~n7221;
  assign n7662 = ~n3881 & n7219;
  assign n7663 = n3574 & ~n3824;
  assign n7664 = ~n7661 & ~n7662;
  assign n7665 = ~n7663 & n7664;
  assign n7666 = ~n3881 & ~n7217;
  assign n7667 = n7665 & ~n7666;
  assign n7668 = ~n7660 & n7667;
  assign n7669 = n7645 & ~n7651;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n3869 & ~n7221;
  assign n7672 = ~n3824 & n7219;
  assign n7673 = n3574 & ~n3759;
  assign n7674 = ~n7671 & ~n7672;
  assign n7675 = ~n7673 & n7674;
  assign n7676 = ~n3824 & ~n7217;
  assign n7677 = n7675 & ~n7676;
  assign n7678 = ~n3869 & ~n7213;
  assign n7679 = ~n3824 & n7203;
  assign n7680 = ~n3574 & ~n7679;
  assign n7681 = ~n3824 & ~n7199;
  assign n7682 = n7680 & ~n7681;
  assign n7683 = ~n7678 & n7682;
  assign n7684 = ~n7677 & n7683;
  assign n7685 = n7660 & ~n7667;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = ~n3813 & ~n7213;
  assign n7688 = ~n3759 & n7203;
  assign n7689 = ~n3574 & ~n7688;
  assign n7690 = ~n3759 & ~n7199;
  assign n7691 = n7689 & ~n7690;
  assign n7692 = ~n7687 & n7691;
  assign n7693 = ~n3813 & ~n7221;
  assign n7694 = ~n3759 & n7219;
  assign n7695 = n3574 & ~n3767;
  assign n7696 = ~n7693 & ~n7694;
  assign n7697 = ~n7695 & n7696;
  assign n7698 = ~n3759 & ~n7217;
  assign n7699 = n7697 & ~n7698;
  assign n7700 = ~n7692 & n7699;
  assign n7701 = n7677 & ~n7683;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = ~n3733 & ~n7213;
  assign n7704 = ~n3767 & n7203;
  assign n7705 = ~n3574 & ~n7704;
  assign n7706 = ~n3767 & ~n7199;
  assign n7707 = n7705 & ~n7706;
  assign n7708 = ~n7703 & n7707;
  assign n7709 = ~n3646 & n3649;
  assign n7710 = ~n3574 & ~n7709;
  assign n7711 = n7221 & n7710;
  assign n7712 = n7708 & n7711;
  assign n7713 = n7692 & ~n7699;
  assign n7714 = ~n3733 & ~n7221;
  assign n7715 = ~n3767 & n7219;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = ~n3767 & ~n7217;
  assign n7718 = n7716 & ~n7717;
  assign n7719 = ~n7708 & ~n7711;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = ~n7712 & ~n7713;
  assign n7722 = ~n7720 & n7721;
  assign n7723 = n7702 & ~n7722;
  assign n7724 = n7686 & ~n7723;
  assign n7725 = n7670 & ~n7724;
  assign n7726 = n7654 & ~n7725;
  assign n7727 = n7638 & ~n7726;
  assign n7728 = n7622 & ~n7727;
  assign n7729 = n7606 & ~n7728;
  assign n7730 = n7590 & ~n7729;
  assign n7731 = n7574 & ~n7730;
  assign n7732 = n7558 & ~n7731;
  assign n7733 = n7542 & ~n7732;
  assign n7734 = n7526 & ~n7733;
  assign n7735 = n7510 & ~n7734;
  assign n7736 = n7494 & ~n7735;
  assign n7737 = n7478 & ~n7736;
  assign n7738 = n7462 & ~n7737;
  assign n7739 = n7446 & ~n7738;
  assign n7740 = n7430 & ~n7739;
  assign n7741 = n7414 & ~n7740;
  assign n7742 = n7398 & ~n7741;
  assign n7743 = n7382 & ~n7742;
  assign n7744 = n7366 & ~n7743;
  assign n7745 = n7350 & ~n7744;
  assign n7746 = n7334 & ~n7745;
  assign n7747 = n7318 & ~n7746;
  assign n7748 = n7302 & ~n7747;
  assign n7749 = n7286 & ~n7748;
  assign n7750 = n5537 & ~n7213;
  assign n7751 = ~n5493 & n7203;
  assign n7752 = ~n5493 & ~n7199;
  assign n7753 = ~n3574 & ~n7752;
  assign n7754 = ~n7750 & ~n7751;
  assign n7755 = n7753 & n7754;
  assign n7756 = ~n7285 & n7755;
  assign n7757 = n7252 & ~n7259;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = ~n7278 & n7755;
  assign n7760 = ~n7748 & n7759;
  assign n7761 = n7260 & ~n7749;
  assign n7762 = n7758 & n7761;
  assign n7763 = ~n7760 & n7762;
  assign n7764 = n7264 & ~n7763;
  assign n7765 = n3587 & n7188;
  assign n7766 = n7764 & n7765;
  assign n7767 = ~n7193 & ~n7766;
  assign n7768 = n5376 & ~n5418;
  assign n7769 = ~n5437 & ~n7768;
  assign n7770 = ~n5387 & ~n7769;
  assign n7771 = ~n5256 & ~n5257;
  assign n7772 = ~n5194 & ~n5198;
  assign n7773 = ~n5315 & ~n5316;
  assign n7774 = ~n7771 & ~n7772;
  assign n7775 = ~n7773 & n7774;
  assign n7776 = ~n5325 & n7775;
  assign n7777 = n7770 & n7776;
  assign n7778 = ~n4084 & ~n4085;
  assign n7779 = ~n3886 & ~n3958;
  assign n7780 = ~n7778 & n7779;
  assign n7781 = ~n4222 & ~n4223;
  assign n7782 = ~n4165 & ~n7781;
  assign n7783 = ~n4552 & n7782;
  assign n7784 = n7780 & n7783;
  assign n7785 = ~n4826 & n7784;
  assign n7786 = n3733 & n3767;
  assign n7787 = ~n3830 & ~n7786;
  assign n7788 = ~n4755 & ~n4756;
  assign n7789 = ~n3829 & ~n7787;
  assign n7790 = ~n7788 & n7789;
  assign n7791 = ~n4615 & ~n4616;
  assign n7792 = ~n4302 & ~n4366;
  assign n7793 = ~n7791 & n7792;
  assign n7794 = ~n4819 & ~n4820;
  assign n7795 = n7790 & n7793;
  assign n7796 = ~n7794 & n7795;
  assign n7797 = ~n4867 & ~n4869;
  assign n7798 = ~n5553 & ~n5559;
  assign n7799 = n7785 & n7796;
  assign n7800 = ~n7797 & n7799;
  assign n7801 = ~n4948 & n7800;
  assign n7802 = ~n7798 & n7801;
  assign n7803 = ~n4426 & ~n4427;
  assign n7804 = n5550 & ~n5601;
  assign n7805 = ~n5550 & n5601;
  assign n7806 = ~n7804 & ~n7805;
  assign n7807 = ~n4025 & ~n7803;
  assign n7808 = ~n4491 & n7807;
  assign n7809 = ~n5024 & n7808;
  assign n7810 = ~n7806 & n7809;
  assign n7811 = ~n5076 & ~n5078;
  assign n7812 = n5668 & ~n5679;
  assign n7813 = ~n5668 & n5679;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = n5648 & ~n5662;
  assign n7816 = ~n5648 & n5662;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = ~n7811 & ~n7814;
  assign n7819 = ~n7817 & n7818;
  assign n7820 = n5493 & ~n5537;
  assign n7821 = ~n5609 & ~n7820;
  assign n7822 = n7810 & n7819;
  assign n7823 = ~n7821 & n7822;
  assign n7824 = n7777 & n7802;
  assign n7825 = n7823 & n7824;
  assign n7826 = n3736 & n7825;
  assign n7827 = n3734 & ~n7825;
  assign n7828 = n3741 & ~n7764;
  assign n7829 = n3643 & ~n3646;
  assign n7830 = n7764 & n7829;
  assign n7831 = ~n7828 & ~n7830;
  assign n7832 = ~n7826 & ~n7827;
  assign n7833 = n7831 & n7832;
  assign n7834 = ~n3649 & ~n7833;
  assign n7835 = ~n3652 & ~n5812;
  assign n7836 = n7764 & ~n7835;
  assign n7837 = n3649 & n7836;
  assign n7838 = ~n3775_1 & ~n3784;
  assign n7839 = ~n7764 & ~n7838;
  assign n7840 = ~n7834 & ~n7837;
  assign n7841 = ~n7839 & n7840;
  assign n7842 = n6206 & ~n7841;
  assign n1170 = ~n7767 | n7842;
  assign n7844 = ~n6206 & ~n1330;
  assign n7845 = n3646 & n3790;
  assign n7846 = ~n5798 & ~n7195;
  assign n7847 = ~n3646 & ~n7846;
  assign n7848 = ~n3779 & ~n5788;
  assign n7849 = n3643 & n5812;
  assign n7850 = ~n3785 & ~n7207;
  assign n7851 = ~n7849 & n7850;
  assign n7852 = ~n7845 & ~n7847;
  assign n7853 = n7848 & n7852;
  assign n7854 = n7851 & n7853;
  assign n7855 = ~n3636 & ~n3640_1;
  assign n7856 = n3718 & n7855;
  assign n7857 = ~n7854 & ~n7856;
  assign n7858 = ~n5790 & ~n7857;
  assign n7859 = n3587 & ~n7858;
  assign n7860 = n7844 & ~n7859;
  assign n7861 = n3587 & ~n5800;
  assign n7862 = ~n7856 & n7861;
  assign n7863 = n7860 & ~n7862;
  assign n7864 = ~n4699 & ~n7863;
  assign n7865 = n7856 & n7861;
  assign n7866 = n3587 & n5789;
  assign n7867 = ~n7865 & ~n7866;
  assign n7868 = ~n4737 & ~n7867;
  assign n7869 = P1_STATE_REG & ~n3586;
  assign n7870 = n7240 & n7869;
  assign n7871 = ~n4699 & ~n7856;
  assign n7872 = ~n3726 & n7856;
  assign n7873 = ~n4639 & n7872;
  assign n7874 = n3726 & n7856;
  assign n7875 = ~n4752 & n7874;
  assign n7876 = ~n7871 & ~n7873;
  assign n7877 = ~n7875 & n7876;
  assign n7878 = n7870 & ~n7877;
  assign n7879 = ~n4639 & ~n6945;
  assign n7880 = ~n4673 & n6938;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = ~n4639 & n6938;
  assign n7883 = ~n4673 & ~n6954;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = ~n6935 & ~n7884;
  assign n7886 = n6935 & n7884;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = ~n7881 & ~n7887;
  assign n7889 = n7881 & n7887;
  assign n7890 = ~n4570 & n6938;
  assign n7891 = ~n4609 & ~n6954;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = ~n6935 & ~n7892;
  assign n7894 = n6935 & n7892;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = ~n4570 & ~n6945;
  assign n7897 = ~n4609 & n6938;
  assign n7898 = ~n7896 & ~n7897;
  assign n7899 = n7895 & n7898;
  assign n7900 = ~n7895 & ~n7898;
  assign n7901 = ~n4505 & ~n6945;
  assign n7902 = ~n4542 & n6938;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = ~n4505 & n6938;
  assign n7905 = ~n4542 & ~n6954;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = ~n6935 & ~n7906;
  assign n7908 = n6935 & n7906;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~n7903 & ~n7909;
  assign n7911 = ~n7900 & ~n7910;
  assign n7912 = ~n4423 & ~n6945;
  assign n7913 = ~n4472 & n6938;
  assign n7914 = ~n7912 & ~n7913;
  assign n7915 = ~n4423 & n6938;
  assign n7916 = ~n4472 & ~n6954;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = ~n6935 & ~n7917;
  assign n7919 = n6935 & n7917;
  assign n7920 = ~n7918 & ~n7919;
  assign n7921 = ~n7914 & ~n7920;
  assign n7922 = n7903 & n7909;
  assign n7923 = ~n7899 & ~n7922;
  assign n7924 = n7921 & n7923;
  assign n7925 = n7911 & ~n7924;
  assign n7926 = ~n7899 & ~n7925;
  assign n7927 = n7914 & n7920;
  assign n7928 = n7923 & ~n7927;
  assign n7929 = ~n4355 & ~n6945;
  assign n7930 = ~n4407 & n6938;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = ~n4355 & n6938;
  assign n7933 = ~n4407 & ~n6954;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = ~n6935 & ~n7934;
  assign n7936 = n6935 & n7934;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = ~n7931 & ~n7937;
  assign n7939 = n7931 & n7937;
  assign n7940 = ~n4287 & ~n6945;
  assign n7941 = ~n4340 & n6938;
  assign n7942 = ~n7940 & ~n7941;
  assign n7943 = ~n4219 & ~n6945;
  assign n7944 = ~n4272 & n6938;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = ~n4219 & n6938;
  assign n7947 = ~n4272 & ~n6954;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n6935 & ~n7948;
  assign n7950 = n6935 & n7948;
  assign n7951 = ~n7949 & ~n7950;
  assign n7952 = ~n7945 & ~n7951;
  assign n7953 = n7945 & n7951;
  assign n7954 = ~n4146 & ~n6945;
  assign n7955 = ~n4204 & n6938;
  assign n7956 = ~n7954 & ~n7955;
  assign n7957 = ~n4081 & ~n6945;
  assign n7958 = ~n4130 & n6938;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = ~n4081 & n6938;
  assign n7961 = ~n4130 & ~n6954;
  assign n7962 = ~n7960 & ~n7961;
  assign n7963 = ~n6935 & ~n7962;
  assign n7964 = n6935 & n7962;
  assign n7965 = ~n7963 & ~n7964;
  assign n7966 = ~n7959 & ~n7965;
  assign n7967 = ~n7956 & n7966;
  assign n7968 = ~n4146 & n6938;
  assign n7969 = ~n4204 & ~n6954;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = ~n6935 & ~n7970;
  assign n7972 = n6935 & n7970;
  assign n7973 = ~n7971 & ~n7972;
  assign n7974 = n7956 & ~n7966;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = ~n7967 & ~n7975;
  assign n7977 = n7959 & n7965;
  assign n7978 = n7956 & n7973;
  assign n7979 = ~n7977 & ~n7978;
  assign n7980 = ~n4011 & ~n6945;
  assign n7981 = ~n4066 & n6938;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = ~n4011 & n6938;
  assign n7984 = ~n4066 & ~n6954;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = ~n6935 & ~n7985;
  assign n7987 = n6935 & n7985;
  assign n7988 = ~n7986 & ~n7987;
  assign n7989 = ~n7982 & ~n7988;
  assign n7990 = n7982 & n7988;
  assign n7991 = ~n3945 & ~n6945;
  assign n7992 = ~n3996 & n6938;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = ~n3881 & ~n6945;
  assign n7995 = ~n3931 & n6938;
  assign n7996 = ~n7994 & ~n7995;
  assign n7997 = ~n3824 & ~n6945;
  assign n7998 = ~n3869 & n6938;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = ~n3824 & n6938;
  assign n8001 = ~n3869 & ~n6954;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = ~n6935 & ~n8002;
  assign n8004 = n6935 & n8002;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = ~n7999 & ~n8005;
  assign n8007 = ~n7996 & n8006;
  assign n8008 = ~n3881 & n6938;
  assign n8009 = ~n3931 & ~n6954;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = ~n6935 & ~n8010;
  assign n8012 = n6935 & n8010;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = n7996 & ~n8006;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~n8007 & ~n8015;
  assign n8017 = n7999 & n8005;
  assign n8018 = n7996 & n8013;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~n3759 & ~n6945;
  assign n8021 = ~n3813 & n6938;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = ~n3759 & n6938;
  assign n8024 = ~n3813 & ~n6954;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n6935 & ~n8025;
  assign n8027 = n6935 & n8025;
  assign n8028 = ~n8026 & ~n8027;
  assign n8029 = ~n8022 & ~n8028;
  assign n8030 = n8022 & n8028;
  assign n8031 = n6935 & ~n6947;
  assign n8032 = ~n6935 & n6947;
  assign n8033 = ~n6959 & ~n8032;
  assign n8034 = ~n8031 & ~n8033;
  assign n8035 = ~n8030 & ~n8034;
  assign n8036 = ~n8029 & ~n8035;
  assign n8037 = n8019 & ~n8036;
  assign n8038 = n8016 & ~n8037;
  assign n8039 = ~n7993 & ~n8038;
  assign n8040 = ~n3945 & n6938;
  assign n8041 = ~n3996 & ~n6954;
  assign n8042 = ~n8040 & ~n8041;
  assign n8043 = ~n6935 & ~n8042;
  assign n8044 = n6935 & n8042;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = n7993 & n8038;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = ~n8039 & ~n8047;
  assign n8049 = ~n7990 & ~n8048;
  assign n8050 = ~n7989 & ~n8049;
  assign n8051 = n7979 & ~n8050;
  assign n8052 = n7976 & ~n8051;
  assign n8053 = ~n7953 & ~n8052;
  assign n8054 = ~n7952 & ~n8053;
  assign n8055 = ~n7942 & ~n8054;
  assign n8056 = ~n4287 & n6938;
  assign n8057 = ~n4340 & ~n6954;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = ~n6935 & ~n8058;
  assign n8060 = n6935 & n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = n7942 & n8054;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n8055 & ~n8063;
  assign n8065 = ~n7939 & ~n8064;
  assign n8066 = ~n7938 & ~n8065;
  assign n8067 = n7928 & ~n8066;
  assign n8068 = ~n7926 & ~n8067;
  assign n8069 = ~n7889 & ~n8068;
  assign n8070 = ~n7888 & ~n8069;
  assign n8071 = ~n4703 & n6938;
  assign n8072 = ~n4737 & ~n6954;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n6935 & ~n8073;
  assign n8075 = n6935 & n8073;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~n4703 & ~n6945;
  assign n8078 = ~n4737 & n6938;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = ~n8076 & n8079;
  assign n8081 = n8076 & ~n8079;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = n8070 & ~n8082;
  assign n8084 = ~n8070 & n8082;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = n3587 & ~n7854;
  assign n8087 = n7856 & n8086;
  assign n8088 = ~n8085 & n8087;
  assign n8089 = ~n7864 & ~n7868;
  assign n8090 = ~n6536 & n8089;
  assign n8091 = ~n7878 & n8090;
  assign n1175 = n8088 | ~n8091;
  assign n8093 = ~n5372 & ~n7863;
  assign n8094 = ~n5800 & n7856;
  assign n8095 = ~n5789 & ~n8094;
  assign n8096 = n3587 & ~n8095;
  assign n8097 = n5418 & n8096;
  assign n8098 = P1_REG3_REG_26_ & ~P1_STATE_REG;
  assign n8099 = ~n5372 & ~n7856;
  assign n8100 = ~n5312 & n7872;
  assign n8101 = ~n5433 & n7874;
  assign n8102 = ~n8099 & ~n8100;
  assign n8103 = ~n8101 & n8102;
  assign n8104 = n7870 & ~n8103;
  assign n8105 = ~n5253 & ~n6945;
  assign n8106 = n5297 & n6938;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = ~n5253 & n6938;
  assign n8109 = n5297 & ~n6954;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = ~n6935 & ~n8110;
  assign n8112 = n6935 & n8110;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = ~n8107 & ~n8113;
  assign n8115 = n8107 & n8113;
  assign n8116 = ~n5191 & ~n6945;
  assign n8117 = n5238 & n6938;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = ~n5191 & n6938;
  assign n8120 = n5238 & ~n6954;
  assign n8121 = ~n8119 & ~n8120;
  assign n8122 = ~n6935 & ~n8121;
  assign n8123 = n6935 & n8121;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~n8118 & ~n8124;
  assign n8126 = n8118 & n8124;
  assign n8127 = ~n5132 & ~n6945;
  assign n8128 = n5176 & n6938;
  assign n8129 = ~n8127 & ~n8128;
  assign n8130 = ~n5132 & n6938;
  assign n8131 = n5176 & ~n6954;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~n6935 & ~n8132;
  assign n8134 = n6935 & n8132;
  assign n8135 = ~n8133 & ~n8134;
  assign n8136 = ~n8129 & ~n8135;
  assign n8137 = n8129 & n8135;
  assign n8138 = ~n4967 & n6938;
  assign n8139 = ~n4998 & ~n6954;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n6935 & ~n8140;
  assign n8142 = n6935 & n8140;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~n4967 & ~n6945;
  assign n8145 = ~n4998 & n6938;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = n8143 & n8146;
  assign n8148 = ~n4895 & ~n6945;
  assign n8149 = ~n4934 & n6938;
  assign n8150 = ~n8148 & ~n8149;
  assign n8151 = ~n4895 & n6938;
  assign n8152 = ~n4934 & ~n6954;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = ~n6935 & ~n8153;
  assign n8155 = n6935 & n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n8150 & ~n8156;
  assign n8158 = n8150 & n8156;
  assign n8159 = ~n4813 & ~n6945;
  assign n8160 = ~n4865 & n6938;
  assign n8161 = ~n8159 & ~n8160;
  assign n8162 = ~n4752 & ~n6945;
  assign n8163 = ~n4798 & n6938;
  assign n8164 = ~n8162 & ~n8163;
  assign n8165 = ~n4752 & n6938;
  assign n8166 = ~n4798 & ~n6954;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n6935 & ~n8167;
  assign n8169 = n6935 & n8167;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = ~n8164 & ~n8170;
  assign n8172 = ~n8161 & n8171;
  assign n8173 = ~n4813 & n6938;
  assign n8174 = ~n4865 & ~n6954;
  assign n8175 = ~n8173 & ~n8174;
  assign n8176 = ~n6935 & ~n8175;
  assign n8177 = n6935 & n8175;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = n8161 & ~n8171;
  assign n8180 = ~n8178 & ~n8179;
  assign n8181 = ~n8172 & ~n8180;
  assign n8182 = n8164 & n8170;
  assign n8183 = n8161 & n8178;
  assign n8184 = ~n8182 & ~n8183;
  assign n8185 = ~n8076 & ~n8079;
  assign n8186 = n8076 & n8079;
  assign n8187 = ~n8070 & ~n8186;
  assign n8188 = ~n8185 & ~n8187;
  assign n8189 = n8184 & ~n8188;
  assign n8190 = n8181 & ~n8189;
  assign n8191 = ~n8158 & ~n8190;
  assign n8192 = ~n8157 & ~n8191;
  assign n8193 = ~n5013 & n6938;
  assign n8194 = n5057 & ~n6954;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n6935 & ~n8195;
  assign n8197 = n6935 & n8195;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = ~n5013 & ~n6945;
  assign n8200 = n5057 & n6938;
  assign n8201 = ~n8199 & ~n8200;
  assign n8202 = n8198 & n8201;
  assign n8203 = ~n5073 & n6938;
  assign n8204 = n5117 & ~n6954;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~n6935 & ~n8205;
  assign n8207 = n6935 & n8205;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = ~n5073 & ~n6945;
  assign n8210 = n5117 & n6938;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = n8208 & n8211;
  assign n8213 = ~n8202 & ~n8212;
  assign n8214 = ~n8147 & ~n8192;
  assign n8215 = n8213 & n8214;
  assign n8216 = ~n8208 & ~n8211;
  assign n8217 = ~n8198 & ~n8201;
  assign n8218 = ~n8143 & ~n8146;
  assign n8219 = n8213 & n8218;
  assign n8220 = ~n8217 & ~n8219;
  assign n8221 = ~n8212 & ~n8220;
  assign n8222 = ~n8215 & ~n8216;
  assign n8223 = ~n8221 & n8222;
  assign n8224 = ~n8137 & ~n8223;
  assign n8225 = ~n8136 & ~n8224;
  assign n8226 = ~n8126 & ~n8225;
  assign n8227 = ~n8125 & ~n8226;
  assign n8228 = ~n8115 & ~n8227;
  assign n8229 = ~n8114 & ~n8228;
  assign n8230 = ~n5312 & ~n6945;
  assign n8231 = n5361 & n6938;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = ~n5312 & n6938;
  assign n8234 = n5361 & ~n6954;
  assign n8235 = ~n8233 & ~n8234;
  assign n8236 = ~n6935 & ~n8235;
  assign n8237 = n6935 & n8235;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n8232 & ~n8238;
  assign n8240 = n8229 & ~n8239;
  assign n8241 = ~n5376 & ~n6945;
  assign n8242 = n5418 & n6938;
  assign n8243 = ~n8241 & ~n8242;
  assign n8244 = ~n5376 & n6938;
  assign n8245 = n5418 & ~n6954;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~n6935 & ~n8246;
  assign n8248 = n6935 & n8246;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = ~n8243 & ~n8249;
  assign n8251 = n8232 & n8238;
  assign n8252 = ~n8243 & ~n8251;
  assign n8253 = ~n8249 & ~n8251;
  assign n8254 = ~n8252 & ~n8253;
  assign n8255 = ~n8240 & ~n8250;
  assign n8256 = ~n8254 & n8255;
  assign n8257 = n8243 & ~n8249;
  assign n8258 = ~n8243 & n8249;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~n8239 & n8259;
  assign n8261 = ~n8229 & ~n8251;
  assign n8262 = n8260 & ~n8261;
  assign n8263 = ~n8256 & ~n8262;
  assign n8264 = n8087 & n8263;
  assign n8265 = ~n8093 & ~n8097;
  assign n8266 = ~n8098 & n8265;
  assign n8267 = ~n8104 & n8266;
  assign n1180 = n8264 | ~n8267;
  assign n8269 = ~n4074 & ~n7863;
  assign n8270 = ~n4130 & ~n7867;
  assign n8271 = ~n4146 & n7874;
  assign n8272 = ~n4011 & n7872;
  assign n8273 = ~n4074 & ~n7856;
  assign n8274 = ~n8271 & ~n8272;
  assign n8275 = ~n8273 & n8274;
  assign n8276 = n7870 & ~n8275;
  assign n8277 = ~n6831 & ~n8276;
  assign n8278 = n7959 & ~n7965;
  assign n8279 = ~n7959 & n7965;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = n8050 & ~n8280;
  assign n8282 = ~n7966 & ~n7977;
  assign n8283 = ~n8050 & ~n8282;
  assign n8284 = ~n8281 & ~n8283;
  assign n8285 = n8087 & ~n8284;
  assign n8286 = ~n8269 & ~n8270;
  assign n8287 = n8277 & n8286;
  assign n1185 = n8285 | ~n8287;
  assign n8289 = ~n4891 & ~n7863;
  assign n8290 = ~n4934 & ~n7867;
  assign n8291 = ~n4891 & ~n7856;
  assign n8292 = ~n4813 & n7872;
  assign n8293 = ~n4967 & n7874;
  assign n8294 = ~n8291 & ~n8292;
  assign n8295 = ~n8293 & n8294;
  assign n8296 = n7870 & ~n8295;
  assign n8297 = n8150 & ~n8156;
  assign n8298 = ~n8150 & n8156;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = n8190 & ~n8299;
  assign n8301 = ~n8190 & n8299;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = n8087 & ~n8302;
  assign n8304 = ~n8289 & ~n8290;
  assign n8305 = ~n6440 & n8304;
  assign n8306 = ~n8296 & n8305;
  assign n1190 = n8303 | ~n8306;
  assign n8308 = n7999 & ~n8005;
  assign n8309 = ~n7999 & n8005;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = n8036 & ~n8310;
  assign n8312 = ~n8006 & ~n8017;
  assign n8313 = ~n8036 & ~n8312;
  assign n8314 = ~n8311 & ~n8313;
  assign n8315 = n8087 & ~n8314;
  assign n8316 = ~n3869 & ~n7867;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = P1_REG3_REG_2_ & ~n7863;
  assign n8319 = ~n3881 & n7874;
  assign n8320 = ~n3759 & n7872;
  assign n8321 = P1_REG3_REG_2_ & ~n7856;
  assign n8322 = ~n8319 & ~n8320;
  assign n8323 = ~n8321 & n8322;
  assign n8324 = n7870 & ~n8323;
  assign n8325 = ~n7033 & ~n8324;
  assign n8326 = n8317 & ~n8318;
  assign n1195 = ~n8325 | ~n8326;
  assign n8328 = ~n4419 & ~n7863;
  assign n8329 = ~n4472 & ~n7867;
  assign n8330 = ~n4505 & n7874;
  assign n8331 = ~n4355 & n7872;
  assign n8332 = ~n4419 & ~n7856;
  assign n8333 = ~n8330 & ~n8331;
  assign n8334 = ~n8332 & n8333;
  assign n8335 = n7870 & ~n8334;
  assign n8336 = ~n6663 & ~n8335;
  assign n8337 = n7914 & ~n7920;
  assign n8338 = ~n7914 & n7920;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = n8066 & ~n8339;
  assign n8341 = ~n7921 & ~n7927;
  assign n8342 = ~n8066 & ~n8341;
  assign n8343 = ~n8340 & ~n8342;
  assign n8344 = n8087 & ~n8343;
  assign n8345 = ~n8328 & ~n8329;
  assign n8346 = n8336 & n8345;
  assign n1200 = n8344 | ~n8346;
  assign n8348 = ~n5128 & ~n7863;
  assign n8349 = n5176 & n8096;
  assign n8350 = P1_REG3_REG_22_ & ~P1_STATE_REG;
  assign n8351 = ~n5128 & ~n7856;
  assign n8352 = ~n5073 & n7872;
  assign n8353 = ~n5191 & n7874;
  assign n8354 = ~n8351 & ~n8352;
  assign n8355 = ~n8353 & n8354;
  assign n8356 = n7870 & ~n8355;
  assign n8357 = n8129 & ~n8135;
  assign n8358 = ~n8129 & n8135;
  assign n8359 = ~n8357 & ~n8358;
  assign n8360 = n8223 & ~n8359;
  assign n8361 = ~n8223 & n8359;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = n8087 & ~n8362;
  assign n8364 = ~n8348 & ~n8349;
  assign n8365 = ~n8350 & n8364;
  assign n8366 = ~n8356 & n8365;
  assign n1205 = n8363 | ~n8366;
  assign n8368 = ~n4566 & ~n7863;
  assign n8369 = ~n4609 & ~n7867;
  assign n8370 = ~n4566 & ~n7856;
  assign n8371 = ~n4505 & n7872;
  assign n8372 = ~n4639 & n7874;
  assign n8373 = ~n8370 & ~n8371;
  assign n8374 = ~n8372 & n8373;
  assign n8375 = n7870 & ~n8374;
  assign n8376 = ~n6598 & ~n8375;
  assign n8377 = ~n7900 & n7923;
  assign n8378 = ~n7927 & ~n8066;
  assign n8379 = ~n7921 & ~n8378;
  assign n8380 = ~n7910 & n8379;
  assign n8381 = n8377 & ~n8380;
  assign n8382 = ~n7895 & n7898;
  assign n8383 = n7895 & ~n7898;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~n7910 & n8384;
  assign n8386 = ~n7922 & ~n8379;
  assign n8387 = n8385 & ~n8386;
  assign n8388 = ~n8381 & ~n8387;
  assign n8389 = n8087 & n8388;
  assign n8390 = ~n8368 & ~n8369;
  assign n8391 = n8376 & n8390;
  assign n1210 = n8389 | ~n8391;
  assign n8393 = ~n5009 & ~n7863;
  assign n8394 = n5057 & n8096;
  assign n8395 = P1_REG3_REG_20_ & ~P1_STATE_REG;
  assign n8396 = ~n5009 & ~n7856;
  assign n8397 = ~n4967 & n7872;
  assign n8398 = ~n5073 & n7874;
  assign n8399 = ~n8396 & ~n8397;
  assign n8400 = ~n8398 & n8399;
  assign n8401 = n7870 & ~n8400;
  assign n8402 = ~n8198 & n8201;
  assign n8403 = n8198 & ~n8201;
  assign n8404 = ~n8402 & ~n8403;
  assign n8405 = ~n8214 & ~n8218;
  assign n8406 = ~n8404 & n8405;
  assign n8407 = ~n8202 & ~n8217;
  assign n8408 = ~n8405 & ~n8407;
  assign n8409 = ~n8406 & ~n8408;
  assign n8410 = n8087 & ~n8409;
  assign n8411 = ~n8393 & ~n8394;
  assign n8412 = ~n8395 & n8411;
  assign n8413 = ~n8401 & n8412;
  assign n1215 = n8410 | ~n8413;
  assign n8415 = ~n7861 & ~n7870;
  assign n8416 = ~n7856 & ~n8415;
  assign n8417 = n7860 & ~n8416;
  assign n8418 = P1_REG3_REG_0_ & ~n8417;
  assign n8419 = ~n3733 & ~n7867;
  assign n8420 = ~n3759 & n7870;
  assign n8421 = n7874 & n8420;
  assign n8422 = ~n6962 & n8087;
  assign n8423 = ~n7072 & ~n8422;
  assign n8424 = ~n8419 & ~n8421;
  assign n8425 = n8423 & n8424;
  assign n1220 = n8418 | ~n8425;
  assign n8427 = ~n4283 & ~n7863;
  assign n8428 = ~n4340 & ~n7867;
  assign n8429 = ~n4355 & n7874;
  assign n8430 = ~n4219 & n7872;
  assign n8431 = ~n4283 & ~n7856;
  assign n8432 = ~n8429 & ~n8430;
  assign n8433 = ~n8431 & n8432;
  assign n8434 = n7870 & ~n8433;
  assign n8435 = ~n6733 & ~n8434;
  assign n8436 = n7942 & ~n8061;
  assign n8437 = ~n7942 & n8061;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = n8054 & ~n8438;
  assign n8440 = ~n8054 & n8438;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = n8087 & ~n8441;
  assign n8443 = ~n8427 & ~n8428;
  assign n8444 = n8435 & n8443;
  assign n1225 = n8442 | ~n8444;
  assign n8446 = n7993 & ~n8045;
  assign n8447 = ~n7993 & n8045;
  assign n8448 = ~n8446 & ~n8447;
  assign n8449 = n8038 & ~n8448;
  assign n8450 = ~n8038 & n8448;
  assign n8451 = ~n8449 & ~n8450;
  assign n8452 = n8087 & ~n8451;
  assign n8453 = ~n3996 & ~n7867;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = ~n3938 & ~n7863;
  assign n8456 = ~n4011 & n7874;
  assign n8457 = ~n3881 & n7872;
  assign n8458 = ~n3938 & ~n7856;
  assign n8459 = ~n8456 & ~n8457;
  assign n8460 = ~n8458 & n8459;
  assign n8461 = n7870 & ~n8460;
  assign n8462 = ~n6923 & ~n8461;
  assign n8463 = n8454 & ~n8455;
  assign n1230 = ~n8462 | ~n8463;
  assign n8465 = ~n5249 & ~n7863;
  assign n8466 = n5297 & n8096;
  assign n8467 = P1_REG3_REG_24_ & ~P1_STATE_REG;
  assign n8468 = ~n5249 & ~n7856;
  assign n8469 = ~n5191 & n7872;
  assign n8470 = ~n5312 & n7874;
  assign n8471 = ~n8468 & ~n8469;
  assign n8472 = ~n8470 & n8471;
  assign n8473 = n7870 & ~n8472;
  assign n8474 = n8107 & ~n8113;
  assign n8475 = ~n8107 & n8113;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = n8227 & ~n8476;
  assign n8478 = ~n8114 & ~n8115;
  assign n8479 = ~n8227 & ~n8478;
  assign n8480 = ~n8477 & ~n8479;
  assign n8481 = n8087 & ~n8480;
  assign n8482 = ~n8465 & ~n8466;
  assign n8483 = ~n8467 & n8482;
  assign n8484 = ~n8473 & n8483;
  assign n1235 = n8481 | ~n8484;
  assign n8486 = ~n4809 & ~n7863;
  assign n8487 = ~n4865 & ~n7867;
  assign n8488 = ~n4809 & ~n7856;
  assign n8489 = ~n4752 & n7872;
  assign n8490 = ~n4895 & n7874;
  assign n8491 = ~n8488 & ~n8489;
  assign n8492 = ~n8490 & n8491;
  assign n8493 = n7870 & ~n8492;
  assign n8494 = ~n8161 & ~n8178;
  assign n8495 = n8184 & ~n8494;
  assign n8496 = ~n8171 & n8188;
  assign n8497 = n8495 & ~n8496;
  assign n8498 = n8161 & ~n8178;
  assign n8499 = ~n8161 & n8178;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~n8171 & n8500;
  assign n8502 = ~n8182 & ~n8188;
  assign n8503 = n8501 & ~n8502;
  assign n8504 = ~n8497 & ~n8503;
  assign n8505 = n8087 & n8504;
  assign n8506 = ~n8486 & ~n8487;
  assign n8507 = ~n6473 & n8506;
  assign n8508 = ~n8493 & n8507;
  assign n1240 = n8505 | ~n8508;
  assign n8510 = ~n4004 & ~n7863;
  assign n8511 = ~n4066 & ~n7867;
  assign n8512 = n7982 & ~n7988;
  assign n8513 = ~n7982 & n7988;
  assign n8514 = ~n8512 & ~n8513;
  assign n8515 = n8048 & ~n8514;
  assign n8516 = ~n8048 & n8514;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = n8087 & ~n8517;
  assign n8519 = ~n4081 & n7874;
  assign n8520 = ~n3945 & n7872;
  assign n8521 = ~n4004 & ~n7856;
  assign n8522 = ~n8519 & ~n8520;
  assign n8523 = ~n8521 & n8522;
  assign n8524 = n7870 & ~n8523;
  assign n8525 = ~n6871 & ~n8524;
  assign n8526 = ~n8510 & ~n8511;
  assign n8527 = ~n8518 & n8526;
  assign n1245 = ~n8525 | ~n8527;
  assign n8529 = ~n4748 & ~n7863;
  assign n8530 = ~n4798 & ~n7867;
  assign n8531 = ~n4748 & ~n7856;
  assign n8532 = ~n4703 & n7872;
  assign n8533 = ~n4813 & n7874;
  assign n8534 = ~n8531 & ~n8532;
  assign n8535 = ~n8533 & n8534;
  assign n8536 = n7870 & ~n8535;
  assign n8537 = n8164 & ~n8170;
  assign n8538 = ~n8164 & n8170;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = n8188 & ~n8539;
  assign n8541 = ~n8171 & ~n8182;
  assign n8542 = ~n8188 & ~n8541;
  assign n8543 = ~n8540 & ~n8542;
  assign n8544 = n8087 & ~n8543;
  assign n8545 = ~n8529 & ~n8530;
  assign n8546 = ~n6507 & n8545;
  assign n8547 = ~n8536 & n8546;
  assign n1250 = n8544 | ~n8547;
  assign n8549 = ~n5308 & ~n7863;
  assign n8550 = n5361 & n8096;
  assign n8551 = P1_REG3_REG_25_ & ~P1_STATE_REG;
  assign n8552 = ~n5308 & ~n7856;
  assign n8553 = ~n5253 & n7872;
  assign n8554 = ~n5376 & n7874;
  assign n8555 = ~n8552 & ~n8553;
  assign n8556 = ~n8554 & n8555;
  assign n8557 = n7870 & ~n8556;
  assign n8558 = n8232 & ~n8238;
  assign n8559 = ~n8232 & n8238;
  assign n8560 = ~n8558 & ~n8559;
  assign n8561 = n8229 & ~n8560;
  assign n8562 = ~n8239 & ~n8251;
  assign n8563 = ~n8229 & ~n8562;
  assign n8564 = ~n8561 & ~n8563;
  assign n8565 = n8087 & ~n8564;
  assign n8566 = ~n8549 & ~n8550;
  assign n8567 = ~n8551 & n8566;
  assign n8568 = ~n8557 & n8567;
  assign n1255 = n8565 | ~n8568;
  assign n8570 = ~n4501 & ~n7863;
  assign n8571 = ~n4542 & ~n7867;
  assign n8572 = ~n4501 & ~n7856;
  assign n8573 = ~n4423 & n7872;
  assign n8574 = ~n4570 & n7874;
  assign n8575 = ~n8572 & ~n8573;
  assign n8576 = ~n8574 & n8575;
  assign n8577 = n7870 & ~n8576;
  assign n8578 = ~n6633 & ~n8577;
  assign n8579 = n7903 & ~n7909;
  assign n8580 = ~n7903 & n7909;
  assign n8581 = ~n8579 & ~n8580;
  assign n8582 = n8379 & ~n8581;
  assign n8583 = ~n7910 & ~n7922;
  assign n8584 = ~n8379 & ~n8583;
  assign n8585 = ~n8582 & ~n8584;
  assign n8586 = n8087 & ~n8585;
  assign n8587 = ~n8570 & ~n8571;
  assign n8588 = n8578 & n8587;
  assign n1260 = n8586 | ~n8588;
  assign n8590 = ~n5069 & ~n7863;
  assign n8591 = n5117 & n8096;
  assign n8592 = P1_REG3_REG_21_ & ~P1_STATE_REG;
  assign n8593 = ~n5069 & ~n7856;
  assign n8594 = ~n5013 & n7872;
  assign n8595 = ~n5132 & n7874;
  assign n8596 = ~n8593 & ~n8594;
  assign n8597 = ~n8595 & n8596;
  assign n8598 = n7870 & ~n8597;
  assign n8599 = ~n8217 & n8405;
  assign n8600 = ~n8216 & ~n8599;
  assign n8601 = n8213 & n8600;
  assign n8602 = ~n8208 & n8211;
  assign n8603 = n8208 & ~n8211;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8217 & n8604;
  assign n8606 = ~n8202 & ~n8405;
  assign n8607 = n8605 & ~n8606;
  assign n8608 = ~n8601 & ~n8607;
  assign n8609 = n8087 & n8608;
  assign n8610 = ~n8590 & ~n8591;
  assign n8611 = ~n8592 & n8610;
  assign n8612 = ~n8598 & n8611;
  assign n1265 = n8609 | ~n8612;
  assign n8614 = n8022 & ~n8028;
  assign n8615 = ~n8022 & n8028;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = n8034 & ~n8616;
  assign n8618 = ~n8034 & n8616;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = n8087 & ~n8619;
  assign n8621 = ~n3813 & ~n7867;
  assign n8622 = ~n8620 & ~n8621;
  assign n8623 = P1_REG3_REG_1_ & ~n7863;
  assign n8624 = ~n3824 & n7874;
  assign n8625 = ~n3767 & n7872;
  assign n8626 = P1_REG3_REG_1_ & ~n7856;
  assign n8627 = ~n8624 & ~n8625;
  assign n8628 = ~n8626 & n8627;
  assign n8629 = n7870 & ~n8628;
  assign n8630 = ~n7049 & ~n8629;
  assign n8631 = n8622 & ~n8623;
  assign n1270 = ~n8630 | ~n8631;
  assign n8633 = ~n4212 & ~n7863;
  assign n8634 = ~n4272 & ~n7867;
  assign n8635 = ~n4287 & n7874;
  assign n8636 = ~n4146 & n7872;
  assign n8637 = ~n4212 & ~n7856;
  assign n8638 = ~n8635 & ~n8636;
  assign n8639 = ~n8637 & n8638;
  assign n8640 = n7870 & ~n8639;
  assign n8641 = ~n6763 & ~n8640;
  assign n8642 = n7945 & ~n7951;
  assign n8643 = ~n7945 & n7951;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = n8052 & ~n8644;
  assign n8646 = ~n8052 & n8644;
  assign n8647 = ~n8645 & ~n8646;
  assign n8648 = n8087 & ~n8647;
  assign n8649 = ~n8633 & ~n8634;
  assign n8650 = n8641 & n8649;
  assign n1275 = n8648 | ~n8650;
  assign n8652 = ~n5489 & ~n7863;
  assign n8653 = n5537 & n8096;
  assign n8654 = P1_REG3_REG_28_ & ~P1_STATE_REG;
  assign n8655 = ~n5550 & n7874;
  assign n8656 = ~n5433 & n7872;
  assign n8657 = ~n5489 & ~n7856;
  assign n8658 = ~n8655 & ~n8656;
  assign n8659 = ~n8657 & n8658;
  assign n8660 = n7870 & ~n8659;
  assign n8661 = ~n5433 & n6938;
  assign n8662 = n5478 & ~n6954;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = ~n6935 & ~n8663;
  assign n8665 = n6935 & n8663;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~n5433 & ~n6945;
  assign n8668 = n5478 & n6938;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = n8666 & n8669;
  assign n8671 = n8250 & ~n8670;
  assign n8672 = ~n8115 & ~n8670;
  assign n8673 = ~n8227 & ~n8254;
  assign n8674 = n8672 & n8673;
  assign n8675 = ~n8114 & ~n8239;
  assign n8676 = ~n8254 & ~n8675;
  assign n8677 = ~n8670 & n8676;
  assign n8678 = ~n8666 & ~n8669;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = ~n5493 & ~n6945;
  assign n8681 = n5537 & n6938;
  assign n8682 = ~n8680 & ~n8681;
  assign n8683 = ~n6935 & ~n8682;
  assign n8684 = n6935 & n8682;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~n5493 & n6938;
  assign n8687 = n5537 & ~n6954;
  assign n8688 = ~n8686 & ~n8687;
  assign n8689 = ~n8685 & n8688;
  assign n8690 = n8685 & ~n8688;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = ~n8671 & ~n8674;
  assign n8693 = n8679 & n8692;
  assign n8694 = ~n8691 & n8693;
  assign n8695 = n8228 & ~n8254;
  assign n8696 = ~n8250 & ~n8678;
  assign n8697 = ~n8676 & ~n8695;
  assign n8698 = n8696 & n8697;
  assign n8699 = ~n8670 & ~n8698;
  assign n8700 = n8691 & n8699;
  assign n8701 = ~n8694 & ~n8700;
  assign n8702 = n8087 & ~n8701;
  assign n8703 = ~n8652 & ~n8653;
  assign n8704 = ~n8654 & n8703;
  assign n8705 = ~n8660 & n8704;
  assign n1280 = n8702 | ~n8705;
  assign n8707 = ~n4963 & ~n7863;
  assign n8708 = ~n4998 & ~n7867;
  assign n8709 = ~n4963 & ~n7856;
  assign n8710 = ~n4895 & n7872;
  assign n8711 = ~n5013 & n7874;
  assign n8712 = ~n8709 & ~n8710;
  assign n8713 = ~n8711 & n8712;
  assign n8714 = n7870 & ~n8713;
  assign n8715 = ~n8143 & n8146;
  assign n8716 = n8143 & ~n8146;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = n8192 & ~n8717;
  assign n8719 = ~n8147 & ~n8218;
  assign n8720 = ~n8192 & ~n8719;
  assign n8721 = ~n8718 & ~n8720;
  assign n8722 = n8087 & ~n8721;
  assign n8723 = ~n8707 & ~n8708;
  assign n8724 = ~n6309 & n8723;
  assign n8725 = ~n8714 & n8724;
  assign n1285 = n8722 | ~n8725;
  assign n8727 = ~n7996 & ~n8013;
  assign n8728 = n8019 & ~n8727;
  assign n8729 = ~n8006 & n8036;
  assign n8730 = n8728 & ~n8729;
  assign n8731 = n7996 & ~n8013;
  assign n8732 = ~n7996 & n8013;
  assign n8733 = ~n8731 & ~n8732;
  assign n8734 = ~n8006 & n8733;
  assign n8735 = ~n8017 & ~n8036;
  assign n8736 = n8734 & ~n8735;
  assign n8737 = ~n8730 & ~n8736;
  assign n8738 = n8087 & n8737;
  assign n8739 = ~n3931 & ~n7867;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~P1_REG3_REG_3_ & ~n7863;
  assign n8742 = ~n3945 & n7874;
  assign n8743 = ~n3824 & n7872;
  assign n8744 = ~P1_REG3_REG_3_ & ~n7856;
  assign n8745 = ~n8742 & ~n8743;
  assign n8746 = ~n8744 & n8745;
  assign n8747 = n7870 & ~n8746;
  assign n8748 = ~n6988 & ~n8747;
  assign n8749 = n8740 & ~n8741;
  assign n1290 = ~n8748 | ~n8749;
  assign n8751 = ~n4351 & ~n7863;
  assign n8752 = ~n4407 & ~n7867;
  assign n8753 = ~n4423 & n7874;
  assign n8754 = ~n4287 & n7872;
  assign n8755 = ~n4351 & ~n7856;
  assign n8756 = ~n8753 & ~n8754;
  assign n8757 = ~n8755 & n8756;
  assign n8758 = n7870 & ~n8757;
  assign n8759 = ~n6698 & ~n8758;
  assign n8760 = n7931 & ~n7937;
  assign n8761 = ~n7931 & n7937;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = n8064 & ~n8762;
  assign n8764 = ~n8064 & n8762;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = n8087 & ~n8765;
  assign n8767 = ~n8751 & ~n8752;
  assign n8768 = n8759 & n8767;
  assign n1295 = n8766 | ~n8768;
  assign n8770 = ~n5187 & ~n7863;
  assign n8771 = n5238 & n8096;
  assign n8772 = P1_REG3_REG_23_ & ~P1_STATE_REG;
  assign n8773 = ~n5187 & ~n7856;
  assign n8774 = ~n5132 & n7872;
  assign n8775 = ~n5253 & n7874;
  assign n8776 = ~n8773 & ~n8774;
  assign n8777 = ~n8775 & n8776;
  assign n8778 = n7870 & ~n8777;
  assign n8779 = n8118 & ~n8124;
  assign n8780 = ~n8118 & n8124;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = n8225 & ~n8781;
  assign n8783 = ~n8225 & n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = n8087 & ~n8784;
  assign n8786 = ~n8770 & ~n8771;
  assign n8787 = ~n8772 & n8786;
  assign n8788 = ~n8778 & n8787;
  assign n1300 = n8785 | ~n8788;
  assign n8790 = ~n4635 & ~n7863;
  assign n8791 = ~n4673 & ~n7867;
  assign n8792 = ~n4635 & ~n7856;
  assign n8793 = ~n4570 & n7872;
  assign n8794 = ~n4703 & n7874;
  assign n8795 = ~n8792 & ~n8793;
  assign n8796 = ~n8794 & n8795;
  assign n8797 = n7870 & ~n8796;
  assign n8798 = n7881 & ~n7887;
  assign n8799 = ~n7881 & n7887;
  assign n8800 = ~n8798 & ~n8799;
  assign n8801 = n8068 & ~n8800;
  assign n8802 = ~n8068 & n8800;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = n8087 & ~n8803;
  assign n8805 = ~n8790 & ~n8791;
  assign n8806 = ~n6564 & n8805;
  assign n8807 = ~n8797 & n8806;
  assign n1305 = n8804 | ~n8807;
  assign n8809 = ~n5429 & ~n7863;
  assign n8810 = n5478 & n8096;
  assign n8811 = P1_REG3_REG_27_ & ~P1_STATE_REG;
  assign n8812 = ~n5429 & ~n7856;
  assign n8813 = ~n5376 & n7872;
  assign n8814 = ~n5493 & n7874;
  assign n8815 = ~n8812 & ~n8813;
  assign n8816 = ~n8814 & n8815;
  assign n8817 = n7870 & ~n8816;
  assign n8818 = ~n8250 & n8697;
  assign n8819 = ~n8666 & n8669;
  assign n8820 = n8666 & ~n8669;
  assign n8821 = ~n8819 & ~n8820;
  assign n8822 = n8818 & ~n8821;
  assign n8823 = ~n8818 & n8821;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = n8087 & ~n8824;
  assign n8826 = ~n8809 & ~n8810;
  assign n8827 = ~n8811 & n8826;
  assign n8828 = ~n8817 & n8827;
  assign n1310 = n8825 | ~n8828;
  assign n8830 = ~n4139 & ~n7863;
  assign n8831 = ~n4204 & ~n7867;
  assign n8832 = ~n4219 & n7874;
  assign n8833 = ~n4081 & n7872;
  assign n8834 = ~n4139 & ~n7856;
  assign n8835 = ~n8832 & ~n8833;
  assign n8836 = ~n8834 & n8835;
  assign n8837 = n7870 & ~n8836;
  assign n8838 = ~n6797 & ~n8837;
  assign n8839 = ~n7956 & ~n7973;
  assign n8840 = n7979 & ~n8839;
  assign n8841 = ~n7966 & n8050;
  assign n8842 = n8840 & ~n8841;
  assign n8843 = n7956 & ~n7973;
  assign n8844 = ~n7956 & n7973;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n7966 & n8845;
  assign n8847 = ~n7977 & ~n8050;
  assign n8848 = n8846 & ~n8847;
  assign n8849 = ~n8842 & ~n8848;
  assign n8850 = n8087 & n8849;
  assign n8851 = ~n8830 & ~n8831;
  assign n8852 = n8838 & n8851;
  assign n1315 = n8850 | ~n8852;
  assign n8854 = ~P2_IR_REG_31_ & P2_STATE_REG;
  assign n8855 = P2_STATE_REG & ~n8854;
  assign n8856 = P2_IR_REG_0_ & n8855;
  assign n8857 = P2_IR_REG_0_ & n8854;
  assign n8858 = n2615_1 & ~n2622;
  assign n8859 = P1_DATAO_REG_0_ & ~n2615_1;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = ~P2_STATE_REG & ~n8860;
  assign n8862 = ~n8856 & ~n8857;
  assign n1335 = n8861 | ~n8862;
  assign n8864 = P2_IR_REG_0_ & ~P2_IR_REG_1_;
  assign n8865 = ~P2_IR_REG_0_ & P2_IR_REG_1_;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = n8855 & ~n8866;
  assign n8868 = P2_IR_REG_1_ & n8854;
  assign n8869 = n2615_1 & ~n2648;
  assign n8870 = P1_DATAO_REG_1_ & ~n2615_1;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = ~P2_STATE_REG & ~n8871;
  assign n8873 = ~n8867 & ~n8868;
  assign n1340 = n8872 | ~n8873;
  assign n8875 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_;
  assign n8876 = P2_IR_REG_2_ & ~n8875;
  assign n8877 = ~P2_IR_REG_2_ & n8875;
  assign n8878 = ~n8876 & ~n8877;
  assign n8879 = n8855 & n8878;
  assign n8880 = P2_IR_REG_2_ & n8854;
  assign n8881 = n2615_1 & ~n2673;
  assign n8882 = P1_DATAO_REG_2_ & ~n2615_1;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = ~P2_STATE_REG & ~n8883;
  assign n8885 = ~n8879 & ~n8880;
  assign n1345 = n8884 | ~n8885;
  assign n8887 = P2_IR_REG_3_ & ~n8877;
  assign n8888 = ~P2_IR_REG_3_ & n8877;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = n8855 & n8889;
  assign n8891 = P2_IR_REG_3_ & n8854;
  assign n8892 = n2615_1 & ~n2704;
  assign n8893 = P1_DATAO_REG_3_ & ~n2615_1;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 = ~P2_STATE_REG & ~n8894;
  assign n8896 = ~n8890 & ~n8891;
  assign n1350 = n8895 | ~n8896;
  assign n8898 = P2_IR_REG_4_ & ~n8888;
  assign n8899 = ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign n8900 = n8877 & n8899;
  assign n8901 = ~n8898 & ~n8900;
  assign n8902 = n8855 & n8901;
  assign n8903 = P2_IR_REG_4_ & n8854;
  assign n8904 = n2615_1 & ~n2732;
  assign n8905 = P1_DATAO_REG_4_ & ~n2615_1;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = ~P2_STATE_REG & ~n8906;
  assign n8908 = ~n8902 & ~n8903;
  assign n1355 = n8907 | ~n8908;
  assign n8910 = ~P2_IR_REG_5_ & n8900;
  assign n8911 = P2_IR_REG_5_ & ~n8900;
  assign n8912 = ~n8910 & ~n8911;
  assign n8913 = n8855 & n8912;
  assign n8914 = P2_IR_REG_5_ & n8854;
  assign n8915 = n2615_1 & ~n2756;
  assign n8916 = P1_DATAO_REG_5_ & ~n2615_1;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = ~P2_STATE_REG & ~n8917;
  assign n8919 = ~n8913 & ~n8914;
  assign n1360 = n8918 | ~n8919;
  assign n8921 = P2_IR_REG_6_ & ~n8910;
  assign n8922 = ~P2_IR_REG_5_ & ~P2_IR_REG_6_;
  assign n8923 = n8900 & n8922;
  assign n8924 = ~n8921 & ~n8923;
  assign n8925 = n8855 & n8924;
  assign n8926 = P2_IR_REG_6_ & n8854;
  assign n8927 = n2615_1 & ~n2784;
  assign n8928 = P1_DATAO_REG_6_ & ~n2615_1;
  assign n8929 = ~n8927 & ~n8928;
  assign n8930 = ~P2_STATE_REG & ~n8929;
  assign n8931 = ~n8925 & ~n8926;
  assign n1365 = n8930 | ~n8931;
  assign n8933 = P2_IR_REG_7_ & ~n8923;
  assign n8934 = ~P2_IR_REG_7_ & n8923;
  assign n8935 = ~n8933 & ~n8934;
  assign n8936 = n8855 & n8935;
  assign n8937 = P2_IR_REG_7_ & n8854;
  assign n8938 = n2615_1 & ~n2811;
  assign n8939 = P1_DATAO_REG_7_ & ~n2615_1;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = ~P2_STATE_REG & ~n8940;
  assign n8942 = ~n8936 & ~n8937;
  assign n1370 = n8941 | ~n8942;
  assign n8944 = P2_IR_REG_8_ & ~n8934;
  assign n8945 = ~P2_IR_REG_7_ & ~P2_IR_REG_8_;
  assign n8946 = ~P2_IR_REG_5_ & n8899;
  assign n8947 = ~P2_IR_REG_6_ & n8946;
  assign n8948 = n8877 & n8945;
  assign n8949 = n8947 & n8948;
  assign n8950 = ~n8944 & ~n8949;
  assign n8951 = n8855 & n8950;
  assign n8952 = P2_IR_REG_8_ & n8854;
  assign n8953 = n2615_1 & ~n2839;
  assign n8954 = P1_DATAO_REG_8_ & ~n2615_1;
  assign n8955 = ~n8953 & ~n8954;
  assign n8956 = ~P2_STATE_REG & ~n8955;
  assign n8957 = ~n8951 & ~n8952;
  assign n1375 = n8956 | ~n8957;
  assign n8959 = ~P2_IR_REG_9_ & n8949;
  assign n8960 = P2_IR_REG_9_ & ~n8949;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = n8855 & n8961;
  assign n8963 = P2_IR_REG_9_ & n8854;
  assign n8964 = n2615_1 & ~n2866;
  assign n8965 = P1_DATAO_REG_9_ & ~n2615_1;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = ~P2_STATE_REG & ~n8966;
  assign n8968 = ~n8962 & ~n8963;
  assign n1380 = n8967 | ~n8968;
  assign n8970 = P2_IR_REG_10_ & ~n8959;
  assign n8971 = ~P2_IR_REG_9_ & ~P2_IR_REG_10_;
  assign n8972 = n8949 & n8971;
  assign n8973 = ~n8970 & ~n8972;
  assign n8974 = n8855 & n8973;
  assign n8975 = P2_IR_REG_10_ & n8854;
  assign n8976 = n2615_1 & ~n2894;
  assign n8977 = P1_DATAO_REG_10_ & ~n2615_1;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = ~P2_STATE_REG & ~n8978;
  assign n8980 = ~n8974 & ~n8975;
  assign n1385 = n8979 | ~n8980;
  assign n8982 = P2_IR_REG_11_ & ~n8972;
  assign n8983 = ~P2_IR_REG_11_ & n8972;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = n8855 & n8984;
  assign n8986 = P2_IR_REG_11_ & n8854;
  assign n8987 = n2615_1 & ~n2921;
  assign n8988 = P1_DATAO_REG_11_ & ~n2615_1;
  assign n8989 = ~n8987 & ~n8988;
  assign n8990 = ~P2_STATE_REG & ~n8989;
  assign n8991 = ~n8985 & ~n8986;
  assign n1390 = n8990 | ~n8991;
  assign n8993 = P2_IR_REG_12_ & ~n8983;
  assign n8994 = ~P2_IR_REG_10_ & ~P2_IR_REG_11_;
  assign n8995 = ~P2_IR_REG_12_ & n8994;
  assign n8996 = ~P2_IR_REG_9_ & n8995;
  assign n8997 = n8949 & n8996;
  assign n8998 = ~n8993 & ~n8997;
  assign n8999 = n8855 & n8998;
  assign n9000 = P2_IR_REG_12_ & n8854;
  assign n9001 = n2615_1 & ~n2948;
  assign n9002 = P1_DATAO_REG_12_ & ~n2615_1;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = ~P2_STATE_REG & ~n9003;
  assign n9005 = ~n8999 & ~n9000;
  assign n1395 = n9004 | ~n9005;
  assign n9007 = ~P2_IR_REG_13_ & n8997;
  assign n9008 = P2_IR_REG_13_ & ~n8997;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = n8855 & n9009;
  assign n9011 = P2_IR_REG_13_ & n8854;
  assign n9012 = n2615_1 & ~n2975_1;
  assign n9013 = P1_DATAO_REG_13_ & ~n2615_1;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~P2_STATE_REG & ~n9014;
  assign n9016 = ~n9010 & ~n9011;
  assign n1400 = n9015 | ~n9016;
  assign n9018 = P2_IR_REG_14_ & ~n9007;
  assign n9019 = ~P2_IR_REG_13_ & ~P2_IR_REG_14_;
  assign n9020 = n8997 & n9019;
  assign n9021 = ~n9018 & ~n9020;
  assign n9022 = n8855 & n9021;
  assign n9023 = P2_IR_REG_14_ & n8854;
  assign n9024 = n2615_1 & ~n3003;
  assign n9025 = P1_DATAO_REG_14_ & ~n2615_1;
  assign n9026 = ~n9024 & ~n9025;
  assign n9027 = ~P2_STATE_REG & ~n9026;
  assign n9028 = ~n9022 & ~n9023;
  assign n1405 = n9027 | ~n9028;
  assign n9030 = P2_IR_REG_15_ & ~n9020;
  assign n9031 = ~P2_IR_REG_15_ & n9020;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = n8855 & n9032;
  assign n9034 = P2_IR_REG_15_ & n8854;
  assign n9035 = n2615_1 & ~n3030_1;
  assign n9036 = P1_DATAO_REG_15_ & ~n2615_1;
  assign n9037 = ~n9035 & ~n9036;
  assign n9038 = ~P2_STATE_REG & ~n9037;
  assign n9039 = ~n9033 & ~n9034;
  assign n1410 = n9038 | ~n9039;
  assign n9041 = P2_IR_REG_16_ & ~n9031;
  assign n9042 = ~P2_IR_REG_6_ & ~P2_IR_REG_7_;
  assign n9043 = ~P2_IR_REG_8_ & n9042;
  assign n9044 = ~P2_IR_REG_9_ & n9043;
  assign n9045 = ~P2_IR_REG_2_ & ~P2_IR_REG_3_;
  assign n9046 = ~P2_IR_REG_4_ & n9045;
  assign n9047 = ~P2_IR_REG_5_ & n9046;
  assign n9048 = ~P2_IR_REG_15_ & ~P2_IR_REG_16_;
  assign n9049 = ~P2_IR_REG_1_ & n9048;
  assign n9050 = ~P2_IR_REG_0_ & n9049;
  assign n9051 = ~P2_IR_REG_12_ & n9019;
  assign n9052 = ~P2_IR_REG_10_ & n9051;
  assign n9053 = ~P2_IR_REG_11_ & n9052;
  assign n9054 = n9044 & n9047;
  assign n9055 = n9050 & n9054;
  assign n9056 = n9053 & n9055;
  assign n9057 = ~n9041 & ~n9056;
  assign n9058 = n8855 & n9057;
  assign n9059 = P2_IR_REG_16_ & n8854;
  assign n9060 = n2615_1 & ~n3071;
  assign n9061 = P1_DATAO_REG_16_ & ~n2615_1;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~P2_STATE_REG & ~n9062;
  assign n9064 = ~n9058 & ~n9059;
  assign n1415 = n9063 | ~n9064;
  assign n9066 = ~P2_IR_REG_17_ & n9056;
  assign n9067 = P2_IR_REG_17_ & ~n9056;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = n8855 & n9068;
  assign n9070 = P2_IR_REG_17_ & n8854;
  assign n9071 = n2615_1 & ~n3095_1;
  assign n9072 = P1_DATAO_REG_17_ & ~n2615_1;
  assign n9073 = ~n9071 & ~n9072;
  assign n9074 = ~P2_STATE_REG & ~n9073;
  assign n9075 = ~n9069 & ~n9070;
  assign n1420 = n9074 | ~n9075;
  assign n9077 = P2_IR_REG_18_ & ~n9066;
  assign n9078 = ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign n9079 = n9056 & n9078;
  assign n9080 = ~n9077 & ~n9079;
  assign n9081 = n8855 & n9080;
  assign n9082 = P2_IR_REG_18_ & n8854;
  assign n9083 = n2615_1 & ~n3129;
  assign n9084 = P1_DATAO_REG_18_ & ~n2615_1;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~P2_STATE_REG & ~n9085;
  assign n9087 = ~n9081 & ~n9082;
  assign n1425 = n9086 | ~n9087;
  assign n9089 = ~P2_IR_REG_19_ & n9079;
  assign n9090 = P2_IR_REG_19_ & ~n9079;
  assign n9091 = ~n9089 & ~n9090;
  assign n9092 = n8855 & n9091;
  assign n9093 = P2_IR_REG_19_ & n8854;
  assign n9094 = n2615_1 & ~n3166;
  assign n9095 = P1_DATAO_REG_19_ & ~n2615_1;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = ~P2_STATE_REG & ~n9096;
  assign n9098 = ~n9092 & ~n9093;
  assign n1430 = n9097 | ~n9098;
  assign n9100 = ~P2_IR_REG_20_ & n9089;
  assign n9101 = P2_IR_REG_20_ & ~n9089;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 = n8855 & n9102;
  assign n9104 = P2_IR_REG_20_ & n8854;
  assign n9105 = n2615_1 & ~n3203;
  assign n9106 = P1_DATAO_REG_20_ & ~n2615_1;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = ~P2_STATE_REG & ~n9107;
  assign n9109 = ~n9103 & ~n9104;
  assign n1435 = n9108 | ~n9109;
  assign n9111 = ~P2_IR_REG_19_ & n9078;
  assign n9112 = ~P2_IR_REG_20_ & n9111;
  assign n9113 = n9056 & n9112;
  assign n9114 = ~P2_IR_REG_21_ & n9113;
  assign n9115 = P2_IR_REG_21_ & ~n9113;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = n8855 & n9116;
  assign n9118 = P2_IR_REG_21_ & n8854;
  assign n9119 = n2615_1 & ~n3227;
  assign n9120 = P1_DATAO_REG_21_ & ~n2615_1;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = ~P2_STATE_REG & ~n9121;
  assign n9123 = ~n9117 & ~n9118;
  assign n1440 = n9122 | ~n9123;
  assign n9125 = ~P2_IR_REG_22_ & n9114;
  assign n9126 = P2_IR_REG_22_ & ~n9114;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = n8855 & n9127;
  assign n9129 = P2_IR_REG_22_ & n8854;
  assign n9130 = n2615_1 & ~n3264;
  assign n9131 = P1_DATAO_REG_22_ & ~n2615_1;
  assign n9132 = ~n9130 & ~n9131;
  assign n9133 = ~P2_STATE_REG & ~n9132;
  assign n9134 = ~n9128 & ~n9129;
  assign n1445 = n9133 | ~n9134;
  assign n9136 = P2_IR_REG_23_ & ~n9125;
  assign n9137 = ~P2_IR_REG_21_ & ~P2_IR_REG_23_;
  assign n9138 = ~P2_IR_REG_22_ & n9137;
  assign n9139 = n9113 & n9138;
  assign n9140 = ~n9136 & ~n9139;
  assign n9141 = n8855 & n9140;
  assign n9142 = P2_IR_REG_23_ & n8854;
  assign n9143 = n2615_1 & ~n3306;
  assign n9144 = P1_DATAO_REG_23_ & ~n2615_1;
  assign n9145 = ~n9143 & ~n9144;
  assign n9146 = ~P2_STATE_REG & ~n9145;
  assign n9147 = ~n9141 & ~n9142;
  assign n1450 = n9146 | ~n9147;
  assign n9149 = P2_IR_REG_24_ & ~n9139;
  assign n9150 = ~P2_IR_REG_24_ & n9139;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = n8855 & n9151;
  assign n9153 = P2_IR_REG_24_ & n8854;
  assign n9154 = n2615_1 & ~n3346;
  assign n9155 = P1_DATAO_REG_24_ & ~n2615_1;
  assign n9156 = ~n9154 & ~n9155;
  assign n9157 = ~P2_STATE_REG & ~n9156;
  assign n9158 = ~n9152 & ~n9153;
  assign n1455 = n9157 | ~n9158;
  assign n9160 = ~P2_IR_REG_25_ & n9150;
  assign n9161 = P2_IR_REG_25_ & ~n9150;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = n8855 & n9162;
  assign n9164 = P2_IR_REG_25_ & n8854;
  assign n9165 = n2615_1 & ~n3370_1;
  assign n9166 = P1_DATAO_REG_25_ & ~n2615_1;
  assign n9167 = ~n9165 & ~n9166;
  assign n9168 = ~P2_STATE_REG & ~n9167;
  assign n9169 = ~n9163 & ~n9164;
  assign n1460 = n9168 | ~n9169;
  assign n9171 = P2_IR_REG_26_ & ~n9160;
  assign n9172 = ~P2_IR_REG_7_ & ~P2_IR_REG_9_;
  assign n9173 = ~P2_IR_REG_8_ & n9172;
  assign n9174 = ~P2_IR_REG_4_ & ~P2_IR_REG_6_;
  assign n9175 = ~P2_IR_REG_5_ & n9174;
  assign n9176 = ~P2_IR_REG_3_ & ~P2_IR_REG_26_;
  assign n9177 = ~P2_IR_REG_2_ & n9176;
  assign n9178 = ~P2_IR_REG_22_ & ~P2_IR_REG_23_;
  assign n9179 = ~P2_IR_REG_24_ & n9178;
  assign n9180 = ~P2_IR_REG_25_ & n9179;
  assign n9181 = n9173 & n9175;
  assign n9182 = n9177 & n9181;
  assign n9183 = n9180 & n9182;
  assign n9184 = ~P2_IR_REG_0_ & ~P2_IR_REG_21_;
  assign n9185 = ~P2_IR_REG_20_ & n9184;
  assign n9186 = ~P2_IR_REG_1_ & n9111;
  assign n9187 = ~P2_IR_REG_14_ & ~P2_IR_REG_16_;
  assign n9188 = ~P2_IR_REG_15_ & n9187;
  assign n9189 = ~P2_IR_REG_13_ & n8995;
  assign n9190 = n9185 & n9186;
  assign n9191 = n9188 & n9190;
  assign n9192 = n9189 & n9191;
  assign n9193 = n9183 & n9192;
  assign n9194 = ~n9171 & ~n9193;
  assign n9195 = n8855 & n9194;
  assign n9196 = P2_IR_REG_26_ & n8854;
  assign n9197 = n2615_1 & ~n3413;
  assign n9198 = P1_DATAO_REG_26_ & ~n2615_1;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = ~P2_STATE_REG & ~n9199;
  assign n9201 = ~n9195 & ~n9196;
  assign n1465 = n9200 | ~n9201;
  assign n9203 = ~P2_IR_REG_27_ & n9193;
  assign n9204 = P2_IR_REG_27_ & ~n9193;
  assign n9205 = ~n9203 & ~n9204;
  assign n9206 = n8855 & n9205;
  assign n9207 = P2_IR_REG_27_ & n8854;
  assign n9208 = n2615_1 & ~n3437;
  assign n9209 = P1_DATAO_REG_27_ & ~n2615_1;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = ~P2_STATE_REG & ~n9210;
  assign n9212 = ~n9206 & ~n9207;
  assign n1470 = n9211 | ~n9212;
  assign n9214 = ~P2_IR_REG_2_ & ~P2_IR_REG_26_;
  assign n9215 = ~P2_IR_REG_27_ & n9214;
  assign n9216 = n8947 & n9173;
  assign n9217 = n9215 & n9216;
  assign n9218 = n9180 & n9217;
  assign n9219 = n9192 & n9218;
  assign n9220 = ~P2_IR_REG_28_ & n9219;
  assign n9221 = P2_IR_REG_28_ & ~n9219;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = n8855 & n9222;
  assign n9224 = P2_IR_REG_28_ & n8854;
  assign n9225 = n2615_1 & ~n3482;
  assign n9226 = P1_DATAO_REG_28_ & ~n2615_1;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = ~P2_STATE_REG & ~n9227;
  assign n9229 = ~n9223 & ~n9224;
  assign n1475 = n9228 | ~n9229;
  assign n9231 = ~P2_IR_REG_2_ & ~P2_IR_REG_27_;
  assign n9232 = ~P2_IR_REG_28_ & n9231;
  assign n9233 = ~P2_IR_REG_23_ & ~P2_IR_REG_24_;
  assign n9234 = ~P2_IR_REG_25_ & n9233;
  assign n9235 = ~P2_IR_REG_26_ & n9234;
  assign n9236 = n9216 & n9232;
  assign n9237 = n9235 & n9236;
  assign n9238 = ~P2_IR_REG_20_ & ~P2_IR_REG_22_;
  assign n9239 = ~P2_IR_REG_21_ & n9238;
  assign n9240 = ~P2_IR_REG_18_ & ~P2_IR_REG_19_;
  assign n9241 = ~P2_IR_REG_1_ & n9240;
  assign n9242 = ~P2_IR_REG_0_ & n9241;
  assign n9243 = ~P2_IR_REG_14_ & ~P2_IR_REG_15_;
  assign n9244 = ~P2_IR_REG_16_ & n9243;
  assign n9245 = ~P2_IR_REG_17_ & n9244;
  assign n9246 = n9239 & n9242;
  assign n9247 = n9245 & n9246;
  assign n9248 = n9189 & n9247;
  assign n9249 = n9237 & n9248;
  assign n9250 = P2_IR_REG_29_ & ~n9249;
  assign n9251 = ~P2_IR_REG_27_ & ~P2_IR_REG_28_;
  assign n9252 = ~P2_IR_REG_29_ & n9251;
  assign n9253 = ~P2_IR_REG_2_ & n9252;
  assign n9254 = n9216 & n9253;
  assign n9255 = n9235 & n9254;
  assign n9256 = n9248 & n9255;
  assign n9257 = ~n9250 & ~n9256;
  assign n9258 = n8855 & n9257;
  assign n9259 = P2_IR_REG_29_ & n8854;
  assign n9260 = n2615_1 & ~n3511;
  assign n9261 = P1_DATAO_REG_29_ & ~n2615_1;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~P2_STATE_REG & ~n9262;
  assign n9264 = ~n9258 & ~n9259;
  assign n1480 = n9263 | ~n9264;
  assign n9266 = ~P2_IR_REG_30_ & n9256;
  assign n9267 = P2_IR_REG_30_ & ~n9256;
  assign n9268 = ~n9266 & ~n9267;
  assign n9269 = n8855 & n9268;
  assign n9270 = P2_IR_REG_30_ & n8854;
  assign n9271 = n2615_1 & ~n3535_1;
  assign n9272 = P1_DATAO_REG_30_ & ~n2615_1;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = ~P2_STATE_REG & ~n9273;
  assign n9275 = ~n9269 & ~n9270;
  assign n1485 = n9274 | ~n9275;
  assign n9277 = P2_IR_REG_31_ & n9266;
  assign n9278 = ~P2_IR_REG_31_ & ~n9266;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = n8855 & ~n9279;
  assign n9281 = P2_IR_REG_31_ & n8854;
  assign n9282 = n2615_1 & n3566;
  assign n9283 = P1_DATAO_REG_31_ & ~n2615_1;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = ~P2_STATE_REG & ~n9284;
  assign n9286 = ~n9280 & ~n9281;
  assign n1490 = n9285 | ~n9286;
  assign n9288 = P2_IR_REG_31_ & n9140;
  assign n9289 = P2_IR_REG_23_ & ~P2_IR_REG_31_;
  assign n9290 = ~n9288 & ~n9289;
  assign n9291 = P2_IR_REG_31_ & n9162;
  assign n9292 = P2_IR_REG_25_ & ~P2_IR_REG_31_;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = P2_IR_REG_31_ & n9151;
  assign n9295 = P2_IR_REG_24_ & ~P2_IR_REG_31_;
  assign n9296 = ~n9294 & ~n9295;
  assign n9297 = P2_IR_REG_31_ & n9194;
  assign n9298 = P2_IR_REG_26_ & ~P2_IR_REG_31_;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = ~n9293 & ~n9296;
  assign n9301 = ~n9299 & n9300;
  assign n9302 = n9290 & ~n9301;
  assign n9303 = P2_STATE_REG & n9302;
  assign n9304 = n9293 & ~n9299;
  assign n9305 = ~P2_B_REG & ~n9296;
  assign n9306 = P2_B_REG & n9296;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = n9304 & ~n9307;
  assign n9309 = ~n9299 & ~n9308;
  assign n9310 = n9303 & ~n9309;
  assign n9311 = n9296 & ~n9304;
  assign n9312 = n9310 & ~n9311;
  assign n9313 = P2_D_REG_0_ & ~n9310;
  assign n1495 = n9312 | n9313;
  assign n9315 = n9293 & ~n9304;
  assign n9316 = n9310 & ~n9315;
  assign n9317 = P2_D_REG_1_ & ~n9310;
  assign n1500 = n9316 | n9317;
  assign n1505 = P2_D_REG_2_ & ~n9310;
  assign n1510 = P2_D_REG_3_ & ~n9310;
  assign n1515 = P2_D_REG_4_ & ~n9310;
  assign n1520 = P2_D_REG_5_ & ~n9310;
  assign n1525 = P2_D_REG_6_ & ~n9310;
  assign n1530 = P2_D_REG_7_ & ~n9310;
  assign n1535 = P2_D_REG_8_ & ~n9310;
  assign n1540 = P2_D_REG_9_ & ~n9310;
  assign n1545 = P2_D_REG_10_ & ~n9310;
  assign n1550 = P2_D_REG_11_ & ~n9310;
  assign n1555 = P2_D_REG_12_ & ~n9310;
  assign n1560 = P2_D_REG_13_ & ~n9310;
  assign n1565 = P2_D_REG_14_ & ~n9310;
  assign n1570 = P2_D_REG_15_ & ~n9310;
  assign n1575 = P2_D_REG_16_ & ~n9310;
  assign n1580 = P2_D_REG_17_ & ~n9310;
  assign n1585 = P2_D_REG_18_ & ~n9310;
  assign n1590 = P2_D_REG_19_ & ~n9310;
  assign n1595 = P2_D_REG_20_ & ~n9310;
  assign n1600 = P2_D_REG_21_ & ~n9310;
  assign n1605 = P2_D_REG_22_ & ~n9310;
  assign n1610 = P2_D_REG_23_ & ~n9310;
  assign n1615 = P2_D_REG_24_ & ~n9310;
  assign n1620 = P2_D_REG_25_ & ~n9310;
  assign n1625 = P2_D_REG_26_ & ~n9310;
  assign n1630 = P2_D_REG_27_ & ~n9310;
  assign n1635 = P2_D_REG_28_ & ~n9310;
  assign n1640 = P2_D_REG_29_ & ~n9310;
  assign n1645 = P2_D_REG_30_ & ~n9310;
  assign n1650 = P2_D_REG_31_ & ~n9310;
  assign n9349 = P2_D_REG_0_ & n9309;
  assign n9350 = n9296 & n9299;
  assign n9351 = ~n9309 & ~n9350;
  assign n9352 = ~n9349 & ~n9351;
  assign n9353 = n9303 & n9352;
  assign n9354 = ~n9309 & ~n9315;
  assign n9355 = P2_D_REG_1_ & n9309;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = P2_IR_REG_31_ & n9127;
  assign n9358 = P2_IR_REG_22_ & ~P2_IR_REG_31_;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = P2_IR_REG_31_ & n9116;
  assign n9361 = P2_IR_REG_21_ & ~P2_IR_REG_31_;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = P2_IR_REG_31_ & n9102;
  assign n9364 = P2_IR_REG_20_ & ~P2_IR_REG_31_;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = n9362 & n9365;
  assign n9367 = n9359 & ~n9366;
  assign n9368 = ~n9359 & n9362;
  assign n9369 = P2_IR_REG_31_ & n9091;
  assign n9370 = P2_IR_REG_19_ & ~P2_IR_REG_31_;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = n9365 & n9371;
  assign n9373 = ~n9367 & ~n9368;
  assign n9374 = ~n9372 & n9373;
  assign n9375 = n9356 & ~n9374;
  assign n9376 = P2_D_REG_8_ & n9309;
  assign n9377 = P2_D_REG_7_ & n9309;
  assign n9378 = P2_D_REG_9_ & n9309;
  assign n9379 = ~n9376 & ~n9377;
  assign n9380 = ~n9378 & n9379;
  assign n9381 = P2_D_REG_6_ & n9309;
  assign n9382 = P2_D_REG_5_ & n9309;
  assign n9383 = P2_D_REG_4_ & n9309;
  assign n9384 = P2_D_REG_3_ & n9309;
  assign n9385 = ~n9381 & ~n9382;
  assign n9386 = ~n9383 & n9385;
  assign n9387 = ~n9384 & n9386;
  assign n9388 = P2_D_REG_31_ & n9309;
  assign n9389 = P2_D_REG_30_ & n9309;
  assign n9390 = P2_D_REG_2_ & n9309;
  assign n9391 = P2_D_REG_29_ & n9309;
  assign n9392 = ~n9388 & ~n9389;
  assign n9393 = ~n9390 & n9392;
  assign n9394 = ~n9391 & n9393;
  assign n9395 = P2_D_REG_28_ & n9309;
  assign n9396 = P2_D_REG_27_ & n9309;
  assign n9397 = P2_D_REG_26_ & n9309;
  assign n9398 = P2_D_REG_25_ & n9309;
  assign n9399 = ~n9395 & ~n9396;
  assign n9400 = ~n9397 & n9399;
  assign n9401 = ~n9398 & n9400;
  assign n9402 = n9380 & n9387;
  assign n9403 = n9394 & n9402;
  assign n9404 = n9401 & n9403;
  assign n9405 = P2_D_REG_23_ & n9309;
  assign n9406 = P2_D_REG_22_ & n9309;
  assign n9407 = P2_D_REG_24_ & n9309;
  assign n9408 = ~n9405 & ~n9406;
  assign n9409 = ~n9407 & n9408;
  assign n9410 = P2_D_REG_21_ & n9309;
  assign n9411 = P2_D_REG_20_ & n9309;
  assign n9412 = P2_D_REG_19_ & n9309;
  assign n9413 = P2_D_REG_18_ & n9309;
  assign n9414 = ~n9410 & ~n9411;
  assign n9415 = ~n9412 & n9414;
  assign n9416 = ~n9413 & n9415;
  assign n9417 = P2_D_REG_17_ & n9309;
  assign n9418 = P2_D_REG_16_ & n9309;
  assign n9419 = P2_D_REG_15_ & n9309;
  assign n9420 = P2_D_REG_14_ & n9309;
  assign n9421 = ~n9417 & ~n9418;
  assign n9422 = ~n9419 & n9421;
  assign n9423 = ~n9420 & n9422;
  assign n9424 = P2_D_REG_13_ & n9309;
  assign n9425 = P2_D_REG_12_ & n9309;
  assign n9426 = P2_D_REG_11_ & n9309;
  assign n9427 = P2_D_REG_10_ & n9309;
  assign n9428 = ~n9424 & ~n9425;
  assign n9429 = ~n9426 & n9428;
  assign n9430 = ~n9427 & n9429;
  assign n9431 = n9409 & n9416;
  assign n9432 = n9423 & n9431;
  assign n9433 = n9430 & n9432;
  assign n9434 = n9404 & n9433;
  assign n9435 = n9375 & n9434;
  assign n9436 = n9353 & n9435;
  assign n9437 = P2_IR_REG_0_ & P2_IR_REG_31_;
  assign n9438 = P2_IR_REG_0_ & ~P2_IR_REG_31_;
  assign n9439 = ~n9437 & ~n9438;
  assign n9440 = P2_IR_REG_31_ & n9205;
  assign n9441 = P2_IR_REG_27_ & ~P2_IR_REG_31_;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = P2_IR_REG_31_ & n9222;
  assign n9444 = P2_IR_REG_28_ & ~P2_IR_REG_31_;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = n9442 & n9445;
  assign n9447 = ~n9439 & n9446;
  assign n9448 = ~n8860 & ~n9446;
  assign n9449 = ~n9447 & ~n9448;
  assign n9450 = n9359 & n9362;
  assign n9451 = ~n9371 & n9450;
  assign n9452 = ~n9365 & n9371;
  assign n9453 = n9359 & n9452;
  assign n9454 = n9362 & n9453;
  assign n9455 = ~n9451 & ~n9454;
  assign n9456 = ~n9449 & ~n9455;
  assign n9457 = ~n9359 & ~n9362;
  assign n9458 = n9445 & n9457;
  assign n9459 = P2_IR_REG_31_ & n9268;
  assign n9460 = P2_IR_REG_30_ & ~P2_IR_REG_31_;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = P2_IR_REG_31_ & n9257;
  assign n9463 = P2_IR_REG_29_ & ~P2_IR_REG_31_;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = ~n9461 & ~n9464;
  assign n9466 = P2_REG3_REG_1_ & n9465;
  assign n9467 = n9461 & n9464;
  assign n9468 = P2_REG0_REG_1_ & n9467;
  assign n9469 = n9461 & ~n9464;
  assign n9470 = P2_REG1_REG_1_ & n9469;
  assign n9471 = ~n9461 & n9464;
  assign n9472 = P2_REG2_REG_1_ & n9471;
  assign n9473 = ~n9466 & ~n9468;
  assign n9474 = ~n9470 & n9473;
  assign n9475 = ~n9472 & n9474;
  assign n9476 = n9458 & ~n9475;
  assign n9477 = P2_REG3_REG_0_ & n9465;
  assign n9478 = P2_REG0_REG_0_ & n9467;
  assign n9479 = P2_REG1_REG_0_ & n9469;
  assign n9480 = P2_REG2_REG_0_ & n9471;
  assign n9481 = ~n9477 & ~n9478;
  assign n9482 = ~n9479 & n9481;
  assign n9483 = ~n9480 & n9482;
  assign n9484 = ~n9449 & n9483;
  assign n9485 = n9449 & ~n9483;
  assign n9486 = ~n9484 & ~n9485;
  assign n9487 = n9359 & ~n9371;
  assign n9488 = n9365 & n9487;
  assign n9489 = ~n9486 & n9488;
  assign n9490 = n9365 & n9450;
  assign n9491 = ~n9449 & n9490;
  assign n9492 = ~n9489 & ~n9491;
  assign n9493 = n9362 & n9371;
  assign n9494 = ~n9359 & n9493;
  assign n9495 = n9365 & n9494;
  assign n9496 = ~n9486 & n9495;
  assign n9497 = ~n9362 & n9452;
  assign n9498 = ~n9486 & n9497;
  assign n9499 = ~n9496 & ~n9498;
  assign n9500 = ~n9362 & n9372;
  assign n9501 = n9359 & n9500;
  assign n9502 = ~n9486 & n9501;
  assign n9503 = ~n9365 & ~n9371;
  assign n9504 = ~n9362 & n9503;
  assign n9505 = ~n9486 & n9504;
  assign n9506 = ~n9359 & n9452;
  assign n9507 = ~n9486 & n9506;
  assign n9508 = ~n9359 & n9503;
  assign n9509 = ~n9486 & n9508;
  assign n9510 = n9365 & ~n9371;
  assign n9511 = ~n9359 & n9510;
  assign n9512 = ~n9486 & n9511;
  assign n9513 = ~n9505 & ~n9507;
  assign n9514 = ~n9509 & n9513;
  assign n9515 = ~n9512 & n9514;
  assign n9516 = n9499 & ~n9502;
  assign n9517 = n9515 & n9516;
  assign n9518 = ~n9456 & ~n9476;
  assign n9519 = n9492 & n9518;
  assign n9520 = n9517 & n9519;
  assign n9521 = n9436 & ~n9520;
  assign n9522 = P2_REG0_REG_0_ & ~n9436;
  assign n1655 = n9521 | n9522;
  assign n9524 = P2_REG3_REG_2_ & n9465;
  assign n9525 = P2_REG0_REG_2_ & n9467;
  assign n9526 = P2_REG1_REG_2_ & n9469;
  assign n9527 = P2_REG2_REG_2_ & n9471;
  assign n9528 = ~n9524 & ~n9525;
  assign n9529 = ~n9526 & n9528;
  assign n9530 = ~n9527 & n9529;
  assign n9531 = n9458 & ~n9530;
  assign n9532 = P2_IR_REG_31_ & ~n8866;
  assign n9533 = P2_IR_REG_1_ & ~P2_IR_REG_31_;
  assign n9534 = ~n9532 & ~n9533;
  assign n9535 = n9446 & ~n9534;
  assign n9536 = ~n8871 & ~n9446;
  assign n9537 = ~n9535 & ~n9536;
  assign n9538 = ~n9449 & n9537;
  assign n9539 = n9449 & ~n9537;
  assign n9540 = ~n9538 & ~n9539;
  assign n9541 = n9490 & ~n9540;
  assign n9542 = ~n9455 & ~n9537;
  assign n9543 = ~n9475 & ~n9537;
  assign n9544 = n9475 & n9537;
  assign n9545 = ~n9543 & ~n9544;
  assign n9546 = ~n9449 & ~n9483;
  assign n9547 = n9545 & ~n9546;
  assign n9548 = ~n9545 & n9546;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = n9488 & ~n9549;
  assign n9551 = ~n9531 & ~n9541;
  assign n9552 = ~n9542 & n9551;
  assign n9553 = ~n9550 & n9552;
  assign n9554 = ~n9475 & n9537;
  assign n9555 = n9475 & ~n9537;
  assign n9556 = ~n9554 & ~n9555;
  assign n9557 = ~n9484 & ~n9556;
  assign n9558 = n9484 & n9556;
  assign n9559 = ~n9557 & ~n9558;
  assign n9560 = n9511 & ~n9559;
  assign n9561 = ~n9445 & n9457;
  assign n9562 = ~n9483 & n9561;
  assign n9563 = n9506 & ~n9549;
  assign n9564 = n9508 & ~n9559;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = n9501 & ~n9549;
  assign n9567 = n9495 & ~n9549;
  assign n9568 = n9497 & ~n9559;
  assign n9569 = n9504 & ~n9559;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 = ~n9566 & ~n9567;
  assign n9572 = n9570 & n9571;
  assign n9573 = ~n9560 & ~n9562;
  assign n9574 = n9565 & n9573;
  assign n9575 = n9572 & n9574;
  assign n9576 = n9553 & n9575;
  assign n9577 = n9436 & ~n9576;
  assign n9578 = P2_REG0_REG_1_ & ~n9436;
  assign n1660 = n9577 | n9578;
  assign n9580 = ~P2_REG3_REG_3_ & n9465;
  assign n9581 = P2_REG0_REG_3_ & n9467;
  assign n9582 = P2_REG1_REG_3_ & n9469;
  assign n9583 = P2_REG2_REG_3_ & n9471;
  assign n9584 = ~n9580 & ~n9581;
  assign n9585 = ~n9582 & n9584;
  assign n9586 = ~n9583 & n9585;
  assign n9587 = n9458 & ~n9586;
  assign n9588 = P2_IR_REG_31_ & n8878;
  assign n9589 = P2_IR_REG_2_ & ~P2_IR_REG_31_;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = n9446 & ~n9590;
  assign n9592 = ~n8883 & ~n9446;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = n9449 & n9537;
  assign n9595 = ~n9593 & ~n9594;
  assign n9596 = n9593 & n9594;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = n9490 & n9597;
  assign n9599 = ~n9455 & ~n9593;
  assign n9600 = ~n9530 & ~n9593;
  assign n9601 = n9530 & n9593;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = ~n9544 & n9546;
  assign n9604 = ~n9543 & ~n9603;
  assign n9605 = n9602 & ~n9604;
  assign n9606 = n9530 & ~n9593;
  assign n9607 = ~n9530 & n9593;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~n9543 & n9608;
  assign n9610 = ~n9603 & n9609;
  assign n9611 = ~n9605 & ~n9610;
  assign n9612 = n9488 & n9611;
  assign n9613 = ~n9587 & ~n9598;
  assign n9614 = ~n9599 & n9613;
  assign n9615 = ~n9612 & n9614;
  assign n9616 = ~n9475 & ~n9484;
  assign n9617 = ~n9484 & n9537;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = ~n9554 & n9618;
  assign n9620 = n9608 & n9619;
  assign n9621 = ~n9608 & ~n9619;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = n9511 & ~n9622;
  assign n9624 = ~n9475 & n9561;
  assign n9625 = n9506 & n9611;
  assign n9626 = n9508 & ~n9622;
  assign n9627 = ~n9625 & ~n9626;
  assign n9628 = n9501 & n9611;
  assign n9629 = n9495 & n9611;
  assign n9630 = n9497 & ~n9622;
  assign n9631 = n9504 & ~n9622;
  assign n9632 = ~n9630 & ~n9631;
  assign n9633 = ~n9628 & ~n9629;
  assign n9634 = n9632 & n9633;
  assign n9635 = ~n9623 & ~n9624;
  assign n9636 = n9627 & n9635;
  assign n9637 = n9634 & n9636;
  assign n9638 = n9615 & n9637;
  assign n9639 = n9436 & ~n9638;
  assign n9640 = P2_REG0_REG_2_ & ~n9436;
  assign n1665 = n9639 | n9640;
  assign n9642 = ~P2_REG3_REG_4_ & P2_REG3_REG_3_;
  assign n9643 = P2_REG3_REG_4_ & ~P2_REG3_REG_3_;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = n9465 & ~n9644;
  assign n9646 = P2_REG0_REG_4_ & n9467;
  assign n9647 = P2_REG1_REG_4_ & n9469;
  assign n9648 = P2_REG2_REG_4_ & n9471;
  assign n9649 = ~n9645 & ~n9646;
  assign n9650 = ~n9647 & n9649;
  assign n9651 = ~n9648 & n9650;
  assign n9652 = n9458 & ~n9651;
  assign n9653 = P2_IR_REG_31_ & n8889;
  assign n9654 = P2_IR_REG_3_ & ~P2_IR_REG_31_;
  assign n9655 = ~n9653 & ~n9654;
  assign n9656 = n9446 & ~n9655;
  assign n9657 = ~n8894 & ~n9446;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = ~n9596 & ~n9658;
  assign n9660 = n9596 & n9658;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = n9490 & n9661;
  assign n9663 = ~n9455 & ~n9658;
  assign n9664 = n9543 & ~n9601;
  assign n9665 = ~n9600 & ~n9664;
  assign n9666 = ~n9601 & n9603;
  assign n9667 = n9665 & ~n9666;
  assign n9668 = n9586 & ~n9658;
  assign n9669 = ~n9586 & n9658;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = n9667 & ~n9670;
  assign n9672 = ~n9586 & ~n9658;
  assign n9673 = n9586 & n9658;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = ~n9667 & ~n9674;
  assign n9676 = ~n9671 & ~n9675;
  assign n9677 = n9488 & ~n9676;
  assign n9678 = ~n9652 & ~n9662;
  assign n9679 = ~n9663 & n9678;
  assign n9680 = ~n9677 & n9679;
  assign n9681 = ~n9606 & ~n9670;
  assign n9682 = ~n9607 & n9619;
  assign n9683 = n9681 & ~n9682;
  assign n9684 = ~n9607 & n9670;
  assign n9685 = ~n9606 & ~n9619;
  assign n9686 = n9684 & ~n9685;
  assign n9687 = ~n9683 & ~n9686;
  assign n9688 = n9511 & ~n9687;
  assign n9689 = ~n9530 & n9561;
  assign n9690 = n9506 & ~n9676;
  assign n9691 = n9508 & ~n9687;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = n9501 & ~n9676;
  assign n9694 = n9495 & ~n9676;
  assign n9695 = n9497 & ~n9687;
  assign n9696 = n9504 & ~n9687;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n9693 & ~n9694;
  assign n9699 = n9697 & n9698;
  assign n9700 = ~n9688 & ~n9689;
  assign n9701 = n9692 & n9700;
  assign n9702 = n9699 & n9701;
  assign n9703 = n9680 & n9702;
  assign n9704 = n9436 & ~n9703;
  assign n9705 = P2_REG0_REG_3_ & ~n9436;
  assign n1670 = n9704 | n9705;
  assign n9707 = P2_REG3_REG_4_ & P2_REG3_REG_3_;
  assign n9708 = ~P2_REG3_REG_5_ & n9707;
  assign n9709 = P2_REG3_REG_5_ & ~n9707;
  assign n9710 = ~n9708 & ~n9709;
  assign n9711 = n9465 & ~n9710;
  assign n9712 = P2_REG0_REG_5_ & n9467;
  assign n9713 = P2_REG1_REG_5_ & n9469;
  assign n9714 = P2_REG2_REG_5_ & n9471;
  assign n9715 = ~n9711 & ~n9712;
  assign n9716 = ~n9713 & n9715;
  assign n9717 = ~n9714 & n9716;
  assign n9718 = n9458 & ~n9717;
  assign n9719 = P2_IR_REG_31_ & n8901;
  assign n9720 = P2_IR_REG_4_ & ~P2_IR_REG_31_;
  assign n9721 = ~n9719 & ~n9720;
  assign n9722 = n9446 & ~n9721;
  assign n9723 = ~n8906 & ~n9446;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = ~n9660 & ~n9724;
  assign n9726 = n9660 & n9724;
  assign n9727 = ~n9725 & ~n9726;
  assign n9728 = n9490 & n9727;
  assign n9729 = ~n9455 & ~n9724;
  assign n9730 = n9651 & ~n9724;
  assign n9731 = ~n9651 & n9724;
  assign n9732 = ~n9730 & ~n9731;
  assign n9733 = ~n9601 & ~n9673;
  assign n9734 = n9603 & n9733;
  assign n9735 = ~n9672 & ~n9734;
  assign n9736 = ~n9665 & ~n9673;
  assign n9737 = n9735 & ~n9736;
  assign n9738 = ~n9732 & n9737;
  assign n9739 = n9651 & n9724;
  assign n9740 = ~n9651 & ~n9724;
  assign n9741 = ~n9739 & ~n9740;
  assign n9742 = ~n9737 & ~n9741;
  assign n9743 = ~n9738 & ~n9742;
  assign n9744 = n9488 & ~n9743;
  assign n9745 = ~n9718 & ~n9728;
  assign n9746 = ~n9729 & n9745;
  assign n9747 = ~n9744 & n9746;
  assign n9748 = n9586 & ~n9607;
  assign n9749 = n9658 & ~n9748;
  assign n9750 = ~n9586 & n9607;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = ~n9606 & ~n9668;
  assign n9753 = ~n9619 & n9752;
  assign n9754 = n9751 & ~n9753;
  assign n9755 = n9732 & n9754;
  assign n9756 = ~n9732 & ~n9754;
  assign n9757 = ~n9755 & ~n9756;
  assign n9758 = n9511 & ~n9757;
  assign n9759 = n9561 & ~n9586;
  assign n9760 = n9506 & ~n9743;
  assign n9761 = n9508 & ~n9757;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = n9501 & ~n9743;
  assign n9764 = n9495 & ~n9743;
  assign n9765 = n9497 & ~n9757;
  assign n9766 = n9504 & ~n9757;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = ~n9763 & ~n9764;
  assign n9769 = n9767 & n9768;
  assign n9770 = ~n9758 & ~n9759;
  assign n9771 = n9762 & n9770;
  assign n9772 = n9769 & n9771;
  assign n9773 = n9747 & n9772;
  assign n9774 = n9436 & ~n9773;
  assign n9775 = P2_REG0_REG_4_ & ~n9436;
  assign n1675 = n9774 | n9775;
  assign n9777 = P2_REG3_REG_5_ & P2_REG3_REG_3_;
  assign n9778 = P2_REG3_REG_4_ & n9777;
  assign n9779 = ~P2_REG3_REG_6_ & n9778;
  assign n9780 = P2_REG3_REG_6_ & ~n9778;
  assign n9781 = ~n9779 & ~n9780;
  assign n9782 = n9465 & ~n9781;
  assign n9783 = P2_REG0_REG_6_ & n9467;
  assign n9784 = P2_REG1_REG_6_ & n9469;
  assign n9785 = P2_REG2_REG_6_ & n9471;
  assign n9786 = ~n9782 & ~n9783;
  assign n9787 = ~n9784 & n9786;
  assign n9788 = ~n9785 & n9787;
  assign n9789 = n9458 & ~n9788;
  assign n9790 = P2_IR_REG_31_ & n8912;
  assign n9791 = P2_IR_REG_5_ & ~P2_IR_REG_31_;
  assign n9792 = ~n9790 & ~n9791;
  assign n9793 = n9446 & ~n9792;
  assign n9794 = ~n8917 & ~n9446;
  assign n9795 = ~n9793 & ~n9794;
  assign n9796 = n9726 & n9795;
  assign n9797 = ~n9726 & ~n9795;
  assign n9798 = ~n9796 & ~n9797;
  assign n9799 = n9490 & n9798;
  assign n9800 = ~n9455 & ~n9795;
  assign n9801 = ~n9717 & ~n9795;
  assign n9802 = n9717 & n9795;
  assign n9803 = ~n9739 & ~n9802;
  assign n9804 = ~n9801 & n9803;
  assign n9805 = n9737 & ~n9740;
  assign n9806 = n9804 & ~n9805;
  assign n9807 = n9717 & ~n9795;
  assign n9808 = ~n9717 & n9795;
  assign n9809 = ~n9807 & ~n9808;
  assign n9810 = ~n9740 & n9809;
  assign n9811 = ~n9737 & ~n9739;
  assign n9812 = n9810 & ~n9811;
  assign n9813 = ~n9806 & ~n9812;
  assign n9814 = n9488 & n9813;
  assign n9815 = ~n9789 & ~n9799;
  assign n9816 = ~n9800 & n9815;
  assign n9817 = ~n9814 & n9816;
  assign n9818 = ~n9730 & ~n9754;
  assign n9819 = ~n9731 & ~n9818;
  assign n9820 = n9809 & n9819;
  assign n9821 = ~n9809 & ~n9819;
  assign n9822 = ~n9820 & ~n9821;
  assign n9823 = n9511 & ~n9822;
  assign n9824 = n9561 & ~n9651;
  assign n9825 = n9506 & n9813;
  assign n9826 = n9508 & ~n9822;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = n9501 & n9813;
  assign n9829 = n9495 & n9813;
  assign n9830 = n9497 & ~n9822;
  assign n9831 = n9504 & ~n9822;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = ~n9828 & ~n9829;
  assign n9834 = n9832 & n9833;
  assign n9835 = ~n9823 & ~n9824;
  assign n9836 = n9827 & n9835;
  assign n9837 = n9834 & n9836;
  assign n9838 = n9817 & n9837;
  assign n9839 = n9436 & ~n9838;
  assign n9840 = P2_REG0_REG_5_ & ~n9436;
  assign n1680 = n9839 | n9840;
  assign n9842 = P2_REG3_REG_6_ & n9778;
  assign n9843 = ~P2_REG3_REG_7_ & n9842;
  assign n9844 = P2_REG3_REG_7_ & ~n9842;
  assign n9845 = ~n9843 & ~n9844;
  assign n9846 = n9465 & ~n9845;
  assign n9847 = P2_REG0_REG_7_ & n9467;
  assign n9848 = P2_REG1_REG_7_ & n9469;
  assign n9849 = P2_REG2_REG_7_ & n9471;
  assign n9850 = ~n9846 & ~n9847;
  assign n9851 = ~n9848 & n9850;
  assign n9852 = ~n9849 & n9851;
  assign n9853 = n9458 & ~n9852;
  assign n9854 = P2_IR_REG_31_ & n8924;
  assign n9855 = P2_IR_REG_6_ & ~P2_IR_REG_31_;
  assign n9856 = ~n9854 & ~n9855;
  assign n9857 = n9446 & ~n9856;
  assign n9858 = ~n8929 & ~n9446;
  assign n9859 = ~n9857 & ~n9858;
  assign n9860 = ~n9796 & ~n9859;
  assign n9861 = n9795 & n9859;
  assign n9862 = n9726 & n9861;
  assign n9863 = ~n9860 & ~n9862;
  assign n9864 = n9490 & n9863;
  assign n9865 = ~n9455 & ~n9859;
  assign n9866 = n9788 & ~n9859;
  assign n9867 = ~n9788 & n9859;
  assign n9868 = ~n9866 & ~n9867;
  assign n9869 = n9740 & ~n9795;
  assign n9870 = ~n9740 & n9795;
  assign n9871 = ~n9717 & ~n9870;
  assign n9872 = ~n9869 & ~n9871;
  assign n9873 = n9600 & ~n9673;
  assign n9874 = ~n9672 & ~n9873;
  assign n9875 = ~n9604 & n9733;
  assign n9876 = n9874 & ~n9875;
  assign n9877 = n9803 & ~n9876;
  assign n9878 = n9872 & ~n9877;
  assign n9879 = ~n9868 & n9878;
  assign n9880 = n9788 & n9859;
  assign n9881 = ~n9788 & ~n9859;
  assign n9882 = ~n9880 & ~n9881;
  assign n9883 = ~n9878 & ~n9882;
  assign n9884 = ~n9879 & ~n9883;
  assign n9885 = n9488 & ~n9884;
  assign n9886 = ~n9853 & ~n9864;
  assign n9887 = ~n9865 & n9886;
  assign n9888 = ~n9885 & n9887;
  assign n9889 = ~n9807 & ~n9868;
  assign n9890 = ~n9808 & n9819;
  assign n9891 = n9889 & ~n9890;
  assign n9892 = ~n9808 & ~n9867;
  assign n9893 = ~n9866 & n9892;
  assign n9894 = ~n9807 & ~n9819;
  assign n9895 = n9893 & ~n9894;
  assign n9896 = ~n9891 & ~n9895;
  assign n9897 = n9511 & ~n9896;
  assign n9898 = n9561 & ~n9717;
  assign n9899 = ~n9673 & n9803;
  assign n9900 = ~n9600 & ~n9672;
  assign n9901 = ~n9601 & ~n9604;
  assign n9902 = n9900 & ~n9901;
  assign n9903 = n9899 & ~n9902;
  assign n9904 = n9872 & ~n9903;
  assign n9905 = ~n9868 & n9904;
  assign n9906 = ~n9882 & ~n9904;
  assign n9907 = ~n9905 & ~n9906;
  assign n9908 = n9506 & ~n9907;
  assign n9909 = n9508 & ~n9896;
  assign n9910 = ~n9908 & ~n9909;
  assign n9911 = n9501 & ~n9907;
  assign n9912 = n9495 & ~n9907;
  assign n9913 = n9497 & ~n9896;
  assign n9914 = n9504 & ~n9896;
  assign n9915 = ~n9913 & ~n9914;
  assign n9916 = ~n9911 & ~n9912;
  assign n9917 = n9915 & n9916;
  assign n9918 = ~n9897 & ~n9898;
  assign n9919 = n9910 & n9918;
  assign n9920 = n9917 & n9919;
  assign n9921 = n9888 & n9920;
  assign n9922 = n9436 & ~n9921;
  assign n9923 = P2_REG0_REG_6_ & ~n9436;
  assign n1685 = n9922 | n9923;
  assign n9925 = P2_REG3_REG_6_ & P2_REG3_REG_7_;
  assign n9926 = n9778 & n9925;
  assign n9927 = ~P2_REG3_REG_8_ & n9926;
  assign n9928 = P2_REG3_REG_8_ & ~n9926;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = n9465 & ~n9929;
  assign n9931 = P2_REG0_REG_8_ & n9467;
  assign n9932 = P2_REG1_REG_8_ & n9469;
  assign n9933 = P2_REG2_REG_8_ & n9471;
  assign n9934 = ~n9930 & ~n9931;
  assign n9935 = ~n9932 & n9934;
  assign n9936 = ~n9933 & n9935;
  assign n9937 = n9458 & ~n9936;
  assign n9938 = P2_IR_REG_31_ & n8935;
  assign n9939 = P2_IR_REG_7_ & ~P2_IR_REG_31_;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = n9446 & ~n9940;
  assign n9942 = ~n8940 & ~n9446;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = ~n9862 & ~n9943;
  assign n9945 = n9862 & n9943;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = n9490 & n9946;
  assign n9948 = ~n9455 & ~n9943;
  assign n9949 = ~n9852 & ~n9943;
  assign n9950 = n9852 & n9943;
  assign n9951 = ~n9880 & ~n9950;
  assign n9952 = ~n9949 & n9951;
  assign n9953 = n9878 & ~n9881;
  assign n9954 = n9952 & ~n9953;
  assign n9955 = n9852 & ~n9943;
  assign n9956 = ~n9852 & n9943;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~n9881 & n9957;
  assign n9959 = ~n9878 & ~n9880;
  assign n9960 = n9958 & ~n9959;
  assign n9961 = ~n9954 & ~n9960;
  assign n9962 = n9488 & n9961;
  assign n9963 = ~n9937 & ~n9947;
  assign n9964 = ~n9948 & n9963;
  assign n9965 = ~n9962 & n9964;
  assign n9966 = n9731 & ~n9807;
  assign n9967 = n9892 & ~n9966;
  assign n9968 = ~n9866 & ~n9967;
  assign n9969 = ~n9730 & ~n9866;
  assign n9970 = ~n9807 & n9969;
  assign n9971 = ~n9754 & n9970;
  assign n9972 = ~n9968 & ~n9971;
  assign n9973 = n9957 & n9972;
  assign n9974 = ~n9957 & ~n9972;
  assign n9975 = ~n9973 & ~n9974;
  assign n9976 = n9511 & ~n9975;
  assign n9977 = n9561 & ~n9788;
  assign n9978 = ~n9881 & n9904;
  assign n9979 = n9952 & ~n9978;
  assign n9980 = ~n9880 & ~n9904;
  assign n9981 = n9958 & ~n9980;
  assign n9982 = ~n9979 & ~n9981;
  assign n9983 = n9506 & n9982;
  assign n9984 = n9508 & ~n9975;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = n9501 & n9982;
  assign n9987 = n9495 & n9982;
  assign n9988 = n9497 & ~n9975;
  assign n9989 = n9504 & ~n9975;
  assign n9990 = ~n9988 & ~n9989;
  assign n9991 = ~n9986 & ~n9987;
  assign n9992 = n9990 & n9991;
  assign n9993 = ~n9976 & ~n9977;
  assign n9994 = n9985 & n9993;
  assign n9995 = n9992 & n9994;
  assign n9996 = n9965 & n9995;
  assign n9997 = n9436 & ~n9996;
  assign n9998 = P2_REG0_REG_7_ & ~n9436;
  assign n1690 = n9997 | n9998;
  assign n10000 = P2_REG3_REG_8_ & n9926;
  assign n10001 = ~P2_REG3_REG_9_ & n10000;
  assign n10002 = P2_REG3_REG_9_ & ~n10000;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = n9465 & ~n10003;
  assign n10005 = P2_REG0_REG_9_ & n9467;
  assign n10006 = P2_REG1_REG_9_ & n9469;
  assign n10007 = P2_REG2_REG_9_ & n9471;
  assign n10008 = ~n10004 & ~n10005;
  assign n10009 = ~n10006 & n10008;
  assign n10010 = ~n10007 & n10009;
  assign n10011 = n9458 & ~n10010;
  assign n10012 = P2_IR_REG_31_ & n8950;
  assign n10013 = P2_IR_REG_8_ & ~P2_IR_REG_31_;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = n9446 & ~n10014;
  assign n10016 = ~n8955 & ~n9446;
  assign n10017 = ~n10015 & ~n10016;
  assign n10018 = ~n9945 & ~n10017;
  assign n10019 = n9945 & n10017;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = n9490 & n10020;
  assign n10022 = ~n9455 & ~n10017;
  assign n10023 = n9881 & ~n9943;
  assign n10024 = ~n9881 & n9943;
  assign n10025 = ~n9852 & ~n10024;
  assign n10026 = ~n10023 & ~n10025;
  assign n10027 = ~n9878 & n9951;
  assign n10028 = n10026 & ~n10027;
  assign n10029 = n9936 & ~n10017;
  assign n10030 = ~n9936 & n10017;
  assign n10031 = ~n10029 & ~n10030;
  assign n10032 = n10028 & ~n10031;
  assign n10033 = n9936 & n10017;
  assign n10034 = ~n9936 & ~n10017;
  assign n10035 = ~n10033 & ~n10034;
  assign n10036 = ~n10028 & ~n10035;
  assign n10037 = ~n10032 & ~n10036;
  assign n10038 = n9488 & ~n10037;
  assign n10039 = ~n10011 & ~n10021;
  assign n10040 = ~n10022 & n10039;
  assign n10041 = ~n10038 & n10040;
  assign n10042 = ~n9955 & ~n10031;
  assign n10043 = ~n9956 & n9972;
  assign n10044 = n10042 & ~n10043;
  assign n10045 = ~n9956 & n10031;
  assign n10046 = ~n9955 & ~n9972;
  assign n10047 = n10045 & ~n10046;
  assign n10048 = ~n10044 & ~n10047;
  assign n10049 = n9511 & ~n10048;
  assign n10050 = n9561 & ~n9852;
  assign n10051 = ~n9904 & n9951;
  assign n10052 = n10026 & ~n10051;
  assign n10053 = ~n10031 & n10052;
  assign n10054 = ~n10035 & ~n10052;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n9506 & ~n10055;
  assign n10057 = n9508 & ~n10048;
  assign n10058 = ~n10056 & ~n10057;
  assign n10059 = n9501 & ~n10055;
  assign n10060 = n9495 & ~n10055;
  assign n10061 = n9497 & ~n10048;
  assign n10062 = n9504 & ~n10048;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10059 & ~n10060;
  assign n10065 = n10063 & n10064;
  assign n10066 = ~n10049 & ~n10050;
  assign n10067 = n10058 & n10066;
  assign n10068 = n10065 & n10067;
  assign n10069 = n10041 & n10068;
  assign n10070 = n9436 & ~n10069;
  assign n10071 = P2_REG0_REG_8_ & ~n9436;
  assign n1695 = n10070 | n10071;
  assign n10073 = P2_REG3_REG_9_ & P2_REG3_REG_8_;
  assign n10074 = n9926 & n10073;
  assign n10075 = ~P2_REG3_REG_10_ & n10074;
  assign n10076 = P2_REG3_REG_10_ & ~n10074;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = n9465 & ~n10077;
  assign n10079 = P2_REG0_REG_10_ & n9467;
  assign n10080 = P2_REG1_REG_10_ & n9469;
  assign n10081 = P2_REG2_REG_10_ & n9471;
  assign n10082 = ~n10078 & ~n10079;
  assign n10083 = ~n10080 & n10082;
  assign n10084 = ~n10081 & n10083;
  assign n10085 = n9458 & ~n10084;
  assign n10086 = P2_IR_REG_31_ & n8961;
  assign n10087 = P2_IR_REG_9_ & ~P2_IR_REG_31_;
  assign n10088 = ~n10086 & ~n10087;
  assign n10089 = n9446 & ~n10088;
  assign n10090 = ~n8966 & ~n9446;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = n10019 & n10091;
  assign n10093 = ~n10019 & ~n10091;
  assign n10094 = ~n10092 & ~n10093;
  assign n10095 = n9490 & n10094;
  assign n10096 = ~n9455 & ~n10091;
  assign n10097 = n10010 & ~n10091;
  assign n10098 = ~n10010 & n10091;
  assign n10099 = ~n10097 & ~n10098;
  assign n10100 = ~n10028 & ~n10033;
  assign n10101 = ~n10034 & ~n10100;
  assign n10102 = ~n10099 & n10101;
  assign n10103 = n10010 & n10091;
  assign n10104 = ~n10010 & ~n10091;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = ~n10101 & ~n10105;
  assign n10107 = ~n10102 & ~n10106;
  assign n10108 = n9488 & ~n10107;
  assign n10109 = ~n10085 & ~n10095;
  assign n10110 = ~n10096 & n10109;
  assign n10111 = ~n10108 & n10110;
  assign n10112 = n9936 & ~n9956;
  assign n10113 = n10017 & ~n10112;
  assign n10114 = ~n9936 & n9956;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~n9955 & ~n10029;
  assign n10117 = ~n9972 & n10116;
  assign n10118 = n10115 & ~n10117;
  assign n10119 = n10099 & n10118;
  assign n10120 = ~n10099 & ~n10118;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 = n9511 & ~n10121;
  assign n10123 = n9561 & ~n9936;
  assign n10124 = ~n10033 & ~n10052;
  assign n10125 = ~n10034 & ~n10124;
  assign n10126 = ~n10099 & n10125;
  assign n10127 = ~n10105 & ~n10125;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = n9506 & ~n10128;
  assign n10130 = n9508 & ~n10121;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = n9501 & ~n10128;
  assign n10133 = n9495 & ~n10128;
  assign n10134 = n9497 & ~n10121;
  assign n10135 = n9504 & ~n10121;
  assign n10136 = ~n10134 & ~n10135;
  assign n10137 = ~n10132 & ~n10133;
  assign n10138 = n10136 & n10137;
  assign n10139 = ~n10122 & ~n10123;
  assign n10140 = n10131 & n10139;
  assign n10141 = n10138 & n10140;
  assign n10142 = n10111 & n10141;
  assign n10143 = n9436 & ~n10142;
  assign n10144 = P2_REG0_REG_9_ & ~n9436;
  assign n1700 = n10143 | n10144;
  assign n10146 = P2_REG3_REG_10_ & n10074;
  assign n10147 = ~P2_REG3_REG_11_ & n10146;
  assign n10148 = P2_REG3_REG_11_ & ~n10146;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = n9465 & ~n10149;
  assign n10151 = P2_REG0_REG_11_ & n9467;
  assign n10152 = P2_REG1_REG_11_ & n9469;
  assign n10153 = P2_REG2_REG_11_ & n9471;
  assign n10154 = ~n10150 & ~n10151;
  assign n10155 = ~n10152 & n10154;
  assign n10156 = ~n10153 & n10155;
  assign n10157 = n9458 & ~n10156;
  assign n10158 = P2_IR_REG_31_ & n8973;
  assign n10159 = P2_IR_REG_10_ & ~P2_IR_REG_31_;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = n9446 & ~n10160;
  assign n10162 = ~n8978 & ~n9446;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = ~n10092 & ~n10163;
  assign n10165 = n10091 & n10163;
  assign n10166 = n10019 & n10165;
  assign n10167 = ~n10164 & ~n10166;
  assign n10168 = n9490 & n10167;
  assign n10169 = ~n9455 & ~n10163;
  assign n10170 = ~n10084 & ~n10163;
  assign n10171 = n10084 & n10163;
  assign n10172 = ~n10103 & ~n10171;
  assign n10173 = ~n10170 & n10172;
  assign n10174 = n10101 & ~n10104;
  assign n10175 = n10173 & ~n10174;
  assign n10176 = n10084 & ~n10163;
  assign n10177 = ~n10084 & n10163;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10104 & n10178;
  assign n10180 = ~n10101 & ~n10103;
  assign n10181 = n10179 & ~n10180;
  assign n10182 = ~n10175 & ~n10181;
  assign n10183 = n9488 & n10182;
  assign n10184 = ~n10157 & ~n10168;
  assign n10185 = ~n10169 & n10184;
  assign n10186 = ~n10183 & n10185;
  assign n10187 = ~n10097 & ~n10118;
  assign n10188 = ~n10098 & ~n10187;
  assign n10189 = n10178 & n10188;
  assign n10190 = ~n10178 & ~n10188;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = n9511 & ~n10191;
  assign n10193 = n9561 & ~n10010;
  assign n10194 = ~n10104 & n10125;
  assign n10195 = n10173 & ~n10194;
  assign n10196 = ~n10103 & ~n10125;
  assign n10197 = n10179 & ~n10196;
  assign n10198 = ~n10195 & ~n10197;
  assign n10199 = n9506 & n10198;
  assign n10200 = n9508 & ~n10191;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = n9501 & n10198;
  assign n10203 = n9495 & n10198;
  assign n10204 = n9497 & ~n10191;
  assign n10205 = n9504 & ~n10191;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = ~n10202 & ~n10203;
  assign n10208 = n10206 & n10207;
  assign n10209 = ~n10192 & ~n10193;
  assign n10210 = n10201 & n10209;
  assign n10211 = n10208 & n10210;
  assign n10212 = n10186 & n10211;
  assign n10213 = n9436 & ~n10212;
  assign n10214 = P2_REG0_REG_10_ & ~n9436;
  assign n1705 = n10213 | n10214;
  assign n10216 = P2_REG3_REG_11_ & P2_REG3_REG_10_;
  assign n10217 = n10074 & n10216;
  assign n10218 = ~P2_REG3_REG_12_ & n10217;
  assign n10219 = P2_REG3_REG_12_ & ~n10217;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = n9465 & ~n10220;
  assign n10222 = P2_REG0_REG_12_ & n9467;
  assign n10223 = P2_REG1_REG_12_ & n9469;
  assign n10224 = P2_REG2_REG_12_ & n9471;
  assign n10225 = ~n10221 & ~n10222;
  assign n10226 = ~n10223 & n10225;
  assign n10227 = ~n10224 & n10226;
  assign n10228 = n9458 & ~n10227;
  assign n10229 = P2_IR_REG_31_ & n8984;
  assign n10230 = P2_IR_REG_11_ & ~P2_IR_REG_31_;
  assign n10231 = ~n10229 & ~n10230;
  assign n10232 = n9446 & ~n10231;
  assign n10233 = ~n8989 & ~n9446;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = ~n10166 & ~n10234;
  assign n10236 = n10166 & n10234;
  assign n10237 = ~n10235 & ~n10236;
  assign n10238 = n9490 & n10237;
  assign n10239 = ~n9455 & ~n10234;
  assign n10240 = ~n10104 & ~n10170;
  assign n10241 = n10034 & n10172;
  assign n10242 = n10240 & ~n10241;
  assign n10243 = ~n10171 & ~n10242;
  assign n10244 = ~n10033 & n10172;
  assign n10245 = ~n10028 & n10244;
  assign n10246 = ~n10243 & ~n10245;
  assign n10247 = n10156 & ~n10234;
  assign n10248 = ~n10156 & n10234;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = n10246 & ~n10249;
  assign n10251 = n10156 & n10234;
  assign n10252 = ~n10156 & ~n10234;
  assign n10253 = ~n10251 & ~n10252;
  assign n10254 = ~n10246 & ~n10253;
  assign n10255 = ~n10250 & ~n10254;
  assign n10256 = n9488 & ~n10255;
  assign n10257 = ~n10228 & ~n10238;
  assign n10258 = ~n10239 & n10257;
  assign n10259 = ~n10256 & n10258;
  assign n10260 = ~n10176 & ~n10249;
  assign n10261 = ~n10177 & n10188;
  assign n10262 = n10260 & ~n10261;
  assign n10263 = ~n10177 & ~n10248;
  assign n10264 = ~n10247 & n10263;
  assign n10265 = ~n10176 & ~n10188;
  assign n10266 = n10264 & ~n10265;
  assign n10267 = ~n10262 & ~n10266;
  assign n10268 = n9511 & ~n10267;
  assign n10269 = n9561 & ~n10084;
  assign n10270 = ~n10052 & n10244;
  assign n10271 = ~n10243 & ~n10270;
  assign n10272 = ~n10249 & n10271;
  assign n10273 = ~n10253 & ~n10271;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = n9506 & ~n10274;
  assign n10276 = n9508 & ~n10267;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = n9501 & ~n10274;
  assign n10279 = n9495 & ~n10274;
  assign n10280 = n9497 & ~n10267;
  assign n10281 = n9504 & ~n10267;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = ~n10278 & ~n10279;
  assign n10284 = n10282 & n10283;
  assign n10285 = ~n10268 & ~n10269;
  assign n10286 = n10277 & n10285;
  assign n10287 = n10284 & n10286;
  assign n10288 = n10259 & n10287;
  assign n10289 = n9436 & ~n10288;
  assign n10290 = P2_REG0_REG_11_ & ~n9436;
  assign n1710 = n10289 | n10290;
  assign n10292 = P2_REG3_REG_12_ & n10217;
  assign n10293 = ~P2_REG3_REG_13_ & n10292;
  assign n10294 = P2_REG3_REG_13_ & ~n10292;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = n9465 & ~n10295;
  assign n10297 = P2_REG0_REG_13_ & n9467;
  assign n10298 = P2_REG1_REG_13_ & n9469;
  assign n10299 = P2_REG2_REG_13_ & n9471;
  assign n10300 = ~n10296 & ~n10297;
  assign n10301 = ~n10298 & n10300;
  assign n10302 = ~n10299 & n10301;
  assign n10303 = n9458 & ~n10302;
  assign n10304 = P2_IR_REG_31_ & n8998;
  assign n10305 = P2_IR_REG_12_ & ~P2_IR_REG_31_;
  assign n10306 = ~n10304 & ~n10305;
  assign n10307 = n9446 & ~n10306;
  assign n10308 = ~n9003 & ~n9446;
  assign n10309 = ~n10307 & ~n10308;
  assign n10310 = ~n10236 & ~n10309;
  assign n10311 = n10236 & n10309;
  assign n10312 = ~n10310 & ~n10311;
  assign n10313 = n9490 & n10312;
  assign n10314 = ~n9455 & ~n10309;
  assign n10315 = n10227 & ~n10309;
  assign n10316 = ~n10227 & n10309;
  assign n10317 = ~n10315 & ~n10316;
  assign n10318 = ~n10246 & ~n10251;
  assign n10319 = ~n10252 & ~n10318;
  assign n10320 = ~n10317 & n10319;
  assign n10321 = n10227 & n10309;
  assign n10322 = ~n10227 & ~n10309;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n10319 & ~n10323;
  assign n10325 = ~n10320 & ~n10324;
  assign n10326 = n9488 & ~n10325;
  assign n10327 = ~n10303 & ~n10313;
  assign n10328 = ~n10314 & n10327;
  assign n10329 = ~n10326 & n10328;
  assign n10330 = n10098 & ~n10176;
  assign n10331 = n10263 & ~n10330;
  assign n10332 = ~n10247 & ~n10331;
  assign n10333 = ~n10097 & ~n10247;
  assign n10334 = ~n10176 & n10333;
  assign n10335 = ~n10118 & n10334;
  assign n10336 = ~n10332 & ~n10335;
  assign n10337 = ~n10317 & ~n10336;
  assign n10338 = n10317 & n10336;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = n9511 & ~n10339;
  assign n10341 = n9561 & ~n10156;
  assign n10342 = ~n10251 & ~n10271;
  assign n10343 = ~n10252 & ~n10342;
  assign n10344 = ~n10317 & n10343;
  assign n10345 = ~n10323 & ~n10343;
  assign n10346 = ~n10344 & ~n10345;
  assign n10347 = n9506 & ~n10346;
  assign n10348 = n9508 & ~n10339;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = n9501 & ~n10346;
  assign n10351 = n9495 & ~n10346;
  assign n10352 = n9497 & ~n10339;
  assign n10353 = n9504 & ~n10339;
  assign n10354 = ~n10352 & ~n10353;
  assign n10355 = ~n10350 & ~n10351;
  assign n10356 = n10354 & n10355;
  assign n10357 = ~n10340 & ~n10341;
  assign n10358 = n10349 & n10357;
  assign n10359 = n10356 & n10358;
  assign n10360 = n10329 & n10359;
  assign n10361 = n9436 & ~n10360;
  assign n10362 = P2_REG0_REG_12_ & ~n9436;
  assign n1715 = n10361 | n10362;
  assign n10364 = P2_REG3_REG_13_ & n10292;
  assign n10365 = ~P2_REG3_REG_14_ & n10364;
  assign n10366 = P2_REG3_REG_14_ & ~n10364;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = n9465 & ~n10367;
  assign n10369 = P2_REG0_REG_14_ & n9467;
  assign n10370 = P2_REG1_REG_14_ & n9469;
  assign n10371 = P2_REG2_REG_14_ & n9471;
  assign n10372 = ~n10368 & ~n10369;
  assign n10373 = ~n10370 & n10372;
  assign n10374 = ~n10371 & n10373;
  assign n10375 = n9458 & ~n10374;
  assign n10376 = P2_IR_REG_31_ & n9009;
  assign n10377 = P2_IR_REG_13_ & ~P2_IR_REG_31_;
  assign n10378 = ~n10376 & ~n10377;
  assign n10379 = n9446 & ~n10378;
  assign n10380 = ~n9014 & ~n9446;
  assign n10381 = ~n10379 & ~n10380;
  assign n10382 = n10311 & n10381;
  assign n10383 = ~n10311 & ~n10381;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = n9490 & n10384;
  assign n10386 = ~n9455 & ~n10381;
  assign n10387 = ~n10302 & ~n10381;
  assign n10388 = n10302 & n10381;
  assign n10389 = ~n10321 & ~n10388;
  assign n10390 = ~n10387 & n10389;
  assign n10391 = n10319 & ~n10322;
  assign n10392 = n10390 & ~n10391;
  assign n10393 = n10302 & ~n10381;
  assign n10394 = ~n10302 & n10381;
  assign n10395 = ~n10393 & ~n10394;
  assign n10396 = ~n10322 & n10395;
  assign n10397 = ~n10319 & ~n10321;
  assign n10398 = n10396 & ~n10397;
  assign n10399 = ~n10392 & ~n10398;
  assign n10400 = n9488 & n10399;
  assign n10401 = ~n10375 & ~n10385;
  assign n10402 = ~n10386 & n10401;
  assign n10403 = ~n10400 & n10402;
  assign n10404 = ~n10315 & ~n10336;
  assign n10405 = ~n10316 & ~n10404;
  assign n10406 = ~n10395 & ~n10405;
  assign n10407 = n10395 & n10405;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = n9511 & ~n10408;
  assign n10410 = n9561 & ~n10227;
  assign n10411 = ~n10322 & n10343;
  assign n10412 = n10390 & ~n10411;
  assign n10413 = ~n10321 & ~n10343;
  assign n10414 = n10396 & ~n10413;
  assign n10415 = ~n10412 & ~n10414;
  assign n10416 = n9506 & n10415;
  assign n10417 = n9508 & ~n10408;
  assign n10418 = ~n10416 & ~n10417;
  assign n10419 = n9501 & n10415;
  assign n10420 = n9495 & n10415;
  assign n10421 = n9497 & ~n10408;
  assign n10422 = n9504 & ~n10408;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = ~n10419 & ~n10420;
  assign n10425 = n10423 & n10424;
  assign n10426 = ~n10409 & ~n10410;
  assign n10427 = n10418 & n10426;
  assign n10428 = n10425 & n10427;
  assign n10429 = n10403 & n10428;
  assign n10430 = n9436 & ~n10429;
  assign n10431 = P2_REG0_REG_13_ & ~n9436;
  assign n1720 = n10430 | n10431;
  assign n10433 = P2_REG3_REG_14_ & n10364;
  assign n10434 = ~P2_REG3_REG_15_ & n10433;
  assign n10435 = P2_REG3_REG_15_ & ~n10433;
  assign n10436 = ~n10434 & ~n10435;
  assign n10437 = n9465 & ~n10436;
  assign n10438 = P2_REG0_REG_15_ & n9467;
  assign n10439 = P2_REG1_REG_15_ & n9469;
  assign n10440 = P2_REG2_REG_15_ & n9471;
  assign n10441 = ~n10437 & ~n10438;
  assign n10442 = ~n10439 & n10441;
  assign n10443 = ~n10440 & n10442;
  assign n10444 = n9458 & ~n10443;
  assign n10445 = P2_IR_REG_31_ & n9021;
  assign n10446 = P2_IR_REG_14_ & ~P2_IR_REG_31_;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = n9446 & ~n10447;
  assign n10449 = ~n9026 & ~n9446;
  assign n10450 = ~n10448 & ~n10449;
  assign n10451 = ~n10382 & ~n10450;
  assign n10452 = n10381 & n10450;
  assign n10453 = n10311 & n10452;
  assign n10454 = ~n10451 & ~n10453;
  assign n10455 = n9490 & n10454;
  assign n10456 = ~n9455 & ~n10450;
  assign n10457 = ~n10322 & ~n10387;
  assign n10458 = n10252 & n10389;
  assign n10459 = n10457 & ~n10458;
  assign n10460 = ~n10388 & ~n10459;
  assign n10461 = ~n10251 & n10389;
  assign n10462 = ~n10246 & n10461;
  assign n10463 = ~n10460 & ~n10462;
  assign n10464 = n10374 & ~n10450;
  assign n10465 = ~n10374 & n10450;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = n10463 & ~n10466;
  assign n10468 = ~n10463 & n10466;
  assign n10469 = ~n10467 & ~n10468;
  assign n10470 = n9488 & ~n10469;
  assign n10471 = ~n10444 & ~n10455;
  assign n10472 = ~n10456 & n10471;
  assign n10473 = ~n10470 & n10472;
  assign n10474 = ~n10393 & ~n10405;
  assign n10475 = ~n10394 & ~n10474;
  assign n10476 = n10466 & n10475;
  assign n10477 = ~n10466 & ~n10475;
  assign n10478 = ~n10476 & ~n10477;
  assign n10479 = n9511 & ~n10478;
  assign n10480 = n9561 & ~n10302;
  assign n10481 = ~n10271 & n10461;
  assign n10482 = ~n10460 & ~n10481;
  assign n10483 = ~n10466 & n10482;
  assign n10484 = n10466 & ~n10482;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = n9506 & ~n10485;
  assign n10487 = n9508 & ~n10478;
  assign n10488 = ~n10486 & ~n10487;
  assign n10489 = n9501 & ~n10485;
  assign n10490 = n9495 & ~n10485;
  assign n10491 = n9497 & ~n10478;
  assign n10492 = n9504 & ~n10478;
  assign n10493 = ~n10491 & ~n10492;
  assign n10494 = ~n10489 & ~n10490;
  assign n10495 = n10493 & n10494;
  assign n10496 = ~n10479 & ~n10480;
  assign n10497 = n10488 & n10496;
  assign n10498 = n10495 & n10497;
  assign n10499 = n10473 & n10498;
  assign n10500 = n9436 & ~n10499;
  assign n10501 = P2_REG0_REG_14_ & ~n9436;
  assign n1725 = n10500 | n10501;
  assign n10503 = P2_REG3_REG_15_ & n10433;
  assign n10504 = ~P2_REG3_REG_16_ & n10503;
  assign n10505 = P2_REG3_REG_16_ & ~n10503;
  assign n10506 = ~n10504 & ~n10505;
  assign n10507 = n9465 & ~n10506;
  assign n10508 = P2_REG0_REG_16_ & n9467;
  assign n10509 = P2_REG1_REG_16_ & n9469;
  assign n10510 = P2_REG2_REG_16_ & n9471;
  assign n10511 = ~n10507 & ~n10508;
  assign n10512 = ~n10509 & n10511;
  assign n10513 = ~n10510 & n10512;
  assign n10514 = n9458 & ~n10513;
  assign n10515 = P2_IR_REG_31_ & n9032;
  assign n10516 = P2_IR_REG_15_ & ~P2_IR_REG_31_;
  assign n10517 = ~n10515 & ~n10516;
  assign n10518 = n9446 & ~n10517;
  assign n10519 = ~n9037 & ~n9446;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = ~n10453 & ~n10520;
  assign n10522 = n10453 & n10520;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = n9490 & n10523;
  assign n10525 = ~n9455 & ~n10520;
  assign n10526 = ~n10374 & ~n10450;
  assign n10527 = n10374 & n10450;
  assign n10528 = ~n10463 & ~n10527;
  assign n10529 = ~n10526 & ~n10528;
  assign n10530 = n10443 & ~n10520;
  assign n10531 = ~n10443 & n10520;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = n10529 & ~n10532;
  assign n10534 = ~n10529 & n10532;
  assign n10535 = ~n10533 & ~n10534;
  assign n10536 = n9488 & ~n10535;
  assign n10537 = ~n10514 & ~n10524;
  assign n10538 = ~n10525 & n10537;
  assign n10539 = ~n10536 & n10538;
  assign n10540 = ~n10464 & ~n10475;
  assign n10541 = ~n10465 & ~n10540;
  assign n10542 = n10532 & n10541;
  assign n10543 = ~n10532 & ~n10541;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = n9511 & ~n10544;
  assign n10546 = n9561 & ~n10374;
  assign n10547 = ~n10482 & ~n10527;
  assign n10548 = ~n10526 & ~n10547;
  assign n10549 = ~n10532 & n10548;
  assign n10550 = n10532 & ~n10548;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = n9506 & ~n10551;
  assign n10553 = n9508 & ~n10544;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = n9501 & ~n10551;
  assign n10556 = n9495 & ~n10551;
  assign n10557 = n9497 & ~n10544;
  assign n10558 = n9504 & ~n10544;
  assign n10559 = ~n10557 & ~n10558;
  assign n10560 = ~n10555 & ~n10556;
  assign n10561 = n10559 & n10560;
  assign n10562 = ~n10545 & ~n10546;
  assign n10563 = n10554 & n10562;
  assign n10564 = n10561 & n10563;
  assign n10565 = n10539 & n10564;
  assign n10566 = n9436 & ~n10565;
  assign n10567 = P2_REG0_REG_15_ & ~n9436;
  assign n1730 = n10566 | n10567;
  assign n10569 = P2_REG1_REG_17_ & n9469;
  assign n10570 = P2_REG0_REG_17_ & n9467;
  assign n10571 = P2_REG2_REG_17_ & n9471;
  assign n10572 = P2_REG3_REG_16_ & n10503;
  assign n10573 = ~P2_REG3_REG_17_ & n10572;
  assign n10574 = P2_REG3_REG_17_ & ~n10572;
  assign n10575 = ~n10573 & ~n10574;
  assign n10576 = n9465 & ~n10575;
  assign n10577 = ~n10569 & ~n10570;
  assign n10578 = ~n10571 & n10577;
  assign n10579 = ~n10576 & n10578;
  assign n10580 = n9458 & ~n10579;
  assign n10581 = P2_IR_REG_31_ & n9057;
  assign n10582 = P2_IR_REG_16_ & ~P2_IR_REG_31_;
  assign n10583 = ~n10581 & ~n10582;
  assign n10584 = n9446 & ~n10583;
  assign n10585 = ~n9062 & ~n9446;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = ~n10522 & ~n10586;
  assign n10588 = n10522 & n10586;
  assign n10589 = ~n10587 & ~n10588;
  assign n10590 = n9490 & n10589;
  assign n10591 = ~n9455 & ~n10586;
  assign n10592 = n10513 & ~n10586;
  assign n10593 = ~n10513 & n10586;
  assign n10594 = ~n10592 & ~n10593;
  assign n10595 = ~n10443 & ~n10520;
  assign n10596 = n10443 & n10520;
  assign n10597 = ~n10529 & ~n10596;
  assign n10598 = ~n10595 & ~n10597;
  assign n10599 = ~n10594 & n10598;
  assign n10600 = n10513 & n10586;
  assign n10601 = ~n10513 & ~n10586;
  assign n10602 = ~n10600 & ~n10601;
  assign n10603 = ~n10598 & ~n10602;
  assign n10604 = ~n10599 & ~n10603;
  assign n10605 = n9488 & ~n10604;
  assign n10606 = ~n10580 & ~n10590;
  assign n10607 = ~n10591 & n10606;
  assign n10608 = ~n10605 & n10607;
  assign n10609 = ~n10530 & ~n10594;
  assign n10610 = ~n10531 & n10541;
  assign n10611 = n10609 & ~n10610;
  assign n10612 = ~n10531 & ~n10593;
  assign n10613 = ~n10592 & n10612;
  assign n10614 = ~n10530 & ~n10541;
  assign n10615 = n10613 & ~n10614;
  assign n10616 = ~n10611 & ~n10615;
  assign n10617 = n9511 & ~n10616;
  assign n10618 = n9561 & ~n10443;
  assign n10619 = ~n10548 & ~n10596;
  assign n10620 = ~n10595 & ~n10619;
  assign n10621 = ~n10594 & n10620;
  assign n10622 = ~n10602 & ~n10620;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = n9506 & ~n10623;
  assign n10625 = n9508 & ~n10616;
  assign n10626 = ~n10624 & ~n10625;
  assign n10627 = n9501 & ~n10623;
  assign n10628 = n9495 & ~n10623;
  assign n10629 = n9497 & ~n10616;
  assign n10630 = n9504 & ~n10616;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = ~n10627 & ~n10628;
  assign n10633 = n10631 & n10632;
  assign n10634 = ~n10617 & ~n10618;
  assign n10635 = n10626 & n10634;
  assign n10636 = n10633 & n10635;
  assign n10637 = n10608 & n10636;
  assign n10638 = n9436 & ~n10637;
  assign n10639 = P2_REG0_REG_16_ & ~n9436;
  assign n1735 = n10638 | n10639;
  assign n10641 = P2_REG1_REG_18_ & n9469;
  assign n10642 = P2_REG0_REG_18_ & n9467;
  assign n10643 = P2_REG2_REG_18_ & n9471;
  assign n10644 = P2_REG3_REG_17_ & n10572;
  assign n10645 = ~P2_REG3_REG_18_ & n10644;
  assign n10646 = P2_REG3_REG_18_ & ~n10644;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = n9465 & ~n10647;
  assign n10649 = ~n10641 & ~n10642;
  assign n10650 = ~n10643 & n10649;
  assign n10651 = ~n10648 & n10650;
  assign n10652 = n9458 & ~n10651;
  assign n10653 = P2_IR_REG_31_ & n9068;
  assign n10654 = P2_IR_REG_17_ & ~P2_IR_REG_31_;
  assign n10655 = ~n10653 & ~n10654;
  assign n10656 = n9446 & ~n10655;
  assign n10657 = ~n9073 & ~n9446;
  assign n10658 = ~n10656 & ~n10657;
  assign n10659 = n10588 & n10658;
  assign n10660 = ~n10588 & ~n10658;
  assign n10661 = ~n10659 & ~n10660;
  assign n10662 = n9490 & n10661;
  assign n10663 = ~n9455 & ~n10658;
  assign n10664 = ~n10579 & ~n10658;
  assign n10665 = n10579 & n10658;
  assign n10666 = ~n10600 & ~n10665;
  assign n10667 = ~n10664 & n10666;
  assign n10668 = n10598 & ~n10601;
  assign n10669 = n10667 & ~n10668;
  assign n10670 = n10579 & ~n10658;
  assign n10671 = ~n10579 & n10658;
  assign n10672 = ~n10670 & ~n10671;
  assign n10673 = ~n10601 & n10672;
  assign n10674 = ~n10598 & ~n10600;
  assign n10675 = n10673 & ~n10674;
  assign n10676 = ~n10669 & ~n10675;
  assign n10677 = n9488 & n10676;
  assign n10678 = ~n10652 & ~n10662;
  assign n10679 = ~n10663 & n10678;
  assign n10680 = ~n10677 & n10679;
  assign n10681 = ~n10530 & ~n10592;
  assign n10682 = n10465 & n10681;
  assign n10683 = n10612 & ~n10682;
  assign n10684 = ~n10592 & ~n10683;
  assign n10685 = ~n10464 & n10681;
  assign n10686 = ~n10475 & n10685;
  assign n10687 = ~n10684 & ~n10686;
  assign n10688 = ~n10672 & ~n10687;
  assign n10689 = n10672 & n10687;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = n9511 & ~n10690;
  assign n10692 = n9561 & ~n10513;
  assign n10693 = ~n10601 & n10620;
  assign n10694 = n10667 & ~n10693;
  assign n10695 = ~n10600 & ~n10620;
  assign n10696 = n10673 & ~n10695;
  assign n10697 = ~n10694 & ~n10696;
  assign n10698 = n9506 & n10697;
  assign n10699 = n9508 & ~n10690;
  assign n10700 = ~n10698 & ~n10699;
  assign n10701 = n9501 & n10697;
  assign n10702 = n9495 & n10697;
  assign n10703 = n9497 & ~n10690;
  assign n10704 = n9504 & ~n10690;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n10701 & ~n10702;
  assign n10707 = n10705 & n10706;
  assign n10708 = ~n10691 & ~n10692;
  assign n10709 = n10700 & n10708;
  assign n10710 = n10707 & n10709;
  assign n10711 = n10680 & n10710;
  assign n10712 = n9436 & ~n10711;
  assign n10713 = P2_REG0_REG_17_ & ~n9436;
  assign n1740 = n10712 | n10713;
  assign n10715 = P2_REG1_REG_19_ & n9469;
  assign n10716 = P2_REG0_REG_19_ & n9467;
  assign n10717 = P2_REG2_REG_19_ & n9471;
  assign n10718 = P2_REG3_REG_18_ & n10644;
  assign n10719 = ~P2_REG3_REG_19_ & n10718;
  assign n10720 = P2_REG3_REG_19_ & ~n10718;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = n9465 & ~n10721;
  assign n10723 = ~n10715 & ~n10716;
  assign n10724 = ~n10717 & n10723;
  assign n10725 = ~n10722 & n10724;
  assign n10726 = n9458 & ~n10725;
  assign n10727 = P2_IR_REG_31_ & n9080;
  assign n10728 = P2_IR_REG_18_ & ~P2_IR_REG_31_;
  assign n10729 = ~n10727 & ~n10728;
  assign n10730 = n9446 & ~n10729;
  assign n10731 = ~n9085 & ~n9446;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 = ~n10659 & ~n10732;
  assign n10734 = n10658 & n10732;
  assign n10735 = n10588 & n10734;
  assign n10736 = ~n10733 & ~n10735;
  assign n10737 = n9490 & n10736;
  assign n10738 = ~n9455 & ~n10732;
  assign n10739 = n10601 & ~n10658;
  assign n10740 = ~n10601 & n10658;
  assign n10741 = ~n10579 & ~n10740;
  assign n10742 = ~n10739 & ~n10741;
  assign n10743 = ~n10598 & n10666;
  assign n10744 = n10742 & ~n10743;
  assign n10745 = n10651 & ~n10732;
  assign n10746 = ~n10651 & n10732;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = n10744 & ~n10747;
  assign n10749 = n10651 & n10732;
  assign n10750 = ~n10651 & ~n10732;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = ~n10744 & ~n10751;
  assign n10753 = ~n10748 & ~n10752;
  assign n10754 = n9488 & ~n10753;
  assign n10755 = ~n10726 & ~n10737;
  assign n10756 = ~n10738 & n10755;
  assign n10757 = ~n10754 & n10756;
  assign n10758 = ~n10670 & ~n10687;
  assign n10759 = ~n10671 & ~n10758;
  assign n10760 = ~n10747 & ~n10759;
  assign n10761 = n10747 & n10759;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = n9511 & ~n10762;
  assign n10764 = n9561 & ~n10579;
  assign n10765 = ~n10620 & n10666;
  assign n10766 = n10742 & ~n10765;
  assign n10767 = ~n10747 & n10766;
  assign n10768 = ~n10751 & ~n10766;
  assign n10769 = ~n10767 & ~n10768;
  assign n10770 = n9506 & ~n10769;
  assign n10771 = n9508 & ~n10762;
  assign n10772 = ~n10770 & ~n10771;
  assign n10773 = n9501 & ~n10769;
  assign n10774 = n9495 & ~n10769;
  assign n10775 = n9497 & ~n10762;
  assign n10776 = n9504 & ~n10762;
  assign n10777 = ~n10775 & ~n10776;
  assign n10778 = ~n10773 & ~n10774;
  assign n10779 = n10777 & n10778;
  assign n10780 = ~n10763 & ~n10764;
  assign n10781 = n10772 & n10780;
  assign n10782 = n10779 & n10781;
  assign n10783 = n10757 & n10782;
  assign n10784 = n9436 & ~n10783;
  assign n10785 = P2_REG0_REG_18_ & ~n9436;
  assign n1745 = n10784 | n10785;
  assign n10787 = P2_REG1_REG_20_ & n9469;
  assign n10788 = P2_REG0_REG_20_ & n9467;
  assign n10789 = P2_REG2_REG_20_ & n9471;
  assign n10790 = P2_REG3_REG_19_ & n10718;
  assign n10791 = ~P2_REG3_REG_20_ & n10790;
  assign n10792 = P2_REG3_REG_20_ & ~n10790;
  assign n10793 = ~n10791 & ~n10792;
  assign n10794 = n9465 & ~n10793;
  assign n10795 = ~n10787 & ~n10788;
  assign n10796 = ~n10789 & n10795;
  assign n10797 = ~n10794 & n10796;
  assign n10798 = n9458 & ~n10797;
  assign n10799 = ~n9371 & n9446;
  assign n10800 = ~n9096 & ~n9446;
  assign n10801 = ~n10799 & ~n10800;
  assign n10802 = n10735 & n10801;
  assign n10803 = ~n10735 & ~n10801;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = n9490 & n10804;
  assign n10806 = ~n9455 & ~n10801;
  assign n10807 = n10725 & ~n10801;
  assign n10808 = ~n10725 & n10801;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = ~n10744 & ~n10749;
  assign n10811 = ~n10750 & ~n10810;
  assign n10812 = ~n10809 & n10811;
  assign n10813 = n10725 & n10801;
  assign n10814 = ~n10725 & ~n10801;
  assign n10815 = ~n10813 & ~n10814;
  assign n10816 = ~n10811 & ~n10815;
  assign n10817 = ~n10812 & ~n10816;
  assign n10818 = n9488 & ~n10817;
  assign n10819 = ~n10798 & ~n10805;
  assign n10820 = ~n10806 & n10819;
  assign n10821 = ~n10818 & n10820;
  assign n10822 = ~n10651 & ~n10759;
  assign n10823 = n10651 & n10759;
  assign n10824 = n10732 & ~n10823;
  assign n10825 = ~n10822 & ~n10824;
  assign n10826 = ~n10809 & ~n10825;
  assign n10827 = n10809 & n10825;
  assign n10828 = ~n10826 & ~n10827;
  assign n10829 = n9511 & ~n10828;
  assign n10830 = n9561 & ~n10651;
  assign n10831 = ~n10749 & ~n10766;
  assign n10832 = ~n10750 & ~n10831;
  assign n10833 = ~n10809 & n10832;
  assign n10834 = ~n10815 & ~n10832;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = n9506 & ~n10835;
  assign n10837 = n9508 & ~n10828;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = n9501 & ~n10835;
  assign n10840 = n9495 & ~n10835;
  assign n10841 = n9497 & ~n10828;
  assign n10842 = n9504 & ~n10828;
  assign n10843 = ~n10841 & ~n10842;
  assign n10844 = ~n10839 & ~n10840;
  assign n10845 = n10843 & n10844;
  assign n10846 = ~n10829 & ~n10830;
  assign n10847 = n10838 & n10846;
  assign n10848 = n10845 & n10847;
  assign n10849 = n10821 & n10848;
  assign n10850 = n9436 & ~n10849;
  assign n10851 = P2_REG0_REG_19_ & ~n9436;
  assign n1750 = n10850 | n10851;
  assign n10853 = P2_REG1_REG_21_ & n9469;
  assign n10854 = P2_REG0_REG_21_ & n9467;
  assign n10855 = P2_REG2_REG_21_ & n9471;
  assign n10856 = P2_REG3_REG_20_ & n10790;
  assign n10857 = ~P2_REG3_REG_21_ & n10856;
  assign n10858 = P2_REG3_REG_21_ & ~n10856;
  assign n10859 = ~n10857 & ~n10858;
  assign n10860 = n9465 & ~n10859;
  assign n10861 = ~n10853 & ~n10854;
  assign n10862 = ~n10855 & n10861;
  assign n10863 = ~n10860 & n10862;
  assign n10864 = n9458 & ~n10863;
  assign n10865 = ~n9107 & ~n9446;
  assign n10866 = ~n10802 & n10865;
  assign n10867 = n10801 & ~n10865;
  assign n10868 = n10735 & n10867;
  assign n10869 = ~n10866 & ~n10868;
  assign n10870 = n9490 & n10869;
  assign n10871 = ~n9455 & n10865;
  assign n10872 = ~n10797 & n10865;
  assign n10873 = n10797 & ~n10865;
  assign n10874 = ~n10813 & ~n10873;
  assign n10875 = ~n10872 & n10874;
  assign n10876 = n10811 & ~n10814;
  assign n10877 = n10875 & ~n10876;
  assign n10878 = n10797 & n10865;
  assign n10879 = ~n10797 & ~n10865;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = ~n10814 & n10880;
  assign n10882 = ~n10811 & ~n10813;
  assign n10883 = n10881 & ~n10882;
  assign n10884 = ~n10877 & ~n10883;
  assign n10885 = n9488 & n10884;
  assign n10886 = ~n10864 & ~n10870;
  assign n10887 = ~n10871 & n10886;
  assign n10888 = ~n10885 & n10887;
  assign n10889 = ~n10807 & ~n10825;
  assign n10890 = ~n10808 & ~n10889;
  assign n10891 = ~n10880 & ~n10890;
  assign n10892 = n10880 & n10890;
  assign n10893 = ~n10891 & ~n10892;
  assign n10894 = n9511 & ~n10893;
  assign n10895 = n9561 & ~n10725;
  assign n10896 = ~n10814 & n10832;
  assign n10897 = n10875 & ~n10896;
  assign n10898 = ~n10813 & ~n10832;
  assign n10899 = n10881 & ~n10898;
  assign n10900 = ~n10897 & ~n10899;
  assign n10901 = n9506 & n10900;
  assign n10902 = n9508 & ~n10893;
  assign n10903 = ~n10901 & ~n10902;
  assign n10904 = n9501 & n10900;
  assign n10905 = n9495 & n10900;
  assign n10906 = n9497 & ~n10893;
  assign n10907 = n9504 & ~n10893;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = ~n10904 & ~n10905;
  assign n10910 = n10908 & n10909;
  assign n10911 = ~n10894 & ~n10895;
  assign n10912 = n10903 & n10911;
  assign n10913 = n10910 & n10912;
  assign n10914 = n10888 & n10913;
  assign n10915 = n9436 & ~n10914;
  assign n10916 = P2_REG0_REG_20_ & ~n9436;
  assign n1755 = n10915 | n10916;
  assign n10918 = P2_REG1_REG_22_ & n9469;
  assign n10919 = P2_REG0_REG_22_ & n9467;
  assign n10920 = P2_REG2_REG_22_ & n9471;
  assign n10921 = P2_REG3_REG_21_ & n10856;
  assign n10922 = ~P2_REG3_REG_22_ & n10921;
  assign n10923 = P2_REG3_REG_22_ & ~n10921;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = n9465 & ~n10924;
  assign n10926 = ~n10918 & ~n10919;
  assign n10927 = ~n10920 & n10926;
  assign n10928 = ~n10925 & n10927;
  assign n10929 = n9458 & ~n10928;
  assign n10930 = ~n9121 & ~n9446;
  assign n10931 = n10868 & ~n10930;
  assign n10932 = ~n10868 & n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = n9490 & n10933;
  assign n10935 = ~n9455 & n10930;
  assign n10936 = n10863 & n10930;
  assign n10937 = ~n10863 & ~n10930;
  assign n10938 = ~n10936 & ~n10937;
  assign n10939 = ~n10811 & n10874;
  assign n10940 = ~n10814 & ~n10865;
  assign n10941 = n10814 & n10865;
  assign n10942 = n10797 & ~n10941;
  assign n10943 = ~n10940 & ~n10942;
  assign n10944 = ~n10939 & ~n10943;
  assign n10945 = ~n10938 & ~n10944;
  assign n10946 = n10938 & ~n10943;
  assign n10947 = ~n10939 & n10946;
  assign n10948 = ~n10945 & ~n10947;
  assign n10949 = n9488 & n10948;
  assign n10950 = ~n10929 & ~n10934;
  assign n10951 = ~n10935 & n10950;
  assign n10952 = ~n10949 & n10951;
  assign n10953 = ~n10878 & ~n10890;
  assign n10954 = ~n10879 & ~n10953;
  assign n10955 = n10938 & n10954;
  assign n10956 = ~n10938 & ~n10954;
  assign n10957 = ~n10955 & ~n10956;
  assign n10958 = n9511 & ~n10957;
  assign n10959 = n9561 & ~n10797;
  assign n10960 = ~n10832 & n10874;
  assign n10961 = ~n10943 & ~n10960;
  assign n10962 = ~n10938 & ~n10961;
  assign n10963 = n10946 & ~n10960;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = n9506 & n10964;
  assign n10966 = n9508 & ~n10957;
  assign n10967 = ~n10965 & ~n10966;
  assign n10968 = n9501 & n10964;
  assign n10969 = n9495 & n10964;
  assign n10970 = n9497 & ~n10957;
  assign n10971 = n9504 & ~n10957;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = ~n10968 & ~n10969;
  assign n10974 = n10972 & n10973;
  assign n10975 = ~n10958 & ~n10959;
  assign n10976 = n10967 & n10975;
  assign n10977 = n10974 & n10976;
  assign n10978 = n10952 & n10977;
  assign n10979 = n9436 & ~n10978;
  assign n10980 = P2_REG0_REG_21_ & ~n9436;
  assign n1760 = n10979 | n10980;
  assign n10982 = P2_REG1_REG_23_ & n9469;
  assign n10983 = P2_REG0_REG_23_ & n9467;
  assign n10984 = P2_REG2_REG_23_ & n9471;
  assign n10985 = P2_REG3_REG_22_ & n10921;
  assign n10986 = ~P2_REG3_REG_23_ & n10985;
  assign n10987 = P2_REG3_REG_23_ & ~n10985;
  assign n10988 = ~n10986 & ~n10987;
  assign n10989 = n9465 & ~n10988;
  assign n10990 = ~n10982 & ~n10983;
  assign n10991 = ~n10984 & n10990;
  assign n10992 = ~n10989 & n10991;
  assign n10993 = n9458 & ~n10992;
  assign n10994 = ~n9132 & ~n9446;
  assign n10995 = ~n10931 & n10994;
  assign n10996 = ~n10930 & ~n10994;
  assign n10997 = n10868 & n10996;
  assign n10998 = ~n10995 & ~n10997;
  assign n10999 = n9490 & n10998;
  assign n11000 = ~n9455 & n10994;
  assign n11001 = n10863 & ~n10930;
  assign n11002 = n10750 & n10874;
  assign n11003 = ~n10943 & ~n11002;
  assign n11004 = ~n11001 & ~n11003;
  assign n11005 = ~n10863 & n10930;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = ~n10749 & n10874;
  assign n11008 = ~n10744 & ~n11001;
  assign n11009 = n11007 & n11008;
  assign n11010 = n11006 & ~n11009;
  assign n11011 = n10928 & n10994;
  assign n11012 = ~n10928 & ~n10994;
  assign n11013 = ~n11011 & ~n11012;
  assign n11014 = n11010 & ~n11013;
  assign n11015 = ~n11010 & n11013;
  assign n11016 = ~n11014 & ~n11015;
  assign n11017 = n9488 & ~n11016;
  assign n11018 = ~n10993 & ~n10999;
  assign n11019 = ~n11000 & n11018;
  assign n11020 = ~n11017 & n11019;
  assign n11021 = ~n10936 & ~n10954;
  assign n11022 = ~n10937 & ~n11021;
  assign n11023 = n11013 & n11022;
  assign n11024 = ~n11013 & ~n11022;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = n9511 & ~n11025;
  assign n11027 = n9561 & ~n10863;
  assign n11028 = ~n10766 & ~n11001;
  assign n11029 = n11007 & n11028;
  assign n11030 = n11006 & ~n11029;
  assign n11031 = ~n11013 & n11030;
  assign n11032 = n11013 & ~n11030;
  assign n11033 = ~n11031 & ~n11032;
  assign n11034 = n9506 & ~n11033;
  assign n11035 = n9508 & ~n11025;
  assign n11036 = ~n11034 & ~n11035;
  assign n11037 = n9501 & ~n11033;
  assign n11038 = n9495 & ~n11033;
  assign n11039 = n9497 & ~n11025;
  assign n11040 = n9504 & ~n11025;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = ~n11037 & ~n11038;
  assign n11043 = n11041 & n11042;
  assign n11044 = ~n11026 & ~n11027;
  assign n11045 = n11036 & n11044;
  assign n11046 = n11043 & n11045;
  assign n11047 = n11020 & n11046;
  assign n11048 = n9436 & ~n11047;
  assign n11049 = P2_REG0_REG_22_ & ~n9436;
  assign n1765 = n11048 | n11049;
  assign n11051 = P2_REG1_REG_24_ & n9469;
  assign n11052 = P2_REG0_REG_24_ & n9467;
  assign n11053 = P2_REG2_REG_24_ & n9471;
  assign n11054 = P2_REG3_REG_23_ & n10985;
  assign n11055 = ~P2_REG3_REG_24_ & n11054;
  assign n11056 = P2_REG3_REG_24_ & ~n11054;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = n9465 & ~n11057;
  assign n11059 = ~n11051 & ~n11052;
  assign n11060 = ~n11053 & n11059;
  assign n11061 = ~n11058 & n11060;
  assign n11062 = n9458 & ~n11061;
  assign n11063 = ~n9145 & ~n9446;
  assign n11064 = n10997 & ~n11063;
  assign n11065 = ~n10997 & n11063;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = n9490 & n11066;
  assign n11068 = ~n9455 & n11063;
  assign n11069 = ~n10928 & n10994;
  assign n11070 = n10928 & ~n10994;
  assign n11071 = ~n11010 & ~n11070;
  assign n11072 = ~n11069 & ~n11071;
  assign n11073 = n10992 & n11063;
  assign n11074 = ~n10992 & ~n11063;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = n11072 & ~n11075;
  assign n11077 = ~n11072 & n11075;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = n9488 & ~n11078;
  assign n11080 = ~n11062 & ~n11067;
  assign n11081 = ~n11068 & n11080;
  assign n11082 = ~n11079 & n11081;
  assign n11083 = ~n11011 & ~n11075;
  assign n11084 = ~n11012 & n11022;
  assign n11085 = n11083 & ~n11084;
  assign n11086 = ~n11012 & ~n11074;
  assign n11087 = ~n11073 & n11086;
  assign n11088 = ~n11011 & ~n11022;
  assign n11089 = n11087 & ~n11088;
  assign n11090 = ~n11085 & ~n11089;
  assign n11091 = n9511 & ~n11090;
  assign n11092 = n9561 & ~n10928;
  assign n11093 = ~n11030 & ~n11070;
  assign n11094 = ~n11069 & ~n11093;
  assign n11095 = ~n11075 & n11094;
  assign n11096 = n11075 & ~n11094;
  assign n11097 = ~n11095 & ~n11096;
  assign n11098 = n9506 & ~n11097;
  assign n11099 = n9508 & ~n11090;
  assign n11100 = ~n11098 & ~n11099;
  assign n11101 = n9501 & ~n11097;
  assign n11102 = n9495 & ~n11097;
  assign n11103 = n9497 & ~n11090;
  assign n11104 = n9504 & ~n11090;
  assign n11105 = ~n11103 & ~n11104;
  assign n11106 = ~n11101 & ~n11102;
  assign n11107 = n11105 & n11106;
  assign n11108 = ~n11091 & ~n11092;
  assign n11109 = n11100 & n11108;
  assign n11110 = n11107 & n11109;
  assign n11111 = n11082 & n11110;
  assign n11112 = n9436 & ~n11111;
  assign n11113 = P2_REG0_REG_23_ & ~n9436;
  assign n1770 = n11112 | n11113;
  assign n11115 = P2_REG1_REG_25_ & n9469;
  assign n11116 = P2_REG0_REG_25_ & n9467;
  assign n11117 = P2_REG2_REG_25_ & n9471;
  assign n11118 = P2_REG3_REG_24_ & n11054;
  assign n11119 = ~P2_REG3_REG_25_ & n11118;
  assign n11120 = P2_REG3_REG_25_ & ~n11118;
  assign n11121 = ~n11119 & ~n11120;
  assign n11122 = n9465 & ~n11121;
  assign n11123 = ~n11115 & ~n11116;
  assign n11124 = ~n11117 & n11123;
  assign n11125 = ~n11122 & n11124;
  assign n11126 = n9458 & ~n11125;
  assign n11127 = ~n9156 & ~n9446;
  assign n11128 = ~n11064 & n11127;
  assign n11129 = n11064 & ~n11127;
  assign n11130 = ~n11128 & ~n11129;
  assign n11131 = n9490 & n11130;
  assign n11132 = ~n9455 & n11127;
  assign n11133 = ~n10992 & n11063;
  assign n11134 = n10992 & ~n11063;
  assign n11135 = ~n11072 & ~n11134;
  assign n11136 = ~n11133 & ~n11135;
  assign n11137 = n11061 & n11127;
  assign n11138 = ~n11061 & ~n11127;
  assign n11139 = ~n11137 & ~n11138;
  assign n11140 = n11136 & ~n11139;
  assign n11141 = n11061 & ~n11127;
  assign n11142 = ~n11061 & n11127;
  assign n11143 = ~n11141 & ~n11142;
  assign n11144 = ~n11136 & ~n11143;
  assign n11145 = ~n11140 & ~n11144;
  assign n11146 = n9488 & ~n11145;
  assign n11147 = ~n11126 & ~n11131;
  assign n11148 = ~n11132 & n11147;
  assign n11149 = ~n11146 & n11148;
  assign n11150 = ~n11011 & ~n11073;
  assign n11151 = n10937 & n11150;
  assign n11152 = n11086 & ~n11151;
  assign n11153 = ~n11073 & ~n11152;
  assign n11154 = ~n10936 & n11150;
  assign n11155 = ~n10954 & n11154;
  assign n11156 = ~n11153 & ~n11155;
  assign n11157 = ~n11139 & ~n11156;
  assign n11158 = n11139 & n11156;
  assign n11159 = ~n11157 & ~n11158;
  assign n11160 = n9511 & ~n11159;
  assign n11161 = n9561 & ~n10992;
  assign n11162 = ~n11094 & ~n11134;
  assign n11163 = ~n11133 & ~n11162;
  assign n11164 = ~n11139 & n11163;
  assign n11165 = ~n11143 & ~n11163;
  assign n11166 = ~n11164 & ~n11165;
  assign n11167 = n9506 & ~n11166;
  assign n11168 = n9508 & ~n11159;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = n9501 & ~n11166;
  assign n11171 = n9495 & ~n11166;
  assign n11172 = n9497 & ~n11159;
  assign n11173 = n9504 & ~n11159;
  assign n11174 = ~n11172 & ~n11173;
  assign n11175 = ~n11170 & ~n11171;
  assign n11176 = n11174 & n11175;
  assign n11177 = ~n11160 & ~n11161;
  assign n11178 = n11169 & n11177;
  assign n11179 = n11176 & n11178;
  assign n11180 = n11149 & n11179;
  assign n11181 = n9436 & ~n11180;
  assign n11182 = P2_REG0_REG_24_ & ~n9436;
  assign n1775 = n11181 | n11182;
  assign n11184 = P2_REG1_REG_26_ & n9469;
  assign n11185 = P2_REG0_REG_26_ & n9467;
  assign n11186 = P2_REG2_REG_26_ & n9471;
  assign n11187 = P2_REG3_REG_25_ & n11118;
  assign n11188 = ~P2_REG3_REG_26_ & n11187;
  assign n11189 = P2_REG3_REG_26_ & ~n11187;
  assign n11190 = ~n11188 & ~n11189;
  assign n11191 = n9465 & ~n11190;
  assign n11192 = ~n11184 & ~n11185;
  assign n11193 = ~n11186 & n11192;
  assign n11194 = ~n11191 & n11193;
  assign n11195 = n9458 & ~n11194;
  assign n11196 = ~n9167 & ~n9446;
  assign n11197 = n11129 & ~n11196;
  assign n11198 = ~n11129 & n11196;
  assign n11199 = ~n11197 & ~n11198;
  assign n11200 = n9490 & n11199;
  assign n11201 = ~n9455 & n11196;
  assign n11202 = n11125 & n11196;
  assign n11203 = ~n11125 & ~n11196;
  assign n11204 = ~n11202 & ~n11203;
  assign n11205 = ~n11136 & ~n11141;
  assign n11206 = ~n11142 & ~n11205;
  assign n11207 = ~n11204 & n11206;
  assign n11208 = n11125 & ~n11196;
  assign n11209 = ~n11125 & n11196;
  assign n11210 = ~n11208 & ~n11209;
  assign n11211 = ~n11206 & ~n11210;
  assign n11212 = ~n11207 & ~n11211;
  assign n11213 = n9488 & ~n11212;
  assign n11214 = ~n11195 & ~n11200;
  assign n11215 = ~n11201 & n11214;
  assign n11216 = ~n11213 & n11215;
  assign n11217 = ~n11137 & ~n11156;
  assign n11218 = ~n11138 & ~n11217;
  assign n11219 = ~n11204 & ~n11218;
  assign n11220 = n11204 & n11218;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = n9511 & ~n11221;
  assign n11223 = n9561 & ~n11061;
  assign n11224 = ~n11141 & ~n11163;
  assign n11225 = ~n11142 & ~n11224;
  assign n11226 = ~n11204 & n11225;
  assign n11227 = ~n11210 & ~n11225;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = n9506 & ~n11228;
  assign n11230 = n9508 & ~n11221;
  assign n11231 = ~n11229 & ~n11230;
  assign n11232 = n9501 & ~n11228;
  assign n11233 = n9495 & ~n11228;
  assign n11234 = n9497 & ~n11221;
  assign n11235 = n9504 & ~n11221;
  assign n11236 = ~n11234 & ~n11235;
  assign n11237 = ~n11232 & ~n11233;
  assign n11238 = n11236 & n11237;
  assign n11239 = ~n11222 & ~n11223;
  assign n11240 = n11231 & n11239;
  assign n11241 = n11238 & n11240;
  assign n11242 = n11216 & n11241;
  assign n11243 = n9436 & ~n11242;
  assign n11244 = P2_REG0_REG_25_ & ~n9436;
  assign n1780 = n11243 | n11244;
  assign n11246 = P2_REG1_REG_27_ & n9469;
  assign n11247 = P2_REG0_REG_27_ & n9467;
  assign n11248 = P2_REG2_REG_27_ & n9471;
  assign n11249 = P2_REG3_REG_26_ & n11187;
  assign n11250 = ~P2_REG3_REG_27_ & n11249;
  assign n11251 = P2_REG3_REG_27_ & ~n11249;
  assign n11252 = ~n11250 & ~n11251;
  assign n11253 = n9465 & ~n11252;
  assign n11254 = ~n11246 & ~n11247;
  assign n11255 = ~n11248 & n11254;
  assign n11256 = ~n11253 & n11255;
  assign n11257 = n9458 & ~n11256;
  assign n11258 = ~n9199 & ~n9446;
  assign n11259 = ~n11197 & n11258;
  assign n11260 = n11197 & ~n11258;
  assign n11261 = ~n11259 & ~n11260;
  assign n11262 = n9490 & n11261;
  assign n11263 = ~n9455 & n11258;
  assign n11264 = n11206 & ~n11209;
  assign n11265 = ~n11194 & n11258;
  assign n11266 = ~n11208 & n11258;
  assign n11267 = ~n11194 & ~n11208;
  assign n11268 = ~n11266 & ~n11267;
  assign n11269 = ~n11264 & ~n11265;
  assign n11270 = ~n11268 & n11269;
  assign n11271 = ~n11206 & ~n11208;
  assign n11272 = n11194 & n11258;
  assign n11273 = ~n11194 & ~n11258;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~n11209 & ~n11271;
  assign n11276 = n11274 & n11275;
  assign n11277 = ~n11270 & ~n11276;
  assign n11278 = n9488 & n11277;
  assign n11279 = ~n11257 & ~n11262;
  assign n11280 = ~n11263 & n11279;
  assign n11281 = ~n11278 & n11280;
  assign n11282 = ~n11202 & ~n11218;
  assign n11283 = ~n11203 & ~n11282;
  assign n11284 = n11274 & n11283;
  assign n11285 = ~n11274 & ~n11283;
  assign n11286 = ~n11284 & ~n11285;
  assign n11287 = n9511 & ~n11286;
  assign n11288 = n9561 & ~n11125;
  assign n11289 = ~n11209 & n11225;
  assign n11290 = ~n11265 & ~n11289;
  assign n11291 = ~n11268 & n11290;
  assign n11292 = ~n11208 & ~n11225;
  assign n11293 = ~n11209 & ~n11292;
  assign n11294 = n11274 & n11293;
  assign n11295 = ~n11291 & ~n11294;
  assign n11296 = n9506 & n11295;
  assign n11297 = n9508 & ~n11286;
  assign n11298 = ~n11296 & ~n11297;
  assign n11299 = n9501 & n11295;
  assign n11300 = n9495 & n11295;
  assign n11301 = n9497 & ~n11286;
  assign n11302 = n9504 & ~n11286;
  assign n11303 = ~n11301 & ~n11302;
  assign n11304 = ~n11299 & ~n11300;
  assign n11305 = n11303 & n11304;
  assign n11306 = ~n11287 & ~n11288;
  assign n11307 = n11298 & n11306;
  assign n11308 = n11305 & n11307;
  assign n11309 = n11281 & n11308;
  assign n11310 = n9436 & ~n11309;
  assign n11311 = P2_REG0_REG_26_ & ~n9436;
  assign n1785 = n11310 | n11311;
  assign n11313 = P2_REG1_REG_28_ & n9469;
  assign n11314 = P2_REG0_REG_28_ & n9467;
  assign n11315 = P2_REG2_REG_28_ & n9471;
  assign n11316 = P2_REG3_REG_27_ & n11249;
  assign n11317 = ~P2_REG3_REG_28_ & n11316;
  assign n11318 = P2_REG3_REG_28_ & ~n11316;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = n9465 & ~n11319;
  assign n11321 = ~n11313 & ~n11314;
  assign n11322 = ~n11315 & n11321;
  assign n11323 = ~n11320 & n11322;
  assign n11324 = n9458 & ~n11323;
  assign n11325 = ~n9210 & ~n9446;
  assign n11326 = n11260 & ~n11325;
  assign n11327 = ~n11260 & n11325;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = n9490 & n11328;
  assign n11330 = ~n9455 & n11325;
  assign n11331 = ~n11142 & ~n11209;
  assign n11332 = ~n11268 & ~n11331;
  assign n11333 = n11205 & ~n11268;
  assign n11334 = ~n11332 & ~n11333;
  assign n11335 = ~n11265 & n11334;
  assign n11336 = n11256 & n11325;
  assign n11337 = ~n11256 & ~n11325;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = n11335 & ~n11338;
  assign n11340 = ~n11335 & n11338;
  assign n11341 = ~n11339 & ~n11340;
  assign n11342 = n9488 & ~n11341;
  assign n11343 = ~n11324 & ~n11329;
  assign n11344 = ~n11330 & n11343;
  assign n11345 = ~n11342 & n11344;
  assign n11346 = ~n11272 & ~n11338;
  assign n11347 = ~n11273 & n11283;
  assign n11348 = n11346 & ~n11347;
  assign n11349 = ~n11273 & n11338;
  assign n11350 = ~n11272 & ~n11283;
  assign n11351 = n11349 & ~n11350;
  assign n11352 = ~n11348 & ~n11351;
  assign n11353 = n9511 & ~n11352;
  assign n11354 = n9561 & ~n11194;
  assign n11355 = n11224 & ~n11268;
  assign n11356 = ~n11332 & ~n11355;
  assign n11357 = ~n11265 & n11356;
  assign n11358 = ~n11338 & n11357;
  assign n11359 = n11338 & ~n11357;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = n9506 & ~n11360;
  assign n11362 = n9508 & ~n11352;
  assign n11363 = ~n11361 & ~n11362;
  assign n11364 = n9501 & ~n11360;
  assign n11365 = n9495 & ~n11360;
  assign n11366 = n9497 & ~n11352;
  assign n11367 = n9504 & ~n11352;
  assign n11368 = ~n11366 & ~n11367;
  assign n11369 = ~n11364 & ~n11365;
  assign n11370 = n11368 & n11369;
  assign n11371 = ~n11353 & ~n11354;
  assign n11372 = n11363 & n11371;
  assign n11373 = n11370 & n11372;
  assign n11374 = n11345 & n11373;
  assign n11375 = n9436 & ~n11374;
  assign n11376 = P2_REG0_REG_27_ & ~n9436;
  assign n1790 = n11375 | n11376;
  assign n11378 = P2_REG0_REG_29_ & n9467;
  assign n11379 = P2_REG1_REG_29_ & n9469;
  assign n11380 = P2_REG2_REG_29_ & n9471;
  assign n11381 = P2_REG3_REG_28_ & P2_REG3_REG_27_;
  assign n11382 = n11249 & n11381;
  assign n11383 = n9465 & n11382;
  assign n11384 = ~n11378 & ~n11379;
  assign n11385 = ~n11380 & n11384;
  assign n11386 = ~n11383 & n11385;
  assign n11387 = n9458 & ~n11386;
  assign n11388 = ~n9227 & ~n9446;
  assign n11389 = ~n11326 & n11388;
  assign n11390 = n11326 & ~n11388;
  assign n11391 = ~n11389 & ~n11390;
  assign n11392 = n9490 & n11391;
  assign n11393 = ~n9455 & n11388;
  assign n11394 = n11256 & ~n11325;
  assign n11395 = n11265 & ~n11394;
  assign n11396 = ~n11141 & ~n11394;
  assign n11397 = ~n11136 & ~n11268;
  assign n11398 = n11396 & n11397;
  assign n11399 = n11332 & ~n11394;
  assign n11400 = ~n11256 & n11325;
  assign n11401 = ~n11399 & ~n11400;
  assign n11402 = ~n11395 & ~n11398;
  assign n11403 = n11401 & n11402;
  assign n11404 = n11323 & n11388;
  assign n11405 = ~n11323 & ~n11388;
  assign n11406 = ~n11404 & ~n11405;
  assign n11407 = n11403 & ~n11406;
  assign n11408 = ~n11403 & n11406;
  assign n11409 = ~n11407 & ~n11408;
  assign n11410 = n9488 & ~n11409;
  assign n11411 = ~n11387 & ~n11392;
  assign n11412 = ~n11393 & n11411;
  assign n11413 = ~n11410 & n11412;
  assign n11414 = n11256 & ~n11273;
  assign n11415 = ~n11325 & ~n11414;
  assign n11416 = ~n11256 & n11273;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = ~n11336 & n11350;
  assign n11419 = n11417 & ~n11418;
  assign n11420 = ~n11406 & ~n11419;
  assign n11421 = n11406 & n11419;
  assign n11422 = ~n11420 & ~n11421;
  assign n11423 = n9511 & ~n11422;
  assign n11424 = n9561 & ~n11256;
  assign n11425 = n9508 & ~n11422;
  assign n11426 = ~n11163 & ~n11268;
  assign n11427 = n11396 & n11426;
  assign n11428 = ~n11395 & ~n11427;
  assign n11429 = n11401 & n11428;
  assign n11430 = ~n11406 & n11429;
  assign n11431 = n11406 & ~n11429;
  assign n11432 = ~n11430 & ~n11431;
  assign n11433 = n9506 & ~n11432;
  assign n11434 = n9501 & ~n11432;
  assign n11435 = n9495 & ~n11432;
  assign n11436 = n9497 & ~n11422;
  assign n11437 = n9504 & ~n11422;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = ~n11434 & ~n11435;
  assign n11440 = n11438 & n11439;
  assign n11441 = ~n11423 & ~n11424;
  assign n11442 = ~n11425 & n11441;
  assign n11443 = ~n11433 & n11442;
  assign n11444 = n11440 & n11443;
  assign n11445 = n11413 & n11444;
  assign n11446 = n9436 & ~n11445;
  assign n11447 = P2_REG0_REG_28_ & ~n9436;
  assign n1795 = n11446 | n11447;
  assign n11449 = ~n9262 & ~n9446;
  assign n11450 = ~n9455 & n11449;
  assign n11451 = n11390 & ~n11449;
  assign n11452 = ~n11390 & n11449;
  assign n11453 = ~n11451 & ~n11452;
  assign n11454 = n9490 & n11453;
  assign n11455 = n11388 & ~n11403;
  assign n11456 = ~n11323 & ~n11403;
  assign n11457 = ~n11323 & n11388;
  assign n11458 = ~n11455 & ~n11456;
  assign n11459 = ~n11457 & n11458;
  assign n11460 = n11386 & n11449;
  assign n11461 = ~n11386 & ~n11449;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = n11459 & ~n11462;
  assign n11464 = ~n11459 & n11462;
  assign n11465 = ~n11463 & ~n11464;
  assign n11466 = n9488 & ~n11465;
  assign n11467 = ~n11450 & ~n11454;
  assign n11468 = ~n11466 & n11467;
  assign n11469 = n9561 & ~n11323;
  assign n11470 = ~P2_B_REG & n9445;
  assign n11471 = ~n9446 & ~n11470;
  assign n11472 = n9457 & ~n11471;
  assign n11473 = P2_REG1_REG_30_ & n9469;
  assign n11474 = P2_REG0_REG_30_ & n9467;
  assign n11475 = P2_REG2_REG_30_ & n9471;
  assign n11476 = ~n11473 & ~n11474;
  assign n11477 = ~n11475 & n11476;
  assign n11478 = n11472 & ~n11477;
  assign n11479 = ~n11404 & ~n11462;
  assign n11480 = ~n11405 & n11419;
  assign n11481 = n11479 & ~n11480;
  assign n11482 = ~n11405 & n11462;
  assign n11483 = ~n11404 & ~n11419;
  assign n11484 = n11482 & ~n11483;
  assign n11485 = ~n11481 & ~n11484;
  assign n11486 = n9511 & ~n11485;
  assign n11487 = n11388 & ~n11429;
  assign n11488 = ~n11323 & ~n11429;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = ~n11457 & n11489;
  assign n11491 = ~n11462 & n11490;
  assign n11492 = n11462 & ~n11490;
  assign n11493 = ~n11491 & ~n11492;
  assign n11494 = n9506 & ~n11493;
  assign n11495 = n9508 & ~n11485;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = n9501 & ~n11493;
  assign n11498 = n9495 & ~n11493;
  assign n11499 = n9497 & ~n11485;
  assign n11500 = n9504 & ~n11485;
  assign n11501 = ~n11499 & ~n11500;
  assign n11502 = ~n11497 & ~n11498;
  assign n11503 = n11501 & n11502;
  assign n11504 = ~n11469 & ~n11478;
  assign n11505 = ~n11486 & n11504;
  assign n11506 = n11496 & n11505;
  assign n11507 = n11503 & n11506;
  assign n11508 = n11468 & n11507;
  assign n11509 = n9436 & ~n11508;
  assign n11510 = P2_REG0_REG_29_ & ~n9436;
  assign n1800 = n11509 | n11510;
  assign n11512 = ~n9273 & ~n9446;
  assign n11513 = ~n9455 & n11512;
  assign n11514 = P2_REG1_REG_31_ & n9469;
  assign n11515 = P2_REG0_REG_31_ & n9467;
  assign n11516 = P2_REG2_REG_31_ & n9471;
  assign n11517 = ~n11514 & ~n11515;
  assign n11518 = ~n11516 & n11517;
  assign n11519 = n11472 & ~n11518;
  assign n11520 = ~n11451 & n11512;
  assign n11521 = n11451 & ~n11512;
  assign n11522 = ~n11520 & ~n11521;
  assign n11523 = n9490 & n11522;
  assign n11524 = ~n11513 & ~n11519;
  assign n11525 = ~n11523 & n11524;
  assign n11526 = n9436 & ~n11525;
  assign n11527 = P2_REG0_REG_30_ & ~n9436;
  assign n1805 = n11526 | n11527;
  assign n11529 = ~n9284 & ~n9446;
  assign n11530 = ~n9455 & n11529;
  assign n11531 = n11521 & ~n11529;
  assign n11532 = ~n11521 & n11529;
  assign n11533 = ~n11531 & ~n11532;
  assign n11534 = n9490 & n11533;
  assign n11535 = ~n11519 & ~n11530;
  assign n11536 = ~n11534 & n11535;
  assign n11537 = n9436 & ~n11536;
  assign n11538 = P2_REG0_REG_31_ & ~n9436;
  assign n1810 = n11537 | n11538;
  assign n11540 = n9303 & ~n9352;
  assign n11541 = n9435 & n11540;
  assign n11542 = ~n9520 & n11541;
  assign n11543 = P2_REG1_REG_0_ & ~n11541;
  assign n1815 = n11542 | n11543;
  assign n11545 = ~n9576 & n11541;
  assign n11546 = P2_REG1_REG_1_ & ~n11541;
  assign n1820 = n11545 | n11546;
  assign n11548 = ~n9638 & n11541;
  assign n11549 = P2_REG1_REG_2_ & ~n11541;
  assign n1825 = n11548 | n11549;
  assign n11551 = ~n9703 & n11541;
  assign n11552 = P2_REG1_REG_3_ & ~n11541;
  assign n1830 = n11551 | n11552;
  assign n11554 = ~n9773 & n11541;
  assign n11555 = P2_REG1_REG_4_ & ~n11541;
  assign n1835 = n11554 | n11555;
  assign n11557 = ~n9838 & n11541;
  assign n11558 = P2_REG1_REG_5_ & ~n11541;
  assign n1840 = n11557 | n11558;
  assign n11560 = ~n9921 & n11541;
  assign n11561 = P2_REG1_REG_6_ & ~n11541;
  assign n1845 = n11560 | n11561;
  assign n11563 = ~n9996 & n11541;
  assign n11564 = P2_REG1_REG_7_ & ~n11541;
  assign n1850 = n11563 | n11564;
  assign n11566 = ~n10069 & n11541;
  assign n11567 = P2_REG1_REG_8_ & ~n11541;
  assign n1855 = n11566 | n11567;
  assign n11569 = ~n10142 & n11541;
  assign n11570 = P2_REG1_REG_9_ & ~n11541;
  assign n1860 = n11569 | n11570;
  assign n11572 = ~n10212 & n11541;
  assign n11573 = P2_REG1_REG_10_ & ~n11541;
  assign n1865 = n11572 | n11573;
  assign n11575 = ~n10288 & n11541;
  assign n11576 = P2_REG1_REG_11_ & ~n11541;
  assign n1870 = n11575 | n11576;
  assign n11578 = ~n10360 & n11541;
  assign n11579 = P2_REG1_REG_12_ & ~n11541;
  assign n1875 = n11578 | n11579;
  assign n11581 = ~n10429 & n11541;
  assign n11582 = P2_REG1_REG_13_ & ~n11541;
  assign n1880 = n11581 | n11582;
  assign n11584 = ~n10499 & n11541;
  assign n11585 = P2_REG1_REG_14_ & ~n11541;
  assign n1885 = n11584 | n11585;
  assign n11587 = ~n10565 & n11541;
  assign n11588 = P2_REG1_REG_15_ & ~n11541;
  assign n1890 = n11587 | n11588;
  assign n11590 = ~n10637 & n11541;
  assign n11591 = P2_REG1_REG_16_ & ~n11541;
  assign n1895 = n11590 | n11591;
  assign n11593 = ~n10711 & n11541;
  assign n11594 = P2_REG1_REG_17_ & ~n11541;
  assign n1900 = n11593 | n11594;
  assign n11596 = ~n10783 & n11541;
  assign n11597 = P2_REG1_REG_18_ & ~n11541;
  assign n1905 = n11596 | n11597;
  assign n11599 = ~n10849 & n11541;
  assign n11600 = P2_REG1_REG_19_ & ~n11541;
  assign n1910 = n11599 | n11600;
  assign n11602 = ~n10914 & n11541;
  assign n11603 = P2_REG1_REG_20_ & ~n11541;
  assign n1915 = n11602 | n11603;
  assign n11605 = ~n10978 & n11541;
  assign n11606 = P2_REG1_REG_21_ & ~n11541;
  assign n1920 = n11605 | n11606;
  assign n11608 = ~n11047 & n11541;
  assign n11609 = P2_REG1_REG_22_ & ~n11541;
  assign n1925 = n11608 | n11609;
  assign n11611 = ~n11111 & n11541;
  assign n11612 = P2_REG1_REG_23_ & ~n11541;
  assign n1930 = n11611 | n11612;
  assign n11614 = ~n11180 & n11541;
  assign n11615 = P2_REG1_REG_24_ & ~n11541;
  assign n1935 = n11614 | n11615;
  assign n11617 = ~n11242 & n11541;
  assign n11618 = P2_REG1_REG_25_ & ~n11541;
  assign n1940 = n11617 | n11618;
  assign n11620 = ~n11309 & n11541;
  assign n11621 = P2_REG1_REG_26_ & ~n11541;
  assign n1945 = n11620 | n11621;
  assign n11623 = ~n11374 & n11541;
  assign n11624 = P2_REG1_REG_27_ & ~n11541;
  assign n1950 = n11623 | n11624;
  assign n11626 = ~n11445 & n11541;
  assign n11627 = P2_REG1_REG_28_ & ~n11541;
  assign n1955 = n11626 | n11627;
  assign n11629 = ~n11508 & n11541;
  assign n11630 = P2_REG1_REG_29_ & ~n11541;
  assign n1960 = n11629 | n11630;
  assign n11632 = ~n11525 & n11541;
  assign n11633 = P2_REG1_REG_30_ & ~n11541;
  assign n1965 = n11632 | n11633;
  assign n11635 = ~n11536 & n11541;
  assign n11636 = P2_REG1_REG_31_ & ~n11541;
  assign n1970 = n11635 | n11636;
  assign n11638 = n9371 & n9450;
  assign n11639 = n9365 & n11638;
  assign n11640 = n9365 & n9451;
  assign n11641 = ~n9372 & n9457;
  assign n11642 = n9352 & ~n11641;
  assign n11643 = ~n9356 & n11642;
  assign n11644 = n9434 & n11643;
  assign n11645 = ~n11640 & ~n11644;
  assign n11646 = n9303 & ~n11645;
  assign n11647 = n11639 & n11646;
  assign n11648 = ~n9449 & n11647;
  assign n11649 = ~n9365 & n9451;
  assign n11650 = ~n9454 & ~n11649;
  assign n11651 = n11646 & ~n11650;
  assign n11652 = ~n9449 & n11651;
  assign n11653 = ~n9517 & n11646;
  assign n11654 = P2_REG2_REG_0_ & ~n11646;
  assign n11655 = ~n11653 & ~n11654;
  assign n11656 = ~n11648 & ~n11652;
  assign n11657 = n11655 & n11656;
  assign n11658 = ~n9362 & n9510;
  assign n11659 = n11646 & n11658;
  assign n11660 = ~n9486 & n11659;
  assign n11661 = n9458 & n11646;
  assign n11662 = ~n9475 & n11661;
  assign n11663 = n11640 & n11646;
  assign n11664 = P2_REG3_REG_0_ & n11663;
  assign n11665 = ~n11660 & ~n11662;
  assign n11666 = ~n11664 & n11665;
  assign n1975 = ~n11657 | ~n11666;
  assign n11668 = ~n9540 & n11647;
  assign n11669 = ~n9537 & n11651;
  assign n11670 = ~n9575 & n11646;
  assign n11671 = P2_REG2_REG_1_ & ~n11646;
  assign n11672 = ~n11670 & ~n11671;
  assign n11673 = ~n11668 & ~n11669;
  assign n11674 = n11672 & n11673;
  assign n11675 = ~n9549 & n11659;
  assign n11676 = ~n9530 & n11661;
  assign n11677 = P2_REG3_REG_1_ & n11663;
  assign n11678 = ~n11675 & ~n11676;
  assign n11679 = ~n11677 & n11678;
  assign n1980 = ~n11674 | ~n11679;
  assign n11681 = n9597 & n11647;
  assign n11682 = ~n9593 & n11651;
  assign n11683 = ~n9637 & n11646;
  assign n11684 = P2_REG2_REG_2_ & ~n11646;
  assign n11685 = ~n11683 & ~n11684;
  assign n11686 = ~n11681 & ~n11682;
  assign n11687 = n11685 & n11686;
  assign n11688 = n9611 & n11659;
  assign n11689 = ~n9586 & n11661;
  assign n11690 = P2_REG3_REG_2_ & n11663;
  assign n11691 = ~n11688 & ~n11689;
  assign n11692 = ~n11690 & n11691;
  assign n1985 = ~n11687 | ~n11692;
  assign n11694 = n9661 & n11647;
  assign n11695 = ~n9658 & n11651;
  assign n11696 = ~n9702 & n11646;
  assign n11697 = P2_REG2_REG_3_ & ~n11646;
  assign n11698 = ~n11696 & ~n11697;
  assign n11699 = ~n11694 & ~n11695;
  assign n11700 = n11698 & n11699;
  assign n11701 = ~n9676 & n11659;
  assign n11702 = ~n9651 & n11661;
  assign n11703 = ~P2_REG3_REG_3_ & n11663;
  assign n11704 = ~n11701 & ~n11702;
  assign n11705 = ~n11703 & n11704;
  assign n1990 = ~n11700 | ~n11705;
  assign n11707 = n9727 & n11647;
  assign n11708 = ~n9724 & n11651;
  assign n11709 = ~n9772 & n11646;
  assign n11710 = P2_REG2_REG_4_ & ~n11646;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = ~n11707 & ~n11708;
  assign n11713 = n11711 & n11712;
  assign n11714 = ~n9743 & n11659;
  assign n11715 = ~n9717 & n11661;
  assign n11716 = ~n9644 & n11663;
  assign n11717 = ~n11714 & ~n11715;
  assign n11718 = ~n11716 & n11717;
  assign n1995 = ~n11713 | ~n11718;
  assign n11720 = n9798 & n11647;
  assign n11721 = ~n9795 & n11651;
  assign n11722 = ~n9837 & n11646;
  assign n11723 = P2_REG2_REG_5_ & ~n11646;
  assign n11724 = ~n11722 & ~n11723;
  assign n11725 = ~n11720 & ~n11721;
  assign n11726 = n11724 & n11725;
  assign n11727 = n9813 & n11659;
  assign n11728 = ~n9788 & n11661;
  assign n11729 = ~n9710 & n11663;
  assign n11730 = ~n11727 & ~n11728;
  assign n11731 = ~n11729 & n11730;
  assign n2000 = ~n11726 | ~n11731;
  assign n11733 = n9863 & n11647;
  assign n11734 = ~n9859 & n11651;
  assign n11735 = ~n9920 & n11646;
  assign n11736 = P2_REG2_REG_6_ & ~n11646;
  assign n11737 = ~n11735 & ~n11736;
  assign n11738 = ~n11733 & ~n11734;
  assign n11739 = n11737 & n11738;
  assign n11740 = ~n9884 & n11659;
  assign n11741 = ~n9852 & n11661;
  assign n11742 = ~n9781 & n11663;
  assign n11743 = ~n11740 & ~n11741;
  assign n11744 = ~n11742 & n11743;
  assign n2005 = ~n11739 | ~n11744;
  assign n11746 = n9946 & n11647;
  assign n11747 = ~n9943 & n11651;
  assign n11748 = ~n9995 & n11646;
  assign n11749 = P2_REG2_REG_7_ & ~n11646;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = ~n11746 & ~n11747;
  assign n11752 = n11750 & n11751;
  assign n11753 = n9961 & n11659;
  assign n11754 = ~n9936 & n11661;
  assign n11755 = ~n9845 & n11663;
  assign n11756 = ~n11753 & ~n11754;
  assign n11757 = ~n11755 & n11756;
  assign n2010 = ~n11752 | ~n11757;
  assign n11759 = n10020 & n11647;
  assign n11760 = ~n10017 & n11651;
  assign n11761 = ~n10068 & n11646;
  assign n11762 = P2_REG2_REG_8_ & ~n11646;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 = ~n11759 & ~n11760;
  assign n11765 = n11763 & n11764;
  assign n11766 = ~n10037 & n11659;
  assign n11767 = ~n10010 & n11661;
  assign n11768 = ~n9929 & n11663;
  assign n11769 = ~n11766 & ~n11767;
  assign n11770 = ~n11768 & n11769;
  assign n2015 = ~n11765 | ~n11770;
  assign n11772 = n10094 & n11647;
  assign n11773 = ~n10091 & n11651;
  assign n11774 = ~n10141 & n11646;
  assign n11775 = P2_REG2_REG_9_ & ~n11646;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = ~n11772 & ~n11773;
  assign n11778 = n11776 & n11777;
  assign n11779 = ~n10107 & n11659;
  assign n11780 = ~n10084 & n11661;
  assign n11781 = ~n10003 & n11663;
  assign n11782 = ~n11779 & ~n11780;
  assign n11783 = ~n11781 & n11782;
  assign n2020 = ~n11778 | ~n11783;
  assign n11785 = n10167 & n11647;
  assign n11786 = ~n10163 & n11651;
  assign n11787 = ~n11785 & ~n11786;
  assign n11788 = n10182 & n11659;
  assign n11789 = ~n10156 & n11661;
  assign n11790 = ~n10077 & n11663;
  assign n11791 = ~n11788 & ~n11789;
  assign n11792 = ~n11790 & n11791;
  assign n11793 = ~n10211 & n11646;
  assign n11794 = P2_REG2_REG_10_ & ~n11646;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = n11787 & n11792;
  assign n2025 = ~n11795 | ~n11796;
  assign n11798 = n10237 & n11647;
  assign n11799 = ~n10234 & n11651;
  assign n11800 = ~n11798 & ~n11799;
  assign n11801 = ~n10255 & n11659;
  assign n11802 = ~n10227 & n11661;
  assign n11803 = ~n10149 & n11663;
  assign n11804 = ~n11801 & ~n11802;
  assign n11805 = ~n11803 & n11804;
  assign n11806 = ~n10287 & n11646;
  assign n11807 = P2_REG2_REG_11_ & ~n11646;
  assign n11808 = ~n11806 & ~n11807;
  assign n11809 = n11800 & n11805;
  assign n2030 = ~n11808 | ~n11809;
  assign n11811 = n10312 & n11647;
  assign n11812 = ~n10309 & n11651;
  assign n11813 = ~n11811 & ~n11812;
  assign n11814 = ~n10325 & n11659;
  assign n11815 = ~n10302 & n11661;
  assign n11816 = ~n10220 & n11663;
  assign n11817 = ~n11814 & ~n11815;
  assign n11818 = ~n11816 & n11817;
  assign n11819 = ~n10359 & n11646;
  assign n11820 = P2_REG2_REG_12_ & ~n11646;
  assign n11821 = ~n11819 & ~n11820;
  assign n11822 = n11813 & n11818;
  assign n2035 = ~n11821 | ~n11822;
  assign n11824 = n10384 & n11647;
  assign n11825 = ~n10381 & n11651;
  assign n11826 = ~n11824 & ~n11825;
  assign n11827 = ~n10295 & n11663;
  assign n11828 = ~n10374 & n11661;
  assign n11829 = n10399 & n11659;
  assign n11830 = ~n11827 & ~n11828;
  assign n11831 = ~n11829 & n11830;
  assign n11832 = ~n10428 & n11646;
  assign n11833 = P2_REG2_REG_13_ & ~n11646;
  assign n11834 = ~n11832 & ~n11833;
  assign n11835 = n11826 & n11831;
  assign n2040 = ~n11834 | ~n11835;
  assign n11837 = n10454 & n11647;
  assign n11838 = ~n10450 & n11651;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = ~n10469 & n11659;
  assign n11841 = ~n10443 & n11661;
  assign n11842 = ~n10367 & n11663;
  assign n11843 = ~n11840 & ~n11841;
  assign n11844 = ~n11842 & n11843;
  assign n11845 = ~n10498 & n11646;
  assign n11846 = P2_REG2_REG_14_ & ~n11646;
  assign n11847 = ~n11845 & ~n11846;
  assign n11848 = n11839 & n11844;
  assign n2045 = ~n11847 | ~n11848;
  assign n11850 = n10523 & n11647;
  assign n11851 = ~n10520 & n11651;
  assign n11852 = ~n11850 & ~n11851;
  assign n11853 = ~n10436 & n11663;
  assign n11854 = ~n10513 & n11661;
  assign n11855 = ~n10535 & n11659;
  assign n11856 = ~n11853 & ~n11854;
  assign n11857 = ~n11855 & n11856;
  assign n11858 = ~n10564 & n11646;
  assign n11859 = P2_REG2_REG_15_ & ~n11646;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = n11852 & n11857;
  assign n2050 = ~n11860 | ~n11861;
  assign n11863 = ~n10506 & n11663;
  assign n11864 = ~n10579 & n11661;
  assign n11865 = ~n11863 & ~n11864;
  assign n11866 = n10589 & n11647;
  assign n11867 = ~n10586 & n11651;
  assign n11868 = ~n11866 & ~n11867;
  assign n11869 = ~n10604 & n11659;
  assign n11870 = ~n10636 & n11646;
  assign n11871 = P2_REG2_REG_16_ & ~n11646;
  assign n11872 = ~n11870 & ~n11871;
  assign n11873 = n11865 & n11868;
  assign n11874 = ~n11869 & n11873;
  assign n2055 = ~n11872 | ~n11874;
  assign n11876 = ~n10575 & n11663;
  assign n11877 = ~n10651 & n11661;
  assign n11878 = ~n11876 & ~n11877;
  assign n11879 = n10661 & n11647;
  assign n11880 = ~n10658 & n11651;
  assign n11881 = ~n11879 & ~n11880;
  assign n11882 = n10676 & n11659;
  assign n11883 = ~n10710 & n11646;
  assign n11884 = P2_REG2_REG_17_ & ~n11646;
  assign n11885 = ~n11883 & ~n11884;
  assign n11886 = n11878 & n11881;
  assign n11887 = ~n11882 & n11886;
  assign n2060 = ~n11885 | ~n11887;
  assign n11889 = ~n10647 & n11663;
  assign n11890 = ~n10725 & n11661;
  assign n11891 = ~n11889 & ~n11890;
  assign n11892 = n10736 & n11647;
  assign n11893 = ~n10732 & n11651;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = ~n10753 & n11659;
  assign n11896 = ~n10782 & n11646;
  assign n11897 = P2_REG2_REG_18_ & ~n11646;
  assign n11898 = ~n11896 & ~n11897;
  assign n11899 = n11891 & n11894;
  assign n11900 = ~n11895 & n11899;
  assign n2065 = ~n11898 | ~n11900;
  assign n11902 = ~n10721 & n11663;
  assign n11903 = ~n10797 & n11661;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = n10804 & n11647;
  assign n11906 = ~n10801 & n11651;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n10817 & n11659;
  assign n11909 = ~n10848 & n11646;
  assign n11910 = P2_REG2_REG_19_ & ~n11646;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = n11904 & n11907;
  assign n11913 = ~n11908 & n11912;
  assign n2070 = ~n11911 | ~n11913;
  assign n11915 = ~n10793 & n11663;
  assign n11916 = ~n10863 & n11661;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = n10869 & n11647;
  assign n11919 = n10865 & n11651;
  assign n11920 = ~n11918 & ~n11919;
  assign n11921 = n10884 & n11659;
  assign n11922 = ~n10913 & n11646;
  assign n11923 = P2_REG2_REG_20_ & ~n11646;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = n11917 & n11920;
  assign n11926 = ~n11921 & n11925;
  assign n2075 = ~n11924 | ~n11926;
  assign n11928 = ~n10859 & n11663;
  assign n11929 = ~n10928 & n11661;
  assign n11930 = ~n11928 & ~n11929;
  assign n11931 = n10933 & n11647;
  assign n11932 = n10930 & n11651;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = n10948 & n11659;
  assign n11935 = ~n10977 & n11646;
  assign n11936 = P2_REG2_REG_21_ & ~n11646;
  assign n11937 = ~n11935 & ~n11936;
  assign n11938 = n11930 & n11933;
  assign n11939 = ~n11934 & n11938;
  assign n2080 = ~n11937 | ~n11939;
  assign n11941 = ~n10924 & n11663;
  assign n11942 = ~n10992 & n11661;
  assign n11943 = ~n11941 & ~n11942;
  assign n11944 = n10998 & n11647;
  assign n11945 = n10994 & n11651;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11016 & n11659;
  assign n11948 = ~n11046 & n11646;
  assign n11949 = P2_REG2_REG_22_ & ~n11646;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = n11943 & n11946;
  assign n11952 = ~n11947 & n11951;
  assign n2085 = ~n11950 | ~n11952;
  assign n11954 = ~n10988 & n11663;
  assign n11955 = ~n11061 & n11661;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = n11066 & n11647;
  assign n11958 = n11063 & n11651;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = ~n11078 & n11659;
  assign n11961 = ~n11110 & n11646;
  assign n11962 = P2_REG2_REG_23_ & ~n11646;
  assign n11963 = ~n11961 & ~n11962;
  assign n11964 = n11956 & n11959;
  assign n11965 = ~n11960 & n11964;
  assign n2090 = ~n11963 | ~n11965;
  assign n11967 = ~n11057 & n11663;
  assign n11968 = ~n11125 & n11661;
  assign n11969 = ~n11967 & ~n11968;
  assign n11970 = n11130 & n11647;
  assign n11971 = n11127 & n11651;
  assign n11972 = ~n11970 & ~n11971;
  assign n11973 = ~n11145 & n11659;
  assign n11974 = ~n11179 & n11646;
  assign n11975 = P2_REG2_REG_24_ & ~n11646;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = n11969 & n11972;
  assign n11978 = ~n11973 & n11977;
  assign n2095 = ~n11976 | ~n11978;
  assign n11980 = ~n11121 & n11663;
  assign n11981 = ~n11194 & n11661;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = n11199 & n11647;
  assign n11984 = n11196 & n11651;
  assign n11985 = ~n11983 & ~n11984;
  assign n11986 = ~n11212 & n11659;
  assign n11987 = ~n11241 & n11646;
  assign n11988 = P2_REG2_REG_25_ & ~n11646;
  assign n11989 = ~n11987 & ~n11988;
  assign n11990 = n11982 & n11985;
  assign n11991 = ~n11986 & n11990;
  assign n2100 = ~n11989 | ~n11991;
  assign n11993 = ~n11190 & n11663;
  assign n11994 = ~n11256 & n11661;
  assign n11995 = ~n11993 & ~n11994;
  assign n11996 = n11261 & n11647;
  assign n11997 = n11258 & n11651;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = n11277 & n11659;
  assign n12000 = ~n11308 & n11646;
  assign n12001 = P2_REG2_REG_26_ & ~n11646;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = n11995 & n11998;
  assign n12004 = ~n11999 & n12003;
  assign n2105 = ~n12002 | ~n12004;
  assign n12006 = ~n11252 & n11663;
  assign n12007 = ~n11323 & n11661;
  assign n12008 = ~n12006 & ~n12007;
  assign n12009 = n11328 & n11647;
  assign n12010 = n11325 & n11651;
  assign n12011 = ~n12009 & ~n12010;
  assign n12012 = ~n11341 & n11659;
  assign n12013 = ~n11373 & n11646;
  assign n12014 = P2_REG2_REG_27_ & ~n11646;
  assign n12015 = ~n12013 & ~n12014;
  assign n12016 = n12008 & n12011;
  assign n12017 = ~n12012 & n12016;
  assign n2110 = ~n12015 | ~n12017;
  assign n12019 = ~n11319 & n11663;
  assign n12020 = ~n11386 & n11661;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = n11391 & n11647;
  assign n12023 = n11388 & n11651;
  assign n12024 = ~n12022 & ~n12023;
  assign n12025 = ~n11409 & n11659;
  assign n12026 = ~n11444 & n11646;
  assign n12027 = P2_REG2_REG_28_ & ~n11646;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = n12021 & n12024;
  assign n12030 = ~n12025 & n12029;
  assign n2115 = ~n12028 | ~n12030;
  assign n12032 = n11382 & n11663;
  assign n12033 = n11449 & n11651;
  assign n12034 = n11453 & n11647;
  assign n12035 = ~n11465 & n11659;
  assign n12036 = ~n11507 & n11646;
  assign n12037 = P2_REG2_REG_29_ & ~n11646;
  assign n12038 = ~n12036 & ~n12037;
  assign n12039 = ~n12032 & ~n12033;
  assign n12040 = ~n12034 & n12039;
  assign n12041 = ~n12035 & n12040;
  assign n2120 = ~n12038 | ~n12041;
  assign n12043 = n11519 & n11646;
  assign n12044 = P2_REG2_REG_30_ & ~n11646;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046 = n11512 & n11651;
  assign n12047 = n11522 & n11647;
  assign n12048 = n12045 & ~n12046;
  assign n2125 = n12047 | ~n12048;
  assign n12050 = P2_REG2_REG_31_ & ~n11646;
  assign n12051 = ~n12043 & ~n12050;
  assign n12052 = n11529 & n11651;
  assign n12053 = n11533 & n11647;
  assign n12054 = n12051 & ~n12052;
  assign n2130 = n12053 | ~n12054;
  assign n12056 = n9290 & n9301;
  assign n2555 = P2_STATE_REG & n12056;
  assign n12058 = n9442 & ~n9445;
  assign n12059 = ~P2_REG1_REG_18_ & n10729;
  assign n12060 = P2_REG1_REG_19_ & n9371;
  assign n12061 = ~P2_REG1_REG_19_ & ~n9371;
  assign n12062 = ~n12060 & ~n12061;
  assign n12063 = P2_REG1_REG_16_ & ~n10583;
  assign n12064 = P2_REG1_REG_17_ & n12063;
  assign n12065 = ~P2_REG1_REG_17_ & ~n12063;
  assign n12066 = ~n10655 & ~n12065;
  assign n12067 = ~P2_REG1_REG_16_ & n10583;
  assign n12068 = ~P2_REG1_REG_17_ & n10655;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = P2_REG1_REG_15_ & ~n10517;
  assign n12071 = ~P2_REG1_REG_15_ & n10517;
  assign n12072 = P2_REG1_REG_14_ & ~n10447;
  assign n12073 = ~P2_REG1_REG_14_ & n10447;
  assign n12074 = ~P2_REG1_REG_13_ & n10378;
  assign n12075 = P2_REG1_REG_13_ & ~n10378;
  assign n12076 = P2_REG1_REG_12_ & ~n10306;
  assign n12077 = P2_REG1_REG_11_ & ~n10231;
  assign n12078 = ~P2_REG1_REG_12_ & n10306;
  assign n12079 = ~n12074 & ~n12078;
  assign n12080 = n12077 & n12079;
  assign n12081 = ~n12075 & ~n12076;
  assign n12082 = ~n12080 & n12081;
  assign n12083 = ~n12074 & ~n12082;
  assign n12084 = ~P2_REG1_REG_11_ & n10231;
  assign n12085 = ~P2_REG1_REG_10_ & n10160;
  assign n12086 = P2_REG1_REG_10_ & ~n10160;
  assign n12087 = P2_REG1_REG_9_ & ~n10088;
  assign n12088 = P2_REG1_REG_8_ & ~n10014;
  assign n12089 = ~P2_REG1_REG_9_ & n10088;
  assign n12090 = ~n12085 & ~n12089;
  assign n12091 = n12088 & n12090;
  assign n12092 = ~n12086 & ~n12087;
  assign n12093 = ~n12091 & n12092;
  assign n12094 = ~n12085 & ~n12093;
  assign n12095 = ~P2_REG1_REG_8_ & n10014;
  assign n12096 = P2_REG1_REG_6_ & ~n9856;
  assign n12097 = P2_REG1_REG_7_ & n12096;
  assign n12098 = ~P2_REG1_REG_7_ & ~n12096;
  assign n12099 = ~n9940 & ~n12098;
  assign n12100 = ~P2_REG1_REG_6_ & n9856;
  assign n12101 = ~P2_REG1_REG_7_ & n9940;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = P2_REG1_REG_4_ & ~n9721;
  assign n12104 = P2_REG1_REG_5_ & n12103;
  assign n12105 = ~P2_REG1_REG_5_ & ~n12103;
  assign n12106 = ~n9792 & ~n12105;
  assign n12107 = ~P2_REG1_REG_4_ & n9721;
  assign n12108 = ~P2_REG1_REG_5_ & n9792;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = P2_REG1_REG_3_ & ~n9655;
  assign n12111 = ~P2_REG1_REG_3_ & n9655;
  assign n12112 = P2_REG1_REG_2_ & ~n9590;
  assign n12113 = ~n12111 & n12112;
  assign n12114 = ~P2_REG1_REG_2_ & n9590;
  assign n12115 = ~n12111 & ~n12114;
  assign n12116 = P2_REG1_REG_0_ & ~n9439;
  assign n12117 = ~P2_REG1_REG_1_ & n9534;
  assign n12118 = n12116 & ~n12117;
  assign n12119 = P2_REG1_REG_1_ & ~n9534;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = n12115 & ~n12120;
  assign n12122 = ~n12110 & ~n12113;
  assign n12123 = ~n12121 & n12122;
  assign n12124 = n12109 & ~n12123;
  assign n12125 = ~n12104 & ~n12106;
  assign n12126 = ~n12124 & n12125;
  assign n12127 = n12102 & ~n12126;
  assign n12128 = ~n12097 & ~n12099;
  assign n12129 = ~n12127 & n12128;
  assign n12130 = n12090 & ~n12095;
  assign n12131 = ~n12129 & n12130;
  assign n12132 = ~n12094 & ~n12131;
  assign n12133 = n12079 & ~n12084;
  assign n12134 = ~n12132 & n12133;
  assign n12135 = ~n12083 & ~n12134;
  assign n12136 = ~n12073 & ~n12135;
  assign n12137 = ~n12072 & ~n12136;
  assign n12138 = ~n12071 & ~n12137;
  assign n12139 = ~n12070 & ~n12138;
  assign n12140 = n12069 & ~n12139;
  assign n12141 = ~n12064 & ~n12066;
  assign n12142 = ~n12140 & n12141;
  assign n12143 = P2_REG1_REG_18_ & ~n10729;
  assign n12144 = n12142 & ~n12143;
  assign n12145 = ~n12059 & ~n12062;
  assign n12146 = ~n12144 & n12145;
  assign n12147 = ~n12059 & ~n12142;
  assign n12148 = n12062 & ~n12143;
  assign n12149 = ~n12147 & n12148;
  assign n12150 = ~n12146 & ~n12149;
  assign n12151 = n12058 & n12150;
  assign n12152 = ~P2_REG2_REG_18_ & n10729;
  assign n12153 = P2_REG2_REG_19_ & n9371;
  assign n12154 = ~P2_REG2_REG_19_ & ~n9371;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = P2_REG2_REG_16_ & ~n10583;
  assign n12157 = P2_REG2_REG_17_ & n12156;
  assign n12158 = ~P2_REG2_REG_17_ & ~n12156;
  assign n12159 = ~n10655 & ~n12158;
  assign n12160 = ~P2_REG2_REG_16_ & n10583;
  assign n12161 = ~P2_REG2_REG_17_ & n10655;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = P2_REG2_REG_15_ & ~n10517;
  assign n12164 = ~P2_REG2_REG_15_ & n10517;
  assign n12165 = P2_REG2_REG_14_ & ~n10447;
  assign n12166 = ~P2_REG2_REG_14_ & n10447;
  assign n12167 = ~P2_REG2_REG_13_ & n10378;
  assign n12168 = P2_REG2_REG_13_ & ~n10378;
  assign n12169 = P2_REG2_REG_12_ & ~n10306;
  assign n12170 = P2_REG2_REG_11_ & ~n10231;
  assign n12171 = ~P2_REG2_REG_12_ & n10306;
  assign n12172 = ~n12167 & ~n12171;
  assign n12173 = n12170 & n12172;
  assign n12174 = ~n12168 & ~n12169;
  assign n12175 = ~n12173 & n12174;
  assign n12176 = ~n12167 & ~n12175;
  assign n12177 = ~P2_REG2_REG_11_ & n10231;
  assign n12178 = ~P2_REG2_REG_10_ & n10160;
  assign n12179 = P2_REG2_REG_10_ & ~n10160;
  assign n12180 = P2_REG2_REG_9_ & ~n10088;
  assign n12181 = P2_REG2_REG_8_ & ~n10014;
  assign n12182 = ~P2_REG2_REG_9_ & n10088;
  assign n12183 = ~n12178 & ~n12182;
  assign n12184 = n12181 & n12183;
  assign n12185 = ~n12179 & ~n12180;
  assign n12186 = ~n12184 & n12185;
  assign n12187 = ~n12178 & ~n12186;
  assign n12188 = ~P2_REG2_REG_8_ & n10014;
  assign n12189 = P2_REG2_REG_6_ & ~n9856;
  assign n12190 = P2_REG2_REG_7_ & n12189;
  assign n12191 = ~P2_REG2_REG_7_ & ~n12189;
  assign n12192 = ~n9940 & ~n12191;
  assign n12193 = ~P2_REG2_REG_6_ & n9856;
  assign n12194 = ~P2_REG2_REG_7_ & n9940;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = P2_REG2_REG_4_ & ~n9721;
  assign n12197 = P2_REG2_REG_5_ & n12196;
  assign n12198 = ~P2_REG2_REG_5_ & ~n12196;
  assign n12199 = ~n9792 & ~n12198;
  assign n12200 = ~P2_REG2_REG_4_ & n9721;
  assign n12201 = ~P2_REG2_REG_5_ & n9792;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = P2_REG2_REG_3_ & ~n9655;
  assign n12204 = ~P2_REG2_REG_3_ & n9655;
  assign n12205 = P2_REG2_REG_2_ & ~n9590;
  assign n12206 = ~n12204 & n12205;
  assign n12207 = ~P2_REG2_REG_2_ & n9590;
  assign n12208 = ~n12204 & ~n12207;
  assign n12209 = P2_REG2_REG_0_ & ~n9439;
  assign n12210 = ~P2_REG2_REG_1_ & n9534;
  assign n12211 = n12209 & ~n12210;
  assign n12212 = P2_REG2_REG_1_ & ~n9534;
  assign n12213 = ~n12211 & ~n12212;
  assign n12214 = n12208 & ~n12213;
  assign n12215 = ~n12203 & ~n12206;
  assign n12216 = ~n12214 & n12215;
  assign n12217 = n12202 & ~n12216;
  assign n12218 = ~n12197 & ~n12199;
  assign n12219 = ~n12217 & n12218;
  assign n12220 = n12195 & ~n12219;
  assign n12221 = ~n12190 & ~n12192;
  assign n12222 = ~n12220 & n12221;
  assign n12223 = n12183 & ~n12188;
  assign n12224 = ~n12222 & n12223;
  assign n12225 = ~n12187 & ~n12224;
  assign n12226 = n12172 & ~n12177;
  assign n12227 = ~n12225 & n12226;
  assign n12228 = ~n12176 & ~n12227;
  assign n12229 = ~n12166 & ~n12228;
  assign n12230 = ~n12165 & ~n12229;
  assign n12231 = ~n12164 & ~n12230;
  assign n12232 = ~n12163 & ~n12231;
  assign n12233 = n12162 & ~n12232;
  assign n12234 = ~n12157 & ~n12159;
  assign n12235 = ~n12233 & n12234;
  assign n12236 = P2_REG2_REG_18_ & ~n10729;
  assign n12237 = n12235 & ~n12236;
  assign n12238 = ~n12152 & ~n12155;
  assign n12239 = ~n12237 & n12238;
  assign n12240 = ~n12152 & ~n12235;
  assign n12241 = n12155 & ~n12236;
  assign n12242 = ~n12240 & n12241;
  assign n12243 = ~n12239 & ~n12242;
  assign n12244 = ~n9442 & ~n9445;
  assign n12245 = n12243 & n12244;
  assign n12246 = ~n9371 & n9445;
  assign n12247 = ~n12151 & ~n12245;
  assign n12248 = ~n12246 & n12247;
  assign n12249 = n2555 & ~n12248;
  assign n12250 = ~n9290 & ~n9446;
  assign n12251 = ~n9446 & ~n9457;
  assign n12252 = ~n12250 & ~n12251;
  assign n12253 = P2_STATE_REG & ~n12056;
  assign n12254 = n12252 & n12253;
  assign n12255 = n9303 & ~n12254;
  assign n12256 = ~n9506 & ~n9508;
  assign n12257 = ~n9511 & n12256;
  assign n12258 = ~n9359 & n9372;
  assign n12259 = ~n9500 & ~n12258;
  assign n12260 = ~n11658 & n12259;
  assign n12261 = ~n9497 & n12260;
  assign n12262 = ~n9504 & n12261;
  assign n12263 = ~n11639 & n12257;
  assign n12264 = n12262 & n12263;
  assign n12265 = n11650 & n12264;
  assign n12266 = ~n11640 & n12265;
  assign n12267 = n9445 & ~n12266;
  assign n12268 = ~n9371 & n12267;
  assign n12269 = n12244 & ~n12266;
  assign n12270 = n12243 & n12269;
  assign n12271 = n9442 & ~n12266;
  assign n12272 = n12150 & n12271;
  assign n12273 = ~n12268 & ~n12270;
  assign n12274 = ~n12272 & n12273;
  assign n12275 = n12255 & ~n12274;
  assign n12276 = P2_ADDR_REG_19_ & n12254;
  assign n12277 = P2_STATE_REG & ~n9290;
  assign n12278 = ~n12254 & n12277;
  assign n12279 = n9445 & n12278;
  assign n12280 = ~n9371 & n12279;
  assign n12281 = n9442 & n12278;
  assign n12282 = n12150 & n12281;
  assign n12283 = P2_REG3_REG_19_ & ~P2_STATE_REG;
  assign n12284 = n12244 & n12278;
  assign n12285 = n12243 & n12284;
  assign n12286 = ~n12276 & ~n12280;
  assign n12287 = ~n12282 & n12286;
  assign n12288 = ~n12283 & n12287;
  assign n12289 = ~n12285 & n12288;
  assign n12290 = ~n12249 & ~n12275;
  assign n2135 = ~n12289 | ~n12290;
  assign n12292 = P2_REG1_REG_18_ & n10729;
  assign n12293 = ~P2_REG1_REG_18_ & ~n10729;
  assign n12294 = ~n12292 & ~n12293;
  assign n12295 = n12142 & ~n12294;
  assign n12296 = ~n12142 & n12294;
  assign n12297 = ~n12295 & ~n12296;
  assign n12298 = n12058 & ~n12297;
  assign n12299 = P2_REG2_REG_18_ & n10729;
  assign n12300 = ~P2_REG2_REG_18_ & ~n10729;
  assign n12301 = ~n12299 & ~n12300;
  assign n12302 = n12235 & ~n12301;
  assign n12303 = ~n12235 & n12301;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = n12244 & ~n12304;
  assign n12306 = n9445 & ~n10729;
  assign n12307 = ~n12298 & ~n12305;
  assign n12308 = ~n12306 & n12307;
  assign n12309 = n2555 & ~n12308;
  assign n12310 = ~n10729 & n12267;
  assign n12311 = n12269 & ~n12304;
  assign n12312 = n12271 & ~n12297;
  assign n12313 = ~n12310 & ~n12311;
  assign n12314 = ~n12312 & n12313;
  assign n12315 = n12255 & ~n12314;
  assign n12316 = P2_ADDR_REG_18_ & n12254;
  assign n12317 = ~n10729 & n12279;
  assign n12318 = n12281 & ~n12297;
  assign n12319 = P2_REG3_REG_18_ & ~P2_STATE_REG;
  assign n12320 = n12284 & ~n12304;
  assign n12321 = ~n12316 & ~n12317;
  assign n12322 = ~n12318 & n12321;
  assign n12323 = ~n12319 & n12322;
  assign n12324 = ~n12320 & n12323;
  assign n12325 = ~n12309 & ~n12315;
  assign n2140 = ~n12324 | ~n12325;
  assign n12327 = P2_REG1_REG_17_ & ~n10655;
  assign n12328 = ~n12063 & n12139;
  assign n12329 = n12069 & ~n12327;
  assign n12330 = ~n12328 & n12329;
  assign n12331 = P2_REG1_REG_17_ & n10655;
  assign n12332 = ~P2_REG1_REG_17_ & ~n10655;
  assign n12333 = ~n12067 & ~n12139;
  assign n12334 = ~n12331 & ~n12332;
  assign n12335 = ~n12063 & n12334;
  assign n12336 = ~n12333 & n12335;
  assign n12337 = ~n12330 & ~n12336;
  assign n12338 = n12058 & n12337;
  assign n12339 = P2_REG2_REG_17_ & ~n10655;
  assign n12340 = ~n12156 & n12232;
  assign n12341 = n12162 & ~n12339;
  assign n12342 = ~n12340 & n12341;
  assign n12343 = P2_REG2_REG_17_ & n10655;
  assign n12344 = ~P2_REG2_REG_17_ & ~n10655;
  assign n12345 = ~n12160 & ~n12232;
  assign n12346 = ~n12343 & ~n12344;
  assign n12347 = ~n12156 & n12346;
  assign n12348 = ~n12345 & n12347;
  assign n12349 = ~n12342 & ~n12348;
  assign n12350 = n12244 & n12349;
  assign n12351 = n9445 & ~n10655;
  assign n12352 = ~n12338 & ~n12350;
  assign n12353 = ~n12351 & n12352;
  assign n12354 = n2555 & ~n12353;
  assign n12355 = ~n10655 & n12267;
  assign n12356 = n12269 & n12349;
  assign n12357 = n12271 & n12337;
  assign n12358 = ~n12355 & ~n12356;
  assign n12359 = ~n12357 & n12358;
  assign n12360 = n12255 & ~n12359;
  assign n12361 = P2_ADDR_REG_17_ & n12254;
  assign n12362 = ~n10655 & n12279;
  assign n12363 = n12281 & n12337;
  assign n12364 = P2_REG3_REG_17_ & ~P2_STATE_REG;
  assign n12365 = n12284 & n12349;
  assign n12366 = ~n12361 & ~n12362;
  assign n12367 = ~n12363 & n12366;
  assign n12368 = ~n12364 & n12367;
  assign n12369 = ~n12365 & n12368;
  assign n12370 = ~n12354 & ~n12360;
  assign n2145 = ~n12369 | ~n12370;
  assign n12372 = P2_REG1_REG_16_ & n10583;
  assign n12373 = ~P2_REG1_REG_16_ & ~n10583;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = n12139 & ~n12374;
  assign n12376 = ~n12063 & ~n12067;
  assign n12377 = ~n12139 & ~n12376;
  assign n12378 = ~n12375 & ~n12377;
  assign n12379 = n12058 & ~n12378;
  assign n12380 = P2_REG2_REG_16_ & n10583;
  assign n12381 = ~P2_REG2_REG_16_ & ~n10583;
  assign n12382 = ~n12380 & ~n12381;
  assign n12383 = n12232 & ~n12382;
  assign n12384 = ~n12156 & ~n12160;
  assign n12385 = ~n12232 & ~n12384;
  assign n12386 = ~n12383 & ~n12385;
  assign n12387 = n12244 & ~n12386;
  assign n12388 = n9445 & ~n10583;
  assign n12389 = ~n12379 & ~n12387;
  assign n12390 = ~n12388 & n12389;
  assign n12391 = n2555 & ~n12390;
  assign n12392 = ~n10583 & n12267;
  assign n12393 = n12269 & ~n12386;
  assign n12394 = n12271 & ~n12378;
  assign n12395 = ~n12392 & ~n12393;
  assign n12396 = ~n12394 & n12395;
  assign n12397 = n12255 & ~n12396;
  assign n12398 = P2_ADDR_REG_16_ & n12254;
  assign n12399 = ~n10583 & n12279;
  assign n12400 = n12281 & ~n12378;
  assign n12401 = P2_REG3_REG_16_ & ~P2_STATE_REG;
  assign n12402 = n12284 & ~n12386;
  assign n12403 = ~n12398 & ~n12399;
  assign n12404 = ~n12400 & n12403;
  assign n12405 = ~n12401 & n12404;
  assign n12406 = ~n12402 & n12405;
  assign n12407 = ~n12391 & ~n12397;
  assign n2150 = ~n12406 | ~n12407;
  assign n12409 = P2_REG1_REG_15_ & n10517;
  assign n12410 = ~P2_REG1_REG_15_ & ~n10517;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = n12137 & ~n12411;
  assign n12413 = ~n12137 & n12411;
  assign n12414 = ~n12412 & ~n12413;
  assign n12415 = n12058 & ~n12414;
  assign n12416 = P2_REG2_REG_15_ & n10517;
  assign n12417 = ~P2_REG2_REG_15_ & ~n10517;
  assign n12418 = ~n12416 & ~n12417;
  assign n12419 = n12230 & ~n12418;
  assign n12420 = ~n12230 & n12418;
  assign n12421 = ~n12419 & ~n12420;
  assign n12422 = n12244 & ~n12421;
  assign n12423 = n9445 & ~n10517;
  assign n12424 = ~n12415 & ~n12422;
  assign n12425 = ~n12423 & n12424;
  assign n12426 = n2555 & ~n12425;
  assign n12427 = ~n10517 & n12267;
  assign n12428 = n12269 & ~n12421;
  assign n12429 = n12271 & ~n12414;
  assign n12430 = ~n12427 & ~n12428;
  assign n12431 = ~n12429 & n12430;
  assign n12432 = n12255 & ~n12431;
  assign n12433 = P2_ADDR_REG_15_ & n12254;
  assign n12434 = ~n10517 & n12279;
  assign n12435 = n12281 & ~n12414;
  assign n12436 = P2_REG3_REG_15_ & ~P2_STATE_REG;
  assign n12437 = n12284 & ~n12421;
  assign n12438 = ~n12433 & ~n12434;
  assign n12439 = ~n12435 & n12438;
  assign n12440 = ~n12436 & n12439;
  assign n12441 = ~n12437 & n12440;
  assign n12442 = ~n12426 & ~n12432;
  assign n2155 = ~n12441 | ~n12442;
  assign n12444 = P2_REG1_REG_14_ & n10447;
  assign n12445 = ~P2_REG1_REG_14_ & ~n10447;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = n12135 & ~n12446;
  assign n12448 = ~n12135 & n12446;
  assign n12449 = ~n12447 & ~n12448;
  assign n12450 = n12058 & ~n12449;
  assign n12451 = P2_REG2_REG_14_ & n10447;
  assign n12452 = ~P2_REG2_REG_14_ & ~n10447;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = n12228 & ~n12453;
  assign n12455 = ~n12228 & n12453;
  assign n12456 = ~n12454 & ~n12455;
  assign n12457 = n12244 & ~n12456;
  assign n12458 = n9445 & ~n10447;
  assign n12459 = ~n12450 & ~n12457;
  assign n12460 = ~n12458 & n12459;
  assign n12461 = n2555 & ~n12460;
  assign n12462 = ~n10447 & n12267;
  assign n12463 = n12269 & ~n12456;
  assign n12464 = n12271 & ~n12449;
  assign n12465 = ~n12462 & ~n12463;
  assign n12466 = ~n12464 & n12465;
  assign n12467 = n12255 & ~n12466;
  assign n12468 = P2_ADDR_REG_14_ & n12254;
  assign n12469 = ~n10447 & n12279;
  assign n12470 = n12281 & ~n12449;
  assign n12471 = P2_REG3_REG_14_ & ~P2_STATE_REG;
  assign n12472 = n12284 & ~n12456;
  assign n12473 = ~n12468 & ~n12469;
  assign n12474 = ~n12470 & n12473;
  assign n12475 = ~n12471 & n12474;
  assign n12476 = ~n12472 & n12475;
  assign n12477 = ~n12461 & ~n12467;
  assign n2160 = ~n12476 | ~n12477;
  assign n12479 = ~n12084 & ~n12132;
  assign n12480 = ~n12077 & ~n12479;
  assign n12481 = ~n12076 & n12480;
  assign n12482 = ~n12075 & n12079;
  assign n12483 = ~n12481 & n12482;
  assign n12484 = P2_REG1_REG_13_ & n10378;
  assign n12485 = ~P2_REG1_REG_13_ & ~n10378;
  assign n12486 = ~n12078 & ~n12480;
  assign n12487 = ~n12484 & ~n12485;
  assign n12488 = ~n12076 & n12487;
  assign n12489 = ~n12486 & n12488;
  assign n12490 = ~n12483 & ~n12489;
  assign n12491 = n12058 & n12490;
  assign n12492 = ~n12177 & ~n12225;
  assign n12493 = ~n12170 & ~n12492;
  assign n12494 = ~n12169 & n12493;
  assign n12495 = ~n12168 & n12172;
  assign n12496 = ~n12494 & n12495;
  assign n12497 = P2_REG2_REG_13_ & n10378;
  assign n12498 = ~P2_REG2_REG_13_ & ~n10378;
  assign n12499 = ~n12171 & ~n12493;
  assign n12500 = ~n12497 & ~n12498;
  assign n12501 = ~n12169 & n12500;
  assign n12502 = ~n12499 & n12501;
  assign n12503 = ~n12496 & ~n12502;
  assign n12504 = n12244 & n12503;
  assign n12505 = n9445 & ~n10378;
  assign n12506 = ~n12491 & ~n12504;
  assign n12507 = ~n12505 & n12506;
  assign n12508 = n2555 & ~n12507;
  assign n12509 = ~n10378 & n12267;
  assign n12510 = n12269 & n12503;
  assign n12511 = n12271 & n12490;
  assign n12512 = ~n12509 & ~n12510;
  assign n12513 = ~n12511 & n12512;
  assign n12514 = n12255 & ~n12513;
  assign n12515 = P2_ADDR_REG_13_ & n12254;
  assign n12516 = ~n10378 & n12279;
  assign n12517 = n12281 & n12490;
  assign n12518 = P2_REG3_REG_13_ & ~P2_STATE_REG;
  assign n12519 = n12284 & n12503;
  assign n12520 = ~n12515 & ~n12516;
  assign n12521 = ~n12517 & n12520;
  assign n12522 = ~n12518 & n12521;
  assign n12523 = ~n12519 & n12522;
  assign n12524 = ~n12508 & ~n12514;
  assign n2165 = ~n12523 | ~n12524;
  assign n12526 = P2_REG1_REG_12_ & n10306;
  assign n12527 = ~P2_REG1_REG_12_ & ~n10306;
  assign n12528 = ~n12526 & ~n12527;
  assign n12529 = n12480 & ~n12528;
  assign n12530 = ~n12076 & ~n12078;
  assign n12531 = ~n12480 & ~n12530;
  assign n12532 = ~n12529 & ~n12531;
  assign n12533 = n12058 & ~n12532;
  assign n12534 = P2_REG2_REG_12_ & n10306;
  assign n12535 = ~P2_REG2_REG_12_ & ~n10306;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = n12493 & ~n12536;
  assign n12538 = ~n12169 & ~n12171;
  assign n12539 = ~n12493 & ~n12538;
  assign n12540 = ~n12537 & ~n12539;
  assign n12541 = n12244 & ~n12540;
  assign n12542 = n9445 & ~n10306;
  assign n12543 = ~n12533 & ~n12541;
  assign n12544 = ~n12542 & n12543;
  assign n12545 = n2555 & ~n12544;
  assign n12546 = ~n10306 & n12267;
  assign n12547 = n12269 & ~n12540;
  assign n12548 = n12271 & ~n12532;
  assign n12549 = ~n12546 & ~n12547;
  assign n12550 = ~n12548 & n12549;
  assign n12551 = n12255 & ~n12550;
  assign n12552 = P2_ADDR_REG_12_ & n12254;
  assign n12553 = ~n10306 & n12279;
  assign n12554 = n12281 & ~n12532;
  assign n12555 = P2_REG3_REG_12_ & ~P2_STATE_REG;
  assign n12556 = n12284 & ~n12540;
  assign n12557 = ~n12552 & ~n12553;
  assign n12558 = ~n12554 & n12557;
  assign n12559 = ~n12555 & n12558;
  assign n12560 = ~n12556 & n12559;
  assign n12561 = ~n12545 & ~n12551;
  assign n2170 = ~n12560 | ~n12561;
  assign n12563 = P2_REG1_REG_11_ & n10231;
  assign n12564 = ~P2_REG1_REG_11_ & ~n10231;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = n12132 & ~n12565;
  assign n12567 = ~n12077 & ~n12084;
  assign n12568 = ~n12132 & ~n12567;
  assign n12569 = ~n12566 & ~n12568;
  assign n12570 = n12058 & ~n12569;
  assign n12571 = P2_REG2_REG_11_ & n10231;
  assign n12572 = ~P2_REG2_REG_11_ & ~n10231;
  assign n12573 = ~n12571 & ~n12572;
  assign n12574 = n12225 & ~n12573;
  assign n12575 = ~n12170 & ~n12177;
  assign n12576 = ~n12225 & ~n12575;
  assign n12577 = ~n12574 & ~n12576;
  assign n12578 = n12244 & ~n12577;
  assign n12579 = n9445 & ~n10231;
  assign n12580 = ~n12570 & ~n12578;
  assign n12581 = ~n12579 & n12580;
  assign n12582 = n2555 & ~n12581;
  assign n12583 = ~n10231 & n12267;
  assign n12584 = n12269 & ~n12577;
  assign n12585 = n12271 & ~n12569;
  assign n12586 = ~n12583 & ~n12584;
  assign n12587 = ~n12585 & n12586;
  assign n12588 = n12255 & ~n12587;
  assign n12589 = n12281 & ~n12569;
  assign n12590 = ~n10231 & n12279;
  assign n12591 = P2_ADDR_REG_11_ & n12254;
  assign n12592 = P2_REG3_REG_11_ & ~P2_STATE_REG;
  assign n12593 = n12284 & ~n12577;
  assign n12594 = ~n12589 & ~n12590;
  assign n12595 = ~n12591 & n12594;
  assign n12596 = ~n12592 & n12595;
  assign n12597 = ~n12593 & n12596;
  assign n12598 = ~n12582 & ~n12588;
  assign n2175 = ~n12597 | ~n12598;
  assign n12600 = ~n12095 & ~n12129;
  assign n12601 = ~n12088 & ~n12600;
  assign n12602 = ~n12087 & n12601;
  assign n12603 = ~n12086 & n12090;
  assign n12604 = ~n12602 & n12603;
  assign n12605 = P2_REG1_REG_10_ & n10160;
  assign n12606 = ~P2_REG1_REG_10_ & ~n10160;
  assign n12607 = ~n12089 & ~n12601;
  assign n12608 = ~n12605 & ~n12606;
  assign n12609 = ~n12087 & n12608;
  assign n12610 = ~n12607 & n12609;
  assign n12611 = ~n12604 & ~n12610;
  assign n12612 = n12058 & n12611;
  assign n12613 = ~n12188 & ~n12222;
  assign n12614 = ~n12181 & ~n12613;
  assign n12615 = ~n12180 & n12614;
  assign n12616 = ~n12179 & n12183;
  assign n12617 = ~n12615 & n12616;
  assign n12618 = P2_REG2_REG_10_ & n10160;
  assign n12619 = ~P2_REG2_REG_10_ & ~n10160;
  assign n12620 = ~n12182 & ~n12614;
  assign n12621 = ~n12618 & ~n12619;
  assign n12622 = ~n12180 & n12621;
  assign n12623 = ~n12620 & n12622;
  assign n12624 = ~n12617 & ~n12623;
  assign n12625 = n12244 & n12624;
  assign n12626 = n9445 & ~n10160;
  assign n12627 = ~n12612 & ~n12625;
  assign n12628 = ~n12626 & n12627;
  assign n12629 = n2555 & ~n12628;
  assign n12630 = ~n10160 & n12267;
  assign n12631 = n12269 & n12624;
  assign n12632 = n12271 & n12611;
  assign n12633 = ~n12630 & ~n12631;
  assign n12634 = ~n12632 & n12633;
  assign n12635 = n12255 & ~n12634;
  assign n12636 = P2_ADDR_REG_10_ & n12254;
  assign n12637 = ~n10160 & n12279;
  assign n12638 = n12281 & n12611;
  assign n12639 = P2_REG3_REG_10_ & ~P2_STATE_REG;
  assign n12640 = n12284 & n12624;
  assign n12641 = ~n12636 & ~n12637;
  assign n12642 = ~n12638 & n12641;
  assign n12643 = ~n12639 & n12642;
  assign n12644 = ~n12640 & n12643;
  assign n12645 = ~n12629 & ~n12635;
  assign n2180 = ~n12644 | ~n12645;
  assign n12647 = P2_REG1_REG_9_ & n10088;
  assign n12648 = ~P2_REG1_REG_9_ & ~n10088;
  assign n12649 = ~n12647 & ~n12648;
  assign n12650 = n12601 & ~n12649;
  assign n12651 = ~n12087 & ~n12089;
  assign n12652 = ~n12601 & ~n12651;
  assign n12653 = ~n12650 & ~n12652;
  assign n12654 = n12058 & ~n12653;
  assign n12655 = P2_REG2_REG_9_ & n10088;
  assign n12656 = ~P2_REG2_REG_9_ & ~n10088;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = n12614 & ~n12657;
  assign n12659 = ~n12180 & ~n12182;
  assign n12660 = ~n12614 & ~n12659;
  assign n12661 = ~n12658 & ~n12660;
  assign n12662 = n12244 & ~n12661;
  assign n12663 = n9445 & ~n10088;
  assign n12664 = ~n12654 & ~n12662;
  assign n12665 = ~n12663 & n12664;
  assign n12666 = n2555 & ~n12665;
  assign n12667 = ~n10088 & n12267;
  assign n12668 = n12269 & ~n12661;
  assign n12669 = n12271 & ~n12653;
  assign n12670 = ~n12667 & ~n12668;
  assign n12671 = ~n12669 & n12670;
  assign n12672 = n12255 & ~n12671;
  assign n12673 = n12281 & ~n12653;
  assign n12674 = ~n10088 & n12279;
  assign n12675 = P2_ADDR_REG_9_ & n12254;
  assign n12676 = P2_REG3_REG_9_ & ~P2_STATE_REG;
  assign n12677 = n12284 & ~n12661;
  assign n12678 = ~n12673 & ~n12674;
  assign n12679 = ~n12675 & n12678;
  assign n12680 = ~n12676 & n12679;
  assign n12681 = ~n12677 & n12680;
  assign n12682 = ~n12666 & ~n12672;
  assign n2185 = ~n12681 | ~n12682;
  assign n12684 = P2_REG1_REG_8_ & n10014;
  assign n12685 = ~P2_REG1_REG_8_ & ~n10014;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = n12129 & ~n12686;
  assign n12688 = ~n12088 & ~n12095;
  assign n12689 = ~n12129 & ~n12688;
  assign n12690 = ~n12687 & ~n12689;
  assign n12691 = n12058 & ~n12690;
  assign n12692 = P2_REG2_REG_8_ & n10014;
  assign n12693 = ~P2_REG2_REG_8_ & ~n10014;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = n12222 & ~n12694;
  assign n12696 = ~n12181 & ~n12188;
  assign n12697 = ~n12222 & ~n12696;
  assign n12698 = ~n12695 & ~n12697;
  assign n12699 = n12244 & ~n12698;
  assign n12700 = n9445 & ~n10014;
  assign n12701 = ~n12691 & ~n12699;
  assign n12702 = ~n12700 & n12701;
  assign n12703 = n2555 & ~n12702;
  assign n12704 = ~n10014 & n12267;
  assign n12705 = n12269 & ~n12698;
  assign n12706 = n12271 & ~n12690;
  assign n12707 = ~n12704 & ~n12705;
  assign n12708 = ~n12706 & n12707;
  assign n12709 = n12255 & ~n12708;
  assign n12710 = P2_REG3_REG_8_ & ~P2_STATE_REG;
  assign n12711 = n12284 & ~n12698;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = n12281 & ~n12690;
  assign n12714 = ~n10014 & n12279;
  assign n12715 = P2_ADDR_REG_8_ & n12254;
  assign n12716 = ~n12713 & ~n12714;
  assign n12717 = ~n12715 & n12716;
  assign n12718 = ~n12703 & ~n12709;
  assign n12719 = n12712 & n12718;
  assign n2190 = ~n12717 | ~n12719;
  assign n12721 = P2_REG1_REG_7_ & ~n9940;
  assign n12722 = ~n12096 & n12126;
  assign n12723 = n12102 & ~n12721;
  assign n12724 = ~n12722 & n12723;
  assign n12725 = P2_REG1_REG_7_ & n9940;
  assign n12726 = ~P2_REG1_REG_7_ & ~n9940;
  assign n12727 = ~n12100 & ~n12126;
  assign n12728 = ~n12725 & ~n12726;
  assign n12729 = ~n12096 & n12728;
  assign n12730 = ~n12727 & n12729;
  assign n12731 = ~n12724 & ~n12730;
  assign n12732 = n12058 & n12731;
  assign n12733 = P2_REG2_REG_7_ & ~n9940;
  assign n12734 = ~n12189 & n12219;
  assign n12735 = n12195 & ~n12733;
  assign n12736 = ~n12734 & n12735;
  assign n12737 = P2_REG2_REG_7_ & n9940;
  assign n12738 = ~P2_REG2_REG_7_ & ~n9940;
  assign n12739 = ~n12193 & ~n12219;
  assign n12740 = ~n12737 & ~n12738;
  assign n12741 = ~n12189 & n12740;
  assign n12742 = ~n12739 & n12741;
  assign n12743 = ~n12736 & ~n12742;
  assign n12744 = n12244 & n12743;
  assign n12745 = n9445 & ~n9940;
  assign n12746 = ~n12732 & ~n12744;
  assign n12747 = ~n12745 & n12746;
  assign n12748 = n2555 & ~n12747;
  assign n12749 = ~n9940 & n12267;
  assign n12750 = n12269 & n12743;
  assign n12751 = n12271 & n12731;
  assign n12752 = ~n12749 & ~n12750;
  assign n12753 = ~n12751 & n12752;
  assign n12754 = n12255 & ~n12753;
  assign n12755 = P2_REG3_REG_7_ & ~P2_STATE_REG;
  assign n12756 = n12284 & n12743;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = n12281 & n12731;
  assign n12759 = ~n9940 & n12279;
  assign n12760 = P2_ADDR_REG_7_ & n12254;
  assign n12761 = ~n12758 & ~n12759;
  assign n12762 = ~n12760 & n12761;
  assign n12763 = ~n12748 & ~n12754;
  assign n12764 = n12757 & n12763;
  assign n2195 = ~n12762 | ~n12764;
  assign n12766 = P2_REG1_REG_6_ & n9856;
  assign n12767 = ~P2_REG1_REG_6_ & ~n9856;
  assign n12768 = ~n12766 & ~n12767;
  assign n12769 = n12126 & ~n12768;
  assign n12770 = ~n12096 & ~n12100;
  assign n12771 = ~n12126 & ~n12770;
  assign n12772 = ~n12769 & ~n12771;
  assign n12773 = n12058 & ~n12772;
  assign n12774 = P2_REG2_REG_6_ & n9856;
  assign n12775 = ~P2_REG2_REG_6_ & ~n9856;
  assign n12776 = ~n12774 & ~n12775;
  assign n12777 = n12219 & ~n12776;
  assign n12778 = ~n12189 & ~n12193;
  assign n12779 = ~n12219 & ~n12778;
  assign n12780 = ~n12777 & ~n12779;
  assign n12781 = n12244 & ~n12780;
  assign n12782 = n9445 & ~n9856;
  assign n12783 = ~n12773 & ~n12781;
  assign n12784 = ~n12782 & n12783;
  assign n12785 = n2555 & ~n12784;
  assign n12786 = ~n9856 & n12267;
  assign n12787 = n12269 & ~n12780;
  assign n12788 = n12271 & ~n12772;
  assign n12789 = ~n12786 & ~n12787;
  assign n12790 = ~n12788 & n12789;
  assign n12791 = n12255 & ~n12790;
  assign n12792 = P2_REG3_REG_6_ & ~P2_STATE_REG;
  assign n12793 = n12284 & ~n12780;
  assign n12794 = ~n12792 & ~n12793;
  assign n12795 = n12281 & ~n12772;
  assign n12796 = ~n9856 & n12279;
  assign n12797 = P2_ADDR_REG_6_ & n12254;
  assign n12798 = ~n12795 & ~n12796;
  assign n12799 = ~n12797 & n12798;
  assign n12800 = ~n12785 & ~n12791;
  assign n12801 = n12794 & n12800;
  assign n2200 = ~n12799 | ~n12801;
  assign n12803 = P2_REG1_REG_5_ & ~n9792;
  assign n12804 = n12115 & n12118;
  assign n12805 = ~n12114 & n12119;
  assign n12806 = ~n12112 & ~n12805;
  assign n12807 = ~n12111 & ~n12806;
  assign n12808 = ~n12110 & ~n12804;
  assign n12809 = ~n12807 & n12808;
  assign n12810 = ~n12103 & n12809;
  assign n12811 = n12109 & ~n12803;
  assign n12812 = ~n12810 & n12811;
  assign n12813 = P2_REG1_REG_5_ & n9792;
  assign n12814 = ~P2_REG1_REG_5_ & ~n9792;
  assign n12815 = ~n12107 & ~n12809;
  assign n12816 = ~n12813 & ~n12814;
  assign n12817 = ~n12103 & n12816;
  assign n12818 = ~n12815 & n12817;
  assign n12819 = ~n12812 & ~n12818;
  assign n12820 = n12058 & n12819;
  assign n12821 = P2_REG2_REG_5_ & ~n9792;
  assign n12822 = n12208 & n12211;
  assign n12823 = ~n12207 & n12212;
  assign n12824 = ~n12205 & ~n12823;
  assign n12825 = ~n12204 & ~n12824;
  assign n12826 = ~n12203 & ~n12822;
  assign n12827 = ~n12825 & n12826;
  assign n12828 = ~n12196 & n12827;
  assign n12829 = n12202 & ~n12821;
  assign n12830 = ~n12828 & n12829;
  assign n12831 = P2_REG2_REG_5_ & n9792;
  assign n12832 = ~P2_REG2_REG_5_ & ~n9792;
  assign n12833 = ~n12200 & ~n12827;
  assign n12834 = ~n12831 & ~n12832;
  assign n12835 = ~n12196 & n12834;
  assign n12836 = ~n12833 & n12835;
  assign n12837 = ~n12830 & ~n12836;
  assign n12838 = n12244 & n12837;
  assign n12839 = n9445 & ~n9792;
  assign n12840 = ~n12820 & ~n12838;
  assign n12841 = ~n12839 & n12840;
  assign n12842 = n2555 & ~n12841;
  assign n12843 = ~n9792 & n12267;
  assign n12844 = n12269 & n12837;
  assign n12845 = n12271 & n12819;
  assign n12846 = ~n12843 & ~n12844;
  assign n12847 = ~n12845 & n12846;
  assign n12848 = n12255 & ~n12847;
  assign n12849 = P2_REG3_REG_5_ & ~P2_STATE_REG;
  assign n12850 = n12284 & n12837;
  assign n12851 = ~n12849 & ~n12850;
  assign n12852 = n12281 & n12819;
  assign n12853 = ~n9792 & n12279;
  assign n12854 = P2_ADDR_REG_5_ & n12254;
  assign n12855 = ~n12852 & ~n12853;
  assign n12856 = ~n12854 & n12855;
  assign n12857 = ~n12842 & ~n12848;
  assign n12858 = n12851 & n12857;
  assign n2205 = ~n12856 | ~n12858;
  assign n12860 = P2_REG1_REG_4_ & n9721;
  assign n12861 = ~P2_REG1_REG_4_ & ~n9721;
  assign n12862 = ~n12860 & ~n12861;
  assign n12863 = n12809 & ~n12862;
  assign n12864 = ~n12103 & ~n12107;
  assign n12865 = ~n12809 & ~n12864;
  assign n12866 = ~n12863 & ~n12865;
  assign n12867 = n12058 & ~n12866;
  assign n12868 = P2_REG2_REG_4_ & n9721;
  assign n12869 = ~P2_REG2_REG_4_ & ~n9721;
  assign n12870 = ~n12868 & ~n12869;
  assign n12871 = n12827 & ~n12870;
  assign n12872 = ~n12196 & ~n12200;
  assign n12873 = ~n12827 & ~n12872;
  assign n12874 = ~n12871 & ~n12873;
  assign n12875 = n12244 & ~n12874;
  assign n12876 = n9445 & ~n9721;
  assign n12877 = ~n12867 & ~n12875;
  assign n12878 = ~n12876 & n12877;
  assign n12879 = n2555 & ~n12878;
  assign n12880 = ~n9721 & n12267;
  assign n12881 = n12269 & ~n12874;
  assign n12882 = n12271 & ~n12866;
  assign n12883 = ~n12880 & ~n12881;
  assign n12884 = ~n12882 & n12883;
  assign n12885 = n12255 & ~n12884;
  assign n12886 = P2_REG3_REG_4_ & ~P2_STATE_REG;
  assign n12887 = n12284 & ~n12874;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = n12281 & ~n12866;
  assign n12890 = ~n9721 & n12279;
  assign n12891 = P2_ADDR_REG_4_ & n12254;
  assign n12892 = ~n12889 & ~n12890;
  assign n12893 = ~n12891 & n12892;
  assign n12894 = ~n12879 & ~n12885;
  assign n12895 = n12888 & n12894;
  assign n2210 = ~n12893 | ~n12895;
  assign n12897 = ~n12114 & n12118;
  assign n12898 = n12806 & ~n12897;
  assign n12899 = P2_REG1_REG_3_ & n9655;
  assign n12900 = ~P2_REG1_REG_3_ & ~n9655;
  assign n12901 = ~n12899 & ~n12900;
  assign n12902 = n12898 & ~n12901;
  assign n12903 = ~n12110 & ~n12111;
  assign n12904 = ~n12898 & ~n12903;
  assign n12905 = ~n12902 & ~n12904;
  assign n12906 = n12058 & ~n12905;
  assign n12907 = ~n12207 & n12211;
  assign n12908 = n12824 & ~n12907;
  assign n12909 = P2_REG2_REG_3_ & n9655;
  assign n12910 = ~P2_REG2_REG_3_ & ~n9655;
  assign n12911 = ~n12909 & ~n12910;
  assign n12912 = n12908 & ~n12911;
  assign n12913 = ~n12203 & ~n12204;
  assign n12914 = ~n12908 & ~n12913;
  assign n12915 = ~n12912 & ~n12914;
  assign n12916 = n12244 & ~n12915;
  assign n12917 = n9445 & ~n9655;
  assign n12918 = ~n12906 & ~n12916;
  assign n12919 = ~n12917 & n12918;
  assign n12920 = n2555 & ~n12919;
  assign n12921 = ~n9655 & n12267;
  assign n12922 = n12269 & ~n12915;
  assign n12923 = n12271 & ~n12905;
  assign n12924 = ~n12921 & ~n12922;
  assign n12925 = ~n12923 & n12924;
  assign n12926 = n12255 & ~n12925;
  assign n12927 = P2_REG3_REG_3_ & ~P2_STATE_REG;
  assign n12928 = n12284 & ~n12915;
  assign n12929 = ~n12927 & ~n12928;
  assign n12930 = n12281 & ~n12905;
  assign n12931 = ~n9655 & n12279;
  assign n12932 = P2_ADDR_REG_3_ & n12254;
  assign n12933 = ~n12930 & ~n12931;
  assign n12934 = ~n12932 & n12933;
  assign n12935 = ~n12920 & ~n12926;
  assign n12936 = n12929 & n12935;
  assign n2215 = ~n12934 | ~n12936;
  assign n12938 = ~n12112 & ~n12114;
  assign n12939 = ~n12120 & n12938;
  assign n12940 = P2_REG1_REG_2_ & n9590;
  assign n12941 = ~P2_REG1_REG_2_ & ~n9590;
  assign n12942 = ~n12940 & ~n12941;
  assign n12943 = ~n12119 & n12942;
  assign n12944 = ~n12118 & n12943;
  assign n12945 = ~n12939 & ~n12944;
  assign n12946 = n12058 & n12945;
  assign n12947 = ~n12205 & ~n12207;
  assign n12948 = ~n12213 & n12947;
  assign n12949 = P2_REG2_REG_2_ & n9590;
  assign n12950 = ~P2_REG2_REG_2_ & ~n9590;
  assign n12951 = ~n12949 & ~n12950;
  assign n12952 = ~n12212 & n12951;
  assign n12953 = ~n12211 & n12952;
  assign n12954 = ~n12948 & ~n12953;
  assign n12955 = n12244 & n12954;
  assign n12956 = n9445 & ~n9590;
  assign n12957 = ~n12946 & ~n12955;
  assign n12958 = ~n12956 & n12957;
  assign n12959 = n2555 & ~n12958;
  assign n12960 = ~n9590 & n12267;
  assign n12961 = n12269 & n12954;
  assign n12962 = n12271 & n12945;
  assign n12963 = ~n12960 & ~n12961;
  assign n12964 = ~n12962 & n12963;
  assign n12965 = n12255 & ~n12964;
  assign n12966 = P2_REG3_REG_2_ & ~P2_STATE_REG;
  assign n12967 = n12284 & n12954;
  assign n12968 = ~n12966 & ~n12967;
  assign n12969 = n12281 & n12945;
  assign n12970 = ~n9590 & n12279;
  assign n12971 = P2_ADDR_REG_2_ & n12254;
  assign n12972 = ~n12969 & ~n12970;
  assign n12973 = ~n12971 & n12972;
  assign n12974 = ~n12959 & ~n12965;
  assign n12975 = n12968 & n12974;
  assign n2220 = ~n12973 | ~n12975;
  assign n12977 = ~n12117 & ~n12119;
  assign n12978 = ~n12116 & n12977;
  assign n12979 = n12116 & ~n12977;
  assign n12980 = ~n12978 & ~n12979;
  assign n12981 = n12058 & ~n12980;
  assign n12982 = ~n12210 & ~n12212;
  assign n12983 = ~n12209 & n12982;
  assign n12984 = n12209 & ~n12982;
  assign n12985 = ~n12983 & ~n12984;
  assign n12986 = n12244 & ~n12985;
  assign n12987 = n9445 & ~n9534;
  assign n12988 = ~n12981 & ~n12986;
  assign n12989 = ~n12987 & n12988;
  assign n12990 = n2555 & ~n12989;
  assign n12991 = ~n9534 & n12267;
  assign n12992 = n12269 & ~n12985;
  assign n12993 = n12271 & ~n12980;
  assign n12994 = ~n12991 & ~n12992;
  assign n12995 = ~n12993 & n12994;
  assign n12996 = n12255 & ~n12995;
  assign n12997 = P2_REG3_REG_1_ & ~P2_STATE_REG;
  assign n12998 = n12284 & ~n12985;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = n12281 & ~n12980;
  assign n13001 = ~n9534 & n12279;
  assign n13002 = P2_ADDR_REG_1_ & n12254;
  assign n13003 = ~n13000 & ~n13001;
  assign n13004 = ~n13002 & n13003;
  assign n13005 = ~n12990 & ~n12996;
  assign n13006 = n12999 & n13005;
  assign n2225 = ~n13004 | ~n13006;
  assign n13008 = P2_REG1_REG_0_ & n9439;
  assign n13009 = ~P2_REG1_REG_0_ & ~n9439;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = n12058 & ~n13010;
  assign n13012 = P2_REG2_REG_0_ & n9439;
  assign n13013 = ~P2_REG2_REG_0_ & ~n9439;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = n12244 & ~n13014;
  assign n13016 = ~n9439 & n9445;
  assign n13017 = ~n13011 & ~n13015;
  assign n13018 = ~n13016 & n13017;
  assign n13019 = n2555 & ~n13018;
  assign n13020 = ~n9439 & n12267;
  assign n13021 = n12269 & ~n13014;
  assign n13022 = n12271 & ~n13010;
  assign n13023 = ~n13020 & ~n13021;
  assign n13024 = ~n13022 & n13023;
  assign n13025 = n12255 & ~n13024;
  assign n13026 = P2_REG3_REG_0_ & ~P2_STATE_REG;
  assign n13027 = n12284 & ~n13014;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = n12281 & ~n13010;
  assign n13030 = ~n9439 & n12279;
  assign n13031 = P2_ADDR_REG_0_ & n12254;
  assign n13032 = ~n13029 & ~n13030;
  assign n13033 = ~n13031 & n13032;
  assign n13034 = ~n13019 & ~n13025;
  assign n13035 = n13028 & n13034;
  assign n2230 = ~n13033 | ~n13035;
  assign n13037 = ~n9483 & n2555;
  assign n13038 = P2_DATAO_REG_0_ & ~n2555;
  assign n2235 = n13037 | n13038;
  assign n13040 = ~n9475 & n2555;
  assign n13041 = P2_DATAO_REG_1_ & ~n2555;
  assign n2240 = n13040 | n13041;
  assign n13043 = ~n9530 & n2555;
  assign n13044 = P2_DATAO_REG_2_ & ~n2555;
  assign n2245 = n13043 | n13044;
  assign n13046 = ~n9586 & n2555;
  assign n13047 = P2_DATAO_REG_3_ & ~n2555;
  assign n2250 = n13046 | n13047;
  assign n13049 = ~n9651 & n2555;
  assign n13050 = P2_DATAO_REG_4_ & ~n2555;
  assign n2255 = n13049 | n13050;
  assign n13052 = ~n9717 & n2555;
  assign n13053 = P2_DATAO_REG_5_ & ~n2555;
  assign n2260 = n13052 | n13053;
  assign n13055 = ~n9788 & n2555;
  assign n13056 = P2_DATAO_REG_6_ & ~n2555;
  assign n2265 = n13055 | n13056;
  assign n13058 = ~n9852 & n2555;
  assign n13059 = P2_DATAO_REG_7_ & ~n2555;
  assign n2270 = n13058 | n13059;
  assign n13061 = ~n9936 & n2555;
  assign n13062 = P2_DATAO_REG_8_ & ~n2555;
  assign n2275 = n13061 | n13062;
  assign n13064 = ~n10010 & n2555;
  assign n13065 = P2_DATAO_REG_9_ & ~n2555;
  assign n2280 = n13064 | n13065;
  assign n13067 = ~n10084 & n2555;
  assign n13068 = P2_DATAO_REG_10_ & ~n2555;
  assign n2285 = n13067 | n13068;
  assign n13070 = ~n10156 & n2555;
  assign n13071 = P2_DATAO_REG_11_ & ~n2555;
  assign n2290 = n13070 | n13071;
  assign n13073 = ~n10227 & n2555;
  assign n13074 = P2_DATAO_REG_12_ & ~n2555;
  assign n2295 = n13073 | n13074;
  assign n13076 = ~n10302 & n2555;
  assign n13077 = P2_DATAO_REG_13_ & ~n2555;
  assign n2300 = n13076 | n13077;
  assign n13079 = ~n10374 & n2555;
  assign n13080 = P2_DATAO_REG_14_ & ~n2555;
  assign n2305 = n13079 | n13080;
  assign n13082 = ~n10443 & n2555;
  assign n13083 = P2_DATAO_REG_15_ & ~n2555;
  assign n2310 = n13082 | n13083;
  assign n13085 = ~n10513 & n2555;
  assign n13086 = P2_DATAO_REG_16_ & ~n2555;
  assign n2315 = n13085 | n13086;
  assign n13088 = ~n10579 & n2555;
  assign n13089 = P2_DATAO_REG_17_ & ~n2555;
  assign n2320 = n13088 | n13089;
  assign n13091 = ~n10651 & n2555;
  assign n13092 = P2_DATAO_REG_18_ & ~n2555;
  assign n2325 = n13091 | n13092;
  assign n13094 = ~n10725 & n2555;
  assign n13095 = P2_DATAO_REG_19_ & ~n2555;
  assign n2330 = n13094 | n13095;
  assign n13097 = ~n10797 & n2555;
  assign n13098 = P2_DATAO_REG_20_ & ~n2555;
  assign n2335 = n13097 | n13098;
  assign n13100 = ~n10863 & n2555;
  assign n13101 = P2_DATAO_REG_21_ & ~n2555;
  assign n2340 = n13100 | n13101;
  assign n13103 = ~n10928 & n2555;
  assign n13104 = P2_DATAO_REG_22_ & ~n2555;
  assign n2345 = n13103 | n13104;
  assign n13106 = ~n10992 & n2555;
  assign n13107 = P2_DATAO_REG_23_ & ~n2555;
  assign n2350 = n13106 | n13107;
  assign n13109 = ~n11061 & n2555;
  assign n13110 = P2_DATAO_REG_24_ & ~n2555;
  assign n2355 = n13109 | n13110;
  assign n13112 = ~n11125 & n2555;
  assign n13113 = P2_DATAO_REG_25_ & ~n2555;
  assign n2360 = n13112 | n13113;
  assign n13115 = ~n11194 & n2555;
  assign n13116 = P2_DATAO_REG_26_ & ~n2555;
  assign n2365 = n13115 | n13116;
  assign n13118 = ~n11256 & n2555;
  assign n13119 = P2_DATAO_REG_27_ & ~n2555;
  assign n2370 = n13118 | n13119;
  assign n13121 = ~n11323 & n2555;
  assign n13122 = P2_DATAO_REG_28_ & ~n2555;
  assign n2375 = n13121 | n13122;
  assign n13124 = ~n11386 & n2555;
  assign n13125 = P2_DATAO_REG_29_ & ~n2555;
  assign n2380 = n13124 | n13125;
  assign n13127 = ~n11477 & n2555;
  assign n13128 = P2_DATAO_REG_30_ & ~n2555;
  assign n2385 = n13127 | n13128;
  assign n13130 = ~n11518 & n2555;
  assign n13131 = P2_DATAO_REG_31_ & ~n2555;
  assign n2390 = n13130 | n13131;
  assign n13133 = ~n9362 & n12258;
  assign n13134 = n12244 & n13133;
  assign n13135 = n9303 & n13134;
  assign n13136 = n9290 & ~n13135;
  assign n13137 = ~n9290 & ~n9359;
  assign n13138 = n9290 & ~n13134;
  assign n13139 = ~n13137 & ~n13138;
  assign n13140 = n12253 & n13139;
  assign n13141 = P2_B_REG & ~n13140;
  assign n13142 = n13136 & ~n13141;
  assign n13143 = ~P2_STATE_REG & ~n13141;
  assign n13144 = ~n13142 & ~n13143;
  assign n13145 = n9362 & ~n9371;
  assign n13146 = ~n9365 & n13145;
  assign n13147 = ~n10170 & ~n10171;
  assign n13148 = ~n10872 & ~n10873;
  assign n13149 = ~n10253 & ~n13147;
  assign n13150 = ~n9741 & n13149;
  assign n13151 = ~n10815 & n13150;
  assign n13152 = ~n13148 & n13151;
  assign n13153 = ~n10387 & ~n10388;
  assign n13154 = ~n10035 & ~n10105;
  assign n13155 = ~n13153 & n13154;
  assign n13156 = ~n10595 & ~n10596;
  assign n13157 = n9449 & n9483;
  assign n13158 = ~n9546 & ~n13157;
  assign n13159 = ~n10526 & ~n10527;
  assign n13160 = ~n13156 & ~n13158;
  assign n13161 = ~n9545 & n13160;
  assign n13162 = ~n13159 & n13161;
  assign n13163 = ~n9801 & ~n9802;
  assign n13164 = ~n10664 & ~n10665;
  assign n13165 = ~n9674 & ~n13163;
  assign n13166 = ~n9602 & n13165;
  assign n13167 = ~n13164 & n13166;
  assign n13168 = ~n9949 & ~n9950;
  assign n13169 = ~n9882 & ~n13168;
  assign n13170 = ~n10323 & n13169;
  assign n13171 = ~n10602 & n13170;
  assign n13172 = n13155 & n13162;
  assign n13173 = ~n10751 & n13172;
  assign n13174 = n13167 & n13173;
  assign n13175 = n13171 & n13174;
  assign n13176 = n11518 & ~n11529;
  assign n13177 = ~n11518 & n11529;
  assign n13178 = ~n13176 & ~n13177;
  assign n13179 = n11477 & ~n11512;
  assign n13180 = ~n11477 & n11512;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = n11194 & ~n11258;
  assign n13183 = ~n11265 & ~n13182;
  assign n13184 = ~n11210 & ~n13183;
  assign n13185 = ~n11069 & ~n11070;
  assign n13186 = ~n11001 & ~n11005;
  assign n13187 = ~n11133 & ~n11134;
  assign n13188 = ~n13185 & ~n13186;
  assign n13189 = ~n13187 & n13188;
  assign n13190 = ~n11143 & n13189;
  assign n13191 = ~n11394 & ~n11400;
  assign n13192 = n11323 & ~n11388;
  assign n13193 = ~n11457 & ~n13192;
  assign n13194 = n11386 & ~n11449;
  assign n13195 = ~n11386 & n11449;
  assign n13196 = ~n13194 & ~n13195;
  assign n13197 = n13184 & n13190;
  assign n13198 = ~n13191 & n13197;
  assign n13199 = ~n13193 & n13198;
  assign n13200 = ~n13196 & n13199;
  assign n13201 = n13152 & n13175;
  assign n13202 = ~n13178 & n13201;
  assign n13203 = ~n13181 & n13202;
  assign n13204 = n13200 & n13203;
  assign n13205 = n13146 & ~n13204;
  assign n13206 = n9362 & n9452;
  assign n13207 = n13204 & n13206;
  assign n13208 = n9359 & n9365;
  assign n13209 = ~n9371 & ~n13208;
  assign n13210 = ~n9362 & ~n13209;
  assign n13211 = ~n9372 & ~n13210;
  assign n13212 = ~n9359 & n13145;
  assign n13213 = ~n9511 & ~n13212;
  assign n13214 = ~n9290 & n13133;
  assign n13215 = ~n9494 & ~n11638;
  assign n13216 = ~n9451 & ~n9501;
  assign n13217 = n13215 & n13216;
  assign n13218 = n13213 & ~n13214;
  assign n13219 = n13217 & n13218;
  assign n13220 = ~n9365 & n9487;
  assign n13221 = ~n9453 & n12256;
  assign n13222 = ~n13220 & n13221;
  assign n13223 = ~n11477 & n11518;
  assign n13224 = ~n13222 & ~n13223;
  assign n13225 = n13219 & ~n13224;
  assign n13226 = ~n11518 & ~n13225;
  assign n13227 = n11477 & ~n11518;
  assign n13228 = ~n13223 & ~n13227;
  assign n13229 = ~n13222 & n13223;
  assign n13230 = n13228 & n13229;
  assign n13231 = ~n13226 & ~n13230;
  assign n13232 = n9446 & n13231;
  assign n13233 = n9359 & n11658;
  assign n13234 = ~n13230 & ~n13233;
  assign n13235 = ~n13226 & n13234;
  assign n13236 = n9284 & n13231;
  assign n13237 = ~n13232 & ~n13235;
  assign n13238 = ~n13236 & n13237;
  assign n13239 = ~n11518 & n13233;
  assign n13240 = n13219 & n13222;
  assign n13241 = ~n9446 & ~n13240;
  assign n13242 = ~n9284 & n13241;
  assign n13243 = ~n13239 & ~n13242;
  assign n13244 = n13238 & n13243;
  assign n13245 = ~n13238 & ~n13243;
  assign n13246 = ~n13244 & ~n13245;
  assign n13247 = ~n11477 & ~n13225;
  assign n13248 = n11477 & n13229;
  assign n13249 = ~n9446 & n13233;
  assign n13250 = ~n9273 & n13249;
  assign n13251 = ~n13247 & ~n13248;
  assign n13252 = ~n13250 & n13251;
  assign n13253 = ~n11477 & n13233;
  assign n13254 = n11512 & ~n13240;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = n13246 & ~n13252;
  assign n13257 = n13255 & n13256;
  assign n13258 = n9290 & n13133;
  assign n13259 = n13243 & ~n13258;
  assign n13260 = ~n13238 & n13258;
  assign n13261 = n13238 & ~n13243;
  assign n13262 = ~n13259 & ~n13260;
  assign n13263 = ~n13261 & n13262;
  assign n13264 = ~n13257 & ~n13263;
  assign n13265 = ~n10579 & n13233;
  assign n13266 = n9290 & ~n10513;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~n10658 & ~n13240;
  assign n13269 = n13267 & ~n13268;
  assign n13270 = ~n10579 & ~n13225;
  assign n13271 = ~n10579 & n13229;
  assign n13272 = ~n9290 & ~n13271;
  assign n13273 = ~n10658 & n13233;
  assign n13274 = ~n13270 & n13272;
  assign n13275 = ~n13273 & n13274;
  assign n13276 = ~n13269 & n13275;
  assign n13277 = ~n10651 & n13233;
  assign n13278 = n9290 & ~n10579;
  assign n13279 = ~n13277 & ~n13278;
  assign n13280 = ~n10732 & ~n13240;
  assign n13281 = n13279 & ~n13280;
  assign n13282 = ~n10651 & ~n13225;
  assign n13283 = ~n10651 & n13229;
  assign n13284 = ~n9290 & ~n13283;
  assign n13285 = ~n10732 & n13233;
  assign n13286 = ~n13282 & n13284;
  assign n13287 = ~n13285 & n13286;
  assign n13288 = ~n13281 & n13287;
  assign n13289 = ~n10725 & n13233;
  assign n13290 = n9290 & ~n10651;
  assign n13291 = ~n13289 & ~n13290;
  assign n13292 = ~n10801 & ~n13240;
  assign n13293 = n13291 & ~n13292;
  assign n13294 = ~n10725 & ~n13225;
  assign n13295 = ~n10725 & n13229;
  assign n13296 = ~n9290 & ~n13295;
  assign n13297 = ~n10801 & n13233;
  assign n13298 = ~n13294 & n13296;
  assign n13299 = ~n13297 & n13298;
  assign n13300 = ~n13293 & n13299;
  assign n13301 = ~n13276 & ~n13288;
  assign n13302 = ~n13300 & n13301;
  assign n13303 = ~n10928 & n13233;
  assign n13304 = n9290 & ~n10863;
  assign n13305 = ~n13303 & ~n13304;
  assign n13306 = n10994 & ~n13240;
  assign n13307 = n13305 & ~n13306;
  assign n13308 = ~n10928 & ~n13225;
  assign n13309 = ~n10928 & n13229;
  assign n13310 = ~n9290 & ~n13309;
  assign n13311 = n10994 & n13233;
  assign n13312 = ~n13308 & n13310;
  assign n13313 = ~n13311 & n13312;
  assign n13314 = ~n13307 & n13313;
  assign n13315 = ~n10992 & n13233;
  assign n13316 = n9290 & ~n10928;
  assign n13317 = ~n13315 & ~n13316;
  assign n13318 = n11063 & ~n13240;
  assign n13319 = n13317 & ~n13318;
  assign n13320 = ~n10992 & ~n13225;
  assign n13321 = ~n10992 & n13229;
  assign n13322 = ~n9290 & ~n13321;
  assign n13323 = n11063 & n13233;
  assign n13324 = ~n13320 & n13322;
  assign n13325 = ~n13323 & n13324;
  assign n13326 = ~n13319 & n13325;
  assign n13327 = ~n11061 & n13233;
  assign n13328 = n9290 & ~n10992;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = n11127 & ~n13240;
  assign n13331 = n13329 & ~n13330;
  assign n13332 = ~n11061 & ~n13225;
  assign n13333 = ~n11061 & n13229;
  assign n13334 = ~n9290 & ~n13333;
  assign n13335 = n11127 & n13233;
  assign n13336 = ~n13332 & n13334;
  assign n13337 = ~n13335 & n13336;
  assign n13338 = ~n13331 & n13337;
  assign n13339 = ~n13314 & ~n13326;
  assign n13340 = ~n13338 & n13339;
  assign n13341 = ~n10863 & n13233;
  assign n13342 = n9290 & ~n10797;
  assign n13343 = ~n13341 & ~n13342;
  assign n13344 = n10930 & ~n13240;
  assign n13345 = n13343 & ~n13344;
  assign n13346 = ~n10863 & ~n13225;
  assign n13347 = ~n10863 & n13229;
  assign n13348 = ~n9290 & ~n13347;
  assign n13349 = n10930 & n13233;
  assign n13350 = ~n13346 & n13348;
  assign n13351 = ~n13349 & n13350;
  assign n13352 = ~n13345 & n13351;
  assign n13353 = ~n10797 & n13233;
  assign n13354 = n9290 & ~n10725;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = n10865 & ~n13240;
  assign n13357 = n13355 & ~n13356;
  assign n13358 = ~n10797 & ~n13225;
  assign n13359 = ~n10797 & n13229;
  assign n13360 = ~n9290 & ~n13359;
  assign n13361 = n10865 & n13233;
  assign n13362 = ~n13358 & n13360;
  assign n13363 = ~n13361 & n13362;
  assign n13364 = ~n13357 & n13363;
  assign n13365 = ~n13352 & ~n13364;
  assign n13366 = ~n11125 & n13233;
  assign n13367 = n9290 & ~n11061;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = n11196 & ~n13240;
  assign n13370 = n13368 & ~n13369;
  assign n13371 = ~n11125 & ~n13225;
  assign n13372 = ~n11125 & n13229;
  assign n13373 = ~n9290 & ~n13372;
  assign n13374 = n11196 & n13233;
  assign n13375 = ~n13371 & n13373;
  assign n13376 = ~n13374 & n13375;
  assign n13377 = ~n13370 & n13376;
  assign n13378 = n13340 & n13365;
  assign n13379 = ~n13377 & n13378;
  assign n13380 = ~n11194 & n13233;
  assign n13381 = n9290 & ~n11125;
  assign n13382 = ~n13380 & ~n13381;
  assign n13383 = n11258 & ~n13240;
  assign n13384 = n13382 & ~n13383;
  assign n13385 = ~n11194 & ~n13225;
  assign n13386 = ~n11194 & n13229;
  assign n13387 = ~n9290 & ~n13386;
  assign n13388 = n11258 & n13233;
  assign n13389 = ~n13385 & n13387;
  assign n13390 = ~n13388 & n13389;
  assign n13391 = ~n13384 & n13390;
  assign n13392 = ~n10513 & n13233;
  assign n13393 = n9290 & ~n10443;
  assign n13394 = ~n13392 & ~n13393;
  assign n13395 = ~n10586 & ~n13240;
  assign n13396 = n13394 & ~n13395;
  assign n13397 = ~n10513 & ~n13225;
  assign n13398 = ~n10513 & n13229;
  assign n13399 = ~n9290 & ~n13398;
  assign n13400 = ~n10586 & n13233;
  assign n13401 = ~n13397 & n13399;
  assign n13402 = ~n13400 & n13401;
  assign n13403 = ~n13396 & n13402;
  assign n13404 = ~n13391 & ~n13403;
  assign n13405 = ~n11256 & n13233;
  assign n13406 = n9290 & ~n11194;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = n11325 & ~n13240;
  assign n13409 = n13407 & ~n13408;
  assign n13410 = ~n11256 & ~n13225;
  assign n13411 = ~n11256 & n13229;
  assign n13412 = ~n9290 & ~n13411;
  assign n13413 = n11325 & n13233;
  assign n13414 = ~n13410 & n13412;
  assign n13415 = ~n13413 & n13414;
  assign n13416 = ~n13409 & n13415;
  assign n13417 = n13302 & n13379;
  assign n13418 = n13404 & n13417;
  assign n13419 = ~n13416 & n13418;
  assign n13420 = n13246 & n13419;
  assign n13421 = ~n9651 & ~n13225;
  assign n13422 = ~n9724 & n13233;
  assign n13423 = ~n9290 & ~n13422;
  assign n13424 = ~n9651 & n13229;
  assign n13425 = n13423 & ~n13424;
  assign n13426 = ~n13421 & n13425;
  assign n13427 = ~n10010 & n13233;
  assign n13428 = n9290 & ~n9936;
  assign n13429 = ~n13427 & ~n13428;
  assign n13430 = ~n10091 & ~n13240;
  assign n13431 = n13429 & ~n13430;
  assign n13432 = ~n10010 & ~n13225;
  assign n13433 = ~n10010 & n13229;
  assign n13434 = ~n10091 & n13233;
  assign n13435 = ~n9290 & ~n13434;
  assign n13436 = ~n13432 & ~n13433;
  assign n13437 = n13435 & n13436;
  assign n13438 = ~n13431 & n13437;
  assign n13439 = ~n10084 & n13233;
  assign n13440 = n9290 & ~n10010;
  assign n13441 = ~n13439 & ~n13440;
  assign n13442 = ~n10163 & ~n13240;
  assign n13443 = n13441 & ~n13442;
  assign n13444 = ~n10084 & ~n13225;
  assign n13445 = ~n10084 & n13229;
  assign n13446 = ~n10163 & n13233;
  assign n13447 = ~n9290 & ~n13446;
  assign n13448 = ~n13444 & ~n13445;
  assign n13449 = n13447 & n13448;
  assign n13450 = ~n13443 & n13449;
  assign n13451 = ~n9936 & n13233;
  assign n13452 = n9290 & ~n9852;
  assign n13453 = ~n13451 & ~n13452;
  assign n13454 = ~n10017 & ~n13240;
  assign n13455 = n13453 & ~n13454;
  assign n13456 = ~n9936 & ~n13225;
  assign n13457 = ~n9936 & n13229;
  assign n13458 = ~n10017 & n13233;
  assign n13459 = ~n9290 & ~n13458;
  assign n13460 = ~n13456 & ~n13457;
  assign n13461 = n13459 & n13460;
  assign n13462 = ~n13455 & n13461;
  assign n13463 = ~n13438 & ~n13450;
  assign n13464 = ~n13462 & n13463;
  assign n13465 = ~n10156 & n13233;
  assign n13466 = n9290 & ~n10084;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = ~n10234 & ~n13240;
  assign n13469 = n13467 & ~n13468;
  assign n13470 = ~n10156 & ~n13225;
  assign n13471 = ~n10156 & n13229;
  assign n13472 = ~n10234 & n13233;
  assign n13473 = ~n9290 & ~n13472;
  assign n13474 = ~n13470 & ~n13471;
  assign n13475 = n13473 & n13474;
  assign n13476 = ~n13469 & n13475;
  assign n13477 = ~n10302 & n13233;
  assign n13478 = n9290 & ~n10227;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = ~n10381 & ~n13240;
  assign n13481 = n13479 & ~n13480;
  assign n13482 = ~n10302 & ~n13225;
  assign n13483 = ~n10302 & n13229;
  assign n13484 = ~n9290 & ~n13483;
  assign n13485 = ~n10381 & n13233;
  assign n13486 = ~n13482 & n13484;
  assign n13487 = ~n13485 & n13486;
  assign n13488 = ~n13481 & n13487;
  assign n13489 = ~n10227 & n13233;
  assign n13490 = n9290 & ~n10156;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = ~n10309 & ~n13240;
  assign n13493 = n13491 & ~n13492;
  assign n13494 = ~n10227 & ~n13225;
  assign n13495 = ~n10227 & n13229;
  assign n13496 = ~n9290 & ~n13495;
  assign n13497 = ~n10309 & n13233;
  assign n13498 = ~n13494 & n13496;
  assign n13499 = ~n13497 & n13498;
  assign n13500 = ~n13493 & n13499;
  assign n13501 = ~n10374 & n13233;
  assign n13502 = n9290 & ~n10302;
  assign n13503 = ~n13501 & ~n13502;
  assign n13504 = ~n10450 & ~n13240;
  assign n13505 = n13503 & ~n13504;
  assign n13506 = ~n10374 & ~n13225;
  assign n13507 = ~n10374 & n13229;
  assign n13508 = ~n9290 & ~n13507;
  assign n13509 = ~n10450 & n13233;
  assign n13510 = ~n13506 & n13508;
  assign n13511 = ~n13509 & n13510;
  assign n13512 = ~n13505 & n13511;
  assign n13513 = ~n13476 & ~n13488;
  assign n13514 = ~n13500 & n13513;
  assign n13515 = ~n13512 & n13514;
  assign n13516 = n13464 & n13515;
  assign n13517 = ~n10443 & n13233;
  assign n13518 = n9290 & ~n10374;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = ~n10520 & ~n13240;
  assign n13521 = n13519 & ~n13520;
  assign n13522 = ~n10443 & ~n13225;
  assign n13523 = ~n10443 & n13229;
  assign n13524 = ~n9290 & ~n13523;
  assign n13525 = ~n10520 & n13233;
  assign n13526 = ~n13522 & n13524;
  assign n13527 = ~n13525 & n13526;
  assign n13528 = ~n13521 & n13527;
  assign n13529 = n13516 & ~n13528;
  assign n13530 = ~n11323 & n13233;
  assign n13531 = n9290 & ~n11256;
  assign n13532 = ~n13530 & ~n13531;
  assign n13533 = n11388 & ~n13240;
  assign n13534 = n13532 & ~n13533;
  assign n13535 = ~n11323 & ~n13225;
  assign n13536 = ~n11323 & n13229;
  assign n13537 = ~n9290 & ~n13536;
  assign n13538 = n11388 & n13233;
  assign n13539 = ~n13535 & n13537;
  assign n13540 = ~n13538 & n13539;
  assign n13541 = ~n13534 & n13540;
  assign n13542 = ~n11386 & n13233;
  assign n13543 = n9290 & ~n11323;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = n11449 & ~n13240;
  assign n13546 = n13544 & ~n13545;
  assign n13547 = ~n11386 & ~n13225;
  assign n13548 = ~n11386 & n13229;
  assign n13549 = ~n9290 & ~n13548;
  assign n13550 = n11449 & n13233;
  assign n13551 = ~n13547 & n13549;
  assign n13552 = ~n13550 & n13551;
  assign n13553 = ~n13546 & n13552;
  assign n13554 = ~n13426 & n13529;
  assign n13555 = ~n13541 & n13554;
  assign n13556 = ~n13553 & n13555;
  assign n13557 = ~n9852 & n13233;
  assign n13558 = ~n9943 & ~n13240;
  assign n13559 = n9290 & ~n9788;
  assign n13560 = ~n13557 & ~n13558;
  assign n13561 = ~n13559 & n13560;
  assign n13562 = ~n9852 & ~n13225;
  assign n13563 = ~n9852 & n13229;
  assign n13564 = ~n9943 & n13233;
  assign n13565 = ~n9290 & ~n13564;
  assign n13566 = ~n13562 & ~n13563;
  assign n13567 = n13565 & n13566;
  assign n13568 = ~n13561 & n13567;
  assign n13569 = ~n9788 & n13233;
  assign n13570 = ~n9859 & ~n13240;
  assign n13571 = n9290 & ~n9717;
  assign n13572 = ~n13569 & ~n13570;
  assign n13573 = ~n13571 & n13572;
  assign n13574 = ~n9788 & ~n13225;
  assign n13575 = ~n9788 & n13229;
  assign n13576 = ~n9859 & n13233;
  assign n13577 = ~n9290 & ~n13576;
  assign n13578 = ~n13574 & ~n13575;
  assign n13579 = n13577 & n13578;
  assign n13580 = ~n13573 & n13579;
  assign n13581 = ~n9717 & n13233;
  assign n13582 = ~n9795 & ~n13240;
  assign n13583 = n9290 & ~n9651;
  assign n13584 = ~n13581 & ~n13582;
  assign n13585 = ~n13583 & n13584;
  assign n13586 = ~n9717 & ~n13225;
  assign n13587 = ~n9717 & n13229;
  assign n13588 = ~n9795 & n13233;
  assign n13589 = ~n9290 & ~n13588;
  assign n13590 = ~n13586 & ~n13587;
  assign n13591 = n13589 & n13590;
  assign n13592 = ~n13585 & n13591;
  assign n13593 = ~n9651 & n13233;
  assign n13594 = ~n9724 & ~n13240;
  assign n13595 = n9290 & ~n9586;
  assign n13596 = ~n13593 & ~n13594;
  assign n13597 = ~n13595 & n13596;
  assign n13598 = n13252 & ~n13255;
  assign n13599 = ~n13568 & ~n13580;
  assign n13600 = ~n13592 & n13599;
  assign n13601 = n13597 & n13600;
  assign n13602 = ~n13598 & n13601;
  assign n13603 = n13420 & n13556;
  assign n13604 = n13602 & n13603;
  assign n13605 = ~n9530 & ~n13225;
  assign n13606 = ~n9593 & n13233;
  assign n13607 = ~n9290 & ~n13606;
  assign n13608 = ~n9530 & n13229;
  assign n13609 = n13607 & ~n13608;
  assign n13610 = ~n13605 & n13609;
  assign n13611 = n13426 & ~n13597;
  assign n13612 = n13599 & ~n13611;
  assign n13613 = ~n13592 & n13612;
  assign n13614 = ~n13610 & n13613;
  assign n13615 = ~n9530 & n13233;
  assign n13616 = ~n9593 & ~n13240;
  assign n13617 = n9290 & ~n9475;
  assign n13618 = ~n13615 & ~n13616;
  assign n13619 = ~n13617 & n13618;
  assign n13620 = ~n9586 & n13233;
  assign n13621 = ~n9658 & ~n13240;
  assign n13622 = n9290 & ~n9530;
  assign n13623 = ~n13620 & ~n13621;
  assign n13624 = ~n13622 & n13623;
  assign n13625 = ~n9586 & ~n13225;
  assign n13626 = ~n9658 & n13233;
  assign n13627 = ~n9290 & ~n13626;
  assign n13628 = ~n9586 & n13229;
  assign n13629 = n13627 & ~n13628;
  assign n13630 = ~n13625 & n13629;
  assign n13631 = ~n13624 & n13630;
  assign n13632 = ~n13553 & n13619;
  assign n13633 = ~n13631 & n13632;
  assign n13634 = ~n13541 & n13633;
  assign n13635 = n13529 & n13614;
  assign n13636 = n13420 & n13635;
  assign n13637 = ~n13598 & n13636;
  assign n13638 = n13634 & n13637;
  assign n13639 = n13264 & ~n13604;
  assign n13640 = ~n13638 & n13639;
  assign n13641 = ~n13488 & ~n13500;
  assign n13642 = ~n13512 & n13641;
  assign n13643 = ~n13528 & n13642;
  assign n13644 = ~n13461 & n13463;
  assign n13645 = n13643 & n13644;
  assign n13646 = n13455 & ~n13553;
  assign n13647 = ~n13476 & n13646;
  assign n13648 = ~n13541 & n13647;
  assign n13649 = n13420 & n13645;
  assign n13650 = ~n13598 & n13649;
  assign n13651 = n13648 & n13650;
  assign n13652 = ~n13449 & ~n13476;
  assign n13653 = n13643 & n13652;
  assign n13654 = n13443 & ~n13541;
  assign n13655 = ~n13553 & n13654;
  assign n13656 = ~n13598 & n13655;
  assign n13657 = n13420 & n13653;
  assign n13658 = n13656 & n13657;
  assign n13659 = ~n13511 & ~n13528;
  assign n13660 = n13505 & ~n13541;
  assign n13661 = ~n13553 & n13660;
  assign n13662 = ~n13598 & n13661;
  assign n13663 = n13420 & n13659;
  assign n13664 = n13662 & n13663;
  assign n13665 = n13302 & ~n13402;
  assign n13666 = ~n13391 & ~n13416;
  assign n13667 = n13396 & ~n13553;
  assign n13668 = n13246 & ~n13541;
  assign n13669 = n13667 & n13668;
  assign n13670 = n13379 & n13665;
  assign n13671 = n13666 & n13670;
  assign n13672 = ~n13598 & n13671;
  assign n13673 = n13669 & n13672;
  assign n13674 = ~n13651 & ~n13658;
  assign n13675 = ~n13664 & n13674;
  assign n13676 = ~n13673 & n13675;
  assign n13677 = ~n13580 & n13585;
  assign n13678 = ~n13568 & n13677;
  assign n13679 = ~n13553 & n13678;
  assign n13680 = ~n13598 & n13679;
  assign n13681 = n13529 & ~n13591;
  assign n13682 = ~n13541 & n13681;
  assign n13683 = n13420 & n13682;
  assign n13684 = n13680 & n13683;
  assign n13685 = ~n13568 & n13573;
  assign n13686 = ~n13553 & n13685;
  assign n13687 = ~n13598 & n13686;
  assign n13688 = n13529 & ~n13579;
  assign n13689 = ~n13541 & n13688;
  assign n13690 = n13420 & n13689;
  assign n13691 = n13687 & n13690;
  assign n13692 = ~n13512 & ~n13528;
  assign n13693 = ~n13487 & n13692;
  assign n13694 = n13481 & ~n13541;
  assign n13695 = ~n13553 & n13694;
  assign n13696 = ~n13598 & n13695;
  assign n13697 = n13420 & n13693;
  assign n13698 = n13696 & n13697;
  assign n13699 = ~n13299 & n13666;
  assign n13700 = n13293 & ~n13541;
  assign n13701 = ~n13553 & n13700;
  assign n13702 = ~n13598 & n13701;
  assign n13703 = n13246 & n13379;
  assign n13704 = n13699 & n13703;
  assign n13705 = n13702 & n13704;
  assign n13706 = ~n13698 & ~n13705;
  assign n13707 = ~n13377 & ~n13541;
  assign n13708 = n13307 & ~n13326;
  assign n13709 = ~n13338 & n13708;
  assign n13710 = ~n13553 & n13709;
  assign n13711 = ~n13598 & n13710;
  assign n13712 = ~n13313 & n13666;
  assign n13713 = n13246 & n13712;
  assign n13714 = n13707 & n13713;
  assign n13715 = n13711 & n13714;
  assign n13716 = ~n13363 & n13666;
  assign n13717 = ~n13352 & n13357;
  assign n13718 = ~n13541 & n13717;
  assign n13719 = ~n13553 & n13718;
  assign n13720 = ~n13598 & n13719;
  assign n13721 = n13340 & ~n13377;
  assign n13722 = n13246 & n13721;
  assign n13723 = n13716 & n13722;
  assign n13724 = n13720 & n13723;
  assign n13725 = ~n13715 & ~n13724;
  assign n13726 = ~n13541 & n13561;
  assign n13727 = ~n13553 & n13726;
  assign n13728 = ~n13598 & n13727;
  assign n13729 = n13529 & ~n13567;
  assign n13730 = n13420 & n13729;
  assign n13731 = n13728 & n13730;
  assign n13732 = ~n13684 & ~n13691;
  assign n13733 = n13706 & n13732;
  assign n13734 = n13725 & n13733;
  assign n13735 = ~n13731 & n13734;
  assign n13736 = n13331 & ~n13541;
  assign n13737 = ~n13553 & n13736;
  assign n13738 = ~n13598 & n13737;
  assign n13739 = ~n13337 & n13666;
  assign n13740 = n13246 & n13739;
  assign n13741 = ~n13377 & n13740;
  assign n13742 = n13738 & n13741;
  assign n13743 = ~n13437 & ~n13450;
  assign n13744 = n13643 & n13743;
  assign n13745 = n13431 & ~n13553;
  assign n13746 = ~n13476 & n13745;
  assign n13747 = ~n13541 & n13746;
  assign n13748 = n13420 & n13744;
  assign n13749 = ~n13598 & n13748;
  assign n13750 = n13747 & n13749;
  assign n13751 = ~n13351 & n13666;
  assign n13752 = n13345 & ~n13553;
  assign n13753 = ~n13377 & n13752;
  assign n13754 = ~n13541 & n13753;
  assign n13755 = n13246 & n13340;
  assign n13756 = n13751 & n13755;
  assign n13757 = ~n13598 & n13756;
  assign n13758 = n13754 & n13757;
  assign n13759 = n13319 & ~n13338;
  assign n13760 = ~n13541 & n13759;
  assign n13761 = ~n13553 & n13760;
  assign n13762 = ~n13598 & n13761;
  assign n13763 = ~n13325 & n13666;
  assign n13764 = n13246 & n13763;
  assign n13765 = ~n13377 & n13764;
  assign n13766 = n13762 & n13765;
  assign n13767 = ~n13758 & ~n13766;
  assign n13768 = n13269 & ~n13553;
  assign n13769 = ~n13288 & n13768;
  assign n13770 = ~n13541 & n13769;
  assign n13771 = ~n13275 & n13666;
  assign n13772 = ~n13300 & n13379;
  assign n13773 = n13246 & n13772;
  assign n13774 = n13771 & n13773;
  assign n13775 = ~n13598 & n13774;
  assign n13776 = n13770 & n13775;
  assign n13777 = ~n13287 & n13666;
  assign n13778 = n13281 & ~n13553;
  assign n13779 = ~n13300 & n13778;
  assign n13780 = ~n13541 & n13779;
  assign n13781 = n13703 & n13777;
  assign n13782 = ~n13598 & n13781;
  assign n13783 = n13780 & n13782;
  assign n13784 = ~n13776 & ~n13783;
  assign n13785 = ~n13527 & ~n13541;
  assign n13786 = n13521 & ~n13553;
  assign n13787 = ~n13598 & n13786;
  assign n13788 = n13420 & n13785;
  assign n13789 = n13787 & n13788;
  assign n13790 = ~n13742 & ~n13750;
  assign n13791 = n13767 & n13790;
  assign n13792 = n13784 & n13791;
  assign n13793 = ~n13789 & n13792;
  assign n13794 = ~n9475 & ~n13225;
  assign n13795 = ~n9537 & n13233;
  assign n13796 = ~n9290 & ~n13795;
  assign n13797 = ~n9475 & n13229;
  assign n13798 = n13796 & ~n13797;
  assign n13799 = ~n13794 & n13798;
  assign n13800 = n13610 & ~n13619;
  assign n13801 = ~n13631 & ~n13800;
  assign n13802 = ~n13799 & n13801;
  assign n13803 = n13613 & n13802;
  assign n13804 = ~n9475 & n13233;
  assign n13805 = ~n9537 & ~n13240;
  assign n13806 = n9290 & ~n9483;
  assign n13807 = ~n13804 & ~n13805;
  assign n13808 = ~n13806 & n13807;
  assign n13809 = ~n13553 & n13808;
  assign n13810 = ~n13598 & n13809;
  assign n13811 = n13529 & n13803;
  assign n13812 = ~n13541 & n13811;
  assign n13813 = n13420 & n13812;
  assign n13814 = n13810 & n13813;
  assign n13815 = ~n9483 & ~n13225;
  assign n13816 = ~n9449 & n13233;
  assign n13817 = ~n9290 & ~n13816;
  assign n13818 = ~n9483 & n13229;
  assign n13819 = n13817 & ~n13818;
  assign n13820 = ~n13815 & n13819;
  assign n13821 = ~n9362 & n9365;
  assign n13822 = ~n9487 & n13821;
  assign n13823 = ~n9290 & n13822;
  assign n13824 = n13820 & n13823;
  assign n13825 = n13613 & n13801;
  assign n13826 = n13516 & ~n13824;
  assign n13827 = n13825 & n13826;
  assign n13828 = n13799 & ~n13808;
  assign n13829 = ~n13528 & ~n13828;
  assign n13830 = ~n9483 & n13233;
  assign n13831 = ~n9449 & ~n13240;
  assign n13832 = ~n13830 & ~n13831;
  assign n13833 = ~n13820 & ~n13823;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = n13829 & ~n13834;
  assign n13836 = ~n13541 & n13835;
  assign n13837 = ~n13553 & n13836;
  assign n13838 = ~n13598 & n13837;
  assign n13839 = n13420 & n13827;
  assign n13840 = n13838 & n13839;
  assign n13841 = ~n13814 & ~n13840;
  assign n13842 = n13613 & ~n13630;
  assign n13843 = ~n13541 & n13624;
  assign n13844 = ~n13553 & n13843;
  assign n13845 = ~n13598 & n13844;
  assign n13846 = n13529 & n13842;
  assign n13847 = n13420 & n13846;
  assign n13848 = n13845 & n13847;
  assign n13849 = n13246 & ~n13598;
  assign n13850 = n13546 & ~n13552;
  assign n13851 = n13384 & ~n13416;
  assign n13852 = ~n13553 & n13851;
  assign n13853 = ~n13390 & n13852;
  assign n13854 = ~n13541 & n13853;
  assign n13855 = ~n13850 & ~n13854;
  assign n13856 = n13849 & ~n13855;
  assign n13857 = ~n13848 & ~n13856;
  assign n13858 = ~n13475 & n13643;
  assign n13859 = n13469 & ~n13541;
  assign n13860 = ~n13553 & n13859;
  assign n13861 = ~n13598 & n13860;
  assign n13862 = n13420 & n13858;
  assign n13863 = n13861 & n13862;
  assign n13864 = n13409 & ~n13415;
  assign n13865 = n13534 & ~n13540;
  assign n13866 = ~n13864 & ~n13865;
  assign n13867 = n13370 & ~n13376;
  assign n13868 = n13666 & n13867;
  assign n13869 = n13866 & ~n13868;
  assign n13870 = ~n13541 & ~n13553;
  assign n13871 = ~n13598 & n13870;
  assign n13872 = n13246 & ~n13869;
  assign n13873 = n13871 & n13872;
  assign n13874 = ~n13488 & ~n13512;
  assign n13875 = ~n13499 & n13874;
  assign n13876 = n13493 & ~n13553;
  assign n13877 = ~n13528 & n13876;
  assign n13878 = ~n13541 & n13877;
  assign n13879 = n13420 & n13875;
  assign n13880 = ~n13598 & n13879;
  assign n13881 = n13878 & n13880;
  assign n13882 = ~n13863 & ~n13873;
  assign n13883 = ~n13881 & n13882;
  assign n13884 = n13841 & n13857;
  assign n13885 = n13883 & n13884;
  assign n13886 = n13640 & n13676;
  assign n13887 = n13735 & n13886;
  assign n13888 = n13793 & n13887;
  assign n13889 = n13885 & n13888;
  assign n13890 = ~n13211 & n13889;
  assign n13891 = n9365 & n13145;
  assign n13892 = ~n9511 & ~n13891;
  assign n13893 = ~n9504 & n13892;
  assign n13894 = ~n13889 & ~n13893;
  assign n13895 = ~n13890 & ~n13894;
  assign n13896 = ~n13205 & ~n13207;
  assign n13897 = ~n13141 & n13896;
  assign n13898 = n13895 & n13897;
  assign n2395 = n13144 & ~n13898;
  assign n13900 = n9303 & ~n11650;
  assign n13901 = ~n9352 & ~n9356;
  assign n13902 = n9434 & n13901;
  assign n13903 = n13900 & ~n13902;
  assign n13904 = n9290 & ~n11641;
  assign n13905 = ~n12056 & n13904;
  assign n13906 = ~n9494 & ~n13212;
  assign n13907 = ~n9501 & n13906;
  assign n13908 = ~n9453 & ~n13220;
  assign n13909 = ~n9362 & ~n13908;
  assign n13910 = ~n11639 & ~n13233;
  assign n13911 = n13907 & ~n13909;
  assign n13912 = n13910 & n13911;
  assign n13913 = ~n13902 & ~n13912;
  assign n13914 = n13905 & ~n13913;
  assign n13915 = P2_STATE_REG & ~n13914;
  assign n13916 = ~n13903 & ~n13915;
  assign n13917 = ~n10436 & ~n13916;
  assign n13918 = n13900 & n13902;
  assign n13919 = n9303 & n11640;
  assign n13920 = ~n13918 & ~n13919;
  assign n13921 = ~n10520 & ~n13920;
  assign n13922 = P2_STATE_REG & n13258;
  assign n13923 = ~n9301 & n13922;
  assign n13924 = n9445 & n13902;
  assign n13925 = ~n10513 & n13924;
  assign n13926 = ~n9445 & n13902;
  assign n13927 = ~n10374 & n13926;
  assign n13928 = ~n10436 & ~n13902;
  assign n13929 = ~n13925 & ~n13927;
  assign n13930 = ~n13928 & n13929;
  assign n13931 = n13923 & ~n13930;
  assign n13932 = ~n13206 & ~n13891;
  assign n13933 = ~n13146 & n13932;
  assign n13934 = n12262 & n13933;
  assign n13935 = ~n10084 & ~n13934;
  assign n13936 = ~n9362 & ~n9365;
  assign n13937 = ~n13145 & ~n13936;
  assign n13938 = ~n9450 & n13937;
  assign n13939 = ~n10163 & n13938;
  assign n13940 = n10163 & ~n13938;
  assign n13941 = ~n13939 & ~n13940;
  assign n13942 = n13935 & ~n13941;
  assign n13943 = ~n10309 & n13938;
  assign n13944 = n10309 & ~n13938;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = ~n10227 & ~n13934;
  assign n13947 = n13945 & ~n13946;
  assign n13948 = ~n10381 & n13938;
  assign n13949 = n10381 & ~n13938;
  assign n13950 = ~n13948 & ~n13949;
  assign n13951 = ~n10302 & ~n13934;
  assign n13952 = n13950 & ~n13951;
  assign n13953 = ~n13947 & ~n13952;
  assign n13954 = ~n10234 & n13938;
  assign n13955 = n10234 & ~n13938;
  assign n13956 = ~n13954 & ~n13955;
  assign n13957 = ~n10156 & ~n13934;
  assign n13958 = n13956 & ~n13957;
  assign n13959 = n13953 & ~n13958;
  assign n13960 = n13942 & n13959;
  assign n13961 = ~n13950 & n13951;
  assign n13962 = ~n13945 & n13946;
  assign n13963 = ~n13961 & ~n13962;
  assign n13964 = ~n13956 & n13957;
  assign n13965 = n13953 & n13964;
  assign n13966 = n13963 & ~n13965;
  assign n13967 = ~n13952 & ~n13966;
  assign n13968 = ~n13960 & ~n13967;
  assign n13969 = ~n10450 & n13938;
  assign n13970 = n10450 & ~n13938;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = ~n10374 & ~n13934;
  assign n13973 = n13971 & ~n13972;
  assign n13974 = ~n13968 & ~n13973;
  assign n13975 = ~n13971 & n13972;
  assign n13976 = ~n13974 & ~n13975;
  assign n13977 = ~n13935 & n13941;
  assign n13978 = n13959 & ~n13977;
  assign n13979 = ~n13973 & n13978;
  assign n13980 = ~n10010 & ~n13934;
  assign n13981 = ~n9852 & ~n13934;
  assign n13982 = ~n9788 & ~n13934;
  assign n13983 = ~n9859 & n13938;
  assign n13984 = n9859 & ~n13938;
  assign n13985 = ~n13983 & ~n13984;
  assign n13986 = n13982 & ~n13985;
  assign n13987 = n13981 & n13986;
  assign n13988 = ~n9943 & n13938;
  assign n13989 = n9943 & ~n13938;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = ~n13981 & ~n13986;
  assign n13992 = ~n13990 & ~n13991;
  assign n13993 = ~n9717 & ~n13934;
  assign n13994 = ~n9795 & n13938;
  assign n13995 = n9795 & ~n13938;
  assign n13996 = ~n13994 & ~n13995;
  assign n13997 = n13993 & ~n13996;
  assign n13998 = ~n13982 & n13985;
  assign n13999 = ~n13981 & n13990;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = n13997 & n14000;
  assign n14002 = ~n13987 & ~n13992;
  assign n14003 = ~n14001 & n14002;
  assign n14004 = ~n10017 & n13938;
  assign n14005 = n10017 & ~n13938;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = ~n9936 & ~n13934;
  assign n14008 = n14006 & ~n14007;
  assign n14009 = ~n14003 & ~n14008;
  assign n14010 = ~n14006 & n14007;
  assign n14011 = ~n14009 & ~n14010;
  assign n14012 = ~n13993 & n13996;
  assign n14013 = n14000 & ~n14012;
  assign n14014 = ~n14008 & n14013;
  assign n14015 = ~n9651 & ~n13934;
  assign n14016 = ~n9586 & ~n13934;
  assign n14017 = ~n9530 & ~n13934;
  assign n14018 = ~n9593 & n13938;
  assign n14019 = n9593 & ~n13938;
  assign n14020 = ~n14018 & ~n14019;
  assign n14021 = n14017 & ~n14020;
  assign n14022 = n14016 & n14021;
  assign n14023 = ~n9658 & n13938;
  assign n14024 = n9658 & ~n13938;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = ~n14016 & ~n14021;
  assign n14027 = ~n14025 & ~n14026;
  assign n14028 = ~n14022 & ~n14027;
  assign n14029 = ~n14017 & n14020;
  assign n14030 = ~n14016 & n14025;
  assign n14031 = ~n14029 & ~n14030;
  assign n14032 = ~n9449 & n13938;
  assign n14033 = n9449 & ~n13938;
  assign n14034 = ~n14032 & ~n14033;
  assign n14035 = ~n13938 & ~n14034;
  assign n14036 = ~n9537 & n13938;
  assign n14037 = n9537 & ~n13938;
  assign n14038 = ~n14036 & ~n14037;
  assign n14039 = ~n9475 & ~n13934;
  assign n14040 = n14038 & ~n14039;
  assign n14041 = n14035 & ~n14040;
  assign n14042 = ~n14038 & n14039;
  assign n14043 = ~n9483 & ~n13934;
  assign n14044 = n13938 & n14034;
  assign n14045 = n14043 & ~n14044;
  assign n14046 = ~n14040 & n14045;
  assign n14047 = ~n14041 & ~n14042;
  assign n14048 = ~n14046 & n14047;
  assign n14049 = n14031 & ~n14048;
  assign n14050 = n14028 & ~n14049;
  assign n14051 = n14015 & ~n14050;
  assign n14052 = ~n9724 & n13938;
  assign n14053 = n9724 & ~n13938;
  assign n14054 = ~n14052 & ~n14053;
  assign n14055 = ~n14050 & ~n14054;
  assign n14056 = n14015 & ~n14054;
  assign n14057 = ~n14051 & ~n14055;
  assign n14058 = ~n14056 & n14057;
  assign n14059 = n14014 & ~n14058;
  assign n14060 = n14011 & ~n14059;
  assign n14061 = n13980 & ~n14060;
  assign n14062 = ~n10091 & n13938;
  assign n14063 = n10091 & ~n13938;
  assign n14064 = ~n14062 & ~n14063;
  assign n14065 = ~n14060 & ~n14064;
  assign n14066 = n13980 & ~n14064;
  assign n14067 = ~n14061 & ~n14065;
  assign n14068 = ~n14066 & n14067;
  assign n14069 = n13979 & ~n14068;
  assign n14070 = n13976 & ~n14069;
  assign n14071 = ~n10520 & n13938;
  assign n14072 = n10520 & ~n13938;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = ~n10443 & ~n13934;
  assign n14075 = ~n14073 & ~n14074;
  assign n14076 = n14073 & n14074;
  assign n14077 = ~n14075 & ~n14076;
  assign n14078 = n14070 & ~n14077;
  assign n14079 = ~n14070 & n14077;
  assign n14080 = ~n14078 & ~n14079;
  assign n14081 = n9303 & ~n13912;
  assign n14082 = n13902 & n14081;
  assign n14083 = ~n14080 & n14082;
  assign n14084 = ~n13917 & ~n13921;
  assign n14085 = ~n12436 & n14084;
  assign n14086 = ~n13931 & n14085;
  assign n2400 = n14083 | ~n14086;
  assign n14088 = P2_REG3_REG_26_ & ~P2_STATE_REG;
  assign n14089 = ~n11190 & ~n13902;
  assign n14090 = ~n11125 & n13926;
  assign n14091 = ~n11256 & n13924;
  assign n14092 = ~n14089 & ~n14090;
  assign n14093 = ~n14091 & n14092;
  assign n14094 = n13923 & ~n14093;
  assign n14095 = ~n11650 & ~n13902;
  assign n14096 = n13914 & ~n14095;
  assign n14097 = P2_STATE_REG & ~n14096;
  assign n14098 = ~n11190 & n14097;
  assign n14099 = ~n11650 & n13902;
  assign n14100 = ~n11640 & ~n14099;
  assign n14101 = n9303 & ~n14100;
  assign n14102 = n11258 & n14101;
  assign n14103 = ~n11194 & ~n13934;
  assign n14104 = n11258 & n13938;
  assign n14105 = ~n11258 & ~n13938;
  assign n14106 = ~n14104 & ~n14105;
  assign n14107 = n14103 & ~n14106;
  assign n14108 = n11196 & n13938;
  assign n14109 = ~n11196 & ~n13938;
  assign n14110 = ~n14108 & ~n14109;
  assign n14111 = ~n11125 & ~n13934;
  assign n14112 = n14110 & ~n14111;
  assign n14113 = n14103 & ~n14112;
  assign n14114 = ~n14106 & ~n14112;
  assign n14115 = ~n14113 & ~n14114;
  assign n14116 = ~n14107 & ~n14115;
  assign n14117 = ~n11061 & ~n13934;
  assign n14118 = n11127 & n13938;
  assign n14119 = ~n11127 & ~n13938;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = n14117 & ~n14120;
  assign n14122 = ~n14110 & n14111;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = ~n14117 & n14120;
  assign n14125 = ~n10992 & ~n13934;
  assign n14126 = n11063 & n13938;
  assign n14127 = ~n11063 & ~n13938;
  assign n14128 = ~n14126 & ~n14127;
  assign n14129 = n14125 & ~n14128;
  assign n14130 = ~n14125 & n14128;
  assign n14131 = ~n10928 & ~n13934;
  assign n14132 = n10994 & n13938;
  assign n14133 = ~n10994 & ~n13938;
  assign n14134 = ~n14132 & ~n14133;
  assign n14135 = n14131 & ~n14134;
  assign n14136 = ~n14131 & n14134;
  assign n14137 = n10930 & n13938;
  assign n14138 = ~n10930 & ~n13938;
  assign n14139 = ~n14137 & ~n14138;
  assign n14140 = ~n10863 & ~n13934;
  assign n14141 = n14139 & ~n14140;
  assign n14142 = ~n14139 & n14140;
  assign n14143 = ~n10797 & ~n13934;
  assign n14144 = n10865 & n13938;
  assign n14145 = ~n10865 & ~n13938;
  assign n14146 = ~n14144 & ~n14145;
  assign n14147 = n14143 & ~n14146;
  assign n14148 = ~n14142 & ~n14147;
  assign n14149 = ~n10725 & ~n13934;
  assign n14150 = ~n10801 & n13938;
  assign n14151 = n10801 & ~n13938;
  assign n14152 = ~n14150 & ~n14151;
  assign n14153 = n14149 & ~n14152;
  assign n14154 = ~n14143 & n14146;
  assign n14155 = ~n14141 & ~n14154;
  assign n14156 = n14153 & n14155;
  assign n14157 = n14148 & ~n14156;
  assign n14158 = ~n14141 & ~n14157;
  assign n14159 = ~n14149 & n14152;
  assign n14160 = n14155 & ~n14159;
  assign n14161 = ~n10651 & ~n13934;
  assign n14162 = ~n10732 & n13938;
  assign n14163 = n10732 & ~n13938;
  assign n14164 = ~n14162 & ~n14163;
  assign n14165 = n14161 & ~n14164;
  assign n14166 = ~n14161 & n14164;
  assign n14167 = ~n10579 & ~n13934;
  assign n14168 = ~n10513 & ~n13934;
  assign n14169 = ~n10586 & n13938;
  assign n14170 = n10586 & ~n13938;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = n14168 & ~n14171;
  assign n14173 = n14167 & n14172;
  assign n14174 = ~n10658 & n13938;
  assign n14175 = n10658 & ~n13938;
  assign n14176 = ~n14174 & ~n14175;
  assign n14177 = ~n14167 & ~n14172;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = ~n14173 & ~n14178;
  assign n14180 = ~n14168 & n14171;
  assign n14181 = ~n14167 & n14176;
  assign n14182 = ~n14180 & ~n14181;
  assign n14183 = ~n14073 & n14074;
  assign n14184 = n14073 & ~n14074;
  assign n14185 = ~n14070 & ~n14184;
  assign n14186 = ~n14183 & ~n14185;
  assign n14187 = n14182 & ~n14186;
  assign n14188 = n14179 & ~n14187;
  assign n14189 = ~n14166 & ~n14188;
  assign n14190 = ~n14165 & ~n14189;
  assign n14191 = n14160 & ~n14190;
  assign n14192 = ~n14158 & ~n14191;
  assign n14193 = ~n14136 & ~n14192;
  assign n14194 = ~n14135 & ~n14193;
  assign n14195 = ~n14130 & ~n14194;
  assign n14196 = ~n14129 & ~n14195;
  assign n14197 = ~n14124 & ~n14196;
  assign n14198 = n14123 & ~n14197;
  assign n14199 = n14116 & ~n14198;
  assign n14200 = ~n14103 & ~n14106;
  assign n14201 = n14103 & n14106;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = n14112 & n14202;
  assign n14204 = ~n14122 & n14202;
  assign n14205 = ~n14121 & ~n14197;
  assign n14206 = n14204 & n14205;
  assign n14207 = ~n14199 & ~n14203;
  assign n14208 = ~n14206 & n14207;
  assign n14209 = n14082 & n14208;
  assign n14210 = ~n14088 & ~n14094;
  assign n14211 = ~n14098 & n14210;
  assign n14212 = ~n14102 & n14211;
  assign n2405 = n14209 | ~n14212;
  assign n14214 = ~n9852 & n13924;
  assign n14215 = ~n9717 & n13926;
  assign n14216 = ~n9781 & ~n13902;
  assign n14217 = ~n14214 & ~n14215;
  assign n14218 = ~n14216 & n14217;
  assign n14219 = n13923 & ~n14218;
  assign n14220 = ~n13982 & ~n13985;
  assign n14221 = n13982 & n13985;
  assign n14222 = ~n14220 & ~n14221;
  assign n14223 = ~n14012 & ~n14058;
  assign n14224 = ~n13997 & ~n14223;
  assign n14225 = ~n14222 & n14224;
  assign n14226 = ~n13986 & ~n13998;
  assign n14227 = ~n14224 & ~n14226;
  assign n14228 = ~n14225 & ~n14227;
  assign n14229 = n14082 & ~n14228;
  assign n14230 = ~n9859 & ~n13920;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = ~n9781 & ~n13916;
  assign n14233 = ~n12792 & ~n14219;
  assign n14234 = n14231 & n14233;
  assign n2410 = n14232 | ~n14234;
  assign n14236 = ~n10647 & ~n13916;
  assign n14237 = ~n10732 & ~n13920;
  assign n14238 = ~n10725 & n13924;
  assign n14239 = ~n10579 & n13926;
  assign n14240 = ~n10647 & ~n13902;
  assign n14241 = ~n14238 & ~n14239;
  assign n14242 = ~n14240 & n14241;
  assign n14243 = n13923 & ~n14242;
  assign n14244 = ~n14161 & ~n14164;
  assign n14245 = n14161 & n14164;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = n14188 & ~n14246;
  assign n14248 = ~n14188 & n14246;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = n14082 & ~n14249;
  assign n14251 = ~n14236 & ~n14237;
  assign n14252 = ~n12319 & n14251;
  assign n14253 = ~n14243 & n14252;
  assign n2415 = n14250 | ~n14253;
  assign n14255 = ~n9586 & n13924;
  assign n14256 = ~n9475 & n13926;
  assign n14257 = P2_REG3_REG_2_ & ~n13902;
  assign n14258 = ~n14255 & ~n14256;
  assign n14259 = ~n14257 & n14258;
  assign n14260 = n13923 & ~n14259;
  assign n14261 = ~n14017 & ~n14020;
  assign n14262 = n14017 & n14020;
  assign n14263 = ~n14261 & ~n14262;
  assign n14264 = n14048 & ~n14263;
  assign n14265 = ~n14021 & ~n14029;
  assign n14266 = ~n14048 & ~n14265;
  assign n14267 = ~n14264 & ~n14266;
  assign n14268 = n14082 & ~n14267;
  assign n14269 = ~n9593 & ~n13920;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = P2_REG3_REG_2_ & ~n13916;
  assign n14272 = ~n12966 & ~n14260;
  assign n14273 = n14270 & n14272;
  assign n2420 = n14271 | ~n14273;
  assign n14275 = ~n10149 & ~n13916;
  assign n14276 = ~n10234 & ~n13920;
  assign n14277 = ~n13977 & ~n14068;
  assign n14278 = ~n13942 & ~n14277;
  assign n14279 = ~n13956 & ~n13957;
  assign n14280 = n13956 & n13957;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = n14278 & ~n14281;
  assign n14283 = ~n13958 & ~n13964;
  assign n14284 = ~n14278 & ~n14283;
  assign n14285 = ~n14282 & ~n14284;
  assign n14286 = n14082 & ~n14285;
  assign n14287 = ~n10227 & n13924;
  assign n14288 = ~n10084 & n13926;
  assign n14289 = ~n10149 & ~n13902;
  assign n14290 = ~n14287 & ~n14288;
  assign n14291 = ~n14289 & n14290;
  assign n14292 = n13923 & ~n14291;
  assign n14293 = ~n14275 & ~n14276;
  assign n14294 = ~n14286 & n14293;
  assign n14295 = ~n12592 & n14294;
  assign n2425 = n14292 | ~n14295;
  assign n14297 = P2_REG3_REG_22_ & ~P2_STATE_REG;
  assign n14298 = ~n10992 & n13924;
  assign n14299 = ~n10863 & n13926;
  assign n14300 = ~n10924 & ~n13902;
  assign n14301 = ~n14298 & ~n14299;
  assign n14302 = ~n14300 & n14301;
  assign n14303 = n13923 & ~n14302;
  assign n14304 = ~n10924 & n14097;
  assign n14305 = n10994 & n14101;
  assign n14306 = ~n14131 & ~n14134;
  assign n14307 = n14131 & n14134;
  assign n14308 = ~n14306 & ~n14307;
  assign n14309 = n14192 & ~n14308;
  assign n14310 = ~n14192 & n14308;
  assign n14311 = ~n14309 & ~n14310;
  assign n14312 = n14082 & ~n14311;
  assign n14313 = ~n14297 & ~n14303;
  assign n14314 = ~n14304 & n14313;
  assign n14315 = ~n14305 & n14314;
  assign n2430 = n14312 | ~n14315;
  assign n14317 = ~n10295 & ~n13916;
  assign n14318 = ~n10381 & ~n13920;
  assign n14319 = ~n10374 & n13924;
  assign n14320 = ~n10227 & n13926;
  assign n14321 = ~n10295 & ~n13902;
  assign n14322 = ~n14319 & ~n14320;
  assign n14323 = ~n14321 & n14322;
  assign n14324 = n13923 & ~n14323;
  assign n14325 = n13953 & ~n13961;
  assign n14326 = ~n13958 & ~n14278;
  assign n14327 = ~n13964 & ~n14326;
  assign n14328 = ~n13962 & n14327;
  assign n14329 = n14325 & ~n14328;
  assign n14330 = ~n13950 & ~n13951;
  assign n14331 = n13950 & n13951;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = ~n13962 & n14332;
  assign n14334 = ~n13947 & ~n14327;
  assign n14335 = n14333 & ~n14334;
  assign n14336 = ~n14329 & ~n14335;
  assign n14337 = n14082 & n14336;
  assign n14338 = ~n14317 & ~n14318;
  assign n14339 = ~n12518 & n14338;
  assign n14340 = ~n14324 & n14339;
  assign n2435 = n14337 | ~n14340;
  assign n14342 = ~n10793 & n14097;
  assign n14343 = n10865 & n14101;
  assign n14344 = P2_REG3_REG_20_ & ~P2_STATE_REG;
  assign n14345 = ~n10863 & n13924;
  assign n14346 = ~n10725 & n13926;
  assign n14347 = ~n10793 & ~n13902;
  assign n14348 = ~n14345 & ~n14346;
  assign n14349 = ~n14347 & n14348;
  assign n14350 = n13923 & ~n14349;
  assign n14351 = ~n14143 & ~n14146;
  assign n14352 = n14143 & n14146;
  assign n14353 = ~n14351 & ~n14352;
  assign n14354 = ~n14159 & ~n14190;
  assign n14355 = ~n14153 & ~n14354;
  assign n14356 = ~n14353 & n14355;
  assign n14357 = ~n14147 & ~n14154;
  assign n14358 = ~n14355 & ~n14357;
  assign n14359 = ~n14356 & ~n14358;
  assign n14360 = n14082 & ~n14359;
  assign n14361 = ~n14342 & ~n14343;
  assign n14362 = ~n14344 & n14361;
  assign n14363 = ~n14350 & n14362;
  assign n2440 = n14360 | ~n14363;
  assign n14365 = ~n13938 & n14034;
  assign n14366 = n13938 & ~n14034;
  assign n14367 = ~n14365 & ~n14366;
  assign n14368 = ~n14043 & ~n14367;
  assign n14369 = n14043 & n14367;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = n14082 & ~n14370;
  assign n14372 = ~n13026 & ~n14371;
  assign n14373 = ~n13900 & ~n13923;
  assign n14374 = ~n13902 & ~n14373;
  assign n14375 = ~n13915 & ~n14374;
  assign n14376 = P2_REG3_REG_0_ & ~n14375;
  assign n14377 = ~n9449 & ~n13920;
  assign n14378 = ~n9475 & n13923;
  assign n14379 = n13924 & n14378;
  assign n14380 = ~n14377 & ~n14379;
  assign n14381 = n14372 & ~n14376;
  assign n2445 = ~n14380 | ~n14381;
  assign n14383 = ~n10003 & ~n13916;
  assign n14384 = ~n10091 & ~n13920;
  assign n14385 = ~n13980 & ~n14064;
  assign n14386 = n13980 & n14064;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = n14060 & ~n14387;
  assign n14389 = ~n14060 & n14387;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = n14082 & ~n14390;
  assign n14392 = ~n10084 & n13924;
  assign n14393 = ~n9936 & n13926;
  assign n14394 = ~n10003 & ~n13902;
  assign n14395 = ~n14392 & ~n14393;
  assign n14396 = ~n14394 & n14395;
  assign n14397 = n13923 & ~n14396;
  assign n14398 = ~n14383 & ~n14384;
  assign n14399 = ~n14391 & n14398;
  assign n14400 = ~n12676 & n14399;
  assign n2450 = n14397 | ~n14400;
  assign n14402 = ~n9717 & n13924;
  assign n14403 = ~n9586 & n13926;
  assign n14404 = ~n9644 & ~n13902;
  assign n14405 = ~n14402 & ~n14403;
  assign n14406 = ~n14404 & n14405;
  assign n14407 = n13923 & ~n14406;
  assign n14408 = ~n14015 & ~n14054;
  assign n14409 = n14015 & n14054;
  assign n14410 = ~n14408 & ~n14409;
  assign n14411 = n14050 & ~n14410;
  assign n14412 = ~n14050 & n14410;
  assign n14413 = ~n14411 & ~n14412;
  assign n14414 = n14082 & ~n14413;
  assign n14415 = ~n9724 & ~n13920;
  assign n14416 = ~n14414 & ~n14415;
  assign n14417 = ~n9644 & ~n13916;
  assign n14418 = ~n12886 & ~n14407;
  assign n14419 = n14416 & n14418;
  assign n2455 = n14417 | ~n14419;
  assign n14421 = P2_REG3_REG_24_ & ~P2_STATE_REG;
  assign n14422 = ~n11125 & n13924;
  assign n14423 = ~n10992 & n13926;
  assign n14424 = ~n11057 & ~n13902;
  assign n14425 = ~n14422 & ~n14423;
  assign n14426 = ~n14424 & n14425;
  assign n14427 = n13923 & ~n14426;
  assign n14428 = ~n11057 & n14097;
  assign n14429 = n11127 & n14101;
  assign n14430 = ~n14117 & ~n14120;
  assign n14431 = n14117 & n14120;
  assign n14432 = ~n14430 & ~n14431;
  assign n14433 = n14196 & ~n14432;
  assign n14434 = ~n14121 & ~n14124;
  assign n14435 = ~n14196 & ~n14434;
  assign n14436 = ~n14433 & ~n14435;
  assign n14437 = n14082 & ~n14436;
  assign n14438 = ~n14421 & ~n14427;
  assign n14439 = ~n14428 & n14438;
  assign n14440 = ~n14429 & n14439;
  assign n2460 = n14437 | ~n14440;
  assign n14442 = ~n10575 & ~n13916;
  assign n14443 = ~n10658 & ~n13920;
  assign n14444 = ~n10651 & n13924;
  assign n14445 = ~n10513 & n13926;
  assign n14446 = ~n10575 & ~n13902;
  assign n14447 = ~n14444 & ~n14445;
  assign n14448 = ~n14446 & n14447;
  assign n14449 = n13923 & ~n14448;
  assign n14450 = n14167 & ~n14176;
  assign n14451 = n14182 & ~n14450;
  assign n14452 = ~n14172 & n14186;
  assign n14453 = n14451 & ~n14452;
  assign n14454 = ~n14167 & ~n14176;
  assign n14455 = n14167 & n14176;
  assign n14456 = ~n14454 & ~n14455;
  assign n14457 = ~n14172 & n14456;
  assign n14458 = ~n14180 & ~n14186;
  assign n14459 = n14457 & ~n14458;
  assign n14460 = ~n14453 & ~n14459;
  assign n14461 = n14082 & n14460;
  assign n14462 = ~n14442 & ~n14443;
  assign n14463 = ~n12364 & n14462;
  assign n14464 = ~n14449 & n14463;
  assign n2465 = n14461 | ~n14464;
  assign n14466 = ~n9788 & n13924;
  assign n14467 = ~n9651 & n13926;
  assign n14468 = ~n9710 & ~n13902;
  assign n14469 = ~n14466 & ~n14467;
  assign n14470 = ~n14468 & n14469;
  assign n14471 = n13923 & ~n14470;
  assign n14472 = ~n13993 & ~n13996;
  assign n14473 = n13993 & n13996;
  assign n14474 = ~n14472 & ~n14473;
  assign n14475 = n14058 & ~n14474;
  assign n14476 = ~n14058 & n14474;
  assign n14477 = ~n14475 & ~n14476;
  assign n14478 = n14082 & ~n14477;
  assign n14479 = ~n9795 & ~n13920;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481 = ~n9710 & ~n13916;
  assign n14482 = ~n12849 & ~n14471;
  assign n14483 = n14480 & n14482;
  assign n2470 = n14481 | ~n14483;
  assign n14485 = ~n10506 & ~n13916;
  assign n14486 = ~n10586 & ~n13920;
  assign n14487 = ~n10579 & n13924;
  assign n14488 = ~n10443 & n13926;
  assign n14489 = ~n10506 & ~n13902;
  assign n14490 = ~n14487 & ~n14488;
  assign n14491 = ~n14489 & n14490;
  assign n14492 = n13923 & ~n14491;
  assign n14493 = ~n14168 & ~n14171;
  assign n14494 = n14168 & n14171;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = n14186 & ~n14495;
  assign n14497 = ~n14172 & ~n14180;
  assign n14498 = ~n14186 & ~n14497;
  assign n14499 = ~n14496 & ~n14498;
  assign n14500 = n14082 & ~n14499;
  assign n14501 = ~n14485 & ~n14486;
  assign n14502 = ~n12401 & n14501;
  assign n14503 = ~n14492 & n14502;
  assign n2475 = n14500 | ~n14503;
  assign n14505 = P2_REG3_REG_25_ & ~P2_STATE_REG;
  assign n14506 = ~n11194 & n13924;
  assign n14507 = ~n11061 & n13926;
  assign n14508 = ~n11121 & ~n13902;
  assign n14509 = ~n14506 & ~n14507;
  assign n14510 = ~n14508 & n14509;
  assign n14511 = n13923 & ~n14510;
  assign n14512 = ~n11121 & n14097;
  assign n14513 = n11196 & n14101;
  assign n14514 = ~n14110 & ~n14111;
  assign n14515 = n14110 & n14111;
  assign n14516 = ~n14514 & ~n14515;
  assign n14517 = n14205 & ~n14516;
  assign n14518 = ~n14112 & ~n14122;
  assign n14519 = ~n14205 & ~n14518;
  assign n14520 = ~n14517 & ~n14519;
  assign n14521 = n14082 & ~n14520;
  assign n14522 = ~n14505 & ~n14511;
  assign n14523 = ~n14512 & n14522;
  assign n14524 = ~n14513 & n14523;
  assign n2480 = n14521 | ~n14524;
  assign n14526 = ~n10220 & ~n13916;
  assign n14527 = ~n10309 & ~n13920;
  assign n14528 = ~n10302 & n13924;
  assign n14529 = ~n10156 & n13926;
  assign n14530 = ~n10220 & ~n13902;
  assign n14531 = ~n14528 & ~n14529;
  assign n14532 = ~n14530 & n14531;
  assign n14533 = n13923 & ~n14532;
  assign n14534 = ~n13945 & ~n13946;
  assign n14535 = n13945 & n13946;
  assign n14536 = ~n14534 & ~n14535;
  assign n14537 = n14327 & ~n14536;
  assign n14538 = ~n13947 & ~n13962;
  assign n14539 = ~n14327 & ~n14538;
  assign n14540 = ~n14537 & ~n14539;
  assign n14541 = n14082 & ~n14540;
  assign n14542 = ~n14526 & ~n14527;
  assign n14543 = ~n12555 & n14542;
  assign n14544 = ~n14533 & n14543;
  assign n2485 = n14541 | ~n14544;
  assign n14546 = ~n10859 & n14097;
  assign n14547 = n10930 & n14101;
  assign n14548 = P2_REG3_REG_21_ & ~P2_STATE_REG;
  assign n14549 = ~n10928 & n13924;
  assign n14550 = ~n10797 & n13926;
  assign n14551 = ~n10859 & ~n13902;
  assign n14552 = ~n14549 & ~n14550;
  assign n14553 = ~n14551 & n14552;
  assign n14554 = n13923 & ~n14553;
  assign n14555 = ~n14142 & n14155;
  assign n14556 = ~n14147 & n14355;
  assign n14557 = n14555 & ~n14556;
  assign n14558 = ~n14139 & ~n14140;
  assign n14559 = n14139 & n14140;
  assign n14560 = ~n14558 & ~n14559;
  assign n14561 = ~n14147 & n14560;
  assign n14562 = ~n14154 & ~n14355;
  assign n14563 = n14561 & ~n14562;
  assign n14564 = ~n14557 & ~n14563;
  assign n14565 = n14082 & n14564;
  assign n14566 = ~n14546 & ~n14547;
  assign n14567 = ~n14548 & n14566;
  assign n14568 = ~n14554 & n14567;
  assign n2490 = n14565 | ~n14568;
  assign n14570 = ~n9530 & n13924;
  assign n14571 = ~n9483 & n13926;
  assign n14572 = P2_REG3_REG_1_ & ~n13902;
  assign n14573 = ~n14570 & ~n14571;
  assign n14574 = ~n14572 & n14573;
  assign n14575 = n13923 & ~n14574;
  assign n14576 = ~n14035 & ~n14045;
  assign n14577 = ~n14038 & ~n14039;
  assign n14578 = n14038 & n14039;
  assign n14579 = ~n14577 & ~n14578;
  assign n14580 = n14576 & ~n14579;
  assign n14581 = ~n14576 & n14579;
  assign n14582 = ~n14580 & ~n14581;
  assign n14583 = n14082 & ~n14582;
  assign n14584 = ~n9537 & ~n13920;
  assign n14585 = ~n14583 & ~n14584;
  assign n14586 = P2_REG3_REG_1_ & ~n13916;
  assign n14587 = ~n12997 & ~n14575;
  assign n14588 = n14585 & n14587;
  assign n2495 = n14586 | ~n14588;
  assign n14590 = ~n10010 & n13924;
  assign n14591 = ~n9852 & n13926;
  assign n14592 = ~n9929 & ~n13902;
  assign n14593 = ~n14590 & ~n14591;
  assign n14594 = ~n14592 & n14593;
  assign n14595 = n13923 & ~n14594;
  assign n14596 = n14013 & ~n14058;
  assign n14597 = n14003 & ~n14596;
  assign n14598 = ~n14006 & ~n14007;
  assign n14599 = n14006 & n14007;
  assign n14600 = ~n14598 & ~n14599;
  assign n14601 = n14597 & ~n14600;
  assign n14602 = ~n14597 & n14600;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = n14082 & ~n14603;
  assign n14605 = ~n10017 & ~n13920;
  assign n14606 = ~n14604 & ~n14605;
  assign n14607 = ~n9929 & ~n13916;
  assign n14608 = ~n12710 & ~n14595;
  assign n14609 = n14606 & n14608;
  assign n2500 = n14607 | ~n14609;
  assign n14611 = P2_REG3_REG_28_ & ~P2_STATE_REG;
  assign n14612 = ~n11386 & n13924;
  assign n14613 = ~n11319 & ~n13902;
  assign n14614 = ~n11256 & n13926;
  assign n14615 = ~n14612 & ~n14613;
  assign n14616 = ~n14614 & n14615;
  assign n14617 = n13923 & ~n14616;
  assign n14618 = ~n11319 & n14097;
  assign n14619 = n11388 & n14101;
  assign n14620 = n11325 & n13938;
  assign n14621 = ~n11325 & ~n13938;
  assign n14622 = ~n14620 & ~n14621;
  assign n14623 = ~n11256 & ~n13934;
  assign n14624 = n14622 & ~n14623;
  assign n14625 = ~n14107 & n14123;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = ~n14107 & ~n14114;
  assign n14628 = ~n14113 & n14627;
  assign n14629 = n14626 & ~n14628;
  assign n14630 = ~n14622 & n14623;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~n14124 & ~n14624;
  assign n14633 = ~n14115 & ~n14196;
  assign n14634 = n14632 & n14633;
  assign n14635 = n11388 & n13938;
  assign n14636 = ~n11388 & ~n13938;
  assign n14637 = ~n14635 & ~n14636;
  assign n14638 = ~n11323 & ~n13934;
  assign n14639 = ~n14637 & ~n14638;
  assign n14640 = n14637 & n14638;
  assign n14641 = ~n14639 & ~n14640;
  assign n14642 = n14631 & ~n14634;
  assign n14643 = ~n14641 & n14642;
  assign n14644 = ~n14115 & ~n14124;
  assign n14645 = ~n14196 & n14644;
  assign n14646 = ~n14103 & n14106;
  assign n14647 = ~n14112 & ~n14123;
  assign n14648 = ~n14646 & n14647;
  assign n14649 = ~n14630 & ~n14648;
  assign n14650 = ~n14107 & ~n14645;
  assign n14651 = n14649 & n14650;
  assign n14652 = ~n14624 & ~n14651;
  assign n14653 = n14641 & n14652;
  assign n14654 = ~n14643 & ~n14653;
  assign n14655 = n14082 & ~n14654;
  assign n14656 = ~n14611 & ~n14617;
  assign n14657 = ~n14618 & n14656;
  assign n14658 = ~n14619 & n14657;
  assign n2505 = n14655 | ~n14658;
  assign n14660 = ~n10721 & ~n13916;
  assign n14661 = ~n10801 & ~n13920;
  assign n14662 = ~n10797 & n13924;
  assign n14663 = ~n10651 & n13926;
  assign n14664 = ~n10721 & ~n13902;
  assign n14665 = ~n14662 & ~n14663;
  assign n14666 = ~n14664 & n14665;
  assign n14667 = n13923 & ~n14666;
  assign n14668 = ~n14149 & ~n14152;
  assign n14669 = n14149 & n14152;
  assign n14670 = ~n14668 & ~n14669;
  assign n14671 = n14190 & ~n14670;
  assign n14672 = ~n14153 & ~n14159;
  assign n14673 = ~n14190 & ~n14672;
  assign n14674 = ~n14671 & ~n14673;
  assign n14675 = n14082 & ~n14674;
  assign n14676 = ~n14660 & ~n14661;
  assign n14677 = ~n12283 & n14676;
  assign n14678 = ~n14667 & n14677;
  assign n2510 = n14675 | ~n14678;
  assign n14680 = ~n9651 & n13924;
  assign n14681 = ~n9530 & n13926;
  assign n14682 = ~P2_REG3_REG_3_ & ~n13902;
  assign n14683 = ~n14680 & ~n14681;
  assign n14684 = ~n14682 & n14683;
  assign n14685 = n13923 & ~n14684;
  assign n14686 = n14016 & ~n14025;
  assign n14687 = n14031 & ~n14686;
  assign n14688 = ~n14021 & n14048;
  assign n14689 = n14687 & ~n14688;
  assign n14690 = ~n14016 & ~n14025;
  assign n14691 = n14016 & n14025;
  assign n14692 = ~n14690 & ~n14691;
  assign n14693 = ~n14021 & n14692;
  assign n14694 = ~n14029 & ~n14048;
  assign n14695 = n14693 & ~n14694;
  assign n14696 = ~n14689 & ~n14695;
  assign n14697 = n14082 & n14696;
  assign n14698 = ~n9658 & ~n13920;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = ~P2_REG3_REG_3_ & ~n13916;
  assign n14701 = ~n12927 & ~n14685;
  assign n14702 = n14699 & n14701;
  assign n2515 = n14700 | ~n14702;
  assign n14704 = ~n10077 & ~n13916;
  assign n14705 = ~n10163 & ~n13920;
  assign n14706 = ~n13935 & ~n13941;
  assign n14707 = n13935 & n13941;
  assign n14708 = ~n14706 & ~n14707;
  assign n14709 = n14068 & ~n14708;
  assign n14710 = ~n14068 & n14708;
  assign n14711 = ~n14709 & ~n14710;
  assign n14712 = n14082 & ~n14711;
  assign n14713 = ~n10156 & n13924;
  assign n14714 = ~n10010 & n13926;
  assign n14715 = ~n10077 & ~n13902;
  assign n14716 = ~n14713 & ~n14714;
  assign n14717 = ~n14715 & n14716;
  assign n14718 = n13923 & ~n14717;
  assign n14719 = ~n14704 & ~n14705;
  assign n14720 = ~n14712 & n14719;
  assign n14721 = ~n12639 & n14720;
  assign n2520 = n14718 | ~n14721;
  assign n14723 = P2_REG3_REG_23_ & ~P2_STATE_REG;
  assign n14724 = ~n11061 & n13924;
  assign n14725 = ~n10928 & n13926;
  assign n14726 = ~n10988 & ~n13902;
  assign n14727 = ~n14724 & ~n14725;
  assign n14728 = ~n14726 & n14727;
  assign n14729 = n13923 & ~n14728;
  assign n14730 = ~n10988 & n14097;
  assign n14731 = n11063 & n14101;
  assign n14732 = ~n14125 & ~n14128;
  assign n14733 = n14125 & n14128;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = n14194 & ~n14734;
  assign n14736 = ~n14194 & n14734;
  assign n14737 = ~n14735 & ~n14736;
  assign n14738 = n14082 & ~n14737;
  assign n14739 = ~n14723 & ~n14729;
  assign n14740 = ~n14730 & n14739;
  assign n14741 = ~n14731 & n14740;
  assign n2525 = n14738 | ~n14741;
  assign n14743 = ~n10367 & ~n13916;
  assign n14744 = ~n10450 & ~n13920;
  assign n14745 = ~n10443 & n13924;
  assign n14746 = ~n10302 & n13926;
  assign n14747 = ~n10367 & ~n13902;
  assign n14748 = ~n14745 & ~n14746;
  assign n14749 = ~n14747 & n14748;
  assign n14750 = n13923 & ~n14749;
  assign n14751 = n13978 & ~n14068;
  assign n14752 = n13968 & ~n14751;
  assign n14753 = ~n13971 & ~n13972;
  assign n14754 = n13971 & n13972;
  assign n14755 = ~n14753 & ~n14754;
  assign n14756 = n14752 & ~n14755;
  assign n14757 = ~n14752 & n14755;
  assign n14758 = ~n14756 & ~n14757;
  assign n14759 = n14082 & ~n14758;
  assign n14760 = ~n14743 & ~n14744;
  assign n14761 = ~n12471 & n14760;
  assign n14762 = ~n14750 & n14761;
  assign n2530 = n14759 | ~n14762;
  assign n14764 = P2_REG3_REG_27_ & ~P2_STATE_REG;
  assign n14765 = ~n11252 & ~n13902;
  assign n14766 = ~n11194 & n13926;
  assign n14767 = ~n11323 & n13924;
  assign n14768 = ~n14765 & ~n14766;
  assign n14769 = ~n14767 & n14768;
  assign n14770 = n13923 & ~n14769;
  assign n14771 = ~n11252 & n14097;
  assign n14772 = n11325 & n14101;
  assign n14773 = ~n14625 & ~n14628;
  assign n14774 = ~n14645 & ~n14773;
  assign n14775 = ~n14622 & ~n14623;
  assign n14776 = n14622 & n14623;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = n14774 & ~n14777;
  assign n14779 = ~n14774 & n14777;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = n14082 & ~n14780;
  assign n14782 = ~n14764 & ~n14770;
  assign n14783 = ~n14771 & n14782;
  assign n14784 = ~n14772 & n14783;
  assign n2535 = n14781 | ~n14784;
  assign n14786 = ~n9936 & n13924;
  assign n14787 = ~n9788 & n13926;
  assign n14788 = ~n9845 & ~n13902;
  assign n14789 = ~n14786 & ~n14787;
  assign n14790 = ~n14788 & n14789;
  assign n14791 = n13923 & ~n14790;
  assign n14792 = n13981 & ~n13990;
  assign n14793 = n14000 & ~n14792;
  assign n14794 = ~n13986 & n14224;
  assign n14795 = n14793 & ~n14794;
  assign n14796 = ~n13981 & ~n13990;
  assign n14797 = n13981 & n13990;
  assign n14798 = ~n14796 & ~n14797;
  assign n14799 = ~n13986 & n14798;
  assign n14800 = ~n13998 & ~n14224;
  assign n14801 = n14799 & ~n14800;
  assign n14802 = ~n14795 & ~n14801;
  assign n14803 = n14082 & n14802;
  assign n14804 = ~n9943 & ~n13920;
  assign n14805 = ~n14803 & ~n14804;
  assign n14806 = ~n9845 & ~n13916;
  assign n14807 = ~n12755 & ~n14791;
  assign n14808 = n14805 & n14807;
  assign n2540 = n14806 | ~n14808;
  assign n14810 = P2_STATE_REG & ~n12250;
  assign n14811 = n9302 & n12251;
  assign n2550 = ~n14810 | n14811;
  assign n14813 = ~P3_IR_REG_31_ & P3_STATE_REG;
  assign n14814 = P3_STATE_REG & ~n14813;
  assign n14815 = P3_IR_REG_0_ & n14814;
  assign n14816 = P3_IR_REG_0_ & n14813;
  assign n14817 = SI_0_ & n2615_1;
  assign n14818 = ~P1_DATAO_REG_0_ & P2_DATAO_REG_0_;
  assign n14819 = P1_DATAO_REG_0_ & ~P2_DATAO_REG_0_;
  assign n14820 = ~n14818 & ~n14819;
  assign n14821 = ~n2615_1 & ~n14820;
  assign n14822 = ~n14817 & ~n14821;
  assign n14823 = ~P3_STATE_REG & ~n14822;
  assign n14824 = ~n14815 & ~n14816;
  assign n2560 = n14823 | ~n14824;
  assign n14826 = P3_IR_REG_0_ & ~P3_IR_REG_1_;
  assign n14827 = ~P3_IR_REG_0_ & P3_IR_REG_1_;
  assign n14828 = ~n14826 & ~n14827;
  assign n14829 = n14814 & ~n14828;
  assign n14830 = P3_IR_REG_1_ & n14813;
  assign n14831 = SI_1_ & n2615_1;
  assign n14832 = P1_DATAO_REG_1_ & ~P2_DATAO_REG_1_;
  assign n14833 = ~P1_DATAO_REG_1_ & P2_DATAO_REG_1_;
  assign n14834 = ~n14832 & ~n14833;
  assign n14835 = ~n14818 & ~n14834;
  assign n14836 = n14818 & n14834;
  assign n14837 = ~n14835 & ~n14836;
  assign n14838 = ~n2615_1 & ~n14837;
  assign n14839 = ~n14831 & ~n14838;
  assign n14840 = ~P3_STATE_REG & ~n14839;
  assign n14841 = ~n14829 & ~n14830;
  assign n2565 = n14840 | ~n14841;
  assign n14843 = ~P3_IR_REG_0_ & ~P3_IR_REG_1_;
  assign n14844 = P3_IR_REG_2_ & ~n14843;
  assign n14845 = ~P3_IR_REG_2_ & n14843;
  assign n14846 = ~n14844 & ~n14845;
  assign n14847 = n14814 & n14846;
  assign n14848 = P3_IR_REG_2_ & n14813;
  assign n14849 = SI_2_ & n2615_1;
  assign n14850 = P1_DATAO_REG_2_ & ~P2_DATAO_REG_2_;
  assign n14851 = ~P1_DATAO_REG_2_ & P2_DATAO_REG_2_;
  assign n14852 = ~n14850 & ~n14851;
  assign n14853 = P1_DATAO_REG_1_ & ~n14818;
  assign n14854 = ~P2_DATAO_REG_1_ & ~n14818;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = ~n14832 & n14855;
  assign n14857 = ~n14852 & ~n14856;
  assign n14858 = n14852 & n14856;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = ~n2615_1 & ~n14859;
  assign n14861 = ~n14849 & ~n14860;
  assign n14862 = ~P3_STATE_REG & ~n14861;
  assign n14863 = ~n14847 & ~n14848;
  assign n2570 = n14862 | ~n14863;
  assign n14865 = P3_IR_REG_3_ & ~n14845;
  assign n14866 = ~P3_IR_REG_3_ & n14845;
  assign n14867 = ~n14865 & ~n14866;
  assign n14868 = n14814 & n14867;
  assign n14869 = P3_IR_REG_3_ & n14813;
  assign n14870 = SI_3_ & n2615_1;
  assign n14871 = P1_DATAO_REG_3_ & ~P2_DATAO_REG_3_;
  assign n14872 = ~P1_DATAO_REG_3_ & P2_DATAO_REG_3_;
  assign n14873 = ~n14871 & ~n14872;
  assign n14874 = ~n14832 & ~n14853;
  assign n14875 = ~n14854 & n14874;
  assign n14876 = ~n14851 & ~n14875;
  assign n14877 = ~n14850 & ~n14876;
  assign n14878 = ~n14873 & ~n14877;
  assign n14879 = n14873 & n14877;
  assign n14880 = ~n14878 & ~n14879;
  assign n14881 = ~n2615_1 & ~n14880;
  assign n14882 = ~n14870 & ~n14881;
  assign n14883 = ~P3_STATE_REG & ~n14882;
  assign n14884 = ~n14868 & ~n14869;
  assign n2575 = n14883 | ~n14884;
  assign n14886 = P3_IR_REG_4_ & ~n14866;
  assign n14887 = ~P3_IR_REG_3_ & ~P3_IR_REG_4_;
  assign n14888 = n14845 & n14887;
  assign n14889 = ~n14886 & ~n14888;
  assign n14890 = n14814 & n14889;
  assign n14891 = P3_IR_REG_4_ & n14813;
  assign n14892 = SI_4_ & n2615_1;
  assign n14893 = P1_DATAO_REG_4_ & ~P2_DATAO_REG_4_;
  assign n14894 = ~P1_DATAO_REG_4_ & P2_DATAO_REG_4_;
  assign n14895 = ~n14893 & ~n14894;
  assign n14896 = ~n14850 & ~n14871;
  assign n14897 = ~n14872 & ~n14896;
  assign n14898 = ~n14851 & ~n14872;
  assign n14899 = ~n14856 & n14898;
  assign n14900 = ~n14897 & ~n14899;
  assign n14901 = ~n14895 & ~n14900;
  assign n14902 = n14895 & n14900;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n2615_1 & ~n14903;
  assign n14905 = ~n14892 & ~n14904;
  assign n14906 = ~P3_STATE_REG & ~n14905;
  assign n14907 = ~n14890 & ~n14891;
  assign n2580 = n14906 | ~n14907;
  assign n14909 = ~P3_IR_REG_5_ & n14888;
  assign n14910 = P3_IR_REG_5_ & ~n14888;
  assign n14911 = ~n14909 & ~n14910;
  assign n14912 = n14814 & n14911;
  assign n14913 = P3_IR_REG_5_ & n14813;
  assign n14914 = SI_5_ & n2615_1;
  assign n14915 = P1_DATAO_REG_5_ & ~P2_DATAO_REG_5_;
  assign n14916 = ~P1_DATAO_REG_5_ & P2_DATAO_REG_5_;
  assign n14917 = ~n14915 & ~n14916;
  assign n14918 = ~n14872 & ~n14894;
  assign n14919 = ~n14896 & n14918;
  assign n14920 = ~n14893 & ~n14919;
  assign n14921 = ~n14894 & n14898;
  assign n14922 = ~n14856 & n14921;
  assign n14923 = n14920 & ~n14922;
  assign n14924 = ~n14917 & ~n14923;
  assign n14925 = n14917 & n14923;
  assign n14926 = ~n14924 & ~n14925;
  assign n14927 = ~n2615_1 & ~n14926;
  assign n14928 = ~n14914 & ~n14927;
  assign n14929 = ~P3_STATE_REG & ~n14928;
  assign n14930 = ~n14912 & ~n14913;
  assign n2585 = n14929 | ~n14930;
  assign n14932 = P3_IR_REG_6_ & ~n14909;
  assign n14933 = ~P3_IR_REG_5_ & ~P3_IR_REG_6_;
  assign n14934 = n14888 & n14933;
  assign n14935 = ~n14932 & ~n14934;
  assign n14936 = n14814 & n14935;
  assign n14937 = P3_IR_REG_6_ & n14813;
  assign n14938 = SI_6_ & n2615_1;
  assign n14939 = P1_DATAO_REG_6_ & ~P2_DATAO_REG_6_;
  assign n14940 = ~P1_DATAO_REG_6_ & P2_DATAO_REG_6_;
  assign n14941 = ~n14939 & ~n14940;
  assign n14942 = ~n14916 & ~n14923;
  assign n14943 = ~n14915 & ~n14942;
  assign n14944 = ~n14941 & ~n14943;
  assign n14945 = n14941 & n14943;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = ~n2615_1 & ~n14946;
  assign n14948 = ~n14938 & ~n14947;
  assign n14949 = ~P3_STATE_REG & ~n14948;
  assign n14950 = ~n14936 & ~n14937;
  assign n2590 = n14949 | ~n14950;
  assign n14952 = P3_IR_REG_7_ & ~n14934;
  assign n14953 = ~P3_IR_REG_7_ & n14934;
  assign n14954 = ~n14952 & ~n14953;
  assign n14955 = n14814 & n14954;
  assign n14956 = P3_IR_REG_7_ & n14813;
  assign n14957 = SI_7_ & n2615_1;
  assign n14958 = P1_DATAO_REG_7_ & ~P2_DATAO_REG_7_;
  assign n14959 = ~P1_DATAO_REG_7_ & P2_DATAO_REG_7_;
  assign n14960 = ~n14958 & ~n14959;
  assign n14961 = n14915 & ~n14940;
  assign n14962 = ~n14939 & ~n14961;
  assign n14963 = ~n14916 & ~n14940;
  assign n14964 = ~n14923 & n14963;
  assign n14965 = n14962 & ~n14964;
  assign n14966 = ~n14960 & ~n14965;
  assign n14967 = n14960 & n14965;
  assign n14968 = ~n14966 & ~n14967;
  assign n14969 = ~n2615_1 & ~n14968;
  assign n14970 = ~n14957 & ~n14969;
  assign n14971 = ~P3_STATE_REG & ~n14970;
  assign n14972 = ~n14955 & ~n14956;
  assign n2595 = n14971 | ~n14972;
  assign n14974 = P3_IR_REG_8_ & ~n14953;
  assign n14975 = ~P3_IR_REG_7_ & ~P3_IR_REG_8_;
  assign n14976 = ~P3_IR_REG_5_ & n14887;
  assign n14977 = ~P3_IR_REG_6_ & n14976;
  assign n14978 = n14845 & n14975;
  assign n14979 = n14977 & n14978;
  assign n14980 = ~n14974 & ~n14979;
  assign n14981 = n14814 & n14980;
  assign n14982 = P3_IR_REG_8_ & n14813;
  assign n14983 = SI_8_ & n2615_1;
  assign n14984 = P1_DATAO_REG_8_ & ~P2_DATAO_REG_8_;
  assign n14985 = ~P1_DATAO_REG_8_ & P2_DATAO_REG_8_;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = ~n14959 & n14963;
  assign n14988 = ~n14923 & n14987;
  assign n14989 = ~n14939 & ~n14958;
  assign n14990 = ~n14961 & n14989;
  assign n14991 = ~n14959 & ~n14990;
  assign n14992 = ~n14988 & ~n14991;
  assign n14993 = ~n14986 & ~n14992;
  assign n14994 = n14986 & n14992;
  assign n14995 = ~n14993 & ~n14994;
  assign n14996 = ~n2615_1 & ~n14995;
  assign n14997 = ~n14983 & ~n14996;
  assign n14998 = ~P3_STATE_REG & ~n14997;
  assign n14999 = ~n14981 & ~n14982;
  assign n2600 = n14998 | ~n14999;
  assign n15001 = ~P3_IR_REG_9_ & n14979;
  assign n15002 = P3_IR_REG_9_ & ~n14979;
  assign n15003 = ~n15001 & ~n15002;
  assign n15004 = n14814 & n15003;
  assign n15005 = P3_IR_REG_9_ & n14813;
  assign n15006 = SI_9_ & n2615_1;
  assign n15007 = P1_DATAO_REG_9_ & ~P2_DATAO_REG_9_;
  assign n15008 = ~P1_DATAO_REG_9_ & P2_DATAO_REG_9_;
  assign n15009 = ~n15007 & ~n15008;
  assign n15010 = ~n14985 & n14991;
  assign n15011 = ~n14984 & ~n15010;
  assign n15012 = ~n14985 & n14987;
  assign n15013 = ~n14923 & n15012;
  assign n15014 = n15011 & ~n15013;
  assign n15015 = ~n15009 & ~n15014;
  assign n15016 = n15009 & n15014;
  assign n15017 = ~n15015 & ~n15016;
  assign n15018 = ~n2615_1 & ~n15017;
  assign n15019 = ~n15006 & ~n15018;
  assign n15020 = ~P3_STATE_REG & ~n15019;
  assign n15021 = ~n15004 & ~n15005;
  assign n2605 = n15020 | ~n15021;
  assign n15023 = P3_IR_REG_10_ & ~n15001;
  assign n15024 = ~P3_IR_REG_9_ & ~P3_IR_REG_10_;
  assign n15025 = n14979 & n15024;
  assign n15026 = ~n15023 & ~n15025;
  assign n15027 = n14814 & n15026;
  assign n15028 = P3_IR_REG_10_ & n14813;
  assign n15029 = SI_10_ & n2615_1;
  assign n15030 = P1_DATAO_REG_10_ & ~P2_DATAO_REG_10_;
  assign n15031 = ~P1_DATAO_REG_10_ & P2_DATAO_REG_10_;
  assign n15032 = ~n15030 & ~n15031;
  assign n15033 = ~n15008 & ~n15014;
  assign n15034 = ~n15007 & ~n15033;
  assign n15035 = ~n15032 & ~n15034;
  assign n15036 = n15032 & n15034;
  assign n15037 = ~n15035 & ~n15036;
  assign n15038 = ~n2615_1 & ~n15037;
  assign n15039 = ~n15029 & ~n15038;
  assign n15040 = ~P3_STATE_REG & ~n15039;
  assign n15041 = ~n15027 & ~n15028;
  assign n2610 = n15040 | ~n15041;
  assign n15043 = P3_IR_REG_11_ & ~n15025;
  assign n15044 = ~P3_IR_REG_11_ & n15025;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = n14814 & n15045;
  assign n15047 = P3_IR_REG_11_ & n14813;
  assign n15048 = SI_11_ & n2615_1;
  assign n15049 = P1_DATAO_REG_11_ & ~P2_DATAO_REG_11_;
  assign n15050 = ~P1_DATAO_REG_11_ & P2_DATAO_REG_11_;
  assign n15051 = ~n15049 & ~n15050;
  assign n15052 = n15007 & ~n15031;
  assign n15053 = ~n15030 & ~n15052;
  assign n15054 = ~n15008 & ~n15031;
  assign n15055 = ~n15014 & n15054;
  assign n15056 = n15053 & ~n15055;
  assign n15057 = ~n15051 & ~n15056;
  assign n15058 = n15051 & n15056;
  assign n15059 = ~n15057 & ~n15058;
  assign n15060 = ~n2615_1 & ~n15059;
  assign n15061 = ~n15048 & ~n15060;
  assign n15062 = ~P3_STATE_REG & ~n15061;
  assign n15063 = ~n15046 & ~n15047;
  assign n2615 = n15062 | ~n15063;
  assign n15065 = P3_IR_REG_12_ & ~n15044;
  assign n15066 = ~P3_IR_REG_10_ & ~P3_IR_REG_11_;
  assign n15067 = ~P3_IR_REG_12_ & n15066;
  assign n15068 = ~P3_IR_REG_9_ & n15067;
  assign n15069 = n14979 & n15068;
  assign n15070 = ~n15065 & ~n15069;
  assign n15071 = n14814 & n15070;
  assign n15072 = P3_IR_REG_12_ & n14813;
  assign n15073 = SI_12_ & n2615_1;
  assign n15074 = P1_DATAO_REG_12_ & ~P2_DATAO_REG_12_;
  assign n15075 = ~P1_DATAO_REG_12_ & P2_DATAO_REG_12_;
  assign n15076 = ~n15074 & ~n15075;
  assign n15077 = ~n15050 & ~n15053;
  assign n15078 = ~n15049 & ~n15077;
  assign n15079 = ~n15050 & n15054;
  assign n15080 = ~n15014 & n15079;
  assign n15081 = n15078 & ~n15080;
  assign n15082 = ~n15076 & ~n15081;
  assign n15083 = n15076 & n15081;
  assign n15084 = ~n15082 & ~n15083;
  assign n15085 = ~n2615_1 & ~n15084;
  assign n15086 = ~n15073 & ~n15085;
  assign n15087 = ~P3_STATE_REG & ~n15086;
  assign n15088 = ~n15071 & ~n15072;
  assign n2620 = n15087 | ~n15088;
  assign n15090 = ~P3_IR_REG_13_ & n15069;
  assign n15091 = P3_IR_REG_13_ & ~n15069;
  assign n15092 = ~n15090 & ~n15091;
  assign n15093 = n14814 & n15092;
  assign n15094 = P3_IR_REG_13_ & n14813;
  assign n15095 = SI_13_ & n2615_1;
  assign n15096 = P1_DATAO_REG_13_ & ~P2_DATAO_REG_13_;
  assign n15097 = ~P1_DATAO_REG_13_ & P2_DATAO_REG_13_;
  assign n15098 = ~n15096 & ~n15097;
  assign n15099 = ~n15075 & ~n15078;
  assign n15100 = ~n15074 & ~n15099;
  assign n15101 = ~n15075 & n15079;
  assign n15102 = ~n15014 & n15101;
  assign n15103 = n15100 & ~n15102;
  assign n15104 = ~n15098 & ~n15103;
  assign n15105 = n15098 & n15103;
  assign n15106 = ~n15104 & ~n15105;
  assign n15107 = ~n2615_1 & ~n15106;
  assign n15108 = ~n15095 & ~n15107;
  assign n15109 = ~P3_STATE_REG & ~n15108;
  assign n15110 = ~n15093 & ~n15094;
  assign n2625 = n15109 | ~n15110;
  assign n15112 = P3_IR_REG_14_ & ~n15090;
  assign n15113 = ~P3_IR_REG_13_ & ~P3_IR_REG_14_;
  assign n15114 = n15069 & n15113;
  assign n15115 = ~n15112 & ~n15114;
  assign n15116 = n14814 & n15115;
  assign n15117 = P3_IR_REG_14_ & n14813;
  assign n15118 = SI_14_ & n2615_1;
  assign n15119 = P1_DATAO_REG_14_ & ~P2_DATAO_REG_14_;
  assign n15120 = ~P1_DATAO_REG_14_ & P2_DATAO_REG_14_;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = ~n15097 & ~n15103;
  assign n15123 = ~n15096 & ~n15122;
  assign n15124 = ~n15121 & ~n15123;
  assign n15125 = n15121 & n15123;
  assign n15126 = ~n15124 & ~n15125;
  assign n15127 = ~n2615_1 & ~n15126;
  assign n15128 = ~n15118 & ~n15127;
  assign n15129 = ~P3_STATE_REG & ~n15128;
  assign n15130 = ~n15116 & ~n15117;
  assign n2630 = n15129 | ~n15130;
  assign n15132 = P3_IR_REG_15_ & ~n15114;
  assign n15133 = ~P3_IR_REG_15_ & n15114;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = n14814 & n15134;
  assign n15136 = P3_IR_REG_15_ & n14813;
  assign n15137 = SI_15_ & n2615_1;
  assign n15138 = P1_DATAO_REG_15_ & ~P2_DATAO_REG_15_;
  assign n15139 = ~P1_DATAO_REG_15_ & P2_DATAO_REG_15_;
  assign n15140 = ~n15138 & ~n15139;
  assign n15141 = ~n15120 & ~n15123;
  assign n15142 = ~n15119 & ~n15141;
  assign n15143 = ~n15140 & ~n15142;
  assign n15144 = n15140 & n15142;
  assign n15145 = ~n15143 & ~n15144;
  assign n15146 = ~n2615_1 & ~n15145;
  assign n15147 = ~n15137 & ~n15146;
  assign n15148 = ~P3_STATE_REG & ~n15147;
  assign n15149 = ~n15135 & ~n15136;
  assign n2635 = n15148 | ~n15149;
  assign n15151 = P3_IR_REG_16_ & ~n15133;
  assign n15152 = ~P3_IR_REG_6_ & ~P3_IR_REG_7_;
  assign n15153 = ~P3_IR_REG_8_ & n15152;
  assign n15154 = ~P3_IR_REG_9_ & n15153;
  assign n15155 = ~P3_IR_REG_2_ & ~P3_IR_REG_3_;
  assign n15156 = ~P3_IR_REG_4_ & n15155;
  assign n15157 = ~P3_IR_REG_5_ & n15156;
  assign n15158 = ~P3_IR_REG_15_ & ~P3_IR_REG_16_;
  assign n15159 = ~P3_IR_REG_1_ & n15158;
  assign n15160 = ~P3_IR_REG_0_ & n15159;
  assign n15161 = ~P3_IR_REG_12_ & n15113;
  assign n15162 = ~P3_IR_REG_10_ & n15161;
  assign n15163 = ~P3_IR_REG_11_ & n15162;
  assign n15164 = n15154 & n15157;
  assign n15165 = n15160 & n15164;
  assign n15166 = n15163 & n15165;
  assign n15167 = ~n15151 & ~n15166;
  assign n15168 = n14814 & n15167;
  assign n15169 = P3_IR_REG_16_ & n14813;
  assign n15170 = SI_16_ & n2615_1;
  assign n15171 = P1_DATAO_REG_16_ & ~P2_DATAO_REG_16_;
  assign n15172 = ~P1_DATAO_REG_16_ & P2_DATAO_REG_16_;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = ~n15139 & ~n15142;
  assign n15175 = ~n15138 & ~n15174;
  assign n15176 = ~n15173 & ~n15175;
  assign n15177 = n15173 & n15175;
  assign n15178 = ~n15176 & ~n15177;
  assign n15179 = ~n2615_1 & ~n15178;
  assign n15180 = ~n15170 & ~n15179;
  assign n15181 = ~P3_STATE_REG & ~n15180;
  assign n15182 = ~n15168 & ~n15169;
  assign n2640 = n15181 | ~n15182;
  assign n15184 = ~P3_IR_REG_17_ & n15166;
  assign n15185 = P3_IR_REG_17_ & ~n15166;
  assign n15186 = ~n15184 & ~n15185;
  assign n15187 = n14814 & n15186;
  assign n15188 = P3_IR_REG_17_ & n14813;
  assign n15189 = SI_17_ & n2615_1;
  assign n15190 = P1_DATAO_REG_17_ & ~P2_DATAO_REG_17_;
  assign n15191 = ~P1_DATAO_REG_17_ & P2_DATAO_REG_17_;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = ~n15172 & ~n15175;
  assign n15194 = ~n15171 & ~n15193;
  assign n15195 = ~n15192 & ~n15194;
  assign n15196 = n15192 & n15194;
  assign n15197 = ~n15195 & ~n15196;
  assign n15198 = ~n2615_1 & ~n15197;
  assign n15199 = ~n15189 & ~n15198;
  assign n15200 = ~P3_STATE_REG & ~n15199;
  assign n15201 = ~n15187 & ~n15188;
  assign n2645 = n15200 | ~n15201;
  assign n15203 = P3_IR_REG_18_ & ~n15184;
  assign n15204 = ~P3_IR_REG_17_ & ~P3_IR_REG_18_;
  assign n15205 = n15166 & n15204;
  assign n15206 = ~n15203 & ~n15205;
  assign n15207 = n14814 & n15206;
  assign n15208 = P3_IR_REG_18_ & n14813;
  assign n15209 = SI_18_ & n2615_1;
  assign n15210 = P1_DATAO_REG_18_ & ~P2_DATAO_REG_18_;
  assign n15211 = ~P1_DATAO_REG_18_ & P2_DATAO_REG_18_;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = ~n15191 & ~n15194;
  assign n15214 = ~n15190 & ~n15213;
  assign n15215 = ~n15212 & ~n15214;
  assign n15216 = n15212 & n15214;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = ~n2615_1 & ~n15217;
  assign n15219 = ~n15209 & ~n15218;
  assign n15220 = ~P3_STATE_REG & ~n15219;
  assign n15221 = ~n15207 & ~n15208;
  assign n2650 = n15220 | ~n15221;
  assign n15223 = P3_IR_REG_19_ & ~n15205;
  assign n15224 = ~P3_IR_REG_19_ & n15205;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = n14814 & n15225;
  assign n15227 = P3_IR_REG_19_ & n14813;
  assign n15228 = SI_19_ & n2615_1;
  assign n15229 = P1_DATAO_REG_19_ & ~P2_DATAO_REG_19_;
  assign n15230 = ~P1_DATAO_REG_19_ & P2_DATAO_REG_19_;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = ~n15211 & ~n15214;
  assign n15233 = ~n15210 & ~n15232;
  assign n15234 = ~n15231 & ~n15233;
  assign n15235 = n15231 & n15233;
  assign n15236 = ~n15234 & ~n15235;
  assign n15237 = ~n2615_1 & ~n15236;
  assign n15238 = ~n15228 & ~n15237;
  assign n15239 = ~P3_STATE_REG & ~n15238;
  assign n15240 = ~n15226 & ~n15227;
  assign n2655 = n15239 | ~n15240;
  assign n15242 = P3_IR_REG_20_ & ~n15224;
  assign n15243 = ~P3_IR_REG_19_ & ~P3_IR_REG_20_;
  assign n15244 = ~P3_IR_REG_17_ & n15243;
  assign n15245 = ~P3_IR_REG_18_ & n15244;
  assign n15246 = n15166 & n15245;
  assign n15247 = ~n15242 & ~n15246;
  assign n15248 = n14814 & n15247;
  assign n15249 = P3_IR_REG_20_ & n14813;
  assign n15250 = SI_20_ & n2615_1;
  assign n15251 = P1_DATAO_REG_20_ & ~P2_DATAO_REG_20_;
  assign n15252 = ~P1_DATAO_REG_20_ & P2_DATAO_REG_20_;
  assign n15253 = ~n15251 & ~n15252;
  assign n15254 = ~n15230 & ~n15233;
  assign n15255 = ~n15229 & ~n15254;
  assign n15256 = ~n15253 & ~n15255;
  assign n15257 = n15253 & n15255;
  assign n15258 = ~n15256 & ~n15257;
  assign n15259 = ~n2615_1 & ~n15258;
  assign n15260 = ~n15250 & ~n15259;
  assign n15261 = ~P3_STATE_REG & ~n15260;
  assign n15262 = ~n15248 & ~n15249;
  assign n2660 = n15261 | ~n15262;
  assign n15264 = ~P3_IR_REG_21_ & n15246;
  assign n15265 = P3_IR_REG_21_ & ~n15246;
  assign n15266 = ~n15264 & ~n15265;
  assign n15267 = n14814 & n15266;
  assign n15268 = P3_IR_REG_21_ & n14813;
  assign n15269 = SI_21_ & n2615_1;
  assign n15270 = P1_DATAO_REG_21_ & ~P2_DATAO_REG_21_;
  assign n15271 = ~P1_DATAO_REG_21_ & P2_DATAO_REG_21_;
  assign n15272 = ~n15270 & ~n15271;
  assign n15273 = ~n15252 & ~n15255;
  assign n15274 = ~n15251 & ~n15273;
  assign n15275 = ~n15272 & ~n15274;
  assign n15276 = n15272 & n15274;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = ~n2615_1 & ~n15277;
  assign n15279 = ~n15269 & ~n15278;
  assign n15280 = ~P3_STATE_REG & ~n15279;
  assign n15281 = ~n15267 & ~n15268;
  assign n2665 = n15280 | ~n15281;
  assign n15283 = P3_IR_REG_22_ & ~n15264;
  assign n15284 = ~P3_IR_REG_21_ & ~P3_IR_REG_22_;
  assign n15285 = n15246 & n15284;
  assign n15286 = ~n15283 & ~n15285;
  assign n15287 = n14814 & n15286;
  assign n15288 = P3_IR_REG_22_ & n14813;
  assign n15289 = SI_22_ & n2615_1;
  assign n15290 = P1_DATAO_REG_22_ & ~P2_DATAO_REG_22_;
  assign n15291 = ~P1_DATAO_REG_22_ & P2_DATAO_REG_22_;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15271 & ~n15274;
  assign n15294 = ~n15270 & ~n15293;
  assign n15295 = ~n15292 & ~n15294;
  assign n15296 = n15292 & n15294;
  assign n15297 = ~n15295 & ~n15296;
  assign n15298 = ~n2615_1 & ~n15297;
  assign n15299 = ~n15289 & ~n15298;
  assign n15300 = ~P3_STATE_REG & ~n15299;
  assign n15301 = ~n15287 & ~n15288;
  assign n2670 = n15300 | ~n15301;
  assign n15303 = P3_IR_REG_23_ & ~n15285;
  assign n15304 = ~P3_IR_REG_23_ & n15285;
  assign n15305 = ~n15303 & ~n15304;
  assign n15306 = n14814 & n15305;
  assign n15307 = P3_IR_REG_23_ & n14813;
  assign n15308 = SI_23_ & n2615_1;
  assign n15309 = P1_DATAO_REG_23_ & ~P2_DATAO_REG_23_;
  assign n15310 = ~P1_DATAO_REG_23_ & P2_DATAO_REG_23_;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = ~n15291 & ~n15294;
  assign n15313 = ~n15290 & ~n15312;
  assign n15314 = ~n15311 & ~n15313;
  assign n15315 = n15311 & n15313;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = ~n2615_1 & ~n15316;
  assign n15318 = ~n15308 & ~n15317;
  assign n15319 = ~P3_STATE_REG & ~n15318;
  assign n15320 = ~n15306 & ~n15307;
  assign n2675 = n15319 | ~n15320;
  assign n15322 = P3_IR_REG_24_ & ~n15304;
  assign n15323 = ~P3_IR_REG_21_ & ~P3_IR_REG_23_;
  assign n15324 = ~P3_IR_REG_22_ & n15323;
  assign n15325 = ~P3_IR_REG_24_ & n15245;
  assign n15326 = n15324 & n15325;
  assign n15327 = n15166 & n15326;
  assign n15328 = ~n15322 & ~n15327;
  assign n15329 = n14814 & n15328;
  assign n15330 = P3_IR_REG_24_ & n14813;
  assign n15331 = SI_24_ & n2615_1;
  assign n15332 = P1_DATAO_REG_24_ & ~P2_DATAO_REG_24_;
  assign n15333 = ~P1_DATAO_REG_24_ & P2_DATAO_REG_24_;
  assign n15334 = ~n15332 & ~n15333;
  assign n15335 = ~n15310 & ~n15313;
  assign n15336 = ~n15309 & ~n15335;
  assign n15337 = ~n15334 & ~n15336;
  assign n15338 = n15334 & n15336;
  assign n15339 = ~n15337 & ~n15338;
  assign n15340 = ~n2615_1 & ~n15339;
  assign n15341 = ~n15331 & ~n15340;
  assign n15342 = ~P3_STATE_REG & ~n15341;
  assign n15343 = ~n15329 & ~n15330;
  assign n2680 = n15342 | ~n15343;
  assign n15345 = ~P3_IR_REG_25_ & n15327;
  assign n15346 = P3_IR_REG_25_ & ~n15327;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = n14814 & n15347;
  assign n15349 = P3_IR_REG_25_ & n14813;
  assign n15350 = SI_25_ & n2615_1;
  assign n15351 = P1_DATAO_REG_25_ & ~P2_DATAO_REG_25_;
  assign n15352 = ~P1_DATAO_REG_25_ & P2_DATAO_REG_25_;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = ~n15333 & ~n15336;
  assign n15355 = ~n15332 & ~n15354;
  assign n15356 = ~n15353 & ~n15355;
  assign n15357 = n15353 & n15355;
  assign n15358 = ~n15356 & ~n15357;
  assign n15359 = ~n2615_1 & ~n15358;
  assign n15360 = ~n15350 & ~n15359;
  assign n15361 = ~P3_STATE_REG & ~n15360;
  assign n15362 = ~n15348 & ~n15349;
  assign n2685 = n15361 | ~n15362;
  assign n15364 = P3_IR_REG_26_ & ~n15345;
  assign n15365 = ~P3_IR_REG_25_ & ~P3_IR_REG_26_;
  assign n15366 = n15327 & n15365;
  assign n15367 = ~n15364 & ~n15366;
  assign n15368 = n14814 & n15367;
  assign n15369 = P3_IR_REG_26_ & n14813;
  assign n15370 = SI_26_ & n2615_1;
  assign n15371 = P1_DATAO_REG_26_ & ~P2_DATAO_REG_26_;
  assign n15372 = ~P1_DATAO_REG_26_ & P2_DATAO_REG_26_;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = ~n15352 & ~n15355;
  assign n15375 = ~n15351 & ~n15374;
  assign n15376 = ~n15373 & ~n15375;
  assign n15377 = n15373 & n15375;
  assign n15378 = ~n15376 & ~n15377;
  assign n15379 = ~n2615_1 & ~n15378;
  assign n15380 = ~n15370 & ~n15379;
  assign n15381 = ~P3_STATE_REG & ~n15380;
  assign n15382 = ~n15368 & ~n15369;
  assign n2690 = n15381 | ~n15382;
  assign n15384 = ~P3_IR_REG_27_ & n15366;
  assign n15385 = P3_IR_REG_27_ & ~n15366;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = n14814 & n15386;
  assign n15388 = P3_IR_REG_27_ & n14813;
  assign n15389 = SI_27_ & n2615_1;
  assign n15390 = P1_DATAO_REG_27_ & ~P2_DATAO_REG_27_;
  assign n15391 = ~P1_DATAO_REG_27_ & P2_DATAO_REG_27_;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = ~n15372 & ~n15375;
  assign n15394 = ~n15371 & ~n15393;
  assign n15395 = ~n15392 & ~n15394;
  assign n15396 = n15392 & n15394;
  assign n15397 = ~n15395 & ~n15396;
  assign n15398 = ~n2615_1 & ~n15397;
  assign n15399 = ~n15389 & ~n15398;
  assign n15400 = ~P3_STATE_REG & ~n15399;
  assign n15401 = ~n15387 & ~n15388;
  assign n2695 = n15400 | ~n15401;
  assign n15403 = P3_IR_REG_27_ & P3_IR_REG_28_;
  assign n15404 = ~P3_IR_REG_27_ & n15365;
  assign n15405 = ~P3_IR_REG_28_ & n15404;
  assign n15406 = n15327 & n15405;
  assign n15407 = ~n15403 & ~n15406;
  assign n15408 = P3_IR_REG_28_ & ~n15366;
  assign n15409 = n15407 & ~n15408;
  assign n15410 = n14814 & n15409;
  assign n15411 = P3_IR_REG_28_ & n14813;
  assign n15412 = SI_28_ & n2615_1;
  assign n15413 = P1_DATAO_REG_28_ & ~P2_DATAO_REG_28_;
  assign n15414 = ~P1_DATAO_REG_28_ & P2_DATAO_REG_28_;
  assign n15415 = ~n15413 & ~n15414;
  assign n15416 = ~n15391 & ~n15394;
  assign n15417 = ~n15390 & ~n15416;
  assign n15418 = ~n15415 & ~n15417;
  assign n15419 = n15415 & n15417;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = ~n2615_1 & ~n15420;
  assign n15422 = ~n15412 & ~n15421;
  assign n15423 = ~P3_STATE_REG & ~n15422;
  assign n15424 = ~n15410 & ~n15411;
  assign n2700 = n15423 | ~n15424;
  assign n15426 = P3_IR_REG_29_ & ~n15406;
  assign n15427 = ~P3_IR_REG_29_ & n15406;
  assign n15428 = ~n15426 & ~n15427;
  assign n15429 = n14814 & n15428;
  assign n15430 = P3_IR_REG_29_ & n14813;
  assign n15431 = SI_29_ & n2615_1;
  assign n15432 = P1_DATAO_REG_29_ & ~P2_DATAO_REG_29_;
  assign n15433 = ~P1_DATAO_REG_29_ & P2_DATAO_REG_29_;
  assign n15434 = ~n15432 & ~n15433;
  assign n15435 = ~n15414 & ~n15417;
  assign n15436 = ~n15413 & ~n15435;
  assign n15437 = ~n15434 & ~n15436;
  assign n15438 = n15434 & n15436;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = ~n2615_1 & ~n15439;
  assign n15441 = ~n15431 & ~n15440;
  assign n15442 = ~P3_STATE_REG & ~n15441;
  assign n15443 = ~n15429 & ~n15430;
  assign n2705 = n15442 | ~n15443;
  assign n15445 = ~P3_IR_REG_30_ & n15427;
  assign n15446 = P3_IR_REG_30_ & ~n15427;
  assign n15447 = ~n15445 & ~n15446;
  assign n15448 = n14814 & n15447;
  assign n15449 = P3_IR_REG_30_ & n14813;
  assign n15450 = SI_30_ & n2615_1;
  assign n15451 = P1_DATAO_REG_30_ & ~P2_DATAO_REG_30_;
  assign n15452 = ~P1_DATAO_REG_30_ & P2_DATAO_REG_30_;
  assign n15453 = ~n15451 & ~n15452;
  assign n15454 = ~n15433 & ~n15436;
  assign n15455 = ~n15432 & ~n15454;
  assign n15456 = ~n15453 & ~n15455;
  assign n15457 = n15453 & n15455;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = ~n2615_1 & ~n15458;
  assign n15460 = ~n15450 & ~n15459;
  assign n15461 = ~P3_STATE_REG & ~n15460;
  assign n15462 = ~n15448 & ~n15449;
  assign n2710 = n15461 | ~n15462;
  assign n15464 = P3_IR_REG_31_ & n15445;
  assign n15465 = ~P3_IR_REG_31_ & ~n15445;
  assign n15466 = ~n15464 & ~n15465;
  assign n15467 = n14814 & ~n15466;
  assign n15468 = P3_IR_REG_31_ & n14813;
  assign n15469 = SI_31_ & n2615_1;
  assign n15470 = P1_DATAO_REG_31_ & ~P2_DATAO_REG_31_;
  assign n15471 = ~P1_DATAO_REG_31_ & P2_DATAO_REG_31_;
  assign n15472 = ~n15470 & ~n15471;
  assign n15473 = ~P1_DATAO_REG_30_ & n15472;
  assign n15474 = P2_DATAO_REG_30_ & n15473;
  assign n15475 = P1_DATAO_REG_30_ & ~n15472;
  assign n15476 = ~P2_DATAO_REG_30_ & n15475;
  assign n15477 = ~n15474 & ~n15476;
  assign n15478 = ~n15451 & n15472;
  assign n15479 = ~n15432 & n15478;
  assign n15480 = ~n15454 & n15479;
  assign n15481 = n15477 & ~n15480;
  assign n15482 = ~n15452 & ~n15472;
  assign n15483 = ~n15455 & n15482;
  assign n15484 = n15481 & ~n15483;
  assign n15485 = ~n2615_1 & ~n15484;
  assign n15486 = ~n15469 & ~n15485;
  assign n15487 = ~P3_STATE_REG & ~n15486;
  assign n15488 = ~n15467 & ~n15468;
  assign n2715 = n15487 | ~n15488;
  assign n15490 = P3_IR_REG_31_ & n15305;
  assign n15491 = P3_IR_REG_23_ & ~P3_IR_REG_31_;
  assign n15492 = ~n15490 & ~n15491;
  assign n15493 = P3_IR_REG_31_ & n15347;
  assign n15494 = P3_IR_REG_25_ & ~P3_IR_REG_31_;
  assign n15495 = ~n15493 & ~n15494;
  assign n15496 = P3_IR_REG_31_ & n15367;
  assign n15497 = P3_IR_REG_26_ & ~P3_IR_REG_31_;
  assign n15498 = ~n15496 & ~n15497;
  assign n15499 = P3_IR_REG_31_ & n15328;
  assign n15500 = P3_IR_REG_24_ & ~P3_IR_REG_31_;
  assign n15501 = ~n15499 & ~n15500;
  assign n15502 = ~n15495 & ~n15498;
  assign n15503 = ~n15501 & n15502;
  assign n15504 = n15492 & ~n15503;
  assign n15505 = P3_STATE_REG & n15504;
  assign n15506 = n15495 & ~n15498;
  assign n15507 = ~P3_B_REG & ~n15501;
  assign n15508 = P3_B_REG & n15501;
  assign n15509 = ~n15507 & ~n15508;
  assign n15510 = n15506 & ~n15509;
  assign n15511 = ~n15498 & ~n15510;
  assign n15512 = n15505 & ~n15511;
  assign n15513 = n15501 & ~n15506;
  assign n15514 = n15512 & ~n15513;
  assign n15515 = P3_D_REG_0_ & ~n15512;
  assign n2720 = n15514 | n15515;
  assign n15517 = n15495 & ~n15506;
  assign n15518 = n15512 & ~n15517;
  assign n15519 = P3_D_REG_1_ & ~n15512;
  assign n2725 = n15518 | n15519;
  assign n2730 = P3_D_REG_2_ & ~n15512;
  assign n2735 = P3_D_REG_3_ & ~n15512;
  assign n2740 = P3_D_REG_4_ & ~n15512;
  assign n2745 = P3_D_REG_5_ & ~n15512;
  assign n2750 = P3_D_REG_6_ & ~n15512;
  assign n2755 = P3_D_REG_7_ & ~n15512;
  assign n2760 = P3_D_REG_8_ & ~n15512;
  assign n2765 = P3_D_REG_9_ & ~n15512;
  assign n2770 = P3_D_REG_10_ & ~n15512;
  assign n2775 = P3_D_REG_11_ & ~n15512;
  assign n2780 = P3_D_REG_12_ & ~n15512;
  assign n2785 = P3_D_REG_13_ & ~n15512;
  assign n2790 = P3_D_REG_14_ & ~n15512;
  assign n2795 = P3_D_REG_15_ & ~n15512;
  assign n2800 = P3_D_REG_16_ & ~n15512;
  assign n2805 = P3_D_REG_17_ & ~n15512;
  assign n2810 = P3_D_REG_18_ & ~n15512;
  assign n2815 = P3_D_REG_19_ & ~n15512;
  assign n2820 = P3_D_REG_20_ & ~n15512;
  assign n2825 = P3_D_REG_21_ & ~n15512;
  assign n2830 = P3_D_REG_22_ & ~n15512;
  assign n2835 = P3_D_REG_23_ & ~n15512;
  assign n2840 = P3_D_REG_24_ & ~n15512;
  assign n2845 = P3_D_REG_25_ & ~n15512;
  assign n2850 = P3_D_REG_26_ & ~n15512;
  assign n2855 = P3_D_REG_27_ & ~n15512;
  assign n2860 = P3_D_REG_28_ & ~n15512;
  assign n2865 = P3_D_REG_29_ & ~n15512;
  assign n2870 = P3_D_REG_30_ & ~n15512;
  assign n2875 = P3_D_REG_31_ & ~n15512;
  assign n15551 = ~n15511 & ~n15517;
  assign n15552 = P3_D_REG_1_ & n15511;
  assign n15553 = ~n15551 & ~n15552;
  assign n15554 = P3_D_REG_0_ & n15511;
  assign n15555 = n15498 & n15501;
  assign n15556 = ~n15511 & ~n15555;
  assign n15557 = ~n15554 & ~n15556;
  assign n15558 = n15553 & n15557;
  assign n15559 = P3_D_REG_8_ & n15511;
  assign n15560 = P3_D_REG_7_ & n15511;
  assign n15561 = P3_D_REG_9_ & n15511;
  assign n15562 = ~n15559 & ~n15560;
  assign n15563 = ~n15561 & n15562;
  assign n15564 = P3_D_REG_6_ & n15511;
  assign n15565 = P3_D_REG_5_ & n15511;
  assign n15566 = P3_D_REG_4_ & n15511;
  assign n15567 = P3_D_REG_3_ & n15511;
  assign n15568 = ~n15564 & ~n15565;
  assign n15569 = ~n15566 & n15568;
  assign n15570 = ~n15567 & n15569;
  assign n15571 = P3_D_REG_31_ & n15511;
  assign n15572 = P3_D_REG_30_ & n15511;
  assign n15573 = P3_D_REG_2_ & n15511;
  assign n15574 = P3_D_REG_29_ & n15511;
  assign n15575 = ~n15571 & ~n15572;
  assign n15576 = ~n15573 & n15575;
  assign n15577 = ~n15574 & n15576;
  assign n15578 = P3_D_REG_28_ & n15511;
  assign n15579 = P3_D_REG_27_ & n15511;
  assign n15580 = P3_D_REG_26_ & n15511;
  assign n15581 = P3_D_REG_25_ & n15511;
  assign n15582 = ~n15578 & ~n15579;
  assign n15583 = ~n15580 & n15582;
  assign n15584 = ~n15581 & n15583;
  assign n15585 = n15563 & n15570;
  assign n15586 = n15577 & n15585;
  assign n15587 = n15584 & n15586;
  assign n15588 = P3_D_REG_23_ & n15511;
  assign n15589 = P3_D_REG_22_ & n15511;
  assign n15590 = P3_D_REG_24_ & n15511;
  assign n15591 = ~n15588 & ~n15589;
  assign n15592 = ~n15590 & n15591;
  assign n15593 = P3_D_REG_21_ & n15511;
  assign n15594 = P3_D_REG_20_ & n15511;
  assign n15595 = P3_D_REG_19_ & n15511;
  assign n15596 = P3_D_REG_18_ & n15511;
  assign n15597 = ~n15593 & ~n15594;
  assign n15598 = ~n15595 & n15597;
  assign n15599 = ~n15596 & n15598;
  assign n15600 = P3_D_REG_17_ & n15511;
  assign n15601 = P3_D_REG_16_ & n15511;
  assign n15602 = P3_D_REG_15_ & n15511;
  assign n15603 = P3_D_REG_14_ & n15511;
  assign n15604 = ~n15600 & ~n15601;
  assign n15605 = ~n15602 & n15604;
  assign n15606 = ~n15603 & n15605;
  assign n15607 = P3_D_REG_13_ & n15511;
  assign n15608 = P3_D_REG_12_ & n15511;
  assign n15609 = P3_D_REG_11_ & n15511;
  assign n15610 = P3_D_REG_10_ & n15511;
  assign n15611 = ~n15607 & ~n15608;
  assign n15612 = ~n15609 & n15611;
  assign n15613 = ~n15610 & n15612;
  assign n15614 = n15592 & n15599;
  assign n15615 = n15606 & n15614;
  assign n15616 = n15613 & n15615;
  assign n15617 = n15587 & n15616;
  assign n15618 = n15558 & n15617;
  assign n15619 = P3_IR_REG_31_ & n15286;
  assign n15620 = P3_IR_REG_22_ & ~P3_IR_REG_31_;
  assign n15621 = ~n15619 & ~n15620;
  assign n15622 = P3_IR_REG_31_ & n15266;
  assign n15623 = P3_IR_REG_21_ & ~P3_IR_REG_31_;
  assign n15624 = ~n15622 & ~n15623;
  assign n15625 = P3_IR_REG_31_ & n15247;
  assign n15626 = P3_IR_REG_20_ & ~P3_IR_REG_31_;
  assign n15627 = ~n15625 & ~n15626;
  assign n15628 = n15624 & n15627;
  assign n15629 = ~n15621 & ~n15628;
  assign n15630 = n15621 & n15628;
  assign n15631 = ~n15629 & ~n15630;
  assign n15632 = P3_IR_REG_31_ & n15225;
  assign n15633 = P3_IR_REG_19_ & ~P3_IR_REG_31_;
  assign n15634 = ~n15632 & ~n15633;
  assign n15635 = n15624 & n15634;
  assign n15636 = ~n15631 & ~n15635;
  assign n15637 = n15618 & ~n15636;
  assign n15638 = ~n15553 & ~n15557;
  assign n15639 = n15617 & n15638;
  assign n15640 = ~n15621 & ~n15634;
  assign n15641 = n15624 & n15640;
  assign n15642 = ~n15627 & n15641;
  assign n15643 = ~n15621 & n15634;
  assign n15644 = n15627 & n15643;
  assign n15645 = ~n15624 & n15644;
  assign n15646 = ~n15642 & ~n15645;
  assign n15647 = n15639 & ~n15646;
  assign n15648 = ~n15637 & ~n15647;
  assign n15649 = n15505 & ~n15648;
  assign n15650 = P3_IR_REG_31_ & n15386;
  assign n15651 = P3_IR_REG_27_ & ~P3_IR_REG_31_;
  assign n15652 = ~n15650 & ~n15651;
  assign n15653 = P3_IR_REG_31_ & n15409;
  assign n15654 = P3_IR_REG_28_ & ~P3_IR_REG_31_;
  assign n15655 = ~n15653 & ~n15654;
  assign n15656 = n15652 & n15655;
  assign n15657 = P3_IR_REG_0_ & P3_IR_REG_31_;
  assign n15658 = P3_IR_REG_0_ & ~P3_IR_REG_31_;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = n15656 & ~n15659;
  assign n15661 = ~n14822 & ~n15656;
  assign n15662 = ~n15660 & ~n15661;
  assign n15663 = n15621 & n15634;
  assign n15664 = n15624 & n15663;
  assign n15665 = n15621 & ~n15634;
  assign n15666 = n15624 & n15665;
  assign n15667 = ~n15664 & ~n15666;
  assign n15668 = ~n15662 & ~n15667;
  assign n15669 = P3_IR_REG_31_ & n15447;
  assign n15670 = P3_IR_REG_30_ & ~P3_IR_REG_31_;
  assign n15671 = ~n15669 & ~n15670;
  assign n15672 = P3_IR_REG_31_ & n15428;
  assign n15673 = P3_IR_REG_29_ & ~P3_IR_REG_31_;
  assign n15674 = ~n15672 & ~n15673;
  assign n15675 = ~n15671 & ~n15674;
  assign n15676 = P3_REG3_REG_0_ & n15675;
  assign n15677 = ~n15671 & n15674;
  assign n15678 = P3_REG2_REG_0_ & n15677;
  assign n15679 = n15671 & ~n15674;
  assign n15680 = P3_REG1_REG_0_ & n15679;
  assign n15681 = n15671 & n15674;
  assign n15682 = P3_REG0_REG_0_ & n15681;
  assign n15683 = ~n15676 & ~n15678;
  assign n15684 = ~n15680 & n15683;
  assign n15685 = ~n15682 & n15684;
  assign n15686 = ~n15662 & n15685;
  assign n15687 = n15662 & ~n15685;
  assign n15688 = ~n15686 & ~n15687;
  assign n15689 = n15627 & n15665;
  assign n15690 = ~n15688 & n15689;
  assign n15691 = ~n15621 & ~n15624;
  assign n15692 = ~n15652 & ~n15655;
  assign n15693 = ~n15656 & ~n15692;
  assign n15694 = n15691 & ~n15693;
  assign n15695 = P3_REG3_REG_1_ & n15675;
  assign n15696 = P3_REG2_REG_1_ & n15677;
  assign n15697 = P3_REG1_REG_1_ & n15679;
  assign n15698 = P3_REG0_REG_1_ & n15681;
  assign n15699 = ~n15695 & ~n15696;
  assign n15700 = ~n15697 & n15699;
  assign n15701 = ~n15698 & n15700;
  assign n15702 = n15694 & ~n15701;
  assign n15703 = ~n15668 & ~n15690;
  assign n15704 = ~n15702 & n15703;
  assign n15705 = n15624 & n15643;
  assign n15706 = n15627 & n15705;
  assign n15707 = ~n15688 & n15706;
  assign n15708 = ~n15624 & n15634;
  assign n15709 = ~n15627 & n15708;
  assign n15710 = ~n15688 & n15709;
  assign n15711 = ~n15624 & n15663;
  assign n15712 = n15627 & n15711;
  assign n15713 = ~n15688 & n15712;
  assign n15714 = ~n15624 & ~n15634;
  assign n15715 = ~n15627 & n15714;
  assign n15716 = ~n15688 & n15715;
  assign n15717 = ~n15627 & n15643;
  assign n15718 = ~n15688 & n15717;
  assign n15719 = ~n15716 & ~n15718;
  assign n15720 = ~n15627 & n15640;
  assign n15721 = ~n15688 & n15720;
  assign n15722 = n15627 & n15640;
  assign n15723 = ~n15688 & n15722;
  assign n15724 = ~n15721 & ~n15723;
  assign n15725 = ~n15707 & ~n15710;
  assign n15726 = ~n15713 & n15725;
  assign n15727 = n15719 & n15726;
  assign n15728 = n15724 & n15727;
  assign n15729 = n15704 & n15728;
  assign n15730 = n15649 & ~n15729;
  assign n15731 = P3_REG0_REG_0_ & ~n15649;
  assign n2880 = n15730 | n15731;
  assign n15733 = P3_REG3_REG_2_ & n15675;
  assign n15734 = P3_REG2_REG_2_ & n15677;
  assign n15735 = P3_REG1_REG_2_ & n15679;
  assign n15736 = P3_REG0_REG_2_ & n15681;
  assign n15737 = ~n15733 & ~n15734;
  assign n15738 = ~n15735 & n15737;
  assign n15739 = ~n15736 & n15738;
  assign n15740 = n15694 & ~n15739;
  assign n15741 = P3_IR_REG_31_ & ~n14828;
  assign n15742 = P3_IR_REG_1_ & ~P3_IR_REG_31_;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = n15656 & ~n15743;
  assign n15745 = ~n14839 & ~n15656;
  assign n15746 = ~n15744 & ~n15745;
  assign n15747 = ~n15667 & ~n15746;
  assign n15748 = ~n15701 & n15746;
  assign n15749 = n15701 & ~n15746;
  assign n15750 = ~n15748 & ~n15749;
  assign n15751 = ~n15686 & ~n15750;
  assign n15752 = n15686 & n15750;
  assign n15753 = ~n15751 & ~n15752;
  assign n15754 = n15689 & ~n15753;
  assign n15755 = ~n15740 & ~n15747;
  assign n15756 = ~n15754 & n15755;
  assign n15757 = ~n15701 & ~n15746;
  assign n15758 = n15701 & n15746;
  assign n15759 = ~n15757 & ~n15758;
  assign n15760 = ~n15662 & ~n15685;
  assign n15761 = n15759 & ~n15760;
  assign n15762 = ~n15759 & n15760;
  assign n15763 = ~n15761 & ~n15762;
  assign n15764 = n15722 & ~n15763;
  assign n15765 = ~n15652 & n15655;
  assign n15766 = n15652 & ~n15655;
  assign n15767 = ~n15765 & ~n15766;
  assign n15768 = n15691 & ~n15767;
  assign n15769 = ~n15685 & n15768;
  assign n15770 = n15717 & ~n15753;
  assign n15771 = n15720 & ~n15763;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = n15712 & ~n15753;
  assign n15774 = n15706 & ~n15753;
  assign n15775 = n15709 & ~n15763;
  assign n15776 = n15715 & ~n15763;
  assign n15777 = ~n15775 & ~n15776;
  assign n15778 = ~n15773 & ~n15774;
  assign n15779 = n15777 & n15778;
  assign n15780 = ~n15764 & ~n15769;
  assign n15781 = n15772 & n15780;
  assign n15782 = n15779 & n15781;
  assign n15783 = n15756 & n15782;
  assign n15784 = n15649 & ~n15783;
  assign n15785 = P3_REG0_REG_1_ & ~n15649;
  assign n2885 = n15784 | n15785;
  assign n15787 = ~P3_REG3_REG_3_ & n15675;
  assign n15788 = P3_REG2_REG_3_ & n15677;
  assign n15789 = P3_REG1_REG_3_ & n15679;
  assign n15790 = P3_REG0_REG_3_ & n15681;
  assign n15791 = ~n15787 & ~n15788;
  assign n15792 = ~n15789 & n15791;
  assign n15793 = ~n15790 & n15792;
  assign n15794 = n15694 & ~n15793;
  assign n15795 = P3_IR_REG_31_ & n14846;
  assign n15796 = P3_IR_REG_2_ & ~P3_IR_REG_31_;
  assign n15797 = ~n15795 & ~n15796;
  assign n15798 = n15656 & ~n15797;
  assign n15799 = ~n14861 & ~n15656;
  assign n15800 = ~n15798 & ~n15799;
  assign n15801 = ~n15667 & ~n15800;
  assign n15802 = ~n15739 & n15800;
  assign n15803 = n15739 & ~n15800;
  assign n15804 = ~n15802 & ~n15803;
  assign n15805 = ~n15686 & ~n15701;
  assign n15806 = ~n15686 & n15746;
  assign n15807 = ~n15805 & ~n15806;
  assign n15808 = ~n15748 & n15807;
  assign n15809 = n15804 & n15808;
  assign n15810 = ~n15804 & ~n15808;
  assign n15811 = ~n15809 & ~n15810;
  assign n15812 = n15689 & ~n15811;
  assign n15813 = ~n15794 & ~n15801;
  assign n15814 = ~n15812 & n15813;
  assign n15815 = ~n15739 & ~n15800;
  assign n15816 = n15739 & n15800;
  assign n15817 = ~n15815 & ~n15816;
  assign n15818 = ~n15758 & n15760;
  assign n15819 = ~n15757 & ~n15818;
  assign n15820 = n15817 & ~n15819;
  assign n15821 = ~n15757 & n15804;
  assign n15822 = ~n15818 & n15821;
  assign n15823 = ~n15820 & ~n15822;
  assign n15824 = n15722 & n15823;
  assign n15825 = ~n15701 & n15768;
  assign n15826 = n15717 & ~n15811;
  assign n15827 = n15720 & n15823;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = n15712 & ~n15811;
  assign n15830 = n15706 & ~n15811;
  assign n15831 = n15709 & n15823;
  assign n15832 = n15715 & n15823;
  assign n15833 = ~n15831 & ~n15832;
  assign n15834 = ~n15829 & ~n15830;
  assign n15835 = n15833 & n15834;
  assign n15836 = ~n15824 & ~n15825;
  assign n15837 = n15828 & n15836;
  assign n15838 = n15835 & n15837;
  assign n15839 = n15814 & n15838;
  assign n15840 = n15649 & ~n15839;
  assign n15841 = P3_REG0_REG_2_ & ~n15649;
  assign n2890 = n15840 | n15841;
  assign n15843 = ~P3_REG3_REG_4_ & ~P3_REG3_REG_3_;
  assign n15844 = P3_REG3_REG_4_ & P3_REG3_REG_3_;
  assign n15845 = ~n15843 & ~n15844;
  assign n15846 = n15675 & ~n15845;
  assign n15847 = P3_REG2_REG_4_ & n15677;
  assign n15848 = P3_REG1_REG_4_ & n15679;
  assign n15849 = P3_REG0_REG_4_ & n15681;
  assign n15850 = ~n15846 & ~n15847;
  assign n15851 = ~n15848 & n15850;
  assign n15852 = ~n15849 & n15851;
  assign n15853 = n15694 & ~n15852;
  assign n15854 = P3_IR_REG_31_ & n14867;
  assign n15855 = P3_IR_REG_3_ & ~P3_IR_REG_31_;
  assign n15856 = ~n15854 & ~n15855;
  assign n15857 = n15656 & ~n15856;
  assign n15858 = ~n14882 & ~n15656;
  assign n15859 = ~n15857 & ~n15858;
  assign n15860 = ~n15667 & ~n15859;
  assign n15861 = ~n15793 & n15859;
  assign n15862 = n15793 & ~n15859;
  assign n15863 = ~n15861 & ~n15862;
  assign n15864 = ~n15803 & ~n15863;
  assign n15865 = ~n15802 & n15808;
  assign n15866 = n15864 & ~n15865;
  assign n15867 = ~n15802 & n15863;
  assign n15868 = ~n15803 & ~n15808;
  assign n15869 = n15867 & ~n15868;
  assign n15870 = ~n15866 & ~n15869;
  assign n15871 = n15689 & ~n15870;
  assign n15872 = ~n15853 & ~n15860;
  assign n15873 = ~n15871 & n15872;
  assign n15874 = n15757 & ~n15816;
  assign n15875 = ~n15815 & ~n15874;
  assign n15876 = ~n15816 & n15818;
  assign n15877 = n15875 & ~n15876;
  assign n15878 = ~n15863 & n15877;
  assign n15879 = ~n15793 & ~n15859;
  assign n15880 = n15793 & n15859;
  assign n15881 = ~n15879 & ~n15880;
  assign n15882 = ~n15877 & ~n15881;
  assign n15883 = ~n15878 & ~n15882;
  assign n15884 = n15722 & ~n15883;
  assign n15885 = ~n15739 & n15768;
  assign n15886 = n15717 & ~n15870;
  assign n15887 = n15720 & ~n15883;
  assign n15888 = ~n15886 & ~n15887;
  assign n15889 = n15712 & ~n15870;
  assign n15890 = n15706 & ~n15870;
  assign n15891 = n15709 & ~n15883;
  assign n15892 = n15715 & ~n15883;
  assign n15893 = ~n15891 & ~n15892;
  assign n15894 = ~n15889 & ~n15890;
  assign n15895 = n15893 & n15894;
  assign n15896 = ~n15884 & ~n15885;
  assign n15897 = n15888 & n15896;
  assign n15898 = n15895 & n15897;
  assign n15899 = n15873 & n15898;
  assign n15900 = n15649 & ~n15899;
  assign n15901 = P3_REG0_REG_3_ & ~n15649;
  assign n2895 = n15900 | n15901;
  assign n15903 = ~P3_REG3_REG_5_ & n15843;
  assign n15904 = P3_REG3_REG_5_ & ~n15843;
  assign n15905 = ~n15903 & ~n15904;
  assign n15906 = n15675 & ~n15905;
  assign n15907 = P3_REG2_REG_5_ & n15677;
  assign n15908 = P3_REG1_REG_5_ & n15679;
  assign n15909 = P3_REG0_REG_5_ & n15681;
  assign n15910 = ~n15906 & ~n15907;
  assign n15911 = ~n15908 & n15910;
  assign n15912 = ~n15909 & n15911;
  assign n15913 = n15694 & ~n15912;
  assign n15914 = P3_IR_REG_31_ & n14889;
  assign n15915 = P3_IR_REG_4_ & ~P3_IR_REG_31_;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = n15656 & ~n15916;
  assign n15918 = ~n14905 & ~n15656;
  assign n15919 = ~n15917 & ~n15918;
  assign n15920 = ~n15667 & ~n15919;
  assign n15921 = n15793 & ~n15802;
  assign n15922 = n15859 & ~n15921;
  assign n15923 = ~n15793 & n15802;
  assign n15924 = ~n15922 & ~n15923;
  assign n15925 = ~n15803 & ~n15862;
  assign n15926 = ~n15808 & n15925;
  assign n15927 = n15924 & ~n15926;
  assign n15928 = ~n15852 & n15919;
  assign n15929 = n15852 & ~n15919;
  assign n15930 = ~n15928 & ~n15929;
  assign n15931 = n15927 & n15930;
  assign n15932 = ~n15927 & ~n15930;
  assign n15933 = ~n15931 & ~n15932;
  assign n15934 = n15689 & ~n15933;
  assign n15935 = ~n15913 & ~n15920;
  assign n15936 = ~n15934 & n15935;
  assign n15937 = ~n15816 & ~n15880;
  assign n15938 = n15818 & n15937;
  assign n15939 = ~n15879 & ~n15938;
  assign n15940 = ~n15875 & ~n15880;
  assign n15941 = n15939 & ~n15940;
  assign n15942 = ~n15930 & n15941;
  assign n15943 = n15852 & n15919;
  assign n15944 = ~n15852 & ~n15919;
  assign n15945 = ~n15943 & ~n15944;
  assign n15946 = ~n15941 & ~n15945;
  assign n15947 = ~n15942 & ~n15946;
  assign n15948 = n15722 & ~n15947;
  assign n15949 = n15768 & ~n15793;
  assign n15950 = n15720 & ~n15947;
  assign n15951 = n15717 & ~n15933;
  assign n15952 = n15712 & ~n15933;
  assign n15953 = n15706 & ~n15933;
  assign n15954 = n15709 & ~n15947;
  assign n15955 = n15715 & ~n15947;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = ~n15952 & ~n15953;
  assign n15958 = n15956 & n15957;
  assign n15959 = ~n15948 & ~n15949;
  assign n15960 = ~n15950 & n15959;
  assign n15961 = ~n15951 & n15960;
  assign n15962 = n15958 & n15961;
  assign n15963 = n15936 & n15962;
  assign n15964 = n15649 & ~n15963;
  assign n15965 = P3_REG0_REG_4_ & ~n15649;
  assign n2900 = n15964 | n15965;
  assign n15967 = ~P3_REG3_REG_6_ & ~P3_REG3_REG_5_;
  assign n15968 = ~P3_REG3_REG_4_ & n15967;
  assign n15969 = ~P3_REG3_REG_3_ & n15968;
  assign n15970 = P3_REG3_REG_6_ & ~n15903;
  assign n15971 = ~n15969 & ~n15970;
  assign n15972 = n15675 & ~n15971;
  assign n15973 = P3_REG2_REG_6_ & n15677;
  assign n15974 = P3_REG1_REG_6_ & n15679;
  assign n15975 = P3_REG0_REG_6_ & n15681;
  assign n15976 = ~n15972 & ~n15973;
  assign n15977 = ~n15974 & n15976;
  assign n15978 = ~n15975 & n15977;
  assign n15979 = n15694 & ~n15978;
  assign n15980 = P3_IR_REG_31_ & n14911;
  assign n15981 = P3_IR_REG_5_ & ~P3_IR_REG_31_;
  assign n15982 = ~n15980 & ~n15981;
  assign n15983 = n15656 & ~n15982;
  assign n15984 = ~n14928 & ~n15656;
  assign n15985 = ~n15983 & ~n15984;
  assign n15986 = ~n15667 & ~n15985;
  assign n15987 = ~n15912 & n15985;
  assign n15988 = n15912 & ~n15985;
  assign n15989 = ~n15987 & ~n15988;
  assign n15990 = ~n15927 & ~n15929;
  assign n15991 = ~n15928 & ~n15990;
  assign n15992 = n15989 & n15991;
  assign n15993 = ~n15989 & ~n15991;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = n15689 & ~n15994;
  assign n15996 = ~n15979 & ~n15986;
  assign n15997 = ~n15995 & n15996;
  assign n15998 = ~n15912 & ~n15985;
  assign n15999 = n15912 & n15985;
  assign n16000 = ~n15943 & ~n15999;
  assign n16001 = ~n15998 & n16000;
  assign n16002 = n15941 & ~n15944;
  assign n16003 = n16001 & ~n16002;
  assign n16004 = ~n15944 & n15989;
  assign n16005 = ~n15941 & ~n15943;
  assign n16006 = n16004 & ~n16005;
  assign n16007 = ~n16003 & ~n16006;
  assign n16008 = n15722 & n16007;
  assign n16009 = n15768 & ~n15852;
  assign n16010 = n15720 & n16007;
  assign n16011 = n15717 & ~n15994;
  assign n16012 = n15712 & ~n15994;
  assign n16013 = n15706 & ~n15994;
  assign n16014 = n15709 & n16007;
  assign n16015 = n15715 & n16007;
  assign n16016 = ~n16014 & ~n16015;
  assign n16017 = ~n16012 & ~n16013;
  assign n16018 = n16016 & n16017;
  assign n16019 = ~n16008 & ~n16009;
  assign n16020 = ~n16010 & n16019;
  assign n16021 = ~n16011 & n16020;
  assign n16022 = n16018 & n16021;
  assign n16023 = n15997 & n16022;
  assign n16024 = n15649 & ~n16023;
  assign n16025 = P3_REG0_REG_5_ & ~n15649;
  assign n2905 = n16024 | n16025;
  assign n16027 = ~P3_REG3_REG_6_ & n15903;
  assign n16028 = ~P3_REG3_REG_7_ & n16027;
  assign n16029 = P3_REG3_REG_7_ & ~n15969;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = n15675 & ~n16030;
  assign n16032 = P3_REG2_REG_7_ & n15677;
  assign n16033 = P3_REG1_REG_7_ & n15679;
  assign n16034 = P3_REG0_REG_7_ & n15681;
  assign n16035 = ~n16031 & ~n16032;
  assign n16036 = ~n16033 & n16035;
  assign n16037 = ~n16034 & n16036;
  assign n16038 = n15694 & ~n16037;
  assign n16039 = P3_IR_REG_31_ & n14935;
  assign n16040 = P3_IR_REG_6_ & ~P3_IR_REG_31_;
  assign n16041 = ~n16039 & ~n16040;
  assign n16042 = n15656 & ~n16041;
  assign n16043 = ~n14948 & ~n15656;
  assign n16044 = ~n16042 & ~n16043;
  assign n16045 = ~n15667 & ~n16044;
  assign n16046 = ~n15978 & n16044;
  assign n16047 = n15978 & ~n16044;
  assign n16048 = ~n16046 & ~n16047;
  assign n16049 = ~n15988 & ~n16048;
  assign n16050 = ~n15987 & n15991;
  assign n16051 = n16049 & ~n16050;
  assign n16052 = ~n15987 & ~n16046;
  assign n16053 = ~n16047 & n16052;
  assign n16054 = ~n15988 & ~n15991;
  assign n16055 = n16053 & ~n16054;
  assign n16056 = ~n16051 & ~n16055;
  assign n16057 = n15689 & ~n16056;
  assign n16058 = ~n16038 & ~n16045;
  assign n16059 = ~n16057 & n16058;
  assign n16060 = n15944 & ~n15985;
  assign n16061 = ~n15944 & n15985;
  assign n16062 = ~n15912 & ~n16061;
  assign n16063 = ~n16060 & ~n16062;
  assign n16064 = ~n15880 & n16000;
  assign n16065 = ~n15815 & ~n15879;
  assign n16066 = ~n15816 & ~n15819;
  assign n16067 = n16065 & ~n16066;
  assign n16068 = n16064 & ~n16067;
  assign n16069 = n16063 & ~n16068;
  assign n16070 = ~n16048 & n16069;
  assign n16071 = n15978 & n16044;
  assign n16072 = ~n15978 & ~n16044;
  assign n16073 = ~n16071 & ~n16072;
  assign n16074 = ~n16069 & ~n16073;
  assign n16075 = ~n16070 & ~n16074;
  assign n16076 = n15722 & ~n16075;
  assign n16077 = n15768 & ~n15912;
  assign n16078 = n15720 & ~n16075;
  assign n16079 = n15717 & ~n16056;
  assign n16080 = n15712 & ~n16056;
  assign n16081 = n15706 & ~n16056;
  assign n16082 = n15709 & ~n16075;
  assign n16083 = n15715 & ~n16075;
  assign n16084 = ~n16082 & ~n16083;
  assign n16085 = ~n16080 & ~n16081;
  assign n16086 = n16084 & n16085;
  assign n16087 = ~n16076 & ~n16077;
  assign n16088 = ~n16078 & n16087;
  assign n16089 = ~n16079 & n16088;
  assign n16090 = n16086 & n16089;
  assign n16091 = n16059 & n16090;
  assign n16092 = n15649 & ~n16091;
  assign n16093 = P3_REG0_REG_6_ & ~n15649;
  assign n2910 = n16092 | n16093;
  assign n16095 = ~P3_REG3_REG_8_ & n16028;
  assign n16096 = P3_REG3_REG_8_ & ~n16028;
  assign n16097 = ~n16095 & ~n16096;
  assign n16098 = n15675 & ~n16097;
  assign n16099 = P3_REG2_REG_8_ & n15677;
  assign n16100 = P3_REG1_REG_8_ & n15679;
  assign n16101 = P3_REG0_REG_8_ & n15681;
  assign n16102 = ~n16098 & ~n16099;
  assign n16103 = ~n16100 & n16102;
  assign n16104 = ~n16101 & n16103;
  assign n16105 = n15694 & ~n16104;
  assign n16106 = P3_IR_REG_31_ & n14954;
  assign n16107 = P3_IR_REG_7_ & ~P3_IR_REG_31_;
  assign n16108 = ~n16106 & ~n16107;
  assign n16109 = n15656 & ~n16108;
  assign n16110 = ~n14970 & ~n15656;
  assign n16111 = ~n16109 & ~n16110;
  assign n16112 = ~n15667 & ~n16111;
  assign n16113 = ~n16037 & n16111;
  assign n16114 = n16037 & ~n16111;
  assign n16115 = ~n16113 & ~n16114;
  assign n16116 = n15928 & ~n15988;
  assign n16117 = n16052 & ~n16116;
  assign n16118 = ~n16047 & ~n16117;
  assign n16119 = ~n15988 & ~n16047;
  assign n16120 = ~n15929 & n16119;
  assign n16121 = ~n15927 & n16120;
  assign n16122 = ~n16118 & ~n16121;
  assign n16123 = n16115 & n16122;
  assign n16124 = ~n16115 & ~n16122;
  assign n16125 = ~n16123 & ~n16124;
  assign n16126 = n15689 & ~n16125;
  assign n16127 = ~n16105 & ~n16112;
  assign n16128 = ~n16126 & n16127;
  assign n16129 = ~n16037 & ~n16111;
  assign n16130 = n16037 & n16111;
  assign n16131 = ~n16071 & ~n16130;
  assign n16132 = ~n16129 & n16131;
  assign n16133 = n16069 & ~n16072;
  assign n16134 = n16132 & ~n16133;
  assign n16135 = ~n16072 & n16115;
  assign n16136 = ~n16069 & ~n16071;
  assign n16137 = n16135 & ~n16136;
  assign n16138 = ~n16134 & ~n16137;
  assign n16139 = n15722 & n16138;
  assign n16140 = n15768 & ~n15978;
  assign n16141 = n15720 & n16138;
  assign n16142 = n15717 & ~n16125;
  assign n16143 = n15712 & ~n16125;
  assign n16144 = n15706 & ~n16125;
  assign n16145 = n15709 & n16138;
  assign n16146 = n15715 & n16138;
  assign n16147 = ~n16145 & ~n16146;
  assign n16148 = ~n16143 & ~n16144;
  assign n16149 = n16147 & n16148;
  assign n16150 = ~n16139 & ~n16140;
  assign n16151 = ~n16141 & n16150;
  assign n16152 = ~n16142 & n16151;
  assign n16153 = n16149 & n16152;
  assign n16154 = n16128 & n16153;
  assign n16155 = n15649 & ~n16154;
  assign n16156 = P3_REG0_REG_7_ & ~n15649;
  assign n2915 = n16155 | n16156;
  assign n16158 = ~P3_REG3_REG_9_ & ~P3_REG3_REG_8_;
  assign n16159 = n16028 & n16158;
  assign n16160 = P3_REG3_REG_9_ & ~n16095;
  assign n16161 = ~n16159 & ~n16160;
  assign n16162 = n15675 & ~n16161;
  assign n16163 = P3_REG2_REG_9_ & n15677;
  assign n16164 = P3_REG1_REG_9_ & n15679;
  assign n16165 = P3_REG0_REG_9_ & n15681;
  assign n16166 = ~n16162 & ~n16163;
  assign n16167 = ~n16164 & n16166;
  assign n16168 = ~n16165 & n16167;
  assign n16169 = n15694 & ~n16168;
  assign n16170 = P3_IR_REG_31_ & n14980;
  assign n16171 = P3_IR_REG_8_ & ~P3_IR_REG_31_;
  assign n16172 = ~n16170 & ~n16171;
  assign n16173 = n15656 & ~n16172;
  assign n16174 = ~n14997 & ~n15656;
  assign n16175 = ~n16173 & ~n16174;
  assign n16176 = ~n15667 & ~n16175;
  assign n16177 = ~n16104 & n16175;
  assign n16178 = n16104 & ~n16175;
  assign n16179 = ~n16177 & ~n16178;
  assign n16180 = ~n16114 & ~n16179;
  assign n16181 = ~n16113 & n16122;
  assign n16182 = n16180 & ~n16181;
  assign n16183 = ~n16113 & n16179;
  assign n16184 = ~n16114 & ~n16122;
  assign n16185 = n16183 & ~n16184;
  assign n16186 = ~n16182 & ~n16185;
  assign n16187 = n15689 & ~n16186;
  assign n16188 = ~n16169 & ~n16176;
  assign n16189 = ~n16187 & n16188;
  assign n16190 = n16072 & ~n16111;
  assign n16191 = ~n16072 & n16111;
  assign n16192 = ~n16037 & ~n16191;
  assign n16193 = ~n16190 & ~n16192;
  assign n16194 = ~n16069 & n16131;
  assign n16195 = n16193 & ~n16194;
  assign n16196 = ~n16179 & n16195;
  assign n16197 = n16104 & n16175;
  assign n16198 = ~n16104 & ~n16175;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = ~n16195 & ~n16199;
  assign n16201 = ~n16196 & ~n16200;
  assign n16202 = n15722 & ~n16201;
  assign n16203 = n15768 & ~n16037;
  assign n16204 = n15720 & ~n16201;
  assign n16205 = n15717 & ~n16186;
  assign n16206 = n15712 & ~n16186;
  assign n16207 = n15706 & ~n16186;
  assign n16208 = n15709 & ~n16201;
  assign n16209 = n15715 & ~n16201;
  assign n16210 = ~n16208 & ~n16209;
  assign n16211 = ~n16206 & ~n16207;
  assign n16212 = n16210 & n16211;
  assign n16213 = ~n16202 & ~n16203;
  assign n16214 = ~n16204 & n16213;
  assign n16215 = ~n16205 & n16214;
  assign n16216 = n16212 & n16215;
  assign n16217 = n16189 & n16216;
  assign n16218 = n15649 & ~n16217;
  assign n16219 = P3_REG0_REG_8_ & ~n15649;
  assign n2920 = n16218 | n16219;
  assign n16221 = ~P3_REG3_REG_10_ & n16159;
  assign n16222 = P3_REG3_REG_10_ & ~n16159;
  assign n16223 = ~n16221 & ~n16222;
  assign n16224 = n15675 & ~n16223;
  assign n16225 = P3_REG2_REG_10_ & n15677;
  assign n16226 = P3_REG1_REG_10_ & n15679;
  assign n16227 = P3_REG0_REG_10_ & n15681;
  assign n16228 = ~n16224 & ~n16225;
  assign n16229 = ~n16226 & n16228;
  assign n16230 = ~n16227 & n16229;
  assign n16231 = n15694 & ~n16230;
  assign n16232 = P3_IR_REG_31_ & n15003;
  assign n16233 = P3_IR_REG_9_ & ~P3_IR_REG_31_;
  assign n16234 = ~n16232 & ~n16233;
  assign n16235 = n15656 & ~n16234;
  assign n16236 = ~n15019 & ~n15656;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = ~n15667 & ~n16237;
  assign n16239 = ~n16114 & ~n16178;
  assign n16240 = n16118 & n16239;
  assign n16241 = ~n16104 & n16113;
  assign n16242 = ~n16175 & ~n16241;
  assign n16243 = n16104 & ~n16113;
  assign n16244 = ~n16242 & ~n16243;
  assign n16245 = ~n16240 & ~n16244;
  assign n16246 = n16120 & n16239;
  assign n16247 = ~n15927 & n16246;
  assign n16248 = n16245 & ~n16247;
  assign n16249 = ~n16168 & n16237;
  assign n16250 = n16168 & ~n16237;
  assign n16251 = ~n16249 & ~n16250;
  assign n16252 = n16248 & n16251;
  assign n16253 = ~n16248 & ~n16251;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = n15689 & ~n16254;
  assign n16256 = ~n16231 & ~n16238;
  assign n16257 = ~n16255 & n16256;
  assign n16258 = ~n16195 & ~n16197;
  assign n16259 = ~n16198 & ~n16258;
  assign n16260 = ~n16251 & n16259;
  assign n16261 = n16168 & n16237;
  assign n16262 = ~n16168 & ~n16237;
  assign n16263 = ~n16261 & ~n16262;
  assign n16264 = ~n16259 & ~n16263;
  assign n16265 = ~n16260 & ~n16264;
  assign n16266 = n15722 & ~n16265;
  assign n16267 = n15768 & ~n16104;
  assign n16268 = n15717 & ~n16254;
  assign n16269 = n15720 & ~n16265;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = n15712 & ~n16254;
  assign n16272 = n15706 & ~n16254;
  assign n16273 = n15709 & ~n16265;
  assign n16274 = n15715 & ~n16265;
  assign n16275 = ~n16273 & ~n16274;
  assign n16276 = ~n16271 & ~n16272;
  assign n16277 = n16275 & n16276;
  assign n16278 = ~n16266 & ~n16267;
  assign n16279 = n16270 & n16278;
  assign n16280 = n16277 & n16279;
  assign n16281 = n16257 & n16280;
  assign n16282 = n15649 & ~n16281;
  assign n16283 = P3_REG0_REG_9_ & ~n15649;
  assign n2925 = n16282 | n16283;
  assign n16285 = ~P3_REG3_REG_11_ & ~P3_REG3_REG_10_;
  assign n16286 = n16159 & n16285;
  assign n16287 = P3_REG3_REG_11_ & ~n16221;
  assign n16288 = ~n16286 & ~n16287;
  assign n16289 = n15675 & ~n16288;
  assign n16290 = P3_REG2_REG_11_ & n15677;
  assign n16291 = P3_REG1_REG_11_ & n15679;
  assign n16292 = P3_REG0_REG_11_ & n15681;
  assign n16293 = ~n16289 & ~n16290;
  assign n16294 = ~n16291 & n16293;
  assign n16295 = ~n16292 & n16294;
  assign n16296 = n15694 & ~n16295;
  assign n16297 = P3_IR_REG_31_ & n15026;
  assign n16298 = P3_IR_REG_10_ & ~P3_IR_REG_31_;
  assign n16299 = ~n16297 & ~n16298;
  assign n16300 = n15656 & ~n16299;
  assign n16301 = ~n15039 & ~n15656;
  assign n16302 = ~n16300 & ~n16301;
  assign n16303 = ~n15667 & ~n16302;
  assign n16304 = ~n16230 & n16302;
  assign n16305 = n16230 & ~n16302;
  assign n16306 = ~n16304 & ~n16305;
  assign n16307 = ~n16248 & ~n16250;
  assign n16308 = ~n16249 & ~n16307;
  assign n16309 = n16306 & n16308;
  assign n16310 = ~n16306 & ~n16308;
  assign n16311 = ~n16309 & ~n16310;
  assign n16312 = n15689 & ~n16311;
  assign n16313 = ~n16296 & ~n16303;
  assign n16314 = ~n16312 & n16313;
  assign n16315 = ~n16230 & ~n16302;
  assign n16316 = n16230 & n16302;
  assign n16317 = ~n16261 & ~n16316;
  assign n16318 = ~n16315 & n16317;
  assign n16319 = n16259 & ~n16262;
  assign n16320 = n16318 & ~n16319;
  assign n16321 = ~n16262 & n16306;
  assign n16322 = ~n16259 & ~n16261;
  assign n16323 = n16321 & ~n16322;
  assign n16324 = ~n16320 & ~n16323;
  assign n16325 = n15722 & n16324;
  assign n16326 = n15768 & ~n16168;
  assign n16327 = n15717 & ~n16311;
  assign n16328 = n15720 & n16324;
  assign n16329 = ~n16327 & ~n16328;
  assign n16330 = n15712 & ~n16311;
  assign n16331 = n15706 & ~n16311;
  assign n16332 = n15709 & n16324;
  assign n16333 = n15715 & n16324;
  assign n16334 = ~n16332 & ~n16333;
  assign n16335 = ~n16330 & ~n16331;
  assign n16336 = n16334 & n16335;
  assign n16337 = ~n16325 & ~n16326;
  assign n16338 = n16329 & n16337;
  assign n16339 = n16336 & n16338;
  assign n16340 = n16314 & n16339;
  assign n16341 = n15649 & ~n16340;
  assign n16342 = P3_REG0_REG_10_ & ~n15649;
  assign n2930 = n16341 | n16342;
  assign n16344 = ~P3_REG3_REG_12_ & n16286;
  assign n16345 = P3_REG3_REG_12_ & ~n16286;
  assign n16346 = ~n16344 & ~n16345;
  assign n16347 = n15675 & ~n16346;
  assign n16348 = P3_REG2_REG_12_ & n15677;
  assign n16349 = P3_REG1_REG_12_ & n15679;
  assign n16350 = P3_REG0_REG_12_ & n15681;
  assign n16351 = ~n16347 & ~n16348;
  assign n16352 = ~n16349 & n16351;
  assign n16353 = ~n16350 & n16352;
  assign n16354 = n15694 & ~n16353;
  assign n16355 = P3_IR_REG_31_ & n15045;
  assign n16356 = P3_IR_REG_11_ & ~P3_IR_REG_31_;
  assign n16357 = ~n16355 & ~n16356;
  assign n16358 = n15656 & ~n16357;
  assign n16359 = ~n15061 & ~n15656;
  assign n16360 = ~n16358 & ~n16359;
  assign n16361 = ~n15667 & ~n16360;
  assign n16362 = ~n16295 & n16360;
  assign n16363 = n16295 & ~n16360;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = ~n16305 & ~n16364;
  assign n16366 = ~n16304 & n16308;
  assign n16367 = n16365 & ~n16366;
  assign n16368 = ~n16304 & ~n16362;
  assign n16369 = ~n16363 & n16368;
  assign n16370 = ~n16305 & ~n16308;
  assign n16371 = n16369 & ~n16370;
  assign n16372 = ~n16367 & ~n16371;
  assign n16373 = n15689 & ~n16372;
  assign n16374 = ~n16354 & ~n16361;
  assign n16375 = ~n16373 & n16374;
  assign n16376 = ~n16262 & ~n16315;
  assign n16377 = n16198 & n16317;
  assign n16378 = n16376 & ~n16377;
  assign n16379 = ~n16316 & ~n16378;
  assign n16380 = ~n16197 & n16317;
  assign n16381 = ~n16195 & n16380;
  assign n16382 = ~n16379 & ~n16381;
  assign n16383 = ~n16364 & n16382;
  assign n16384 = n16295 & n16360;
  assign n16385 = ~n16295 & ~n16360;
  assign n16386 = ~n16384 & ~n16385;
  assign n16387 = ~n16382 & ~n16386;
  assign n16388 = ~n16383 & ~n16387;
  assign n16389 = n15722 & ~n16388;
  assign n16390 = n15768 & ~n16230;
  assign n16391 = n15720 & ~n16388;
  assign n16392 = n15717 & ~n16372;
  assign n16393 = n15712 & ~n16372;
  assign n16394 = n15706 & ~n16372;
  assign n16395 = ~n16262 & ~n16377;
  assign n16396 = ~n16316 & ~n16395;
  assign n16397 = ~n16315 & ~n16396;
  assign n16398 = ~n16381 & n16397;
  assign n16399 = ~n16364 & n16398;
  assign n16400 = ~n16386 & ~n16398;
  assign n16401 = ~n16399 & ~n16400;
  assign n16402 = n15709 & ~n16401;
  assign n16403 = n15715 & ~n16401;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = ~n16393 & ~n16394;
  assign n16406 = n16404 & n16405;
  assign n16407 = ~n16389 & ~n16390;
  assign n16408 = ~n16391 & n16407;
  assign n16409 = ~n16392 & n16408;
  assign n16410 = n16406 & n16409;
  assign n16411 = n16375 & n16410;
  assign n16412 = n15649 & ~n16411;
  assign n16413 = P3_REG0_REG_11_ & ~n15649;
  assign n2935 = n16412 | n16413;
  assign n16415 = ~P3_REG3_REG_13_ & ~P3_REG3_REG_12_;
  assign n16416 = n16286 & n16415;
  assign n16417 = P3_REG3_REG_13_ & ~n16344;
  assign n16418 = ~n16416 & ~n16417;
  assign n16419 = n15675 & ~n16418;
  assign n16420 = P3_REG2_REG_13_ & n15677;
  assign n16421 = P3_REG1_REG_13_ & n15679;
  assign n16422 = P3_REG0_REG_13_ & n15681;
  assign n16423 = ~n16419 & ~n16420;
  assign n16424 = ~n16421 & n16423;
  assign n16425 = ~n16422 & n16424;
  assign n16426 = n15694 & ~n16425;
  assign n16427 = P3_IR_REG_31_ & n15070;
  assign n16428 = P3_IR_REG_12_ & ~P3_IR_REG_31_;
  assign n16429 = ~n16427 & ~n16428;
  assign n16430 = n15656 & ~n16429;
  assign n16431 = ~n15086 & ~n15656;
  assign n16432 = ~n16430 & ~n16431;
  assign n16433 = ~n15667 & ~n16432;
  assign n16434 = ~n16353 & n16432;
  assign n16435 = n16353 & ~n16432;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = ~n16305 & ~n16363;
  assign n16438 = n16249 & n16437;
  assign n16439 = n16368 & ~n16438;
  assign n16440 = ~n16363 & ~n16439;
  assign n16441 = ~n16250 & n16437;
  assign n16442 = ~n16248 & n16441;
  assign n16443 = ~n16440 & ~n16442;
  assign n16444 = ~n16436 & ~n16443;
  assign n16445 = n16436 & n16443;
  assign n16446 = ~n16444 & ~n16445;
  assign n16447 = n15689 & ~n16446;
  assign n16448 = ~n16426 & ~n16433;
  assign n16449 = ~n16447 & n16448;
  assign n16450 = ~n16382 & ~n16384;
  assign n16451 = ~n16385 & ~n16450;
  assign n16452 = ~n16436 & n16451;
  assign n16453 = n16353 & n16432;
  assign n16454 = ~n16353 & ~n16432;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456 = ~n16451 & ~n16455;
  assign n16457 = ~n16452 & ~n16456;
  assign n16458 = n15722 & ~n16457;
  assign n16459 = n15768 & ~n16295;
  assign n16460 = n15717 & ~n16446;
  assign n16461 = n15720 & ~n16457;
  assign n16462 = ~n16460 & ~n16461;
  assign n16463 = n15712 & ~n16446;
  assign n16464 = n15706 & ~n16446;
  assign n16465 = ~n16384 & ~n16398;
  assign n16466 = ~n16385 & ~n16465;
  assign n16467 = ~n16436 & n16466;
  assign n16468 = ~n16455 & ~n16466;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n15709 & ~n16469;
  assign n16471 = n15715 & ~n16469;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = ~n16463 & ~n16464;
  assign n16474 = n16472 & n16473;
  assign n16475 = ~n16458 & ~n16459;
  assign n16476 = n16462 & n16475;
  assign n16477 = n16474 & n16476;
  assign n16478 = n16449 & n16477;
  assign n16479 = n15649 & ~n16478;
  assign n16480 = P3_REG0_REG_12_ & ~n15649;
  assign n2940 = n16479 | n16480;
  assign n16482 = ~P3_REG3_REG_14_ & n16416;
  assign n16483 = P3_REG3_REG_14_ & ~n16416;
  assign n16484 = ~n16482 & ~n16483;
  assign n16485 = n15675 & ~n16484;
  assign n16486 = P3_REG2_REG_14_ & n15677;
  assign n16487 = P3_REG1_REG_14_ & n15679;
  assign n16488 = P3_REG0_REG_14_ & n15681;
  assign n16489 = ~n16485 & ~n16486;
  assign n16490 = ~n16487 & n16489;
  assign n16491 = ~n16488 & n16490;
  assign n16492 = n15694 & ~n16491;
  assign n16493 = P3_IR_REG_31_ & n15092;
  assign n16494 = P3_IR_REG_13_ & ~P3_IR_REG_31_;
  assign n16495 = ~n16493 & ~n16494;
  assign n16496 = n15656 & ~n16495;
  assign n16497 = ~n15108 & ~n15656;
  assign n16498 = ~n16496 & ~n16497;
  assign n16499 = ~n15667 & ~n16498;
  assign n16500 = ~n16425 & n16498;
  assign n16501 = n16425 & ~n16498;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n16435 & ~n16443;
  assign n16504 = ~n16434 & ~n16503;
  assign n16505 = ~n16502 & ~n16504;
  assign n16506 = n16502 & n16504;
  assign n16507 = ~n16505 & ~n16506;
  assign n16508 = n15689 & ~n16507;
  assign n16509 = ~n16492 & ~n16499;
  assign n16510 = ~n16508 & n16509;
  assign n16511 = ~n16425 & ~n16498;
  assign n16512 = n16425 & n16498;
  assign n16513 = ~n16453 & ~n16512;
  assign n16514 = ~n16511 & n16513;
  assign n16515 = n16451 & ~n16454;
  assign n16516 = n16514 & ~n16515;
  assign n16517 = ~n16454 & n16502;
  assign n16518 = ~n16451 & ~n16453;
  assign n16519 = n16517 & ~n16518;
  assign n16520 = ~n16516 & ~n16519;
  assign n16521 = n15722 & n16520;
  assign n16522 = n15768 & ~n16353;
  assign n16523 = n15717 & ~n16507;
  assign n16524 = n15720 & n16520;
  assign n16525 = ~n16523 & ~n16524;
  assign n16526 = n15712 & ~n16507;
  assign n16527 = n15706 & ~n16507;
  assign n16528 = ~n16454 & n16466;
  assign n16529 = n16514 & ~n16528;
  assign n16530 = ~n16453 & ~n16466;
  assign n16531 = n16517 & ~n16530;
  assign n16532 = ~n16529 & ~n16531;
  assign n16533 = n15709 & n16532;
  assign n16534 = n15715 & n16532;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536 = ~n16526 & ~n16527;
  assign n16537 = n16535 & n16536;
  assign n16538 = ~n16521 & ~n16522;
  assign n16539 = n16525 & n16538;
  assign n16540 = n16537 & n16539;
  assign n16541 = n16510 & n16540;
  assign n16542 = n15649 & ~n16541;
  assign n16543 = P3_REG0_REG_13_ & ~n15649;
  assign n2945 = n16542 | n16543;
  assign n16545 = ~P3_REG3_REG_15_ & ~P3_REG3_REG_14_;
  assign n16546 = n16416 & n16545;
  assign n16547 = P3_REG3_REG_15_ & ~n16482;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = n15675 & ~n16548;
  assign n16550 = P3_REG2_REG_15_ & n15677;
  assign n16551 = P3_REG1_REG_15_ & n15679;
  assign n16552 = P3_REG0_REG_15_ & n15681;
  assign n16553 = ~n16549 & ~n16550;
  assign n16554 = ~n16551 & n16553;
  assign n16555 = ~n16552 & n16554;
  assign n16556 = n15694 & ~n16555;
  assign n16557 = P3_IR_REG_31_ & n15115;
  assign n16558 = P3_IR_REG_14_ & ~P3_IR_REG_31_;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = n15656 & ~n16559;
  assign n16561 = ~n15128 & ~n15656;
  assign n16562 = ~n16560 & ~n16561;
  assign n16563 = ~n15667 & ~n16562;
  assign n16564 = ~n16501 & ~n16504;
  assign n16565 = ~n16500 & ~n16564;
  assign n16566 = ~n16491 & n16562;
  assign n16567 = n16491 & ~n16562;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = n16565 & n16568;
  assign n16570 = ~n16565 & ~n16568;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = n15689 & ~n16571;
  assign n16573 = ~n16556 & ~n16563;
  assign n16574 = ~n16572 & n16573;
  assign n16575 = ~n16454 & ~n16511;
  assign n16576 = n16385 & n16513;
  assign n16577 = n16575 & ~n16576;
  assign n16578 = ~n16512 & ~n16577;
  assign n16579 = ~n16384 & n16513;
  assign n16580 = ~n16382 & n16579;
  assign n16581 = ~n16578 & ~n16580;
  assign n16582 = ~n16568 & n16581;
  assign n16583 = n16568 & ~n16581;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = n15722 & ~n16584;
  assign n16586 = n15768 & ~n16425;
  assign n16587 = n15720 & ~n16584;
  assign n16588 = n15717 & ~n16571;
  assign n16589 = n15712 & ~n16571;
  assign n16590 = n15706 & ~n16571;
  assign n16591 = ~n16398 & n16579;
  assign n16592 = ~n16578 & ~n16591;
  assign n16593 = ~n16568 & n16592;
  assign n16594 = n16568 & ~n16592;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = n15709 & ~n16595;
  assign n16597 = n15715 & ~n16595;
  assign n16598 = ~n16596 & ~n16597;
  assign n16599 = ~n16589 & ~n16590;
  assign n16600 = n16598 & n16599;
  assign n16601 = ~n16585 & ~n16586;
  assign n16602 = ~n16587 & n16601;
  assign n16603 = ~n16588 & n16602;
  assign n16604 = n16600 & n16603;
  assign n16605 = n16574 & n16604;
  assign n16606 = n15649 & ~n16605;
  assign n16607 = P3_REG0_REG_14_ & ~n15649;
  assign n2950 = n16606 | n16607;
  assign n16609 = ~P3_REG3_REG_16_ & n16546;
  assign n16610 = P3_REG3_REG_16_ & ~n16546;
  assign n16611 = ~n16609 & ~n16610;
  assign n16612 = n15675 & ~n16611;
  assign n16613 = P3_REG2_REG_16_ & n15677;
  assign n16614 = P3_REG1_REG_16_ & n15679;
  assign n16615 = P3_REG0_REG_16_ & n15681;
  assign n16616 = ~n16612 & ~n16613;
  assign n16617 = ~n16614 & n16616;
  assign n16618 = ~n16615 & n16617;
  assign n16619 = n15694 & ~n16618;
  assign n16620 = P3_IR_REG_31_ & n15134;
  assign n16621 = P3_IR_REG_15_ & ~P3_IR_REG_31_;
  assign n16622 = ~n16620 & ~n16621;
  assign n16623 = n15656 & ~n16622;
  assign n16624 = ~n15147 & ~n15656;
  assign n16625 = ~n16623 & ~n16624;
  assign n16626 = ~n15667 & ~n16625;
  assign n16627 = ~n16555 & n16625;
  assign n16628 = n16555 & ~n16625;
  assign n16629 = ~n16627 & ~n16628;
  assign n16630 = ~n16565 & ~n16567;
  assign n16631 = ~n16566 & ~n16630;
  assign n16632 = n16629 & n16631;
  assign n16633 = ~n16629 & ~n16631;
  assign n16634 = ~n16632 & ~n16633;
  assign n16635 = n15689 & ~n16634;
  assign n16636 = ~n16619 & ~n16626;
  assign n16637 = ~n16635 & n16636;
  assign n16638 = ~n16491 & ~n16562;
  assign n16639 = n16491 & n16562;
  assign n16640 = ~n16581 & ~n16639;
  assign n16641 = ~n16638 & ~n16640;
  assign n16642 = ~n16629 & n16641;
  assign n16643 = n16629 & ~n16641;
  assign n16644 = ~n16642 & ~n16643;
  assign n16645 = n15722 & ~n16644;
  assign n16646 = n15768 & ~n16491;
  assign n16647 = n15720 & ~n16644;
  assign n16648 = n15717 & ~n16634;
  assign n16649 = n15712 & ~n16634;
  assign n16650 = n15706 & ~n16634;
  assign n16651 = ~n16592 & ~n16639;
  assign n16652 = ~n16638 & ~n16651;
  assign n16653 = ~n16629 & n16652;
  assign n16654 = n16629 & ~n16652;
  assign n16655 = ~n16653 & ~n16654;
  assign n16656 = n15709 & ~n16655;
  assign n16657 = n15715 & ~n16655;
  assign n16658 = ~n16656 & ~n16657;
  assign n16659 = ~n16649 & ~n16650;
  assign n16660 = n16658 & n16659;
  assign n16661 = ~n16645 & ~n16646;
  assign n16662 = ~n16647 & n16661;
  assign n16663 = ~n16648 & n16662;
  assign n16664 = n16660 & n16663;
  assign n16665 = n16637 & n16664;
  assign n16666 = n15649 & ~n16665;
  assign n16667 = P3_REG0_REG_15_ & ~n15649;
  assign n2955 = n16666 | n16667;
  assign n16669 = ~P3_REG3_REG_17_ & ~P3_REG3_REG_16_;
  assign n16670 = n16546 & n16669;
  assign n16671 = P3_REG3_REG_17_ & ~n16609;
  assign n16672 = ~n16670 & ~n16671;
  assign n16673 = n15675 & ~n16672;
  assign n16674 = P3_REG2_REG_17_ & n15677;
  assign n16675 = P3_REG1_REG_17_ & n15679;
  assign n16676 = P3_REG0_REG_17_ & n15681;
  assign n16677 = ~n16673 & ~n16674;
  assign n16678 = ~n16675 & n16677;
  assign n16679 = ~n16676 & n16678;
  assign n16680 = n15694 & ~n16679;
  assign n16681 = P3_IR_REG_31_ & n15167;
  assign n16682 = P3_IR_REG_16_ & ~P3_IR_REG_31_;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = n15656 & ~n16683;
  assign n16685 = ~n15180 & ~n15656;
  assign n16686 = ~n16684 & ~n16685;
  assign n16687 = ~n15667 & ~n16686;
  assign n16688 = ~n16618 & n16686;
  assign n16689 = n16618 & ~n16686;
  assign n16690 = ~n16688 & ~n16689;
  assign n16691 = ~n16628 & ~n16690;
  assign n16692 = ~n16627 & n16631;
  assign n16693 = n16691 & ~n16692;
  assign n16694 = ~n16627 & ~n16688;
  assign n16695 = ~n16689 & n16694;
  assign n16696 = ~n16628 & ~n16631;
  assign n16697 = n16695 & ~n16696;
  assign n16698 = ~n16693 & ~n16697;
  assign n16699 = n15689 & ~n16698;
  assign n16700 = ~n16680 & ~n16687;
  assign n16701 = ~n16699 & n16700;
  assign n16702 = ~n16555 & ~n16625;
  assign n16703 = n16555 & n16625;
  assign n16704 = ~n16641 & ~n16703;
  assign n16705 = ~n16702 & ~n16704;
  assign n16706 = ~n16690 & n16705;
  assign n16707 = n16618 & n16686;
  assign n16708 = ~n16618 & ~n16686;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = ~n16705 & ~n16709;
  assign n16711 = ~n16706 & ~n16710;
  assign n16712 = n15722 & ~n16711;
  assign n16713 = n15768 & ~n16555;
  assign n16714 = n15720 & ~n16711;
  assign n16715 = n15717 & ~n16698;
  assign n16716 = n15712 & ~n16698;
  assign n16717 = n15706 & ~n16698;
  assign n16718 = ~n16652 & ~n16703;
  assign n16719 = ~n16702 & ~n16718;
  assign n16720 = ~n16690 & n16719;
  assign n16721 = ~n16709 & ~n16719;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = n15709 & ~n16722;
  assign n16724 = n15715 & ~n16722;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = ~n16716 & ~n16717;
  assign n16727 = n16725 & n16726;
  assign n16728 = ~n16712 & ~n16713;
  assign n16729 = ~n16714 & n16728;
  assign n16730 = ~n16715 & n16729;
  assign n16731 = n16727 & n16730;
  assign n16732 = n16701 & n16731;
  assign n16733 = n15649 & ~n16732;
  assign n16734 = P3_REG0_REG_16_ & ~n15649;
  assign n2960 = n16733 | n16734;
  assign n16736 = ~P3_REG3_REG_18_ & n16670;
  assign n16737 = P3_REG3_REG_18_ & ~n16670;
  assign n16738 = ~n16736 & ~n16737;
  assign n16739 = n15675 & ~n16738;
  assign n16740 = P3_REG2_REG_18_ & n15677;
  assign n16741 = P3_REG1_REG_18_ & n15679;
  assign n16742 = P3_REG0_REG_18_ & n15681;
  assign n16743 = ~n16739 & ~n16740;
  assign n16744 = ~n16741 & n16743;
  assign n16745 = ~n16742 & n16744;
  assign n16746 = n15694 & ~n16745;
  assign n16747 = P3_IR_REG_31_ & n15186;
  assign n16748 = P3_IR_REG_17_ & ~P3_IR_REG_31_;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = n15656 & ~n16749;
  assign n16751 = ~n15199 & ~n15656;
  assign n16752 = ~n16750 & ~n16751;
  assign n16753 = ~n15667 & ~n16752;
  assign n16754 = ~n16679 & n16752;
  assign n16755 = n16679 & ~n16752;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = ~n16628 & ~n16689;
  assign n16758 = n16566 & n16757;
  assign n16759 = n16694 & ~n16758;
  assign n16760 = ~n16689 & ~n16759;
  assign n16761 = ~n16567 & n16757;
  assign n16762 = ~n16565 & n16761;
  assign n16763 = ~n16760 & ~n16762;
  assign n16764 = ~n16756 & ~n16763;
  assign n16765 = n16756 & n16763;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = n15689 & ~n16766;
  assign n16768 = ~n16746 & ~n16753;
  assign n16769 = ~n16767 & n16768;
  assign n16770 = ~n16679 & ~n16752;
  assign n16771 = n16679 & n16752;
  assign n16772 = ~n16707 & ~n16771;
  assign n16773 = ~n16770 & n16772;
  assign n16774 = n16705 & ~n16708;
  assign n16775 = n16773 & ~n16774;
  assign n16776 = ~n16708 & n16756;
  assign n16777 = ~n16705 & ~n16707;
  assign n16778 = n16776 & ~n16777;
  assign n16779 = ~n16775 & ~n16778;
  assign n16780 = n15722 & n16779;
  assign n16781 = n15768 & ~n16618;
  assign n16782 = n15717 & ~n16766;
  assign n16783 = n15720 & n16779;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = n15712 & ~n16766;
  assign n16786 = n15706 & ~n16766;
  assign n16787 = ~n16708 & n16719;
  assign n16788 = n16773 & ~n16787;
  assign n16789 = ~n16707 & ~n16719;
  assign n16790 = n16776 & ~n16789;
  assign n16791 = ~n16788 & ~n16790;
  assign n16792 = n15709 & n16791;
  assign n16793 = n15715 & n16791;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = ~n16785 & ~n16786;
  assign n16796 = n16794 & n16795;
  assign n16797 = ~n16780 & ~n16781;
  assign n16798 = n16784 & n16797;
  assign n16799 = n16796 & n16798;
  assign n16800 = n16769 & n16799;
  assign n16801 = n15649 & ~n16800;
  assign n16802 = P3_REG0_REG_17_ & ~n15649;
  assign n2965 = n16801 | n16802;
  assign n16804 = ~P3_REG3_REG_18_ & ~P3_REG3_REG_19_;
  assign n16805 = n16670 & n16804;
  assign n16806 = P3_REG3_REG_19_ & ~n16736;
  assign n16807 = ~n16805 & ~n16806;
  assign n16808 = n15675 & ~n16807;
  assign n16809 = P3_REG2_REG_19_ & n15677;
  assign n16810 = P3_REG1_REG_19_ & n15679;
  assign n16811 = P3_REG0_REG_19_ & n15681;
  assign n16812 = ~n16808 & ~n16809;
  assign n16813 = ~n16810 & n16812;
  assign n16814 = ~n16811 & n16813;
  assign n16815 = n15694 & ~n16814;
  assign n16816 = P3_IR_REG_31_ & n15206;
  assign n16817 = P3_IR_REG_18_ & ~P3_IR_REG_31_;
  assign n16818 = ~n16816 & ~n16817;
  assign n16819 = n15656 & ~n16818;
  assign n16820 = ~n15219 & ~n15656;
  assign n16821 = ~n16819 & ~n16820;
  assign n16822 = ~n15667 & ~n16821;
  assign n16823 = ~n16745 & n16821;
  assign n16824 = n16745 & ~n16821;
  assign n16825 = ~n16823 & ~n16824;
  assign n16826 = ~n16755 & ~n16763;
  assign n16827 = ~n16754 & ~n16826;
  assign n16828 = ~n16825 & ~n16827;
  assign n16829 = n16825 & n16827;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = n15689 & ~n16830;
  assign n16832 = ~n16815 & ~n16822;
  assign n16833 = ~n16831 & n16832;
  assign n16834 = n16708 & ~n16752;
  assign n16835 = ~n16708 & n16752;
  assign n16836 = ~n16679 & ~n16835;
  assign n16837 = ~n16834 & ~n16836;
  assign n16838 = ~n16705 & n16772;
  assign n16839 = n16837 & ~n16838;
  assign n16840 = ~n16825 & n16839;
  assign n16841 = n16745 & n16821;
  assign n16842 = ~n16745 & ~n16821;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = ~n16839 & ~n16843;
  assign n16845 = ~n16840 & ~n16844;
  assign n16846 = n15722 & ~n16845;
  assign n16847 = n15768 & ~n16679;
  assign n16848 = n15720 & ~n16845;
  assign n16849 = n15717 & ~n16830;
  assign n16850 = n15712 & ~n16830;
  assign n16851 = n15706 & ~n16830;
  assign n16852 = ~n16719 & n16772;
  assign n16853 = n16837 & ~n16852;
  assign n16854 = ~n16825 & n16853;
  assign n16855 = ~n16843 & ~n16853;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = n15709 & ~n16856;
  assign n16858 = n15715 & ~n16856;
  assign n16859 = ~n16857 & ~n16858;
  assign n16860 = ~n16850 & ~n16851;
  assign n16861 = n16859 & n16860;
  assign n16862 = ~n16846 & ~n16847;
  assign n16863 = ~n16848 & n16862;
  assign n16864 = ~n16849 & n16863;
  assign n16865 = n16861 & n16864;
  assign n16866 = n16833 & n16865;
  assign n16867 = n15649 & ~n16866;
  assign n16868 = P3_REG0_REG_18_ & ~n15649;
  assign n2970 = n16867 | n16868;
  assign n16870 = ~P3_REG3_REG_20_ & n16805;
  assign n16871 = P3_REG3_REG_20_ & ~n16805;
  assign n16872 = ~n16870 & ~n16871;
  assign n16873 = n15675 & ~n16872;
  assign n16874 = P3_REG0_REG_20_ & n15681;
  assign n16875 = P3_REG1_REG_20_ & n15679;
  assign n16876 = P3_REG2_REG_20_ & n15677;
  assign n16877 = ~n16873 & ~n16874;
  assign n16878 = ~n16875 & n16877;
  assign n16879 = ~n16876 & n16878;
  assign n16880 = n15694 & ~n16879;
  assign n16881 = ~n15634 & n15656;
  assign n16882 = ~n15238 & ~n15656;
  assign n16883 = ~n16881 & ~n16882;
  assign n16884 = ~n15667 & ~n16883;
  assign n16885 = ~n16814 & n16883;
  assign n16886 = n16814 & ~n16883;
  assign n16887 = ~n16885 & ~n16886;
  assign n16888 = ~n16745 & ~n16827;
  assign n16889 = n16821 & ~n16827;
  assign n16890 = ~n16888 & ~n16889;
  assign n16891 = ~n16823 & n16890;
  assign n16892 = ~n16887 & ~n16891;
  assign n16893 = n16887 & n16891;
  assign n16894 = ~n16892 & ~n16893;
  assign n16895 = n15689 & ~n16894;
  assign n16896 = ~n16880 & ~n16884;
  assign n16897 = ~n16895 & n16896;
  assign n16898 = ~n16839 & ~n16841;
  assign n16899 = ~n16842 & ~n16898;
  assign n16900 = ~n16887 & n16899;
  assign n16901 = n16814 & n16883;
  assign n16902 = ~n16814 & ~n16883;
  assign n16903 = ~n16901 & ~n16902;
  assign n16904 = ~n16899 & ~n16903;
  assign n16905 = ~n16900 & ~n16904;
  assign n16906 = n15722 & ~n16905;
  assign n16907 = n15768 & ~n16745;
  assign n16908 = n15720 & ~n16905;
  assign n16909 = n15717 & ~n16894;
  assign n16910 = n15712 & ~n16894;
  assign n16911 = n15706 & ~n16894;
  assign n16912 = ~n16841 & ~n16853;
  assign n16913 = ~n16842 & ~n16912;
  assign n16914 = ~n16887 & n16913;
  assign n16915 = ~n16903 & ~n16913;
  assign n16916 = ~n16914 & ~n16915;
  assign n16917 = n15709 & ~n16916;
  assign n16918 = n15715 & ~n16916;
  assign n16919 = ~n16917 & ~n16918;
  assign n16920 = ~n16910 & ~n16911;
  assign n16921 = n16919 & n16920;
  assign n16922 = ~n16906 & ~n16907;
  assign n16923 = ~n16908 & n16922;
  assign n16924 = ~n16909 & n16923;
  assign n16925 = n16921 & n16924;
  assign n16926 = n16897 & n16925;
  assign n16927 = n15649 & ~n16926;
  assign n16928 = P3_REG0_REG_19_ & ~n15649;
  assign n2975 = n16927 | n16928;
  assign n16930 = ~P3_REG3_REG_20_ & ~P3_REG3_REG_21_;
  assign n16931 = n16805 & n16930;
  assign n16932 = P3_REG3_REG_21_ & ~n16870;
  assign n16933 = ~n16931 & ~n16932;
  assign n16934 = n15675 & ~n16933;
  assign n16935 = P3_REG0_REG_21_ & n15681;
  assign n16936 = P3_REG1_REG_21_ & n15679;
  assign n16937 = P3_REG2_REG_21_ & n15677;
  assign n16938 = ~n16934 & ~n16935;
  assign n16939 = ~n16936 & n16938;
  assign n16940 = ~n16937 & n16939;
  assign n16941 = n15694 & ~n16940;
  assign n16942 = ~n15260 & ~n15656;
  assign n16943 = ~n15667 & n16942;
  assign n16944 = ~n16879 & ~n16942;
  assign n16945 = n16879 & n16942;
  assign n16946 = ~n16944 & ~n16945;
  assign n16947 = ~n16886 & ~n16891;
  assign n16948 = ~n16885 & ~n16947;
  assign n16949 = ~n16946 & ~n16948;
  assign n16950 = n16946 & n16948;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = n15689 & ~n16951;
  assign n16953 = ~n16941 & ~n16943;
  assign n16954 = ~n16952 & n16953;
  assign n16955 = ~n16879 & n16942;
  assign n16956 = n16879 & ~n16942;
  assign n16957 = ~n16901 & ~n16956;
  assign n16958 = ~n16955 & n16957;
  assign n16959 = n16899 & ~n16902;
  assign n16960 = n16958 & ~n16959;
  assign n16961 = ~n16902 & n16946;
  assign n16962 = ~n16899 & ~n16901;
  assign n16963 = n16961 & ~n16962;
  assign n16964 = ~n16960 & ~n16963;
  assign n16965 = n15722 & n16964;
  assign n16966 = n15768 & ~n16814;
  assign n16967 = n15720 & n16964;
  assign n16968 = n15717 & ~n16951;
  assign n16969 = n15712 & ~n16951;
  assign n16970 = n15706 & ~n16951;
  assign n16971 = ~n16902 & n16913;
  assign n16972 = n16958 & ~n16971;
  assign n16973 = ~n16901 & ~n16913;
  assign n16974 = n16961 & ~n16973;
  assign n16975 = ~n16972 & ~n16974;
  assign n16976 = n15709 & n16975;
  assign n16977 = n15715 & n16975;
  assign n16978 = ~n16976 & ~n16977;
  assign n16979 = ~n16969 & ~n16970;
  assign n16980 = n16978 & n16979;
  assign n16981 = ~n16965 & ~n16966;
  assign n16982 = ~n16967 & n16981;
  assign n16983 = ~n16968 & n16982;
  assign n16984 = n16980 & n16983;
  assign n16985 = n16954 & n16984;
  assign n16986 = n15649 & ~n16985;
  assign n16987 = P3_REG0_REG_20_ & ~n15649;
  assign n2980 = n16986 | n16987;
  assign n16989 = ~P3_REG3_REG_22_ & n16931;
  assign n16990 = P3_REG3_REG_22_ & ~n16931;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = n15675 & ~n16991;
  assign n16993 = P3_REG0_REG_22_ & n15681;
  assign n16994 = P3_REG1_REG_22_ & n15679;
  assign n16995 = P3_REG2_REG_22_ & n15677;
  assign n16996 = ~n16992 & ~n16993;
  assign n16997 = ~n16994 & n16996;
  assign n16998 = ~n16995 & n16997;
  assign n16999 = n15694 & ~n16998;
  assign n17000 = ~n15279 & ~n15656;
  assign n17001 = ~n15667 & n17000;
  assign n17002 = ~n16945 & ~n16948;
  assign n17003 = ~n16944 & ~n17002;
  assign n17004 = ~n16940 & ~n17000;
  assign n17005 = n16940 & n17000;
  assign n17006 = ~n17004 & ~n17005;
  assign n17007 = n17003 & n17006;
  assign n17008 = ~n17003 & ~n17006;
  assign n17009 = ~n17007 & ~n17008;
  assign n17010 = n15689 & ~n17009;
  assign n17011 = ~n16999 & ~n17001;
  assign n17012 = ~n17010 & n17011;
  assign n17013 = ~n16899 & n16957;
  assign n17014 = ~n16902 & ~n16942;
  assign n17015 = n16902 & n16942;
  assign n17016 = n16879 & ~n17015;
  assign n17017 = ~n17014 & ~n17016;
  assign n17018 = ~n17013 & ~n17017;
  assign n17019 = ~n17006 & ~n17018;
  assign n17020 = n17006 & ~n17017;
  assign n17021 = ~n17013 & n17020;
  assign n17022 = ~n17019 & ~n17021;
  assign n17023 = n15722 & n17022;
  assign n17024 = n15768 & ~n16879;
  assign n17025 = n15720 & n17022;
  assign n17026 = n15717 & ~n17009;
  assign n17027 = n15712 & ~n17009;
  assign n17028 = n15706 & ~n17009;
  assign n17029 = ~n16913 & n16957;
  assign n17030 = ~n17017 & ~n17029;
  assign n17031 = ~n17006 & ~n17030;
  assign n17032 = n17020 & ~n17029;
  assign n17033 = ~n17031 & ~n17032;
  assign n17034 = n15709 & n17033;
  assign n17035 = n15715 & n17033;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = ~n17027 & ~n17028;
  assign n17038 = n17036 & n17037;
  assign n17039 = ~n17023 & ~n17024;
  assign n17040 = ~n17025 & n17039;
  assign n17041 = ~n17026 & n17040;
  assign n17042 = n17038 & n17041;
  assign n17043 = n17012 & n17042;
  assign n17044 = n15649 & ~n17043;
  assign n17045 = P3_REG0_REG_21_ & ~n15649;
  assign n2985 = n17044 | n17045;
  assign n17047 = ~P3_REG3_REG_22_ & ~P3_REG3_REG_23_;
  assign n17048 = n16931 & n17047;
  assign n17049 = P3_REG3_REG_23_ & ~n16989;
  assign n17050 = ~n17048 & ~n17049;
  assign n17051 = n15675 & ~n17050;
  assign n17052 = P3_REG0_REG_23_ & n15681;
  assign n17053 = P3_REG1_REG_23_ & n15679;
  assign n17054 = P3_REG2_REG_23_ & n15677;
  assign n17055 = ~n17051 & ~n17052;
  assign n17056 = ~n17053 & n17055;
  assign n17057 = ~n17054 & n17056;
  assign n17058 = n15694 & ~n17057;
  assign n17059 = ~n15299 & ~n15656;
  assign n17060 = ~n15667 & n17059;
  assign n17061 = ~n16998 & ~n17059;
  assign n17062 = n16998 & n17059;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = ~n17003 & ~n17005;
  assign n17065 = ~n17004 & ~n17064;
  assign n17066 = n17063 & n17065;
  assign n17067 = ~n17063 & ~n17065;
  assign n17068 = ~n17066 & ~n17067;
  assign n17069 = n15689 & ~n17068;
  assign n17070 = ~n17058 & ~n17060;
  assign n17071 = ~n17069 & n17070;
  assign n17072 = n16940 & ~n17000;
  assign n17073 = n16842 & n16957;
  assign n17074 = ~n17017 & ~n17073;
  assign n17075 = ~n17072 & ~n17074;
  assign n17076 = ~n16940 & n17000;
  assign n17077 = ~n17075 & ~n17076;
  assign n17078 = ~n16841 & n16957;
  assign n17079 = ~n17072 & n17078;
  assign n17080 = ~n16839 & n17079;
  assign n17081 = n17077 & ~n17080;
  assign n17082 = ~n17063 & n17081;
  assign n17083 = n17063 & ~n17081;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = n15722 & ~n17084;
  assign n17086 = n15768 & ~n16940;
  assign n17087 = n15720 & ~n17084;
  assign n17088 = n15717 & ~n17068;
  assign n17089 = n15712 & ~n17068;
  assign n17090 = n15706 & ~n17068;
  assign n17091 = ~n16853 & n17079;
  assign n17092 = n17077 & ~n17091;
  assign n17093 = ~n17063 & n17092;
  assign n17094 = n17063 & ~n17092;
  assign n17095 = ~n17093 & ~n17094;
  assign n17096 = n15709 & ~n17095;
  assign n17097 = n15715 & ~n17095;
  assign n17098 = ~n17096 & ~n17097;
  assign n17099 = ~n17089 & ~n17090;
  assign n17100 = n17098 & n17099;
  assign n17101 = ~n17085 & ~n17086;
  assign n17102 = ~n17087 & n17101;
  assign n17103 = ~n17088 & n17102;
  assign n17104 = n17100 & n17103;
  assign n17105 = n17071 & n17104;
  assign n17106 = n15649 & ~n17105;
  assign n17107 = P3_REG0_REG_22_ & ~n15649;
  assign n2990 = n17106 | n17107;
  assign n17109 = ~P3_REG3_REG_24_ & n17048;
  assign n17110 = P3_REG3_REG_24_ & ~n17048;
  assign n17111 = ~n17109 & ~n17110;
  assign n17112 = n15675 & ~n17111;
  assign n17113 = P3_REG0_REG_24_ & n15681;
  assign n17114 = P3_REG1_REG_24_ & n15679;
  assign n17115 = P3_REG2_REG_24_ & n15677;
  assign n17116 = ~n17112 & ~n17113;
  assign n17117 = ~n17114 & n17116;
  assign n17118 = ~n17115 & n17117;
  assign n17119 = n15694 & ~n17118;
  assign n17120 = ~n15318 & ~n15656;
  assign n17121 = ~n15667 & n17120;
  assign n17122 = ~n17057 & ~n17120;
  assign n17123 = n17057 & n17120;
  assign n17124 = ~n17122 & ~n17123;
  assign n17125 = ~n17062 & ~n17124;
  assign n17126 = ~n17061 & n17065;
  assign n17127 = n17125 & ~n17126;
  assign n17128 = ~n17061 & ~n17122;
  assign n17129 = ~n17123 & n17128;
  assign n17130 = ~n17062 & ~n17065;
  assign n17131 = n17129 & ~n17130;
  assign n17132 = ~n17127 & ~n17131;
  assign n17133 = n15689 & ~n17132;
  assign n17134 = ~n17119 & ~n17121;
  assign n17135 = ~n17133 & n17134;
  assign n17136 = ~n16998 & n17059;
  assign n17137 = n16998 & ~n17059;
  assign n17138 = ~n17081 & ~n17137;
  assign n17139 = ~n17136 & ~n17138;
  assign n17140 = ~n17124 & n17139;
  assign n17141 = n17124 & ~n17139;
  assign n17142 = ~n17140 & ~n17141;
  assign n17143 = n15722 & ~n17142;
  assign n17144 = n15768 & ~n16998;
  assign n17145 = n15720 & ~n17142;
  assign n17146 = n15717 & ~n17132;
  assign n17147 = n15712 & ~n17132;
  assign n17148 = n15706 & ~n17132;
  assign n17149 = ~n17092 & ~n17137;
  assign n17150 = ~n17136 & ~n17149;
  assign n17151 = ~n17124 & n17150;
  assign n17152 = n17124 & ~n17150;
  assign n17153 = ~n17151 & ~n17152;
  assign n17154 = n15709 & ~n17153;
  assign n17155 = n15715 & ~n17153;
  assign n17156 = ~n17154 & ~n17155;
  assign n17157 = ~n17147 & ~n17148;
  assign n17158 = n17156 & n17157;
  assign n17159 = ~n17143 & ~n17144;
  assign n17160 = ~n17145 & n17159;
  assign n17161 = ~n17146 & n17160;
  assign n17162 = n17158 & n17161;
  assign n17163 = n17135 & n17162;
  assign n17164 = n15649 & ~n17163;
  assign n17165 = P3_REG0_REG_23_ & ~n15649;
  assign n2995 = n17164 | n17165;
  assign n17167 = ~P3_REG3_REG_24_ & ~P3_REG3_REG_25_;
  assign n17168 = n17048 & n17167;
  assign n17169 = P3_REG3_REG_25_ & ~n17109;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = n15675 & ~n17170;
  assign n17172 = P3_REG0_REG_25_ & n15681;
  assign n17173 = P3_REG1_REG_25_ & n15679;
  assign n17174 = P3_REG2_REG_25_ & n15677;
  assign n17175 = ~n17171 & ~n17172;
  assign n17176 = ~n17173 & n17175;
  assign n17177 = ~n17174 & n17176;
  assign n17178 = n15694 & ~n17177;
  assign n17179 = ~n15341 & ~n15656;
  assign n17180 = ~n15667 & n17179;
  assign n17181 = ~n17118 & ~n17179;
  assign n17182 = n17118 & n17179;
  assign n17183 = ~n17181 & ~n17182;
  assign n17184 = ~n17062 & ~n17123;
  assign n17185 = n17004 & n17184;
  assign n17186 = n17128 & ~n17185;
  assign n17187 = ~n17123 & ~n17186;
  assign n17188 = ~n17005 & n17184;
  assign n17189 = ~n17003 & n17188;
  assign n17190 = ~n17187 & ~n17189;
  assign n17191 = ~n17183 & ~n17190;
  assign n17192 = n17183 & n17190;
  assign n17193 = ~n17191 & ~n17192;
  assign n17194 = n15689 & ~n17193;
  assign n17195 = ~n17178 & ~n17180;
  assign n17196 = ~n17194 & n17195;
  assign n17197 = ~n17057 & n17120;
  assign n17198 = n17057 & ~n17120;
  assign n17199 = ~n17139 & ~n17198;
  assign n17200 = ~n17197 & ~n17199;
  assign n17201 = ~n17183 & n17200;
  assign n17202 = n17118 & ~n17179;
  assign n17203 = ~n17118 & n17179;
  assign n17204 = ~n17202 & ~n17203;
  assign n17205 = ~n17200 & ~n17204;
  assign n17206 = ~n17201 & ~n17205;
  assign n17207 = n15722 & ~n17206;
  assign n17208 = n15768 & ~n17057;
  assign n17209 = n15717 & ~n17193;
  assign n17210 = n15720 & ~n17206;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = n15712 & ~n17193;
  assign n17213 = n15706 & ~n17193;
  assign n17214 = ~n17150 & ~n17198;
  assign n17215 = ~n17197 & ~n17214;
  assign n17216 = ~n17183 & n17215;
  assign n17217 = ~n17204 & ~n17215;
  assign n17218 = ~n17216 & ~n17217;
  assign n17219 = n15709 & ~n17218;
  assign n17220 = n15715 & ~n17218;
  assign n17221 = ~n17219 & ~n17220;
  assign n17222 = ~n17212 & ~n17213;
  assign n17223 = n17221 & n17222;
  assign n17224 = ~n17207 & ~n17208;
  assign n17225 = n17211 & n17224;
  assign n17226 = n17223 & n17225;
  assign n17227 = n17196 & n17226;
  assign n17228 = n15649 & ~n17227;
  assign n17229 = P3_REG0_REG_24_ & ~n15649;
  assign n3000 = n17228 | n17229;
  assign n17231 = ~P3_REG3_REG_26_ & n17168;
  assign n17232 = P3_REG3_REG_26_ & ~n17168;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = n15675 & ~n17233;
  assign n17235 = P3_REG0_REG_26_ & n15681;
  assign n17236 = P3_REG1_REG_26_ & n15679;
  assign n17237 = P3_REG2_REG_26_ & n15677;
  assign n17238 = ~n17234 & ~n17235;
  assign n17239 = ~n17236 & n17238;
  assign n17240 = ~n17237 & n17239;
  assign n17241 = n15694 & ~n17240;
  assign n17242 = ~n15360 & ~n15656;
  assign n17243 = ~n15667 & n17242;
  assign n17244 = ~n17177 & ~n17242;
  assign n17245 = n17177 & n17242;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = ~n17182 & ~n17190;
  assign n17248 = ~n17181 & ~n17247;
  assign n17249 = ~n17246 & ~n17248;
  assign n17250 = n17246 & n17248;
  assign n17251 = ~n17249 & ~n17250;
  assign n17252 = n15689 & ~n17251;
  assign n17253 = ~n17241 & ~n17243;
  assign n17254 = ~n17252 & n17253;
  assign n17255 = ~n17200 & ~n17202;
  assign n17256 = ~n17203 & ~n17255;
  assign n17257 = ~n17246 & n17256;
  assign n17258 = n17177 & ~n17242;
  assign n17259 = ~n17177 & n17242;
  assign n17260 = ~n17258 & ~n17259;
  assign n17261 = ~n17256 & ~n17260;
  assign n17262 = ~n17257 & ~n17261;
  assign n17263 = n15722 & ~n17262;
  assign n17264 = n15768 & ~n17118;
  assign n17265 = n15717 & ~n17251;
  assign n17266 = n15720 & ~n17262;
  assign n17267 = ~n17265 & ~n17266;
  assign n17268 = n15712 & ~n17251;
  assign n17269 = n15706 & ~n17251;
  assign n17270 = ~n17202 & ~n17215;
  assign n17271 = ~n17203 & ~n17270;
  assign n17272 = ~n17246 & n17271;
  assign n17273 = ~n17260 & ~n17271;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = n15709 & ~n17274;
  assign n17276 = n15715 & ~n17274;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = ~n17268 & ~n17269;
  assign n17279 = n17277 & n17278;
  assign n17280 = ~n17263 & ~n17264;
  assign n17281 = n17267 & n17280;
  assign n17282 = n17279 & n17281;
  assign n17283 = n17254 & n17282;
  assign n17284 = n15649 & ~n17283;
  assign n17285 = P3_REG0_REG_25_ & ~n15649;
  assign n3005 = n17284 | n17285;
  assign n17287 = P3_REG1_REG_27_ & n15679;
  assign n17288 = P3_REG0_REG_27_ & n15681;
  assign n17289 = P3_REG2_REG_27_ & n15677;
  assign n17290 = ~P3_REG3_REG_26_ & ~P3_REG3_REG_27_;
  assign n17291 = n17168 & n17290;
  assign n17292 = P3_REG3_REG_27_ & ~n17231;
  assign n17293 = ~n17291 & ~n17292;
  assign n17294 = n15675 & ~n17293;
  assign n17295 = ~n17287 & ~n17288;
  assign n17296 = ~n17289 & n17295;
  assign n17297 = ~n17294 & n17296;
  assign n17298 = n15694 & ~n17297;
  assign n17299 = ~n15380 & ~n15656;
  assign n17300 = ~n15667 & n17299;
  assign n17301 = ~n17240 & ~n17299;
  assign n17302 = n17240 & n17299;
  assign n17303 = ~n17301 & ~n17302;
  assign n17304 = ~n17245 & ~n17248;
  assign n17305 = ~n17244 & ~n17304;
  assign n17306 = n17303 & n17305;
  assign n17307 = ~n17303 & ~n17305;
  assign n17308 = ~n17306 & ~n17307;
  assign n17309 = n15689 & ~n17308;
  assign n17310 = ~n17298 & ~n17300;
  assign n17311 = ~n17309 & n17310;
  assign n17312 = n17256 & ~n17259;
  assign n17313 = ~n17240 & n17299;
  assign n17314 = ~n17258 & n17299;
  assign n17315 = ~n17240 & ~n17258;
  assign n17316 = ~n17314 & ~n17315;
  assign n17317 = ~n17312 & ~n17313;
  assign n17318 = ~n17316 & n17317;
  assign n17319 = ~n17256 & ~n17258;
  assign n17320 = ~n17259 & ~n17319;
  assign n17321 = n17303 & n17320;
  assign n17322 = ~n17318 & ~n17321;
  assign n17323 = n15722 & n17322;
  assign n17324 = n15768 & ~n17177;
  assign n17325 = n15717 & ~n17308;
  assign n17326 = n15720 & n17322;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = n15712 & ~n17308;
  assign n17329 = n15706 & ~n17308;
  assign n17330 = ~n17259 & n17271;
  assign n17331 = ~n17313 & ~n17330;
  assign n17332 = ~n17316 & n17331;
  assign n17333 = ~n17258 & ~n17271;
  assign n17334 = ~n17259 & ~n17333;
  assign n17335 = n17303 & n17334;
  assign n17336 = ~n17332 & ~n17335;
  assign n17337 = n15709 & n17336;
  assign n17338 = n15715 & n17336;
  assign n17339 = ~n17337 & ~n17338;
  assign n17340 = ~n17328 & ~n17329;
  assign n17341 = n17339 & n17340;
  assign n17342 = ~n17323 & ~n17324;
  assign n17343 = n17327 & n17342;
  assign n17344 = n17341 & n17343;
  assign n17345 = n17311 & n17344;
  assign n17346 = n15649 & ~n17345;
  assign n17347 = P3_REG0_REG_26_ & ~n15649;
  assign n3010 = n17346 | n17347;
  assign n17349 = ~P3_REG3_REG_28_ & n17291;
  assign n17350 = P3_REG3_REG_28_ & ~n17291;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = n15675 & ~n17351;
  assign n17353 = P3_REG0_REG_28_ & n15681;
  assign n17354 = P3_REG1_REG_28_ & n15679;
  assign n17355 = P3_REG2_REG_28_ & n15677;
  assign n17356 = ~n17352 & ~n17353;
  assign n17357 = ~n17354 & n17356;
  assign n17358 = ~n17355 & n17357;
  assign n17359 = n15694 & ~n17358;
  assign n17360 = ~n15399 & ~n15656;
  assign n17361 = ~n15667 & n17360;
  assign n17362 = ~n17297 & ~n17360;
  assign n17363 = n17297 & n17360;
  assign n17364 = ~n17362 & ~n17363;
  assign n17365 = ~n17302 & ~n17364;
  assign n17366 = ~n17301 & n17305;
  assign n17367 = n17365 & ~n17366;
  assign n17368 = ~n17301 & n17364;
  assign n17369 = ~n17302 & ~n17305;
  assign n17370 = n17368 & ~n17369;
  assign n17371 = ~n17367 & ~n17370;
  assign n17372 = n15689 & ~n17371;
  assign n17373 = ~n17359 & ~n17361;
  assign n17374 = ~n17372 & n17373;
  assign n17375 = ~n17203 & ~n17259;
  assign n17376 = ~n17316 & ~n17375;
  assign n17377 = n17255 & ~n17316;
  assign n17378 = ~n17376 & ~n17377;
  assign n17379 = ~n17313 & n17378;
  assign n17380 = ~n17364 & n17379;
  assign n17381 = n17364 & ~n17379;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = n15722 & ~n17382;
  assign n17384 = n15768 & ~n17240;
  assign n17385 = n15717 & ~n17371;
  assign n17386 = n15720 & ~n17382;
  assign n17387 = ~n17385 & ~n17386;
  assign n17388 = n15712 & ~n17371;
  assign n17389 = n15706 & ~n17371;
  assign n17390 = n17270 & ~n17316;
  assign n17391 = ~n17376 & ~n17390;
  assign n17392 = ~n17313 & n17391;
  assign n17393 = ~n17364 & n17392;
  assign n17394 = n17364 & ~n17392;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = n15709 & ~n17395;
  assign n17397 = n15715 & ~n17395;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~n17388 & ~n17389;
  assign n17400 = n17398 & n17399;
  assign n17401 = ~n17383 & ~n17384;
  assign n17402 = n17387 & n17401;
  assign n17403 = n17400 & n17402;
  assign n17404 = n17374 & n17403;
  assign n17405 = n15649 & ~n17404;
  assign n17406 = P3_REG0_REG_27_ & ~n15649;
  assign n3015 = n17405 | n17406;
  assign n17408 = P3_REG0_REG_29_ & n15681;
  assign n17409 = P3_REG1_REG_29_ & n15679;
  assign n17410 = P3_REG2_REG_29_ & n15677;
  assign n17411 = n15675 & n17349;
  assign n17412 = ~n17408 & ~n17409;
  assign n17413 = ~n17410 & n17412;
  assign n17414 = ~n17411 & n17413;
  assign n17415 = n15694 & ~n17414;
  assign n17416 = ~n15422 & ~n15656;
  assign n17417 = ~n15667 & n17416;
  assign n17418 = ~n17358 & ~n17416;
  assign n17419 = n17358 & n17416;
  assign n17420 = ~n17418 & ~n17419;
  assign n17421 = n17297 & ~n17301;
  assign n17422 = ~n17360 & ~n17421;
  assign n17423 = ~n17297 & n17301;
  assign n17424 = ~n17422 & ~n17423;
  assign n17425 = ~n17302 & ~n17363;
  assign n17426 = ~n17305 & n17425;
  assign n17427 = n17424 & ~n17426;
  assign n17428 = ~n17420 & ~n17427;
  assign n17429 = n17420 & n17427;
  assign n17430 = ~n17428 & ~n17429;
  assign n17431 = n15689 & ~n17430;
  assign n17432 = ~n17415 & ~n17417;
  assign n17433 = ~n17431 & n17432;
  assign n17434 = n17297 & ~n17360;
  assign n17435 = n17313 & ~n17434;
  assign n17436 = ~n17202 & ~n17434;
  assign n17437 = ~n17200 & ~n17316;
  assign n17438 = n17436 & n17437;
  assign n17439 = n17376 & ~n17434;
  assign n17440 = ~n17297 & n17360;
  assign n17441 = ~n17439 & ~n17440;
  assign n17442 = ~n17435 & ~n17438;
  assign n17443 = n17441 & n17442;
  assign n17444 = ~n17420 & n17443;
  assign n17445 = n17420 & ~n17443;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = n15722 & ~n17446;
  assign n17448 = n15768 & ~n17297;
  assign n17449 = n15717 & ~n17430;
  assign n17450 = n15720 & ~n17446;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = n15712 & ~n17430;
  assign n17453 = n15706 & ~n17430;
  assign n17454 = ~n17215 & ~n17316;
  assign n17455 = n17436 & n17454;
  assign n17456 = ~n17435 & ~n17455;
  assign n17457 = n17441 & n17456;
  assign n17458 = ~n17420 & n17457;
  assign n17459 = n17420 & ~n17457;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = n15709 & ~n17460;
  assign n17462 = n15715 & ~n17460;
  assign n17463 = ~n17461 & ~n17462;
  assign n17464 = ~n17452 & ~n17453;
  assign n17465 = n17463 & n17464;
  assign n17466 = ~n17447 & ~n17448;
  assign n17467 = n17451 & n17466;
  assign n17468 = n17465 & n17467;
  assign n17469 = n17433 & n17468;
  assign n17470 = n15649 & ~n17469;
  assign n17471 = P3_REG0_REG_28_ & ~n15649;
  assign n3020 = n17470 | n17471;
  assign n17473 = ~n15441 & ~n15656;
  assign n17474 = ~n15667 & n17473;
  assign n17475 = ~n17414 & ~n17473;
  assign n17476 = n17414 & n17473;
  assign n17477 = ~n17475 & ~n17476;
  assign n17478 = n17358 & n17477;
  assign n17479 = n17416 & n17478;
  assign n17480 = ~n17358 & ~n17477;
  assign n17481 = ~n17416 & n17480;
  assign n17482 = ~n17479 & ~n17481;
  assign n17483 = ~n17419 & ~n17477;
  assign n17484 = ~n17427 & n17483;
  assign n17485 = ~n17418 & n17477;
  assign n17486 = n17427 & n17485;
  assign n17487 = n17482 & ~n17484;
  assign n17488 = ~n17486 & n17487;
  assign n17489 = n15689 & ~n17488;
  assign n17490 = ~n17474 & ~n17489;
  assign n17491 = n15768 & ~n17358;
  assign n17492 = ~P3_B_REG & n15692;
  assign n17493 = ~n15656 & ~n17492;
  assign n17494 = P3_REG0_REG_30_ & n15681;
  assign n17495 = P3_REG1_REG_30_ & n15679;
  assign n17496 = P3_REG2_REG_30_ & n15677;
  assign n17497 = ~n17411 & ~n17494;
  assign n17498 = ~n17495 & n17497;
  assign n17499 = ~n17496 & n17498;
  assign n17500 = n15691 & ~n17493;
  assign n17501 = ~n17499 & n17500;
  assign n17502 = n17416 & ~n17443;
  assign n17503 = ~n17358 & ~n17443;
  assign n17504 = ~n17358 & n17416;
  assign n17505 = ~n17502 & ~n17503;
  assign n17506 = ~n17504 & n17505;
  assign n17507 = ~n17477 & n17506;
  assign n17508 = n17477 & ~n17506;
  assign n17509 = ~n17507 & ~n17508;
  assign n17510 = n15722 & ~n17509;
  assign n17511 = n15717 & ~n17488;
  assign n17512 = n15720 & ~n17509;
  assign n17513 = ~n17511 & ~n17512;
  assign n17514 = n15712 & ~n17488;
  assign n17515 = n15706 & ~n17488;
  assign n17516 = n17416 & ~n17457;
  assign n17517 = ~n17358 & ~n17457;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~n17504 & n17518;
  assign n17520 = ~n17477 & n17519;
  assign n17521 = n17477 & ~n17519;
  assign n17522 = ~n17520 & ~n17521;
  assign n17523 = n15709 & ~n17522;
  assign n17524 = n15715 & ~n17522;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = ~n17514 & ~n17515;
  assign n17527 = n17525 & n17526;
  assign n17528 = ~n17491 & ~n17501;
  assign n17529 = ~n17510 & n17528;
  assign n17530 = n17513 & n17529;
  assign n17531 = n17527 & n17530;
  assign n17532 = n17490 & n17531;
  assign n17533 = n15649 & ~n17532;
  assign n17534 = P3_REG0_REG_29_ & ~n15649;
  assign n3025 = n17533 | n17534;
  assign n17536 = P3_REG0_REG_31_ & n15681;
  assign n17537 = P3_REG1_REG_31_ & n15679;
  assign n17538 = P3_REG2_REG_31_ & n15677;
  assign n17539 = ~n17536 & ~n17537;
  assign n17540 = ~n17538 & n17539;
  assign n17541 = ~n17411 & n17540;
  assign n17542 = n17500 & ~n17541;
  assign n17543 = ~n15460 & ~n15656;
  assign n17544 = ~n15667 & n17543;
  assign n17545 = ~n17542 & ~n17544;
  assign n17546 = n15649 & ~n17545;
  assign n17547 = P3_REG0_REG_30_ & ~n15649;
  assign n3030 = n17546 | n17547;
  assign n17549 = ~n15486 & ~n15656;
  assign n17550 = ~n15667 & n17549;
  assign n17551 = ~n17542 & ~n17550;
  assign n17552 = n15649 & ~n17551;
  assign n17553 = P3_REG0_REG_31_ & ~n15649;
  assign n3035 = n17552 | n17553;
  assign n17555 = n15553 & ~n15557;
  assign n17556 = n15617 & n17555;
  assign n17557 = n15628 & n15634;
  assign n17558 = n15621 & ~n15628;
  assign n17559 = ~n17557 & ~n17558;
  assign n17560 = ~n15641 & n17559;
  assign n17561 = n17556 & ~n17560;
  assign n17562 = ~n15553 & n15557;
  assign n17563 = n15617 & n17562;
  assign n17564 = ~n15627 & n15705;
  assign n17565 = ~n15645 & ~n17564;
  assign n17566 = n17563 & ~n17565;
  assign n17567 = ~n17561 & ~n17566;
  assign n17568 = n15505 & ~n17567;
  assign n17569 = ~n15729 & n17568;
  assign n17570 = P3_REG1_REG_0_ & ~n17568;
  assign n3040 = n17569 | n17570;
  assign n17572 = ~n15783 & n17568;
  assign n17573 = P3_REG1_REG_1_ & ~n17568;
  assign n3045 = n17572 | n17573;
  assign n17575 = ~n15839 & n17568;
  assign n17576 = P3_REG1_REG_2_ & ~n17568;
  assign n3050 = n17575 | n17576;
  assign n17578 = ~n15899 & n17568;
  assign n17579 = P3_REG1_REG_3_ & ~n17568;
  assign n3055 = n17578 | n17579;
  assign n17581 = ~n15963 & n17568;
  assign n17582 = P3_REG1_REG_4_ & ~n17568;
  assign n3060 = n17581 | n17582;
  assign n17584 = ~n16023 & n17568;
  assign n17585 = P3_REG1_REG_5_ & ~n17568;
  assign n3065 = n17584 | n17585;
  assign n17587 = ~n16091 & n17568;
  assign n17588 = P3_REG1_REG_6_ & ~n17568;
  assign n3070 = n17587 | n17588;
  assign n17590 = ~n16154 & n17568;
  assign n17591 = P3_REG1_REG_7_ & ~n17568;
  assign n3075 = n17590 | n17591;
  assign n17593 = ~n16217 & n17568;
  assign n17594 = P3_REG1_REG_8_ & ~n17568;
  assign n3080 = n17593 | n17594;
  assign n17596 = ~n16281 & n17568;
  assign n17597 = P3_REG1_REG_9_ & ~n17568;
  assign n3085 = n17596 | n17597;
  assign n17599 = ~n16340 & n17568;
  assign n17600 = P3_REG1_REG_10_ & ~n17568;
  assign n3090 = n17599 | n17600;
  assign n17602 = ~n16411 & n17568;
  assign n17603 = P3_REG1_REG_11_ & ~n17568;
  assign n3095 = n17602 | n17603;
  assign n17605 = ~n16478 & n17568;
  assign n17606 = P3_REG1_REG_12_ & ~n17568;
  assign n3100 = n17605 | n17606;
  assign n17608 = ~n16541 & n17568;
  assign n17609 = P3_REG1_REG_13_ & ~n17568;
  assign n3105 = n17608 | n17609;
  assign n17611 = ~n16605 & n17568;
  assign n17612 = P3_REG1_REG_14_ & ~n17568;
  assign n3110 = n17611 | n17612;
  assign n17614 = ~n16665 & n17568;
  assign n17615 = P3_REG1_REG_15_ & ~n17568;
  assign n3115 = n17614 | n17615;
  assign n17617 = ~n16732 & n17568;
  assign n17618 = P3_REG1_REG_16_ & ~n17568;
  assign n3120 = n17617 | n17618;
  assign n17620 = ~n16800 & n17568;
  assign n17621 = P3_REG1_REG_17_ & ~n17568;
  assign n3125 = n17620 | n17621;
  assign n17623 = ~n16866 & n17568;
  assign n17624 = P3_REG1_REG_18_ & ~n17568;
  assign n3130 = n17623 | n17624;
  assign n17626 = ~n16926 & n17568;
  assign n17627 = P3_REG1_REG_19_ & ~n17568;
  assign n3135 = n17626 | n17627;
  assign n17629 = ~n16985 & n17568;
  assign n17630 = P3_REG1_REG_20_ & ~n17568;
  assign n3140 = n17629 | n17630;
  assign n17632 = ~n17043 & n17568;
  assign n17633 = P3_REG1_REG_21_ & ~n17568;
  assign n3145 = n17632 | n17633;
  assign n17635 = ~n17105 & n17568;
  assign n17636 = P3_REG1_REG_22_ & ~n17568;
  assign n3150 = n17635 | n17636;
  assign n17638 = ~n17163 & n17568;
  assign n17639 = P3_REG1_REG_23_ & ~n17568;
  assign n3155 = n17638 | n17639;
  assign n17641 = ~n17227 & n17568;
  assign n17642 = P3_REG1_REG_24_ & ~n17568;
  assign n3160 = n17641 | n17642;
  assign n17644 = ~n17283 & n17568;
  assign n17645 = P3_REG1_REG_25_ & ~n17568;
  assign n3165 = n17644 | n17645;
  assign n17647 = ~n17345 & n17568;
  assign n17648 = P3_REG1_REG_26_ & ~n17568;
  assign n3170 = n17647 | n17648;
  assign n17650 = ~n17404 & n17568;
  assign n17651 = P3_REG1_REG_27_ & ~n17568;
  assign n3175 = n17650 | n17651;
  assign n17653 = ~n17469 & n17568;
  assign n17654 = P3_REG1_REG_28_ & ~n17568;
  assign n3180 = n17653 | n17654;
  assign n17656 = ~n17532 & n17568;
  assign n17657 = P3_REG1_REG_29_ & ~n17568;
  assign n3185 = n17656 | n17657;
  assign n17659 = ~n17545 & n17568;
  assign n17660 = P3_REG1_REG_30_ & ~n17568;
  assign n3190 = n17659 | n17660;
  assign n17662 = ~n17551 & n17568;
  assign n17663 = P3_REG1_REG_31_ & ~n17568;
  assign n3195 = n17662 | n17663;
  assign n17665 = ~n15624 & n15627;
  assign n17666 = ~n15634 & n17665;
  assign n17667 = n15624 & ~n15634;
  assign n17668 = ~n15621 & ~n17667;
  assign n17669 = ~n15628 & n17668;
  assign n17670 = n17563 & ~n17669;
  assign n17671 = n15627 & n15666;
  assign n17672 = n17556 & ~n17565;
  assign n17673 = ~n17670 & ~n17671;
  assign n17674 = ~n17672 & n17673;
  assign n17675 = n15505 & ~n17674;
  assign n17676 = n17666 & n17675;
  assign n17677 = ~n15688 & n17676;
  assign n17678 = n15694 & n17675;
  assign n17679 = ~n15701 & n17678;
  assign n17680 = ~n15627 & n15666;
  assign n17681 = ~n15664 & ~n17680;
  assign n17682 = n17675 & ~n17681;
  assign n17683 = ~n15662 & n17682;
  assign n17684 = ~n15728 & n17675;
  assign n17685 = P3_REG2_REG_0_ & ~n17675;
  assign n17686 = ~n17684 & ~n17685;
  assign n17687 = n17671 & n17675;
  assign n17688 = P3_REG3_REG_0_ & n17687;
  assign n17689 = ~n17677 & ~n17679;
  assign n17690 = ~n17683 & n17689;
  assign n17691 = n17686 & n17690;
  assign n3200 = n17688 | ~n17691;
  assign n17693 = ~n15753 & n17676;
  assign n17694 = ~n15739 & n17678;
  assign n17695 = ~n15746 & n17682;
  assign n17696 = ~n15782 & n17675;
  assign n17697 = P3_REG2_REG_1_ & ~n17675;
  assign n17698 = ~n17696 & ~n17697;
  assign n17699 = P3_REG3_REG_1_ & n17687;
  assign n17700 = ~n17693 & ~n17694;
  assign n17701 = ~n17695 & n17700;
  assign n17702 = n17698 & n17701;
  assign n3205 = n17699 | ~n17702;
  assign n17704 = ~n15811 & n17676;
  assign n17705 = ~n15793 & n17678;
  assign n17706 = ~n15800 & n17682;
  assign n17707 = ~n15838 & n17675;
  assign n17708 = P3_REG2_REG_2_ & ~n17675;
  assign n17709 = ~n17707 & ~n17708;
  assign n17710 = P3_REG3_REG_2_ & n17687;
  assign n17711 = ~n17704 & ~n17705;
  assign n17712 = ~n17706 & n17711;
  assign n17713 = n17709 & n17712;
  assign n3210 = n17710 | ~n17713;
  assign n17715 = ~n15870 & n17676;
  assign n17716 = ~n15852 & n17678;
  assign n17717 = ~n15859 & n17682;
  assign n17718 = ~n15898 & n17675;
  assign n17719 = P3_REG2_REG_3_ & ~n17675;
  assign n17720 = ~n17718 & ~n17719;
  assign n17721 = ~P3_REG3_REG_3_ & n17687;
  assign n17722 = ~n17715 & ~n17716;
  assign n17723 = ~n17717 & n17722;
  assign n17724 = n17720 & n17723;
  assign n3215 = n17721 | ~n17724;
  assign n17726 = ~n15933 & n17676;
  assign n17727 = ~n15912 & n17678;
  assign n17728 = ~n15919 & n17682;
  assign n17729 = ~n15962 & n17675;
  assign n17730 = P3_REG2_REG_4_ & ~n17675;
  assign n17731 = ~n17729 & ~n17730;
  assign n17732 = ~n15845 & n17687;
  assign n17733 = ~n17726 & ~n17727;
  assign n17734 = ~n17728 & n17733;
  assign n17735 = n17731 & n17734;
  assign n3220 = n17732 | ~n17735;
  assign n17737 = ~n15994 & n17676;
  assign n17738 = ~n15978 & n17678;
  assign n17739 = ~n15985 & n17682;
  assign n17740 = ~n16022 & n17675;
  assign n17741 = P3_REG2_REG_5_ & ~n17675;
  assign n17742 = ~n17740 & ~n17741;
  assign n17743 = ~n15905 & n17687;
  assign n17744 = ~n17737 & ~n17738;
  assign n17745 = ~n17739 & n17744;
  assign n17746 = n17742 & n17745;
  assign n3225 = n17743 | ~n17746;
  assign n17748 = ~n16056 & n17676;
  assign n17749 = ~n16037 & n17678;
  assign n17750 = ~n16044 & n17682;
  assign n17751 = ~n16090 & n17675;
  assign n17752 = P3_REG2_REG_6_ & ~n17675;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = ~n15971 & n17687;
  assign n17755 = ~n17748 & ~n17749;
  assign n17756 = ~n17750 & n17755;
  assign n17757 = n17753 & n17756;
  assign n3230 = n17754 | ~n17757;
  assign n17759 = ~n16125 & n17676;
  assign n17760 = ~n16104 & n17678;
  assign n17761 = ~n16111 & n17682;
  assign n17762 = ~n16153 & n17675;
  assign n17763 = P3_REG2_REG_7_ & ~n17675;
  assign n17764 = ~n17762 & ~n17763;
  assign n17765 = ~n16030 & n17687;
  assign n17766 = ~n17759 & ~n17760;
  assign n17767 = ~n17761 & n17766;
  assign n17768 = n17764 & n17767;
  assign n3235 = n17765 | ~n17768;
  assign n17770 = ~n16186 & n17676;
  assign n17771 = ~n16168 & n17678;
  assign n17772 = ~n16175 & n17682;
  assign n17773 = ~n16216 & n17675;
  assign n17774 = P3_REG2_REG_8_ & ~n17675;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = ~n16097 & n17687;
  assign n17777 = ~n17770 & ~n17771;
  assign n17778 = ~n17772 & n17777;
  assign n17779 = n17775 & n17778;
  assign n3240 = n17776 | ~n17779;
  assign n17781 = ~n16254 & n17676;
  assign n17782 = ~n16230 & n17678;
  assign n17783 = ~n16237 & n17682;
  assign n17784 = ~n16280 & n17675;
  assign n17785 = P3_REG2_REG_9_ & ~n17675;
  assign n17786 = ~n17784 & ~n17785;
  assign n17787 = ~n16161 & n17687;
  assign n17788 = ~n17781 & ~n17782;
  assign n17789 = ~n17783 & n17788;
  assign n17790 = n17786 & n17789;
  assign n3245 = n17787 | ~n17790;
  assign n17792 = ~n16223 & n17687;
  assign n17793 = ~n16302 & n17682;
  assign n17794 = ~n16311 & n17676;
  assign n17795 = ~n16295 & n17678;
  assign n17796 = ~n16339 & n17675;
  assign n17797 = P3_REG2_REG_10_ & ~n17675;
  assign n17798 = ~n17796 & ~n17797;
  assign n17799 = ~n17792 & ~n17793;
  assign n17800 = ~n17794 & n17799;
  assign n17801 = ~n17795 & n17800;
  assign n3250 = ~n17798 | ~n17801;
  assign n17803 = ~n16288 & n17687;
  assign n17804 = ~n16372 & n17676;
  assign n17805 = ~n16360 & n17682;
  assign n17806 = ~n16353 & n17678;
  assign n17807 = ~n16410 & n17675;
  assign n17808 = P3_REG2_REG_11_ & ~n17675;
  assign n17809 = ~n17807 & ~n17808;
  assign n17810 = ~n17803 & ~n17804;
  assign n17811 = ~n17805 & n17810;
  assign n17812 = ~n17806 & n17811;
  assign n3255 = ~n17809 | ~n17812;
  assign n17814 = ~n16346 & n17687;
  assign n17815 = ~n16432 & n17682;
  assign n17816 = ~n16446 & n17676;
  assign n17817 = ~n16425 & n17678;
  assign n17818 = ~n16477 & n17675;
  assign n17819 = P3_REG2_REG_12_ & ~n17675;
  assign n17820 = ~n17818 & ~n17819;
  assign n17821 = ~n17814 & ~n17815;
  assign n17822 = ~n17816 & n17821;
  assign n17823 = ~n17817 & n17822;
  assign n3260 = ~n17820 | ~n17823;
  assign n17825 = ~n16418 & n17687;
  assign n17826 = ~n16507 & n17676;
  assign n17827 = ~n16498 & n17682;
  assign n17828 = ~n16491 & n17678;
  assign n17829 = ~n16540 & n17675;
  assign n17830 = P3_REG2_REG_13_ & ~n17675;
  assign n17831 = ~n17829 & ~n17830;
  assign n17832 = ~n17825 & ~n17826;
  assign n17833 = ~n17827 & n17832;
  assign n17834 = ~n17828 & n17833;
  assign n3265 = ~n17831 | ~n17834;
  assign n17836 = ~n16562 & n17682;
  assign n17837 = ~n16555 & n17678;
  assign n17838 = ~n16484 & n17687;
  assign n17839 = ~n16571 & n17676;
  assign n17840 = ~n16604 & n17675;
  assign n17841 = P3_REG2_REG_14_ & ~n17675;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = ~n17836 & ~n17837;
  assign n17844 = ~n17838 & n17843;
  assign n17845 = ~n17839 & n17844;
  assign n3270 = ~n17842 | ~n17845;
  assign n17847 = ~n16625 & n17682;
  assign n17848 = ~n16618 & n17678;
  assign n17849 = ~n16548 & n17687;
  assign n17850 = ~n16634 & n17676;
  assign n17851 = ~n16664 & n17675;
  assign n17852 = P3_REG2_REG_15_ & ~n17675;
  assign n17853 = ~n17851 & ~n17852;
  assign n17854 = ~n17847 & ~n17848;
  assign n17855 = ~n17849 & n17854;
  assign n17856 = ~n17850 & n17855;
  assign n3275 = ~n17853 | ~n17856;
  assign n17858 = ~n16686 & n17682;
  assign n17859 = ~n16679 & n17678;
  assign n17860 = ~n16611 & n17687;
  assign n17861 = ~n16698 & n17676;
  assign n17862 = ~n16731 & n17675;
  assign n17863 = P3_REG2_REG_16_ & ~n17675;
  assign n17864 = ~n17862 & ~n17863;
  assign n17865 = ~n17858 & ~n17859;
  assign n17866 = ~n17860 & n17865;
  assign n17867 = ~n17861 & n17866;
  assign n3280 = ~n17864 | ~n17867;
  assign n17869 = ~n16752 & n17682;
  assign n17870 = ~n16745 & n17678;
  assign n17871 = ~n16672 & n17687;
  assign n17872 = ~n16766 & n17676;
  assign n17873 = ~n16799 & n17675;
  assign n17874 = P3_REG2_REG_17_ & ~n17675;
  assign n17875 = ~n17873 & ~n17874;
  assign n17876 = ~n17869 & ~n17870;
  assign n17877 = ~n17871 & n17876;
  assign n17878 = ~n17872 & n17877;
  assign n3285 = ~n17875 | ~n17878;
  assign n17880 = ~n16821 & n17682;
  assign n17881 = ~n16814 & n17678;
  assign n17882 = ~n16738 & n17687;
  assign n17883 = ~n16830 & n17676;
  assign n17884 = ~n16865 & n17675;
  assign n17885 = P3_REG2_REG_18_ & ~n17675;
  assign n17886 = ~n17884 & ~n17885;
  assign n17887 = ~n17880 & ~n17881;
  assign n17888 = ~n17882 & n17887;
  assign n17889 = ~n17883 & n17888;
  assign n3290 = ~n17886 | ~n17889;
  assign n17891 = ~n16883 & n17682;
  assign n17892 = ~n16879 & n17678;
  assign n17893 = ~n16807 & n17687;
  assign n17894 = ~n16894 & n17676;
  assign n17895 = ~n16925 & n17675;
  assign n17896 = P3_REG2_REG_19_ & ~n17675;
  assign n17897 = ~n17895 & ~n17896;
  assign n17898 = ~n17891 & ~n17892;
  assign n17899 = ~n17893 & n17898;
  assign n17900 = ~n17894 & n17899;
  assign n3295 = ~n17897 | ~n17900;
  assign n17902 = n16942 & n17682;
  assign n17903 = ~n16940 & n17678;
  assign n17904 = ~n16872 & n17687;
  assign n17905 = ~n16951 & n17676;
  assign n17906 = ~n16984 & n17675;
  assign n17907 = P3_REG2_REG_20_ & ~n17675;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n17902 & ~n17903;
  assign n17910 = ~n17904 & n17909;
  assign n17911 = ~n17905 & n17910;
  assign n3300 = ~n17908 | ~n17911;
  assign n17913 = n17000 & n17682;
  assign n17914 = ~n16998 & n17678;
  assign n17915 = ~n16933 & n17687;
  assign n17916 = ~n17009 & n17676;
  assign n17917 = ~n17042 & n17675;
  assign n17918 = P3_REG2_REG_21_ & ~n17675;
  assign n17919 = ~n17917 & ~n17918;
  assign n17920 = ~n17913 & ~n17914;
  assign n17921 = ~n17915 & n17920;
  assign n17922 = ~n17916 & n17921;
  assign n3305 = ~n17919 | ~n17922;
  assign n17924 = n17059 & n17682;
  assign n17925 = ~n17057 & n17678;
  assign n17926 = ~n16991 & n17687;
  assign n17927 = ~n17068 & n17676;
  assign n17928 = ~n17104 & n17675;
  assign n17929 = P3_REG2_REG_22_ & ~n17675;
  assign n17930 = ~n17928 & ~n17929;
  assign n17931 = ~n17924 & ~n17925;
  assign n17932 = ~n17926 & n17931;
  assign n17933 = ~n17927 & n17932;
  assign n3310 = ~n17930 | ~n17933;
  assign n17935 = n17120 & n17682;
  assign n17936 = ~n17118 & n17678;
  assign n17937 = ~n17050 & n17687;
  assign n17938 = ~n17132 & n17676;
  assign n17939 = ~n17162 & n17675;
  assign n17940 = P3_REG2_REG_23_ & ~n17675;
  assign n17941 = ~n17939 & ~n17940;
  assign n17942 = ~n17935 & ~n17936;
  assign n17943 = ~n17937 & n17942;
  assign n17944 = ~n17938 & n17943;
  assign n3315 = ~n17941 | ~n17944;
  assign n17946 = n17179 & n17682;
  assign n17947 = ~n17177 & n17678;
  assign n17948 = ~n17111 & n17687;
  assign n17949 = ~n17193 & n17676;
  assign n17950 = ~n17226 & n17675;
  assign n17951 = P3_REG2_REG_24_ & ~n17675;
  assign n17952 = ~n17950 & ~n17951;
  assign n17953 = ~n17946 & ~n17947;
  assign n17954 = ~n17948 & n17953;
  assign n17955 = ~n17949 & n17954;
  assign n3320 = ~n17952 | ~n17955;
  assign n17957 = n17242 & n17682;
  assign n17958 = ~n17240 & n17678;
  assign n17959 = ~n17170 & n17687;
  assign n17960 = ~n17251 & n17676;
  assign n17961 = ~n17282 & n17675;
  assign n17962 = P3_REG2_REG_25_ & ~n17675;
  assign n17963 = ~n17961 & ~n17962;
  assign n17964 = ~n17957 & ~n17958;
  assign n17965 = ~n17959 & n17964;
  assign n17966 = ~n17960 & n17965;
  assign n3325 = ~n17963 | ~n17966;
  assign n17968 = n17299 & n17682;
  assign n17969 = ~n17297 & n17678;
  assign n17970 = ~n17233 & n17687;
  assign n17971 = ~n17308 & n17676;
  assign n17972 = ~n17344 & n17675;
  assign n17973 = P3_REG2_REG_26_ & ~n17675;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~n17968 & ~n17969;
  assign n17976 = ~n17970 & n17975;
  assign n17977 = ~n17971 & n17976;
  assign n3330 = ~n17974 | ~n17977;
  assign n17979 = n17360 & n17682;
  assign n17980 = ~n17358 & n17678;
  assign n17981 = ~n17293 & n17687;
  assign n17982 = ~n17371 & n17676;
  assign n17983 = ~n17403 & n17675;
  assign n17984 = P3_REG2_REG_27_ & ~n17675;
  assign n17985 = ~n17983 & ~n17984;
  assign n17986 = ~n17979 & ~n17980;
  assign n17987 = ~n17981 & n17986;
  assign n17988 = ~n17982 & n17987;
  assign n3335 = ~n17985 | ~n17988;
  assign n17990 = n17416 & n17682;
  assign n17991 = ~n17414 & n17678;
  assign n17992 = ~n17351 & n17687;
  assign n17993 = ~n17430 & n17676;
  assign n17994 = ~n17468 & n17675;
  assign n17995 = P3_REG2_REG_28_ & ~n17675;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = ~n17990 & ~n17991;
  assign n17998 = ~n17992 & n17997;
  assign n17999 = ~n17993 & n17998;
  assign n3340 = ~n17996 | ~n17999;
  assign n18001 = n17473 & n17682;
  assign n18002 = n17349 & n17687;
  assign n18003 = ~n17488 & n17676;
  assign n18004 = ~n17531 & n17675;
  assign n18005 = P3_REG2_REG_29_ & ~n17675;
  assign n18006 = ~n18004 & ~n18005;
  assign n18007 = ~n18001 & ~n18002;
  assign n18008 = ~n18003 & n18007;
  assign n3345 = ~n18006 | ~n18008;
  assign n18010 = P3_REG2_REG_30_ & ~n17675;
  assign n18011 = n17542 & n17675;
  assign n18012 = ~n18002 & ~n18011;
  assign n18013 = n17543 & n17682;
  assign n18014 = ~n18010 & n18012;
  assign n3350 = n18013 | ~n18014;
  assign n18016 = P3_REG2_REG_31_ & ~n17675;
  assign n18017 = n17549 & n17682;
  assign n18018 = n18012 & ~n18016;
  assign n3355 = n18017 | ~n18018;
  assign n18020 = ~n15492 & ~n15656;
  assign n18021 = ~n15656 & ~n15691;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = n15492 & n15503;
  assign n18024 = P3_STATE_REG & ~n18023;
  assign n18025 = n18022 & n18024;
  assign n18026 = n15505 & ~n18025;
  assign n18027 = ~n15709 & ~n17671;
  assign n18028 = ~n15644 & ~n15715;
  assign n18029 = ~n15722 & n18028;
  assign n18030 = ~n15720 & n18029;
  assign n18031 = ~n15717 & n18030;
  assign n18032 = ~n17665 & n17681;
  assign n18033 = n18027 & n18032;
  assign n18034 = n18031 & n18033;
  assign n18035 = n15655 & ~n18034;
  assign n18036 = ~n15634 & n18035;
  assign n18037 = P3_REG2_REG_18_ & n16818;
  assign n18038 = ~P3_REG2_REG_19_ & ~n15634;
  assign n18039 = P3_REG2_REG_19_ & n15634;
  assign n18040 = ~n18038 & ~n18039;
  assign n18041 = ~n18037 & ~n18040;
  assign n18042 = ~P3_REG2_REG_17_ & ~n16749;
  assign n18043 = P3_REG2_REG_17_ & n16749;
  assign n18044 = ~P3_REG2_REG_16_ & ~n16683;
  assign n18045 = P3_REG2_REG_16_ & n16683;
  assign n18046 = ~P3_REG2_REG_14_ & ~n16559;
  assign n18047 = P3_REG2_REG_14_ & n16559;
  assign n18048 = ~P3_REG2_REG_13_ & ~n16495;
  assign n18049 = P3_REG2_REG_13_ & n16495;
  assign n18050 = ~P3_REG2_REG_12_ & ~n16429;
  assign n18051 = P3_REG2_REG_12_ & n16429;
  assign n18052 = ~P3_REG2_REG_11_ & ~n16357;
  assign n18053 = P3_REG2_REG_11_ & n16357;
  assign n18054 = ~P3_REG2_REG_10_ & ~n16299;
  assign n18055 = P3_REG2_REG_10_ & n16299;
  assign n18056 = ~P3_REG2_REG_9_ & ~n16234;
  assign n18057 = P3_REG2_REG_9_ & n16234;
  assign n18058 = ~P3_REG2_REG_8_ & ~n16172;
  assign n18059 = P3_REG2_REG_8_ & n16172;
  assign n18060 = ~P3_REG2_REG_7_ & ~n16108;
  assign n18061 = P3_REG2_REG_7_ & n16108;
  assign n18062 = ~P3_REG2_REG_6_ & ~n16041;
  assign n18063 = P3_REG2_REG_6_ & n16041;
  assign n18064 = ~P3_REG2_REG_5_ & ~n15982;
  assign n18065 = P3_REG2_REG_5_ & n15982;
  assign n18066 = ~P3_REG2_REG_4_ & ~n15916;
  assign n18067 = P3_REG2_REG_4_ & n15916;
  assign n18068 = ~P3_REG2_REG_3_ & ~n15856;
  assign n18069 = P3_REG2_REG_3_ & n15856;
  assign n18070 = ~P3_REG2_REG_2_ & ~n15797;
  assign n18071 = P3_REG2_REG_2_ & n15797;
  assign n18072 = P3_REG2_REG_0_ & n15659;
  assign n18073 = ~P3_REG2_REG_1_ & ~n18072;
  assign n18074 = P3_REG2_REG_1_ & n18072;
  assign n18075 = ~n15743 & ~n18074;
  assign n18076 = ~n18073 & ~n18075;
  assign n18077 = ~n18071 & ~n18076;
  assign n18078 = ~n18070 & ~n18077;
  assign n18079 = ~n18069 & ~n18078;
  assign n18080 = ~n18068 & ~n18079;
  assign n18081 = ~n18067 & ~n18080;
  assign n18082 = ~n18066 & ~n18081;
  assign n18083 = ~n18065 & ~n18082;
  assign n18084 = ~n18064 & ~n18083;
  assign n18085 = ~n18063 & ~n18084;
  assign n18086 = ~n18062 & ~n18085;
  assign n18087 = ~n18061 & ~n18086;
  assign n18088 = ~n18060 & ~n18087;
  assign n18089 = ~n18059 & ~n18088;
  assign n18090 = ~n18058 & ~n18089;
  assign n18091 = ~n18057 & ~n18090;
  assign n18092 = ~n18056 & ~n18091;
  assign n18093 = ~n18055 & ~n18092;
  assign n18094 = ~n18054 & ~n18093;
  assign n18095 = ~n18053 & ~n18094;
  assign n18096 = ~n18052 & ~n18095;
  assign n18097 = ~n18051 & ~n18096;
  assign n18098 = ~n18050 & ~n18097;
  assign n18099 = ~n18049 & ~n18098;
  assign n18100 = ~n18048 & ~n18099;
  assign n18101 = ~n18047 & ~n18100;
  assign n18102 = ~n18046 & ~n18101;
  assign n18103 = ~P3_REG2_REG_15_ & ~n18102;
  assign n18104 = P3_REG2_REG_15_ & n18102;
  assign n18105 = ~n16622 & ~n18104;
  assign n18106 = ~n18103 & ~n18105;
  assign n18107 = ~n18045 & ~n18106;
  assign n18108 = ~n18044 & ~n18107;
  assign n18109 = ~n18043 & ~n18108;
  assign n18110 = ~n18042 & ~n18109;
  assign n18111 = ~P3_REG2_REG_18_ & ~n16818;
  assign n18112 = n18110 & ~n18111;
  assign n18113 = n18041 & ~n18112;
  assign n18114 = n18040 & ~n18111;
  assign n18115 = ~n18037 & ~n18110;
  assign n18116 = n18114 & ~n18115;
  assign n18117 = ~n18113 & ~n18116;
  assign n18118 = n15692 & ~n18034;
  assign n18119 = ~n18117 & n18118;
  assign n18120 = P3_REG1_REG_18_ & n16818;
  assign n18121 = ~P3_REG1_REG_19_ & ~n15634;
  assign n18122 = P3_REG1_REG_19_ & n15634;
  assign n18123 = ~n18121 & ~n18122;
  assign n18124 = ~n18120 & ~n18123;
  assign n18125 = ~P3_REG1_REG_17_ & ~n16749;
  assign n18126 = P3_REG1_REG_17_ & n16749;
  assign n18127 = ~P3_REG1_REG_16_ & ~n16683;
  assign n18128 = P3_REG1_REG_16_ & n16683;
  assign n18129 = ~P3_REG1_REG_14_ & ~n16559;
  assign n18130 = P3_REG1_REG_14_ & n16559;
  assign n18131 = ~P3_REG1_REG_13_ & ~n16495;
  assign n18132 = P3_REG1_REG_13_ & n16495;
  assign n18133 = ~P3_REG1_REG_12_ & ~n16429;
  assign n18134 = P3_REG1_REG_12_ & n16429;
  assign n18135 = ~P3_REG1_REG_11_ & ~n16357;
  assign n18136 = P3_REG1_REG_11_ & n16357;
  assign n18137 = ~P3_REG1_REG_10_ & ~n16299;
  assign n18138 = P3_REG1_REG_10_ & n16299;
  assign n18139 = ~P3_REG1_REG_9_ & ~n16234;
  assign n18140 = P3_REG1_REG_9_ & n16234;
  assign n18141 = ~P3_REG1_REG_8_ & ~n16172;
  assign n18142 = P3_REG1_REG_8_ & n16172;
  assign n18143 = ~P3_REG1_REG_7_ & ~n16108;
  assign n18144 = P3_REG1_REG_7_ & n16108;
  assign n18145 = ~P3_REG1_REG_6_ & ~n16041;
  assign n18146 = P3_REG1_REG_6_ & n16041;
  assign n18147 = ~P3_REG1_REG_5_ & ~n15982;
  assign n18148 = P3_REG1_REG_5_ & n15982;
  assign n18149 = ~P3_REG1_REG_4_ & ~n15916;
  assign n18150 = P3_REG1_REG_4_ & n15916;
  assign n18151 = ~P3_REG1_REG_3_ & ~n15856;
  assign n18152 = P3_REG1_REG_3_ & n15856;
  assign n18153 = ~P3_REG1_REG_2_ & ~n15797;
  assign n18154 = P3_REG1_REG_2_ & n15797;
  assign n18155 = P3_REG1_REG_0_ & n15659;
  assign n18156 = ~P3_REG1_REG_1_ & ~n18155;
  assign n18157 = P3_REG1_REG_1_ & n18155;
  assign n18158 = ~n15743 & ~n18157;
  assign n18159 = ~n18156 & ~n18158;
  assign n18160 = ~n18154 & ~n18159;
  assign n18161 = ~n18153 & ~n18160;
  assign n18162 = ~n18152 & ~n18161;
  assign n18163 = ~n18151 & ~n18162;
  assign n18164 = ~n18150 & ~n18163;
  assign n18165 = ~n18149 & ~n18164;
  assign n18166 = ~n18148 & ~n18165;
  assign n18167 = ~n18147 & ~n18166;
  assign n18168 = ~n18146 & ~n18167;
  assign n18169 = ~n18145 & ~n18168;
  assign n18170 = ~n18144 & ~n18169;
  assign n18171 = ~n18143 & ~n18170;
  assign n18172 = ~n18142 & ~n18171;
  assign n18173 = ~n18141 & ~n18172;
  assign n18174 = ~n18140 & ~n18173;
  assign n18175 = ~n18139 & ~n18174;
  assign n18176 = ~n18138 & ~n18175;
  assign n18177 = ~n18137 & ~n18176;
  assign n18178 = ~n18136 & ~n18177;
  assign n18179 = ~n18135 & ~n18178;
  assign n18180 = ~n18134 & ~n18179;
  assign n18181 = ~n18133 & ~n18180;
  assign n18182 = ~n18132 & ~n18181;
  assign n18183 = ~n18131 & ~n18182;
  assign n18184 = ~n18130 & ~n18183;
  assign n18185 = ~n18129 & ~n18184;
  assign n18186 = ~P3_REG1_REG_15_ & ~n18185;
  assign n18187 = P3_REG1_REG_15_ & n18185;
  assign n18188 = ~n16622 & ~n18187;
  assign n18189 = ~n18186 & ~n18188;
  assign n18190 = ~n18128 & ~n18189;
  assign n18191 = ~n18127 & ~n18190;
  assign n18192 = ~n18126 & ~n18191;
  assign n18193 = ~n18125 & ~n18192;
  assign n18194 = ~P3_REG1_REG_18_ & ~n16818;
  assign n18195 = n18193 & ~n18194;
  assign n18196 = n18124 & ~n18195;
  assign n18197 = n18123 & ~n18194;
  assign n18198 = ~n18120 & ~n18193;
  assign n18199 = n18197 & ~n18198;
  assign n18200 = ~n18196 & ~n18199;
  assign n18201 = n15652 & ~n18034;
  assign n18202 = ~n18200 & n18201;
  assign n18203 = ~n18036 & ~n18119;
  assign n18204 = ~n18202 & n18203;
  assign n18205 = n18026 & ~n18204;
  assign n18206 = P3_STATE_REG & n15492;
  assign n3780 = n15503 & n18206;
  assign n18208 = ~n15655 & n3780;
  assign n18209 = P3_STATE_REG & ~n15492;
  assign n18210 = ~n18025 & n18209;
  assign n18211 = n15655 & n18210;
  assign n18212 = ~n18208 & ~n18211;
  assign n18213 = ~n15634 & ~n18212;
  assign n18214 = P3_REG2_REG_19_ & ~n15652;
  assign n18215 = P3_REG1_REG_19_ & n15652;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = n15634 & ~n18216;
  assign n18218 = ~n15634 & n18216;
  assign n18219 = ~n18217 & ~n18218;
  assign n18220 = P3_REG2_REG_18_ & ~n15652;
  assign n18221 = P3_REG1_REG_18_ & n15652;
  assign n18222 = ~n18220 & ~n18221;
  assign n18223 = P3_REG2_REG_17_ & ~n15652;
  assign n18224 = P3_REG1_REG_17_ & n15652;
  assign n18225 = ~n18223 & ~n18224;
  assign n18226 = n16749 & ~n18225;
  assign n18227 = ~n16749 & n18225;
  assign n18228 = P3_REG2_REG_16_ & ~n15652;
  assign n18229 = P3_REG1_REG_16_ & n15652;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = ~n16683 & n18230;
  assign n18232 = P3_REG2_REG_15_ & ~n15652;
  assign n18233 = P3_REG1_REG_15_ & n15652;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = n16622 & ~n18234;
  assign n18236 = n16683 & ~n18230;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = P3_REG2_REG_14_ & ~n15652;
  assign n18239 = P3_REG1_REG_14_ & n15652;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = n16559 & ~n18240;
  assign n18242 = ~n16622 & n18234;
  assign n18243 = ~n18231 & ~n18242;
  assign n18244 = n18241 & n18243;
  assign n18245 = n18237 & ~n18244;
  assign n18246 = ~n18231 & ~n18245;
  assign n18247 = ~n16559 & n18240;
  assign n18248 = P3_REG2_REG_13_ & ~n15652;
  assign n18249 = P3_REG1_REG_13_ & n15652;
  assign n18250 = ~n18248 & ~n18249;
  assign n18251 = n16495 & ~n18250;
  assign n18252 = ~n16495 & n18250;
  assign n18253 = P3_REG2_REG_12_ & ~n15652;
  assign n18254 = P3_REG1_REG_12_ & n15652;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = n16429 & ~n18255;
  assign n18257 = ~n16429 & n18255;
  assign n18258 = P3_REG2_REG_11_ & ~n15652;
  assign n18259 = P3_REG1_REG_11_ & n15652;
  assign n18260 = ~n18258 & ~n18259;
  assign n18261 = ~n16357 & n18260;
  assign n18262 = P3_REG2_REG_10_ & ~n15652;
  assign n18263 = P3_REG1_REG_10_ & n15652;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = n16299 & ~n18264;
  assign n18266 = n16357 & ~n18260;
  assign n18267 = ~n18265 & ~n18266;
  assign n18268 = P3_REG2_REG_9_ & ~n15652;
  assign n18269 = P3_REG1_REG_9_ & n15652;
  assign n18270 = ~n18268 & ~n18269;
  assign n18271 = n16234 & ~n18270;
  assign n18272 = ~n16299 & n18264;
  assign n18273 = ~n18261 & ~n18272;
  assign n18274 = n18271 & n18273;
  assign n18275 = n18267 & ~n18274;
  assign n18276 = ~n18261 & ~n18275;
  assign n18277 = ~n16234 & n18270;
  assign n18278 = P3_REG2_REG_8_ & ~n15652;
  assign n18279 = P3_REG1_REG_8_ & n15652;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = P3_REG2_REG_7_ & ~n15652;
  assign n18282 = P3_REG1_REG_7_ & n15652;
  assign n18283 = ~n18281 & ~n18282;
  assign n18284 = n16108 & ~n18283;
  assign n18285 = n18280 & ~n18284;
  assign n18286 = n16172 & ~n18285;
  assign n18287 = ~n18280 & n18284;
  assign n18288 = ~n16172 & n18280;
  assign n18289 = ~n16108 & n18283;
  assign n18290 = P3_REG2_REG_6_ & ~n15652;
  assign n18291 = P3_REG1_REG_6_ & n15652;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~n16041 & n18292;
  assign n18294 = P3_REG2_REG_5_ & ~n15652;
  assign n18295 = P3_REG1_REG_5_ & n15652;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = n15982 & ~n18296;
  assign n18298 = n16041 & ~n18292;
  assign n18299 = ~n18297 & ~n18298;
  assign n18300 = P3_REG2_REG_4_ & ~n15652;
  assign n18301 = P3_REG1_REG_4_ & n15652;
  assign n18302 = ~n18300 & ~n18301;
  assign n18303 = n15916 & ~n18302;
  assign n18304 = ~n15982 & n18296;
  assign n18305 = ~n18293 & ~n18304;
  assign n18306 = n18303 & n18305;
  assign n18307 = n18299 & ~n18306;
  assign n18308 = ~n18293 & ~n18307;
  assign n18309 = ~n15916 & n18302;
  assign n18310 = P3_REG2_REG_3_ & ~n15652;
  assign n18311 = P3_REG1_REG_3_ & n15652;
  assign n18312 = ~n18310 & ~n18311;
  assign n18313 = P3_REG2_REG_2_ & ~n15652;
  assign n18314 = P3_REG1_REG_2_ & n15652;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = n15797 & ~n18315;
  assign n18317 = n18312 & ~n18316;
  assign n18318 = n15856 & ~n18317;
  assign n18319 = ~n18312 & n18316;
  assign n18320 = ~n15856 & n18312;
  assign n18321 = ~n15797 & n18315;
  assign n18322 = P3_REG2_REG_1_ & ~n15652;
  assign n18323 = P3_REG1_REG_1_ & n15652;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = P3_REG2_REG_0_ & ~n15652;
  assign n18326 = P3_REG1_REG_0_ & n15652;
  assign n18327 = ~n18325 & ~n18326;
  assign n18328 = ~n15659 & n18327;
  assign n18329 = ~n18324 & ~n18328;
  assign n18330 = n18324 & n18328;
  assign n18331 = n15743 & ~n18330;
  assign n18332 = ~n18329 & ~n18331;
  assign n18333 = ~n18320 & ~n18321;
  assign n18334 = ~n18332 & n18333;
  assign n18335 = ~n18318 & ~n18319;
  assign n18336 = ~n18334 & n18335;
  assign n18337 = n18305 & ~n18309;
  assign n18338 = ~n18336 & n18337;
  assign n18339 = ~n18308 & ~n18338;
  assign n18340 = ~n18288 & ~n18289;
  assign n18341 = ~n18339 & n18340;
  assign n18342 = ~n18286 & ~n18287;
  assign n18343 = ~n18341 & n18342;
  assign n18344 = n18273 & ~n18277;
  assign n18345 = ~n18343 & n18344;
  assign n18346 = ~n18276 & ~n18345;
  assign n18347 = ~n18257 & ~n18346;
  assign n18348 = ~n18256 & ~n18347;
  assign n18349 = ~n18252 & ~n18348;
  assign n18350 = ~n18251 & ~n18349;
  assign n18351 = n18243 & ~n18247;
  assign n18352 = ~n18350 & n18351;
  assign n18353 = ~n18246 & ~n18352;
  assign n18354 = ~n18227 & ~n18353;
  assign n18355 = ~n18226 & ~n18354;
  assign n18356 = ~n18222 & ~n18355;
  assign n18357 = n18222 & n18355;
  assign n18358 = n16818 & ~n18357;
  assign n18359 = ~n18356 & ~n18358;
  assign n18360 = ~n18219 & ~n18359;
  assign n18361 = n18219 & n18359;
  assign n18362 = ~n18360 & ~n18361;
  assign n18363 = ~n15656 & ~n15765;
  assign n18364 = n3780 & ~n18363;
  assign n18365 = ~n18362 & n18364;
  assign n18366 = n15692 & n18210;
  assign n18367 = ~n18117 & n18366;
  assign n18368 = P3_ADDR_REG_19_ & n18025;
  assign n18369 = P3_REG3_REG_19_ & ~P3_STATE_REG;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = n15652 & n18210;
  assign n18372 = ~n18200 & n18371;
  assign n18373 = n18370 & ~n18372;
  assign n18374 = ~n18213 & ~n18365;
  assign n18375 = ~n18367 & n18374;
  assign n18376 = n18373 & n18375;
  assign n3360 = n18205 | ~n18376;
  assign n18378 = ~n16818 & n18035;
  assign n18379 = ~n18037 & ~n18111;
  assign n18380 = ~n18110 & ~n18379;
  assign n18381 = n18110 & n18379;
  assign n18382 = ~n18380 & ~n18381;
  assign n18383 = n18118 & ~n18382;
  assign n18384 = ~n18120 & ~n18194;
  assign n18385 = ~n18193 & ~n18384;
  assign n18386 = n18193 & n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = n18201 & ~n18387;
  assign n18389 = ~n18378 & ~n18383;
  assign n18390 = ~n18388 & n18389;
  assign n18391 = n18026 & ~n18390;
  assign n18392 = ~n16818 & ~n18212;
  assign n18393 = n16818 & ~n18222;
  assign n18394 = ~n16818 & n18222;
  assign n18395 = ~n18393 & ~n18394;
  assign n18396 = ~n18355 & ~n18395;
  assign n18397 = n18355 & n18395;
  assign n18398 = ~n18396 & ~n18397;
  assign n18399 = n18364 & ~n18398;
  assign n18400 = n18366 & ~n18382;
  assign n18401 = P3_ADDR_REG_18_ & n18025;
  assign n18402 = P3_REG3_REG_18_ & ~P3_STATE_REG;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = n18371 & ~n18387;
  assign n18405 = n18403 & ~n18404;
  assign n18406 = ~n18392 & ~n18399;
  assign n18407 = ~n18400 & n18406;
  assign n18408 = n18405 & n18407;
  assign n3365 = n18391 | ~n18408;
  assign n18410 = ~n16749 & n18035;
  assign n18411 = ~n18042 & ~n18043;
  assign n18412 = ~n18108 & ~n18411;
  assign n18413 = n18108 & n18411;
  assign n18414 = ~n18412 & ~n18413;
  assign n18415 = n18118 & ~n18414;
  assign n18416 = ~n18125 & ~n18126;
  assign n18417 = ~n18191 & ~n18416;
  assign n18418 = n18191 & n18416;
  assign n18419 = ~n18417 & ~n18418;
  assign n18420 = n18201 & ~n18419;
  assign n18421 = ~n18410 & ~n18415;
  assign n18422 = ~n18420 & n18421;
  assign n18423 = n18026 & ~n18422;
  assign n18424 = ~n16749 & ~n18212;
  assign n18425 = ~n18226 & ~n18227;
  assign n18426 = ~n18353 & ~n18425;
  assign n18427 = n18353 & n18425;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = n18364 & ~n18428;
  assign n18430 = n18366 & ~n18414;
  assign n18431 = P3_ADDR_REG_17_ & n18025;
  assign n18432 = P3_REG3_REG_17_ & ~P3_STATE_REG;
  assign n18433 = ~n18431 & ~n18432;
  assign n18434 = n18371 & ~n18419;
  assign n18435 = n18433 & ~n18434;
  assign n18436 = ~n18424 & ~n18429;
  assign n18437 = ~n18430 & n18436;
  assign n18438 = n18435 & n18437;
  assign n3370 = n18423 | ~n18438;
  assign n18440 = ~n16683 & n18035;
  assign n18441 = ~n18044 & ~n18045;
  assign n18442 = ~n18106 & ~n18441;
  assign n18443 = n18106 & n18441;
  assign n18444 = ~n18442 & ~n18443;
  assign n18445 = n18118 & ~n18444;
  assign n18446 = ~n18127 & ~n18128;
  assign n18447 = ~n18189 & ~n18446;
  assign n18448 = n18189 & n18446;
  assign n18449 = ~n18447 & ~n18448;
  assign n18450 = n18201 & ~n18449;
  assign n18451 = ~n18440 & ~n18445;
  assign n18452 = ~n18450 & n18451;
  assign n18453 = n18026 & ~n18452;
  assign n18454 = ~n16683 & ~n18212;
  assign n18455 = ~n18231 & ~n18236;
  assign n18456 = ~n18247 & ~n18350;
  assign n18457 = ~n18241 & ~n18456;
  assign n18458 = ~n18235 & n18457;
  assign n18459 = ~n18242 & ~n18455;
  assign n18460 = ~n18458 & n18459;
  assign n18461 = ~n18242 & ~n18457;
  assign n18462 = ~n18231 & n18237;
  assign n18463 = ~n18461 & n18462;
  assign n18464 = ~n18460 & ~n18463;
  assign n18465 = n18364 & ~n18464;
  assign n18466 = n18366 & ~n18444;
  assign n18467 = P3_ADDR_REG_16_ & n18025;
  assign n18468 = P3_REG3_REG_16_ & ~P3_STATE_REG;
  assign n18469 = ~n18467 & ~n18468;
  assign n18470 = n18371 & ~n18449;
  assign n18471 = n18469 & ~n18470;
  assign n18472 = ~n18454 & ~n18465;
  assign n18473 = ~n18466 & n18472;
  assign n18474 = n18471 & n18473;
  assign n3375 = n18453 | ~n18474;
  assign n18476 = ~n16622 & n18035;
  assign n18477 = P3_REG2_REG_15_ & n16622;
  assign n18478 = ~P3_REG2_REG_15_ & ~n16622;
  assign n18479 = ~n18477 & ~n18478;
  assign n18480 = ~n18102 & ~n18479;
  assign n18481 = n18102 & n18479;
  assign n18482 = ~n18480 & ~n18481;
  assign n18483 = n18118 & ~n18482;
  assign n18484 = P3_REG1_REG_15_ & n16622;
  assign n18485 = ~P3_REG1_REG_15_ & ~n16622;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = ~n18185 & ~n18486;
  assign n18488 = n18185 & n18486;
  assign n18489 = ~n18487 & ~n18488;
  assign n18490 = n18201 & ~n18489;
  assign n18491 = ~n18476 & ~n18483;
  assign n18492 = ~n18490 & n18491;
  assign n18493 = n18026 & ~n18492;
  assign n18494 = ~n16622 & ~n18212;
  assign n18495 = ~n18235 & ~n18242;
  assign n18496 = n18457 & n18495;
  assign n18497 = ~n18457 & ~n18495;
  assign n18498 = ~n18496 & ~n18497;
  assign n18499 = n18364 & ~n18498;
  assign n18500 = n18366 & ~n18482;
  assign n18501 = P3_ADDR_REG_15_ & n18025;
  assign n18502 = P3_REG3_REG_15_ & ~P3_STATE_REG;
  assign n18503 = ~n18501 & ~n18502;
  assign n18504 = n18371 & ~n18489;
  assign n18505 = n18503 & ~n18504;
  assign n18506 = ~n18494 & ~n18499;
  assign n18507 = ~n18500 & n18506;
  assign n18508 = n18505 & n18507;
  assign n3380 = n18493 | ~n18508;
  assign n18510 = ~n16559 & n18035;
  assign n18511 = ~n18046 & ~n18047;
  assign n18512 = ~n18100 & ~n18511;
  assign n18513 = n18100 & n18511;
  assign n18514 = ~n18512 & ~n18513;
  assign n18515 = n18118 & ~n18514;
  assign n18516 = ~n18129 & ~n18130;
  assign n18517 = ~n18183 & ~n18516;
  assign n18518 = n18183 & n18516;
  assign n18519 = ~n18517 & ~n18518;
  assign n18520 = n18201 & ~n18519;
  assign n18521 = ~n18510 & ~n18515;
  assign n18522 = ~n18520 & n18521;
  assign n18523 = n18026 & ~n18522;
  assign n18524 = ~n16559 & ~n18212;
  assign n18525 = ~n18241 & ~n18247;
  assign n18526 = n18350 & n18525;
  assign n18527 = ~n18350 & ~n18525;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = n18364 & ~n18528;
  assign n18530 = n18366 & ~n18514;
  assign n18531 = P3_ADDR_REG_14_ & n18025;
  assign n18532 = P3_REG3_REG_14_ & ~P3_STATE_REG;
  assign n18533 = ~n18531 & ~n18532;
  assign n18534 = n18371 & ~n18519;
  assign n18535 = n18533 & ~n18534;
  assign n18536 = ~n18524 & ~n18529;
  assign n18537 = ~n18530 & n18536;
  assign n18538 = n18535 & n18537;
  assign n3385 = n18523 | ~n18538;
  assign n18540 = ~n16495 & n18035;
  assign n18541 = ~n18048 & ~n18049;
  assign n18542 = ~n18098 & ~n18541;
  assign n18543 = n18098 & n18541;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = n18118 & ~n18544;
  assign n18546 = ~n18131 & ~n18132;
  assign n18547 = ~n18181 & ~n18546;
  assign n18548 = n18181 & n18546;
  assign n18549 = ~n18547 & ~n18548;
  assign n18550 = n18201 & ~n18549;
  assign n18551 = ~n18540 & ~n18545;
  assign n18552 = ~n18550 & n18551;
  assign n18553 = n18026 & ~n18552;
  assign n18554 = ~n16495 & ~n18212;
  assign n18555 = ~n18251 & ~n18252;
  assign n18556 = ~n18348 & ~n18555;
  assign n18557 = n18348 & n18555;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = n18364 & ~n18558;
  assign n18560 = n18366 & ~n18544;
  assign n18561 = P3_ADDR_REG_13_ & n18025;
  assign n18562 = P3_REG3_REG_13_ & ~P3_STATE_REG;
  assign n18563 = ~n18561 & ~n18562;
  assign n18564 = n18371 & ~n18549;
  assign n18565 = n18563 & ~n18564;
  assign n18566 = ~n18554 & ~n18559;
  assign n18567 = ~n18560 & n18566;
  assign n18568 = n18565 & n18567;
  assign n3390 = n18553 | ~n18568;
  assign n18570 = ~n16429 & n18035;
  assign n18571 = ~n18050 & ~n18051;
  assign n18572 = ~n18096 & ~n18571;
  assign n18573 = n18096 & n18571;
  assign n18574 = ~n18572 & ~n18573;
  assign n18575 = n18118 & ~n18574;
  assign n18576 = ~n18133 & ~n18134;
  assign n18577 = ~n18179 & ~n18576;
  assign n18578 = n18179 & n18576;
  assign n18579 = ~n18577 & ~n18578;
  assign n18580 = n18201 & ~n18579;
  assign n18581 = ~n18570 & ~n18575;
  assign n18582 = ~n18580 & n18581;
  assign n18583 = n18026 & ~n18582;
  assign n18584 = ~n16429 & ~n18212;
  assign n18585 = ~n18256 & ~n18257;
  assign n18586 = ~n18346 & ~n18585;
  assign n18587 = n18346 & n18585;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = n18364 & ~n18588;
  assign n18590 = n18366 & ~n18574;
  assign n18591 = P3_ADDR_REG_12_ & n18025;
  assign n18592 = P3_REG3_REG_12_ & ~P3_STATE_REG;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = n18371 & ~n18579;
  assign n18595 = n18593 & ~n18594;
  assign n18596 = ~n18584 & ~n18589;
  assign n18597 = ~n18590 & n18596;
  assign n18598 = n18595 & n18597;
  assign n3395 = n18583 | ~n18598;
  assign n18600 = ~n16357 & n18035;
  assign n18601 = ~n18052 & ~n18053;
  assign n18602 = ~n18094 & ~n18601;
  assign n18603 = n18094 & n18601;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = n18118 & ~n18604;
  assign n18606 = ~n18135 & ~n18136;
  assign n18607 = ~n18177 & ~n18606;
  assign n18608 = n18177 & n18606;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = n18201 & ~n18609;
  assign n18611 = ~n18600 & ~n18605;
  assign n18612 = ~n18610 & n18611;
  assign n18613 = n18026 & ~n18612;
  assign n18614 = ~n16357 & ~n18212;
  assign n18615 = ~n18261 & ~n18266;
  assign n18616 = ~n18277 & ~n18343;
  assign n18617 = ~n18271 & ~n18616;
  assign n18618 = ~n18265 & n18617;
  assign n18619 = ~n18272 & ~n18615;
  assign n18620 = ~n18618 & n18619;
  assign n18621 = ~n18272 & ~n18617;
  assign n18622 = ~n18261 & n18267;
  assign n18623 = ~n18621 & n18622;
  assign n18624 = ~n18620 & ~n18623;
  assign n18625 = n18364 & ~n18624;
  assign n18626 = n18366 & ~n18604;
  assign n18627 = P3_ADDR_REG_11_ & n18025;
  assign n18628 = P3_REG3_REG_11_ & ~P3_STATE_REG;
  assign n18629 = ~n18627 & ~n18628;
  assign n18630 = n18371 & ~n18609;
  assign n18631 = n18629 & ~n18630;
  assign n18632 = ~n18614 & ~n18625;
  assign n18633 = ~n18626 & n18632;
  assign n18634 = n18631 & n18633;
  assign n3400 = n18613 | ~n18634;
  assign n18636 = ~n16299 & n18035;
  assign n18637 = ~n18054 & ~n18055;
  assign n18638 = ~n18092 & ~n18637;
  assign n18639 = n18092 & n18637;
  assign n18640 = ~n18638 & ~n18639;
  assign n18641 = n18118 & ~n18640;
  assign n18642 = ~n18137 & ~n18138;
  assign n18643 = ~n18175 & ~n18642;
  assign n18644 = n18175 & n18642;
  assign n18645 = ~n18643 & ~n18644;
  assign n18646 = n18201 & ~n18645;
  assign n18647 = ~n18636 & ~n18641;
  assign n18648 = ~n18646 & n18647;
  assign n18649 = n18026 & ~n18648;
  assign n18650 = ~n16299 & ~n18212;
  assign n18651 = ~n18265 & ~n18272;
  assign n18652 = n18617 & n18651;
  assign n18653 = ~n18617 & ~n18651;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = n18364 & ~n18654;
  assign n18656 = n18366 & ~n18640;
  assign n18657 = P3_ADDR_REG_10_ & n18025;
  assign n18658 = P3_REG3_REG_10_ & ~P3_STATE_REG;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 = n18371 & ~n18645;
  assign n18661 = n18659 & ~n18660;
  assign n18662 = ~n18650 & ~n18655;
  assign n18663 = ~n18656 & n18662;
  assign n18664 = n18661 & n18663;
  assign n3405 = n18649 | ~n18664;
  assign n18666 = ~n16234 & n18035;
  assign n18667 = ~n18056 & ~n18057;
  assign n18668 = ~n18090 & ~n18667;
  assign n18669 = n18090 & n18667;
  assign n18670 = ~n18668 & ~n18669;
  assign n18671 = n18118 & ~n18670;
  assign n18672 = ~n18139 & ~n18140;
  assign n18673 = ~n18173 & ~n18672;
  assign n18674 = n18173 & n18672;
  assign n18675 = ~n18673 & ~n18674;
  assign n18676 = n18201 & ~n18675;
  assign n18677 = ~n18666 & ~n18671;
  assign n18678 = ~n18676 & n18677;
  assign n18679 = n18026 & ~n18678;
  assign n18680 = ~n16234 & ~n18212;
  assign n18681 = ~n18271 & ~n18277;
  assign n18682 = n18343 & n18681;
  assign n18683 = ~n18343 & ~n18681;
  assign n18684 = ~n18682 & ~n18683;
  assign n18685 = n18364 & ~n18684;
  assign n18686 = n18366 & ~n18670;
  assign n18687 = P3_ADDR_REG_9_ & n18025;
  assign n18688 = P3_REG3_REG_9_ & ~P3_STATE_REG;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = n18371 & ~n18675;
  assign n18691 = n18689 & ~n18690;
  assign n18692 = ~n18680 & ~n18685;
  assign n18693 = ~n18686 & n18692;
  assign n18694 = n18691 & n18693;
  assign n3410 = n18679 | ~n18694;
  assign n18696 = ~n16172 & n18035;
  assign n18697 = ~n18058 & ~n18059;
  assign n18698 = ~n18088 & ~n18697;
  assign n18699 = n18088 & n18697;
  assign n18700 = ~n18698 & ~n18699;
  assign n18701 = n18118 & ~n18700;
  assign n18702 = ~n18141 & ~n18142;
  assign n18703 = ~n18171 & ~n18702;
  assign n18704 = n18171 & n18702;
  assign n18705 = ~n18703 & ~n18704;
  assign n18706 = n18201 & ~n18705;
  assign n18707 = ~n18696 & ~n18701;
  assign n18708 = ~n18706 & n18707;
  assign n18709 = n18026 & ~n18708;
  assign n18710 = ~n16172 & ~n18212;
  assign n18711 = n18366 & ~n18700;
  assign n18712 = n16172 & ~n18280;
  assign n18713 = ~n18288 & ~n18712;
  assign n18714 = ~n18284 & n18339;
  assign n18715 = ~n18289 & ~n18713;
  assign n18716 = ~n18714 & n18715;
  assign n18717 = ~n18289 & ~n18339;
  assign n18718 = ~n18284 & n18713;
  assign n18719 = ~n18717 & n18718;
  assign n18720 = ~n18716 & ~n18719;
  assign n18721 = n18364 & ~n18720;
  assign n18722 = P3_ADDR_REG_8_ & n18025;
  assign n18723 = P3_REG3_REG_8_ & ~P3_STATE_REG;
  assign n18724 = ~n18722 & ~n18723;
  assign n18725 = n18371 & ~n18705;
  assign n18726 = n18724 & ~n18725;
  assign n18727 = ~n18710 & ~n18711;
  assign n18728 = ~n18721 & n18727;
  assign n18729 = n18726 & n18728;
  assign n3415 = n18709 | ~n18729;
  assign n18731 = ~n16108 & n18035;
  assign n18732 = ~n18060 & ~n18061;
  assign n18733 = ~n18086 & ~n18732;
  assign n18734 = n18086 & n18732;
  assign n18735 = ~n18733 & ~n18734;
  assign n18736 = n18118 & ~n18735;
  assign n18737 = ~n18143 & ~n18144;
  assign n18738 = ~n18169 & ~n18737;
  assign n18739 = n18169 & n18737;
  assign n18740 = ~n18738 & ~n18739;
  assign n18741 = n18201 & ~n18740;
  assign n18742 = ~n18731 & ~n18736;
  assign n18743 = ~n18741 & n18742;
  assign n18744 = n18026 & ~n18743;
  assign n18745 = ~n16108 & ~n18212;
  assign n18746 = n18366 & ~n18735;
  assign n18747 = ~n18284 & ~n18289;
  assign n18748 = n18339 & n18747;
  assign n18749 = ~n18339 & ~n18747;
  assign n18750 = ~n18748 & ~n18749;
  assign n18751 = n18364 & ~n18750;
  assign n18752 = P3_ADDR_REG_7_ & n18025;
  assign n18753 = P3_REG3_REG_7_ & ~P3_STATE_REG;
  assign n18754 = ~n18752 & ~n18753;
  assign n18755 = n18371 & ~n18740;
  assign n18756 = n18754 & ~n18755;
  assign n18757 = ~n18745 & ~n18746;
  assign n18758 = ~n18751 & n18757;
  assign n18759 = n18756 & n18758;
  assign n3420 = n18744 | ~n18759;
  assign n18761 = ~n16041 & n18035;
  assign n18762 = ~n18062 & ~n18063;
  assign n18763 = ~n18084 & ~n18762;
  assign n18764 = n18084 & n18762;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = n18118 & ~n18765;
  assign n18767 = ~n18145 & ~n18146;
  assign n18768 = ~n18167 & ~n18767;
  assign n18769 = n18167 & n18767;
  assign n18770 = ~n18768 & ~n18769;
  assign n18771 = n18201 & ~n18770;
  assign n18772 = ~n18761 & ~n18766;
  assign n18773 = ~n18771 & n18772;
  assign n18774 = n18026 & ~n18773;
  assign n18775 = n18366 & ~n18765;
  assign n18776 = ~n16041 & ~n18212;
  assign n18777 = P3_ADDR_REG_6_ & n18025;
  assign n18778 = P3_REG3_REG_6_ & ~P3_STATE_REG;
  assign n18779 = ~n18777 & ~n18778;
  assign n18780 = n18371 & ~n18770;
  assign n18781 = n18779 & ~n18780;
  assign n18782 = ~n18775 & ~n18776;
  assign n18783 = n18781 & n18782;
  assign n18784 = ~n18293 & ~n18298;
  assign n18785 = ~n18309 & ~n18336;
  assign n18786 = ~n18303 & ~n18785;
  assign n18787 = ~n18297 & n18786;
  assign n18788 = ~n18304 & ~n18784;
  assign n18789 = ~n18787 & n18788;
  assign n18790 = ~n18304 & ~n18786;
  assign n18791 = ~n18293 & n18299;
  assign n18792 = ~n18790 & n18791;
  assign n18793 = ~n18789 & ~n18792;
  assign n18794 = n18364 & ~n18793;
  assign n18795 = ~n18774 & n18783;
  assign n3425 = n18794 | ~n18795;
  assign n18797 = ~n15982 & n18035;
  assign n18798 = ~n18064 & ~n18065;
  assign n18799 = ~n18082 & ~n18798;
  assign n18800 = n18082 & n18798;
  assign n18801 = ~n18799 & ~n18800;
  assign n18802 = n18118 & ~n18801;
  assign n18803 = ~n18147 & ~n18148;
  assign n18804 = ~n18165 & ~n18803;
  assign n18805 = n18165 & n18803;
  assign n18806 = ~n18804 & ~n18805;
  assign n18807 = n18201 & ~n18806;
  assign n18808 = ~n18797 & ~n18802;
  assign n18809 = ~n18807 & n18808;
  assign n18810 = n18026 & ~n18809;
  assign n18811 = n18366 & ~n18801;
  assign n18812 = ~n15982 & ~n18212;
  assign n18813 = ~n18811 & ~n18812;
  assign n18814 = P3_ADDR_REG_5_ & n18025;
  assign n18815 = P3_REG3_REG_5_ & ~P3_STATE_REG;
  assign n18816 = ~n18814 & ~n18815;
  assign n18817 = n18371 & ~n18806;
  assign n18818 = n18816 & ~n18817;
  assign n18819 = ~n18297 & ~n18304;
  assign n18820 = n18786 & n18819;
  assign n18821 = ~n18786 & ~n18819;
  assign n18822 = ~n18820 & ~n18821;
  assign n18823 = n18364 & ~n18822;
  assign n18824 = ~n18810 & n18813;
  assign n18825 = n18818 & n18824;
  assign n3430 = n18823 | ~n18825;
  assign n18827 = ~n18066 & ~n18067;
  assign n18828 = ~n18080 & ~n18827;
  assign n18829 = n18080 & n18827;
  assign n18830 = ~n18828 & ~n18829;
  assign n18831 = n18366 & ~n18830;
  assign n18832 = ~n15916 & n18035;
  assign n18833 = n18118 & ~n18830;
  assign n18834 = ~n18149 & ~n18150;
  assign n18835 = ~n18163 & ~n18834;
  assign n18836 = n18163 & n18834;
  assign n18837 = ~n18835 & ~n18836;
  assign n18838 = n18201 & ~n18837;
  assign n18839 = ~n18832 & ~n18833;
  assign n18840 = ~n18838 & n18839;
  assign n18841 = n18026 & ~n18840;
  assign n18842 = ~n15916 & ~n18212;
  assign n18843 = P3_ADDR_REG_4_ & n18025;
  assign n18844 = P3_REG3_REG_4_ & ~P3_STATE_REG;
  assign n18845 = ~n18843 & ~n18844;
  assign n18846 = n18371 & ~n18837;
  assign n18847 = n18845 & ~n18846;
  assign n18848 = ~n18303 & ~n18309;
  assign n18849 = n18336 & n18848;
  assign n18850 = ~n18336 & ~n18848;
  assign n18851 = ~n18849 & ~n18850;
  assign n18852 = n18364 & ~n18851;
  assign n18853 = ~n18842 & n18847;
  assign n18854 = ~n18852 & n18853;
  assign n18855 = ~n18831 & ~n18841;
  assign n3435 = ~n18854 | ~n18855;
  assign n18857 = ~n18068 & ~n18069;
  assign n18858 = ~n18078 & ~n18857;
  assign n18859 = n18078 & n18857;
  assign n18860 = ~n18858 & ~n18859;
  assign n18861 = n18366 & ~n18860;
  assign n18862 = ~n15856 & n18035;
  assign n18863 = n18118 & ~n18860;
  assign n18864 = ~n18151 & ~n18152;
  assign n18865 = ~n18161 & ~n18864;
  assign n18866 = n18161 & n18864;
  assign n18867 = ~n18865 & ~n18866;
  assign n18868 = n18201 & ~n18867;
  assign n18869 = ~n18862 & ~n18863;
  assign n18870 = ~n18868 & n18869;
  assign n18871 = n18026 & ~n18870;
  assign n18872 = ~n15856 & ~n18212;
  assign n18873 = P3_ADDR_REG_3_ & n18025;
  assign n18874 = P3_REG3_REG_3_ & ~P3_STATE_REG;
  assign n18875 = ~n18873 & ~n18874;
  assign n18876 = n18371 & ~n18867;
  assign n18877 = n18875 & ~n18876;
  assign n18878 = n15856 & ~n18312;
  assign n18879 = ~n18320 & ~n18878;
  assign n18880 = ~n18316 & n18332;
  assign n18881 = ~n18321 & ~n18879;
  assign n18882 = ~n18880 & n18881;
  assign n18883 = ~n18321 & ~n18332;
  assign n18884 = ~n18316 & n18879;
  assign n18885 = ~n18883 & n18884;
  assign n18886 = ~n18882 & ~n18885;
  assign n18887 = n18364 & ~n18886;
  assign n18888 = ~n18872 & n18877;
  assign n18889 = ~n18887 & n18888;
  assign n18890 = ~n18861 & ~n18871;
  assign n3440 = ~n18889 | ~n18890;
  assign n18892 = ~n15797 & n18035;
  assign n18893 = ~n18070 & ~n18071;
  assign n18894 = ~n18076 & ~n18893;
  assign n18895 = n18076 & n18893;
  assign n18896 = ~n18894 & ~n18895;
  assign n18897 = n18118 & ~n18896;
  assign n18898 = ~n18153 & ~n18154;
  assign n18899 = ~n18159 & ~n18898;
  assign n18900 = n18159 & n18898;
  assign n18901 = ~n18899 & ~n18900;
  assign n18902 = n18201 & ~n18901;
  assign n18903 = ~n18892 & ~n18897;
  assign n18904 = ~n18902 & n18903;
  assign n18905 = n18026 & ~n18904;
  assign n18906 = ~n15797 & ~n18212;
  assign n18907 = n18366 & ~n18896;
  assign n18908 = ~n18316 & ~n18321;
  assign n18909 = n18332 & n18908;
  assign n18910 = ~n18332 & ~n18908;
  assign n18911 = ~n18909 & ~n18910;
  assign n18912 = n18364 & ~n18911;
  assign n18913 = P3_ADDR_REG_2_ & n18025;
  assign n18914 = P3_REG3_REG_2_ & ~P3_STATE_REG;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = n18371 & ~n18901;
  assign n18917 = n18915 & ~n18916;
  assign n18918 = ~n18906 & ~n18907;
  assign n18919 = ~n18912 & n18918;
  assign n18920 = n18917 & n18919;
  assign n3445 = n18905 | ~n18920;
  assign n18922 = ~n15743 & n18035;
  assign n18923 = P3_REG2_REG_1_ & ~n18072;
  assign n18924 = ~P3_REG2_REG_1_ & n18072;
  assign n18925 = ~n18923 & ~n18924;
  assign n18926 = n15743 & ~n18925;
  assign n18927 = ~n15743 & n18925;
  assign n18928 = ~n18926 & ~n18927;
  assign n18929 = n18118 & ~n18928;
  assign n18930 = P3_REG1_REG_1_ & ~n18155;
  assign n18931 = ~P3_REG1_REG_1_ & n18155;
  assign n18932 = ~n18930 & ~n18931;
  assign n18933 = n15743 & ~n18932;
  assign n18934 = ~n15743 & n18932;
  assign n18935 = ~n18933 & ~n18934;
  assign n18936 = n18201 & ~n18935;
  assign n18937 = ~n18922 & ~n18929;
  assign n18938 = ~n18936 & n18937;
  assign n18939 = n18026 & ~n18938;
  assign n18940 = ~n15743 & ~n18212;
  assign n18941 = n15743 & ~n18324;
  assign n18942 = ~n15743 & n18324;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = ~n18328 & ~n18943;
  assign n18945 = n18328 & n18943;
  assign n18946 = ~n18944 & ~n18945;
  assign n18947 = n18364 & ~n18946;
  assign n18948 = n18366 & ~n18928;
  assign n18949 = P3_ADDR_REG_1_ & n18025;
  assign n18950 = P3_REG3_REG_1_ & ~P3_STATE_REG;
  assign n18951 = ~n18949 & ~n18950;
  assign n18952 = n18371 & ~n18935;
  assign n18953 = n18951 & ~n18952;
  assign n18954 = ~n18940 & ~n18947;
  assign n18955 = ~n18948 & n18954;
  assign n18956 = n18953 & n18955;
  assign n3450 = n18939 | ~n18956;
  assign n18958 = ~n15659 & n18035;
  assign n18959 = ~P3_REG2_REG_0_ & ~n15659;
  assign n18960 = ~n18072 & ~n18959;
  assign n18961 = n18118 & ~n18960;
  assign n18962 = ~P3_REG1_REG_0_ & ~n15659;
  assign n18963 = ~n18155 & ~n18962;
  assign n18964 = n18201 & ~n18963;
  assign n18965 = ~n18958 & ~n18961;
  assign n18966 = ~n18964 & n18965;
  assign n18967 = n18026 & ~n18966;
  assign n18968 = ~n15659 & ~n18212;
  assign n18969 = n15659 & ~n18327;
  assign n18970 = ~n18328 & ~n18969;
  assign n18971 = n18364 & ~n18970;
  assign n18972 = n18366 & ~n18960;
  assign n18973 = P3_ADDR_REG_0_ & n18025;
  assign n18974 = P3_REG3_REG_0_ & ~P3_STATE_REG;
  assign n18975 = ~n18973 & ~n18974;
  assign n18976 = n18371 & ~n18963;
  assign n18977 = n18975 & ~n18976;
  assign n18978 = ~n18968 & ~n18971;
  assign n18979 = ~n18972 & n18978;
  assign n18980 = n18977 & n18979;
  assign n3455 = n18967 | ~n18980;
  assign n18982 = ~n15685 & n3780;
  assign n18983 = P3_DATAO_REG_0_ & ~n3780;
  assign n3460 = n18982 | n18983;
  assign n18985 = ~n15701 & n3780;
  assign n18986 = P3_DATAO_REG_1_ & ~n3780;
  assign n3465 = n18985 | n18986;
  assign n18988 = ~n15739 & n3780;
  assign n18989 = P3_DATAO_REG_2_ & ~n3780;
  assign n3470 = n18988 | n18989;
  assign n18991 = ~n15793 & n3780;
  assign n18992 = P3_DATAO_REG_3_ & ~n3780;
  assign n3475 = n18991 | n18992;
  assign n18994 = ~n15852 & n3780;
  assign n18995 = P3_DATAO_REG_4_ & ~n3780;
  assign n3480 = n18994 | n18995;
  assign n18997 = ~n15912 & n3780;
  assign n18998 = P3_DATAO_REG_5_ & ~n3780;
  assign n3485 = n18997 | n18998;
  assign n19000 = ~n15978 & n3780;
  assign n19001 = P3_DATAO_REG_6_ & ~n3780;
  assign n3490 = n19000 | n19001;
  assign n19003 = ~n16037 & n3780;
  assign n19004 = P3_DATAO_REG_7_ & ~n3780;
  assign n3495 = n19003 | n19004;
  assign n19006 = ~n16104 & n3780;
  assign n19007 = P3_DATAO_REG_8_ & ~n3780;
  assign n3500 = n19006 | n19007;
  assign n19009 = ~n16168 & n3780;
  assign n19010 = P3_DATAO_REG_9_ & ~n3780;
  assign n3505 = n19009 | n19010;
  assign n19012 = ~n16230 & n3780;
  assign n19013 = P3_DATAO_REG_10_ & ~n3780;
  assign n3510 = n19012 | n19013;
  assign n19015 = ~n16295 & n3780;
  assign n19016 = P3_DATAO_REG_11_ & ~n3780;
  assign n3515 = n19015 | n19016;
  assign n19018 = ~n16353 & n3780;
  assign n19019 = P3_DATAO_REG_12_ & ~n3780;
  assign n3520 = n19018 | n19019;
  assign n19021 = ~n16425 & n3780;
  assign n19022 = P3_DATAO_REG_13_ & ~n3780;
  assign n3525 = n19021 | n19022;
  assign n19024 = ~n16491 & n3780;
  assign n19025 = P3_DATAO_REG_14_ & ~n3780;
  assign n3530 = n19024 | n19025;
  assign n19027 = ~n16555 & n3780;
  assign n19028 = P3_DATAO_REG_15_ & ~n3780;
  assign n3535 = n19027 | n19028;
  assign n19030 = ~n16618 & n3780;
  assign n19031 = P3_DATAO_REG_16_ & ~n3780;
  assign n3540 = n19030 | n19031;
  assign n19033 = ~n16679 & n3780;
  assign n19034 = P3_DATAO_REG_17_ & ~n3780;
  assign n3545 = n19033 | n19034;
  assign n19036 = ~n16745 & n3780;
  assign n19037 = P3_DATAO_REG_18_ & ~n3780;
  assign n3550 = n19036 | n19037;
  assign n19039 = ~n16814 & n3780;
  assign n19040 = P3_DATAO_REG_19_ & ~n3780;
  assign n3555 = n19039 | n19040;
  assign n19042 = ~n16879 & n3780;
  assign n19043 = P3_DATAO_REG_20_ & ~n3780;
  assign n3560 = n19042 | n19043;
  assign n19045 = ~n16940 & n3780;
  assign n19046 = P3_DATAO_REG_21_ & ~n3780;
  assign n3565 = n19045 | n19046;
  assign n19048 = ~n16998 & n3780;
  assign n19049 = P3_DATAO_REG_22_ & ~n3780;
  assign n3570 = n19048 | n19049;
  assign n19051 = ~n17057 & n3780;
  assign n19052 = P3_DATAO_REG_23_ & ~n3780;
  assign n3575 = n19051 | n19052;
  assign n19054 = ~n17118 & n3780;
  assign n19055 = P3_DATAO_REG_24_ & ~n3780;
  assign n3580 = n19054 | n19055;
  assign n19057 = ~n17177 & n3780;
  assign n19058 = P3_DATAO_REG_25_ & ~n3780;
  assign n3585 = n19057 | n19058;
  assign n19060 = ~n17240 & n3780;
  assign n19061 = P3_DATAO_REG_26_ & ~n3780;
  assign n3590 = n19060 | n19061;
  assign n19063 = ~n17297 & n3780;
  assign n19064 = P3_DATAO_REG_27_ & ~n3780;
  assign n3595 = n19063 | n19064;
  assign n19066 = ~n17358 & n3780;
  assign n19067 = P3_DATAO_REG_28_ & ~n3780;
  assign n3600 = n19066 | n19067;
  assign n19069 = ~n17414 & n3780;
  assign n19070 = P3_DATAO_REG_29_ & ~n3780;
  assign n3605 = n19069 | n19070;
  assign n19072 = ~n17499 & n3780;
  assign n19073 = P3_DATAO_REG_30_ & ~n3780;
  assign n3610 = n19072 | n19073;
  assign n19075 = ~n17541 & n3780;
  assign n19076 = P3_DATAO_REG_31_ & ~n3780;
  assign n3615 = n19075 | n19076;
  assign n19078 = ~n15492 & ~n15621;
  assign n19079 = n15645 & n15766;
  assign n19080 = n15492 & ~n19079;
  assign n19081 = ~n19078 & ~n19080;
  assign n19082 = n18024 & n19081;
  assign n19083 = P3_B_REG & ~n19082;
  assign n19084 = n15492 & ~n15624;
  assign n19085 = n15643 & n19084;
  assign n19086 = n15667 & ~n15705;
  assign n19087 = ~n15624 & n15665;
  assign n19088 = ~n15711 & ~n19087;
  assign n19089 = ~n15641 & n19088;
  assign n19090 = n19086 & n19089;
  assign n19091 = ~n17541 & ~n19090;
  assign n19092 = ~n15624 & n15640;
  assign n19093 = ~n15492 & ~n15624;
  assign n19094 = n15643 & n19093;
  assign n19095 = ~n19092 & ~n19094;
  assign n19096 = n17549 & ~n19095;
  assign n19097 = ~n19091 & ~n19096;
  assign n19098 = n17549 & ~n19090;
  assign n19099 = ~n17541 & ~n19095;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = ~n19085 & n19097;
  assign n19102 = ~n19100 & n19101;
  assign n19103 = n19085 & ~n19097;
  assign n19104 = n19100 & n19103;
  assign n19105 = ~n19102 & ~n19104;
  assign n19106 = ~n19097 & n19100;
  assign n19107 = n19097 & ~n19100;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = n17543 & ~n19090;
  assign n19110 = ~n17499 & ~n19095;
  assign n19111 = ~n19109 & ~n19110;
  assign n19112 = n19108 & n19111;
  assign n19113 = ~n17499 & ~n19090;
  assign n19114 = n17543 & ~n19095;
  assign n19115 = ~n19113 & ~n19114;
  assign n19116 = n19108 & ~n19115;
  assign n19117 = ~n19112 & ~n19116;
  assign n19118 = ~n16940 & ~n19090;
  assign n19119 = n17000 & ~n19095;
  assign n19120 = ~n15492 & ~n19118;
  assign n19121 = ~n19119 & n19120;
  assign n19122 = n15492 & ~n16879;
  assign n19123 = ~n16940 & ~n19095;
  assign n19124 = n17000 & ~n19090;
  assign n19125 = ~n19122 & ~n19123;
  assign n19126 = ~n19124 & n19125;
  assign n19127 = ~n19121 & n19126;
  assign n19128 = ~n16879 & ~n19090;
  assign n19129 = n16942 & ~n19095;
  assign n19130 = ~n15492 & ~n19128;
  assign n19131 = ~n19129 & n19130;
  assign n19132 = n15492 & ~n16814;
  assign n19133 = ~n16879 & ~n19095;
  assign n19134 = n16942 & ~n19090;
  assign n19135 = ~n19132 & ~n19133;
  assign n19136 = ~n19134 & n19135;
  assign n19137 = ~n19131 & n19136;
  assign n19138 = ~n16814 & ~n19090;
  assign n19139 = ~n16883 & ~n19095;
  assign n19140 = ~n15492 & ~n19138;
  assign n19141 = ~n19139 & n19140;
  assign n19142 = ~n16814 & ~n19095;
  assign n19143 = n15492 & ~n16745;
  assign n19144 = ~n16883 & ~n19090;
  assign n19145 = ~n19142 & ~n19143;
  assign n19146 = ~n19144 & n19145;
  assign n19147 = ~n19141 & n19146;
  assign n19148 = n19131 & ~n19136;
  assign n19149 = n19147 & ~n19148;
  assign n19150 = ~n19137 & ~n19149;
  assign n19151 = n19121 & ~n19126;
  assign n19152 = ~n19150 & ~n19151;
  assign n19153 = ~n16998 & ~n19090;
  assign n19154 = n17059 & ~n19095;
  assign n19155 = ~n15492 & ~n19153;
  assign n19156 = ~n19154 & n19155;
  assign n19157 = n15492 & ~n16940;
  assign n19158 = ~n16998 & ~n19095;
  assign n19159 = n17059 & ~n19090;
  assign n19160 = ~n19157 & ~n19158;
  assign n19161 = ~n19159 & n19160;
  assign n19162 = ~n19156 & n19161;
  assign n19163 = ~n17057 & ~n19090;
  assign n19164 = n17120 & ~n19095;
  assign n19165 = ~n15492 & ~n19163;
  assign n19166 = ~n19164 & n19165;
  assign n19167 = n15492 & ~n16998;
  assign n19168 = ~n17057 & ~n19095;
  assign n19169 = n17120 & ~n19090;
  assign n19170 = ~n19167 & ~n19168;
  assign n19171 = ~n19169 & n19170;
  assign n19172 = ~n19166 & n19171;
  assign n19173 = ~n19127 & ~n19152;
  assign n19174 = ~n19162 & n19173;
  assign n19175 = ~n19172 & n19174;
  assign n19176 = ~n19148 & ~n19151;
  assign n19177 = ~n16745 & ~n19095;
  assign n19178 = n15492 & ~n16679;
  assign n19179 = ~n16821 & ~n19090;
  assign n19180 = ~n19177 & ~n19178;
  assign n19181 = ~n19179 & n19180;
  assign n19182 = ~n16745 & ~n19090;
  assign n19183 = ~n16821 & ~n19095;
  assign n19184 = ~n15492 & ~n19182;
  assign n19185 = ~n19183 & n19184;
  assign n19186 = ~n16679 & ~n19095;
  assign n19187 = n15492 & ~n16618;
  assign n19188 = ~n16752 & ~n19090;
  assign n19189 = ~n19186 & ~n19187;
  assign n19190 = ~n19188 & n19189;
  assign n19191 = ~n16679 & ~n19090;
  assign n19192 = ~n16752 & ~n19095;
  assign n19193 = ~n15492 & ~n19191;
  assign n19194 = ~n19192 & n19193;
  assign n19195 = ~n19190 & n19194;
  assign n19196 = ~n16618 & ~n19095;
  assign n19197 = n15492 & ~n16555;
  assign n19198 = ~n16686 & ~n19090;
  assign n19199 = ~n19196 & ~n19197;
  assign n19200 = ~n19198 & n19199;
  assign n19201 = ~n16618 & ~n19090;
  assign n19202 = ~n16686 & ~n19095;
  assign n19203 = ~n15492 & ~n19201;
  assign n19204 = ~n19202 & n19203;
  assign n19205 = ~n19200 & n19204;
  assign n19206 = ~n16175 & ~n19095;
  assign n19207 = ~n15492 & ~n19206;
  assign n19208 = ~n16104 & ~n19090;
  assign n19209 = n19207 & ~n19208;
  assign n19210 = ~n16104 & ~n19095;
  assign n19211 = ~n16175 & ~n19090;
  assign n19212 = n15492 & ~n16037;
  assign n19213 = ~n19210 & ~n19211;
  assign n19214 = ~n19212 & n19213;
  assign n19215 = ~n19209 & n19214;
  assign n19216 = ~n16111 & ~n19095;
  assign n19217 = ~n15492 & ~n19216;
  assign n19218 = ~n16037 & ~n19090;
  assign n19219 = n19217 & ~n19218;
  assign n19220 = ~n16037 & ~n19095;
  assign n19221 = ~n16111 & ~n19090;
  assign n19222 = n15492 & ~n15978;
  assign n19223 = ~n19220 & ~n19221;
  assign n19224 = ~n19222 & n19223;
  assign n19225 = ~n19219 & n19224;
  assign n19226 = ~n15739 & ~n19095;
  assign n19227 = ~n15800 & ~n19090;
  assign n19228 = n15492 & ~n15701;
  assign n19229 = ~n19226 & ~n19227;
  assign n19230 = ~n19228 & n19229;
  assign n19231 = ~n15800 & ~n19095;
  assign n19232 = ~n15492 & ~n19231;
  assign n19233 = ~n15739 & ~n19090;
  assign n19234 = n19232 & ~n19233;
  assign n19235 = ~n19230 & n19234;
  assign n19236 = ~n15793 & ~n19095;
  assign n19237 = ~n15859 & ~n19090;
  assign n19238 = n15492 & ~n15739;
  assign n19239 = ~n19236 & ~n19237;
  assign n19240 = ~n19238 & n19239;
  assign n19241 = ~n15859 & ~n19095;
  assign n19242 = ~n15492 & ~n19241;
  assign n19243 = ~n15793 & ~n19090;
  assign n19244 = n19242 & ~n19243;
  assign n19245 = ~n19240 & n19244;
  assign n19246 = ~n19235 & ~n19245;
  assign n19247 = n19230 & ~n19234;
  assign n19248 = ~n15746 & ~n19095;
  assign n19249 = ~n15492 & ~n19248;
  assign n19250 = ~n15701 & ~n19090;
  assign n19251 = n19249 & ~n19250;
  assign n19252 = ~n15701 & ~n19095;
  assign n19253 = ~n15746 & ~n19090;
  assign n19254 = n15492 & ~n15685;
  assign n19255 = ~n19252 & ~n19253;
  assign n19256 = ~n19254 & n19255;
  assign n19257 = ~n19251 & n19256;
  assign n19258 = ~n19247 & ~n19257;
  assign n19259 = n19246 & ~n19258;
  assign n19260 = n19240 & ~n19244;
  assign n19261 = ~n15685 & ~n19095;
  assign n19262 = ~n15662 & ~n19090;
  assign n19263 = ~n19261 & ~n19262;
  assign n19264 = ~n15662 & ~n19095;
  assign n19265 = ~n15492 & ~n19264;
  assign n19266 = ~n15685 & ~n19090;
  assign n19267 = n19265 & ~n19266;
  assign n19268 = n15621 & ~n15624;
  assign n19269 = ~n15492 & n19268;
  assign n19270 = ~n19267 & ~n19269;
  assign n19271 = ~n19263 & ~n19270;
  assign n19272 = n19251 & ~n19256;
  assign n19273 = n19267 & n19269;
  assign n19274 = n19246 & ~n19271;
  assign n19275 = ~n19272 & n19274;
  assign n19276 = ~n19273 & n19275;
  assign n19277 = ~n16044 & ~n19095;
  assign n19278 = ~n15492 & ~n19277;
  assign n19279 = ~n15978 & ~n19090;
  assign n19280 = n19278 & ~n19279;
  assign n19281 = ~n15978 & ~n19095;
  assign n19282 = ~n16044 & ~n19090;
  assign n19283 = n15492 & ~n15912;
  assign n19284 = ~n19281 & ~n19282;
  assign n19285 = ~n19283 & n19284;
  assign n19286 = ~n19280 & n19285;
  assign n19287 = ~n15985 & ~n19095;
  assign n19288 = ~n15492 & ~n19287;
  assign n19289 = ~n15912 & ~n19090;
  assign n19290 = n19288 & ~n19289;
  assign n19291 = ~n15912 & ~n19095;
  assign n19292 = ~n15985 & ~n19090;
  assign n19293 = n15492 & ~n15852;
  assign n19294 = ~n19291 & ~n19292;
  assign n19295 = ~n19293 & n19294;
  assign n19296 = ~n19290 & n19295;
  assign n19297 = ~n19286 & ~n19296;
  assign n19298 = ~n15919 & ~n19095;
  assign n19299 = ~n15492 & ~n19298;
  assign n19300 = ~n15852 & ~n19090;
  assign n19301 = n19299 & ~n19300;
  assign n19302 = ~n15852 & ~n19095;
  assign n19303 = ~n15919 & ~n19090;
  assign n19304 = n15492 & ~n15793;
  assign n19305 = ~n19302 & ~n19303;
  assign n19306 = ~n19304 & n19305;
  assign n19307 = ~n19301 & n19306;
  assign n19308 = n19297 & ~n19307;
  assign n19309 = ~n19259 & ~n19260;
  assign n19310 = ~n19276 & n19309;
  assign n19311 = n19308 & n19310;
  assign n19312 = n19301 & ~n19306;
  assign n19313 = n19297 & n19312;
  assign n19314 = n19280 & ~n19285;
  assign n19315 = n19219 & ~n19224;
  assign n19316 = n19290 & ~n19295;
  assign n19317 = ~n19286 & n19316;
  assign n19318 = ~n19315 & ~n19317;
  assign n19319 = ~n19313 & ~n19314;
  assign n19320 = n19318 & n19319;
  assign n19321 = ~n19311 & n19320;
  assign n19322 = ~n19225 & ~n19321;
  assign n19323 = n19209 & ~n19214;
  assign n19324 = ~n19322 & ~n19323;
  assign n19325 = ~n19215 & ~n19324;
  assign n19326 = ~n16168 & ~n19095;
  assign n19327 = ~n16237 & ~n19090;
  assign n19328 = n15492 & ~n16104;
  assign n19329 = ~n19326 & ~n19327;
  assign n19330 = ~n19328 & n19329;
  assign n19331 = ~n16237 & ~n19095;
  assign n19332 = ~n15492 & ~n19331;
  assign n19333 = ~n16168 & ~n19090;
  assign n19334 = n19332 & ~n19333;
  assign n19335 = ~n19330 & n19334;
  assign n19336 = ~n19325 & ~n19335;
  assign n19337 = ~n16432 & ~n19095;
  assign n19338 = ~n15492 & ~n19337;
  assign n19339 = ~n16353 & ~n19090;
  assign n19340 = n19338 & ~n19339;
  assign n19341 = ~n16353 & ~n19095;
  assign n19342 = ~n16432 & ~n19090;
  assign n19343 = n15492 & ~n16295;
  assign n19344 = ~n19341 & ~n19342;
  assign n19345 = ~n19343 & n19344;
  assign n19346 = ~n19340 & n19345;
  assign n19347 = ~n16360 & ~n19095;
  assign n19348 = ~n15492 & ~n19347;
  assign n19349 = ~n16295 & ~n19090;
  assign n19350 = n19348 & ~n19349;
  assign n19351 = ~n16295 & ~n19095;
  assign n19352 = ~n16360 & ~n19090;
  assign n19353 = n15492 & ~n16230;
  assign n19354 = ~n19351 & ~n19352;
  assign n19355 = ~n19353 & n19354;
  assign n19356 = ~n19350 & n19355;
  assign n19357 = ~n19346 & ~n19356;
  assign n19358 = n19330 & ~n19334;
  assign n19359 = ~n16302 & ~n19095;
  assign n19360 = ~n15492 & ~n19359;
  assign n19361 = ~n16230 & ~n19090;
  assign n19362 = n19360 & ~n19361;
  assign n19363 = ~n16230 & ~n19095;
  assign n19364 = ~n16302 & ~n19090;
  assign n19365 = n15492 & ~n16168;
  assign n19366 = ~n19363 & ~n19364;
  assign n19367 = ~n19365 & n19366;
  assign n19368 = ~n19362 & n19367;
  assign n19369 = ~n19358 & ~n19368;
  assign n19370 = n19357 & n19369;
  assign n19371 = ~n19336 & n19370;
  assign n19372 = n19350 & ~n19355;
  assign n19373 = ~n19346 & n19372;
  assign n19374 = n19362 & ~n19367;
  assign n19375 = n19357 & n19374;
  assign n19376 = ~n16425 & ~n19095;
  assign n19377 = ~n16498 & ~n19090;
  assign n19378 = n15492 & ~n16353;
  assign n19379 = ~n19376 & ~n19377;
  assign n19380 = ~n19378 & n19379;
  assign n19381 = ~n16498 & ~n19095;
  assign n19382 = ~n15492 & ~n19381;
  assign n19383 = ~n16425 & ~n19090;
  assign n19384 = n19382 & ~n19383;
  assign n19385 = ~n19380 & n19384;
  assign n19386 = n19340 & ~n19345;
  assign n19387 = ~n19385 & ~n19386;
  assign n19388 = ~n16555 & ~n19095;
  assign n19389 = n15492 & ~n16491;
  assign n19390 = ~n16625 & ~n19090;
  assign n19391 = ~n19388 & ~n19389;
  assign n19392 = ~n19390 & n19391;
  assign n19393 = ~n16555 & ~n19090;
  assign n19394 = ~n16625 & ~n19095;
  assign n19395 = ~n15492 & ~n19393;
  assign n19396 = ~n19394 & n19395;
  assign n19397 = ~n19392 & n19396;
  assign n19398 = ~n16491 & ~n19095;
  assign n19399 = n15492 & ~n16425;
  assign n19400 = ~n16562 & ~n19090;
  assign n19401 = ~n19398 & ~n19399;
  assign n19402 = ~n19400 & n19401;
  assign n19403 = ~n16491 & ~n19090;
  assign n19404 = ~n16562 & ~n19095;
  assign n19405 = ~n15492 & ~n19403;
  assign n19406 = ~n19404 & n19405;
  assign n19407 = ~n19402 & n19406;
  assign n19408 = ~n19397 & ~n19407;
  assign n19409 = n19387 & n19408;
  assign n19410 = ~n19373 & ~n19375;
  assign n19411 = n19409 & n19410;
  assign n19412 = ~n19371 & n19411;
  assign n19413 = n19380 & ~n19384;
  assign n19414 = n19408 & n19413;
  assign n19415 = n19402 & ~n19406;
  assign n19416 = ~n19397 & n19415;
  assign n19417 = n19200 & ~n19204;
  assign n19418 = n19392 & ~n19396;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = ~n19414 & ~n19416;
  assign n19421 = n19419 & n19420;
  assign n19422 = ~n19412 & n19421;
  assign n19423 = ~n19205 & ~n19422;
  assign n19424 = n19190 & ~n19194;
  assign n19425 = ~n19423 & ~n19424;
  assign n19426 = ~n19195 & ~n19425;
  assign n19427 = ~n19185 & n19426;
  assign n19428 = ~n19181 & ~n19427;
  assign n19429 = n19141 & ~n19146;
  assign n19430 = n19185 & ~n19426;
  assign n19431 = ~n19429 & ~n19430;
  assign n19432 = n19176 & ~n19428;
  assign n19433 = n19431 & n19432;
  assign n19434 = ~n17118 & ~n19090;
  assign n19435 = n17179 & ~n19095;
  assign n19436 = ~n15492 & ~n19434;
  assign n19437 = ~n19435 & n19436;
  assign n19438 = n15492 & ~n17057;
  assign n19439 = ~n17118 & ~n19095;
  assign n19440 = n17179 & ~n19090;
  assign n19441 = ~n19438 & ~n19439;
  assign n19442 = ~n19440 & n19441;
  assign n19443 = ~n19437 & n19442;
  assign n19444 = n19175 & ~n19433;
  assign n19445 = ~n19443 & n19444;
  assign n19446 = n15492 & ~n17240;
  assign n19447 = ~n17297 & ~n19095;
  assign n19448 = n17360 & ~n19090;
  assign n19449 = ~n19446 & ~n19447;
  assign n19450 = ~n19448 & n19449;
  assign n19451 = ~n17297 & ~n19090;
  assign n19452 = n17360 & ~n19095;
  assign n19453 = ~n15492 & ~n19451;
  assign n19454 = ~n19452 & n19453;
  assign n19455 = ~n19450 & n19454;
  assign n19456 = n15492 & ~n17177;
  assign n19457 = ~n17240 & ~n19095;
  assign n19458 = n17299 & ~n19090;
  assign n19459 = ~n19456 & ~n19457;
  assign n19460 = ~n19458 & n19459;
  assign n19461 = ~n17240 & ~n19090;
  assign n19462 = n17299 & ~n19095;
  assign n19463 = ~n15492 & ~n19461;
  assign n19464 = ~n19462 & n19463;
  assign n19465 = ~n19460 & n19464;
  assign n19466 = ~n19455 & ~n19465;
  assign n19467 = n15492 & ~n17297;
  assign n19468 = ~n17358 & ~n19095;
  assign n19469 = n17416 & ~n19090;
  assign n19470 = ~n19467 & ~n19468;
  assign n19471 = ~n19469 & n19470;
  assign n19472 = ~n17358 & ~n19090;
  assign n19473 = n17416 & ~n19095;
  assign n19474 = ~n15492 & ~n19472;
  assign n19475 = ~n19473 & n19474;
  assign n19476 = ~n19471 & n19475;
  assign n19477 = n19437 & ~n19442;
  assign n19478 = n19166 & ~n19171;
  assign n19479 = n19156 & ~n19161;
  assign n19480 = ~n19478 & ~n19479;
  assign n19481 = ~n19172 & ~n19480;
  assign n19482 = ~n19443 & n19481;
  assign n19483 = n15492 & ~n17118;
  assign n19484 = ~n17177 & ~n19095;
  assign n19485 = n17242 & ~n19090;
  assign n19486 = ~n19483 & ~n19484;
  assign n19487 = ~n19485 & n19486;
  assign n19488 = ~n17177 & ~n19090;
  assign n19489 = n17242 & ~n19095;
  assign n19490 = ~n15492 & ~n19488;
  assign n19491 = ~n19489 & n19490;
  assign n19492 = ~n19487 & n19491;
  assign n19493 = ~n19477 & ~n19482;
  assign n19494 = ~n19492 & n19493;
  assign n19495 = n15492 & ~n17358;
  assign n19496 = ~n17414 & ~n19095;
  assign n19497 = n17473 & ~n19090;
  assign n19498 = ~n19495 & ~n19496;
  assign n19499 = ~n19497 & n19498;
  assign n19500 = ~n17414 & ~n19090;
  assign n19501 = n17473 & ~n19095;
  assign n19502 = ~n15492 & ~n19500;
  assign n19503 = ~n19501 & n19502;
  assign n19504 = ~n19499 & n19503;
  assign n19505 = ~n19445 & n19466;
  assign n19506 = ~n19476 & n19505;
  assign n19507 = n19494 & n19506;
  assign n19508 = ~n19504 & n19507;
  assign n19509 = ~n19117 & n19508;
  assign n19510 = n19487 & ~n19491;
  assign n19511 = n19460 & ~n19464;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = n19466 & ~n19512;
  assign n19514 = ~n19476 & n19513;
  assign n19515 = ~n19504 & n19514;
  assign n19516 = n19471 & ~n19475;
  assign n19517 = n19450 & ~n19454;
  assign n19518 = ~n19476 & n19517;
  assign n19519 = ~n19516 & ~n19518;
  assign n19520 = n19503 & n19519;
  assign n19521 = n19499 & ~n19520;
  assign n19522 = n19111 & ~n19115;
  assign n19523 = ~n19503 & ~n19519;
  assign n19524 = ~n19522 & ~n19523;
  assign n19525 = ~n19515 & ~n19521;
  assign n19526 = n19524 & n19525;
  assign n19527 = ~n19117 & ~n19526;
  assign n19528 = n19105 & ~n19509;
  assign n19529 = ~n19527 & n19528;
  assign n19530 = n15505 & n19079;
  assign n19531 = n19529 & n19530;
  assign n19532 = n15492 & ~n19083;
  assign n19533 = ~n19531 & n19532;
  assign n19534 = ~P3_STATE_REG & ~n19083;
  assign n19535 = ~n19533 & ~n19534;
  assign n19536 = n15662 & n15685;
  assign n19537 = ~n15760 & ~n19536;
  assign n19538 = ~n15759 & ~n19537;
  assign n19539 = ~n16638 & ~n16639;
  assign n19540 = ~n16511 & ~n16512;
  assign n19541 = ~n19539 & ~n19540;
  assign n19542 = ~n16199 & ~n16263;
  assign n19543 = n19538 & n19541;
  assign n19544 = n19542 & n19543;
  assign n19545 = ~n16843 & n19544;
  assign n19546 = ~n15998 & ~n15999;
  assign n19547 = ~n16129 & ~n16130;
  assign n19548 = ~n15817 & ~n19546;
  assign n19549 = ~n19547 & n19548;
  assign n19550 = ~n16702 & ~n16703;
  assign n19551 = ~n16073 & ~n16455;
  assign n19552 = ~n19550 & n19551;
  assign n19553 = ~n16770 & ~n16771;
  assign n19554 = n19549 & n19552;
  assign n19555 = ~n16709 & n19554;
  assign n19556 = ~n19553 & n19555;
  assign n19557 = ~n17197 & ~n17198;
  assign n19558 = n17240 & ~n17299;
  assign n19559 = ~n17313 & ~n19558;
  assign n19560 = ~n17204 & ~n19557;
  assign n19561 = ~n17260 & n19560;
  assign n19562 = ~n19559 & n19561;
  assign n19563 = n17499 & ~n17543;
  assign n19564 = ~n17499 & n17543;
  assign n19565 = ~n19563 & ~n19564;
  assign n19566 = n19545 & n19556;
  assign n19567 = ~n16903 & n19566;
  assign n19568 = n19562 & n19567;
  assign n19569 = ~n19565 & n19568;
  assign n19570 = ~n16315 & ~n16316;
  assign n19571 = ~n15945 & ~n19570;
  assign n19572 = ~n16386 & n19571;
  assign n19573 = ~n15881 & n19572;
  assign n19574 = ~n16955 & ~n16956;
  assign n19575 = ~n17072 & ~n17076;
  assign n19576 = ~n19574 & ~n19575;
  assign n19577 = ~n17136 & ~n17137;
  assign n19578 = n17414 & ~n17473;
  assign n19579 = ~n17414 & n17473;
  assign n19580 = ~n19578 & ~n19579;
  assign n19581 = n17358 & ~n17416;
  assign n19582 = ~n17504 & ~n19581;
  assign n19583 = ~n17434 & ~n17440;
  assign n19584 = n17541 & ~n17549;
  assign n19585 = ~n17541 & n17549;
  assign n19586 = ~n19584 & ~n19585;
  assign n19587 = ~n19582 & ~n19583;
  assign n19588 = ~n19586 & n19587;
  assign n19589 = n19573 & n19576;
  assign n19590 = ~n19577 & n19589;
  assign n19591 = ~n19580 & n19590;
  assign n19592 = n19588 & n19591;
  assign n19593 = n19569 & n19592;
  assign n19594 = ~n15634 & ~n19593;
  assign n19595 = n15634 & n19593;
  assign n19596 = ~n19594 & ~n19595;
  assign n19597 = n15624 & ~n19596;
  assign n19598 = ~n15627 & n19597;
  assign n19599 = n15634 & n15691;
  assign n19600 = ~n15634 & ~n15691;
  assign n19601 = ~n19599 & ~n19600;
  assign n19602 = n19529 & ~n19601;
  assign n19603 = ~n19529 & n19601;
  assign n19604 = ~n19602 & ~n19603;
  assign n19605 = n15627 & n19604;
  assign n19606 = ~n17499 & n17541;
  assign n19607 = ~n17541 & ~n19606;
  assign n19608 = n17499 & ~n17541;
  assign n19609 = ~n19606 & ~n19608;
  assign n19610 = n19606 & n19609;
  assign n19611 = ~n19607 & ~n19610;
  assign n19612 = ~n17549 & ~n19611;
  assign n19613 = ~n17499 & ~n19606;
  assign n19614 = n17499 & n19606;
  assign n19615 = ~n19613 & ~n19614;
  assign n19616 = ~n19612 & ~n19615;
  assign n19617 = ~n17543 & n19616;
  assign n19618 = ~n16555 & ~n19606;
  assign n19619 = ~n16555 & n19606;
  assign n19620 = ~n19618 & ~n19619;
  assign n19621 = n16625 & ~n19620;
  assign n19622 = ~n16491 & ~n19606;
  assign n19623 = ~n16491 & n19606;
  assign n19624 = ~n19622 & ~n19623;
  assign n19625 = n16562 & ~n19624;
  assign n19626 = ~n15978 & ~n19606;
  assign n19627 = ~n15978 & n19606;
  assign n19628 = ~n19626 & ~n19627;
  assign n19629 = ~n16044 & n19628;
  assign n19630 = ~n16037 & ~n19606;
  assign n19631 = ~n16037 & n19606;
  assign n19632 = ~n19630 & ~n19631;
  assign n19633 = n16111 & ~n19632;
  assign n19634 = n19629 & ~n19633;
  assign n19635 = ~n15912 & ~n19606;
  assign n19636 = ~n15912 & n19606;
  assign n19637 = ~n19635 & ~n19636;
  assign n19638 = ~n15985 & n19637;
  assign n19639 = n16044 & ~n19628;
  assign n19640 = ~n19633 & ~n19639;
  assign n19641 = n19638 & n19640;
  assign n19642 = ~n16104 & ~n19606;
  assign n19643 = ~n16104 & n19606;
  assign n19644 = ~n19642 & ~n19643;
  assign n19645 = ~n16175 & n19644;
  assign n19646 = ~n16111 & n19632;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = ~n16230 & ~n19606;
  assign n19649 = ~n16230 & n19606;
  assign n19650 = ~n19648 & ~n19649;
  assign n19651 = ~n16302 & n19650;
  assign n19652 = ~n16168 & ~n19606;
  assign n19653 = ~n16168 & n19606;
  assign n19654 = ~n19652 & ~n19653;
  assign n19655 = ~n16237 & n19654;
  assign n19656 = ~n19651 & ~n19655;
  assign n19657 = n19647 & n19656;
  assign n19658 = ~n19634 & ~n19641;
  assign n19659 = n19657 & n19658;
  assign n19660 = ~n15852 & ~n19606;
  assign n19661 = ~n15852 & n19606;
  assign n19662 = ~n19660 & ~n19661;
  assign n19663 = n15919 & ~n19662;
  assign n19664 = ~n15919 & n19662;
  assign n19665 = ~n15793 & ~n19606;
  assign n19666 = ~n15793 & n19606;
  assign n19667 = ~n19665 & ~n19666;
  assign n19668 = ~n15859 & n19667;
  assign n19669 = ~n19664 & ~n19668;
  assign n19670 = n15859 & ~n19667;
  assign n19671 = ~n15739 & ~n19606;
  assign n19672 = ~n15739 & n19606;
  assign n19673 = ~n19671 & ~n19672;
  assign n19674 = n15800 & ~n19673;
  assign n19675 = ~n19670 & ~n19674;
  assign n19676 = n19669 & ~n19675;
  assign n19677 = n15985 & ~n19637;
  assign n19678 = n19640 & ~n19677;
  assign n19679 = ~n19663 & ~n19676;
  assign n19680 = n19678 & n19679;
  assign n19681 = n19659 & ~n19680;
  assign n19682 = ~n15701 & ~n19606;
  assign n19683 = ~n15701 & n19606;
  assign n19684 = ~n19682 & ~n19683;
  assign n19685 = ~n15746 & n19684;
  assign n19686 = ~n15800 & n19673;
  assign n19687 = ~n15685 & ~n19606;
  assign n19688 = ~n15685 & n19606;
  assign n19689 = ~n19687 & ~n19688;
  assign n19690 = ~n15662 & n19689;
  assign n19691 = n15746 & ~n19684;
  assign n19692 = n19690 & ~n19691;
  assign n19693 = ~n19686 & ~n19692;
  assign n19694 = ~n19634 & n19669;
  assign n19695 = n19657 & ~n19685;
  assign n19696 = n19693 & n19695;
  assign n19697 = ~n19641 & n19696;
  assign n19698 = n19694 & n19697;
  assign n19699 = n16175 & ~n19644;
  assign n19700 = n19656 & n19699;
  assign n19701 = n16237 & ~n19654;
  assign n19702 = ~n19651 & n19701;
  assign n19703 = ~n16295 & ~n19606;
  assign n19704 = ~n16295 & n19606;
  assign n19705 = ~n19703 & ~n19704;
  assign n19706 = n16360 & ~n19705;
  assign n19707 = n16302 & ~n19650;
  assign n19708 = ~n19706 & ~n19707;
  assign n19709 = ~n16425 & ~n19606;
  assign n19710 = ~n16425 & n19606;
  assign n19711 = ~n19709 & ~n19710;
  assign n19712 = n16498 & ~n19711;
  assign n19713 = ~n16353 & ~n19606;
  assign n19714 = ~n16353 & n19606;
  assign n19715 = ~n19713 & ~n19714;
  assign n19716 = n16432 & ~n19715;
  assign n19717 = ~n19712 & ~n19716;
  assign n19718 = n19708 & n19717;
  assign n19719 = ~n19700 & ~n19702;
  assign n19720 = n19718 & n19719;
  assign n19721 = ~n19681 & ~n19698;
  assign n19722 = n19720 & n19721;
  assign n19723 = ~n16432 & n19715;
  assign n19724 = ~n19712 & n19723;
  assign n19725 = ~n16498 & n19711;
  assign n19726 = ~n16562 & n19624;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = ~n19724 & n19727;
  assign n19729 = ~n16360 & n19705;
  assign n19730 = n19717 & n19729;
  assign n19731 = n19728 & ~n19730;
  assign n19732 = ~n19722 & n19731;
  assign n19733 = ~n19625 & ~n19732;
  assign n19734 = ~n16625 & n19620;
  assign n19735 = ~n19733 & ~n19734;
  assign n19736 = ~n19621 & ~n19735;
  assign n19737 = ~n16618 & ~n19606;
  assign n19738 = ~n16618 & n19606;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = ~n16686 & n19739;
  assign n19741 = ~n16814 & ~n19606;
  assign n19742 = ~n16814 & n19606;
  assign n19743 = ~n19741 & ~n19742;
  assign n19744 = ~n16883 & n19743;
  assign n19745 = ~n16745 & ~n19606;
  assign n19746 = ~n16745 & n19606;
  assign n19747 = ~n19745 & ~n19746;
  assign n19748 = ~n16821 & n19747;
  assign n19749 = n16883 & ~n19743;
  assign n19750 = n19748 & ~n19749;
  assign n19751 = ~n19744 & ~n19750;
  assign n19752 = ~n16679 & ~n19606;
  assign n19753 = ~n16679 & n19606;
  assign n19754 = ~n19752 & ~n19753;
  assign n19755 = ~n16752 & n19754;
  assign n19756 = n16821 & ~n19747;
  assign n19757 = ~n19749 & ~n19756;
  assign n19758 = n19755 & n19757;
  assign n19759 = ~n16879 & ~n19606;
  assign n19760 = ~n16879 & n19606;
  assign n19761 = ~n19759 & ~n19760;
  assign n19762 = n16942 & n19761;
  assign n19763 = ~n16998 & ~n19606;
  assign n19764 = ~n16998 & n19606;
  assign n19765 = ~n19763 & ~n19764;
  assign n19766 = n17059 & n19765;
  assign n19767 = ~n16940 & ~n19606;
  assign n19768 = ~n16940 & n19606;
  assign n19769 = ~n19767 & ~n19768;
  assign n19770 = n17000 & n19769;
  assign n19771 = ~n19766 & ~n19770;
  assign n19772 = n19751 & ~n19758;
  assign n19773 = ~n19762 & n19772;
  assign n19774 = n19771 & n19773;
  assign n19775 = ~n19736 & ~n19740;
  assign n19776 = n19774 & n19775;
  assign n19777 = n16686 & ~n19739;
  assign n19778 = n16752 & ~n19754;
  assign n19779 = ~n19777 & ~n19778;
  assign n19780 = n19757 & n19779;
  assign n19781 = n19774 & ~n19780;
  assign n19782 = ~n17057 & ~n19606;
  assign n19783 = ~n17057 & n19606;
  assign n19784 = ~n19782 & ~n19783;
  assign n19785 = ~n17120 & ~n19784;
  assign n19786 = ~n17059 & ~n19765;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = ~n16942 & ~n19761;
  assign n19789 = n19771 & n19788;
  assign n19790 = ~n17000 & ~n19769;
  assign n19791 = ~n19766 & n19790;
  assign n19792 = ~n17118 & ~n19606;
  assign n19793 = ~n17118 & n19606;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = ~n17179 & ~n19794;
  assign n19796 = ~n17177 & ~n19606;
  assign n19797 = ~n17177 & n19606;
  assign n19798 = ~n19796 & ~n19797;
  assign n19799 = ~n17242 & ~n19798;
  assign n19800 = ~n19789 & ~n19791;
  assign n19801 = ~n19795 & n19800;
  assign n19802 = ~n19799 & n19801;
  assign n19803 = ~n19776 & ~n19781;
  assign n19804 = n19787 & n19803;
  assign n19805 = n19802 & n19804;
  assign n19806 = n17179 & n19794;
  assign n19807 = n17120 & n19784;
  assign n19808 = ~n19806 & ~n19807;
  assign n19809 = ~n19795 & ~n19808;
  assign n19810 = ~n19799 & n19809;
  assign n19811 = ~n17543 & ~n19612;
  assign n19812 = ~n19616 & ~n19811;
  assign n19813 = ~n17240 & ~n19606;
  assign n19814 = ~n17240 & n19606;
  assign n19815 = ~n19813 & ~n19814;
  assign n19816 = n17299 & n19815;
  assign n19817 = n17242 & n19798;
  assign n19818 = ~n19816 & ~n19817;
  assign n19819 = ~n17297 & ~n19606;
  assign n19820 = ~n17297 & n19606;
  assign n19821 = ~n19819 & ~n19820;
  assign n19822 = n17360 & n19821;
  assign n19823 = ~n17358 & ~n19606;
  assign n19824 = ~n17358 & n19606;
  assign n19825 = ~n19823 & ~n19824;
  assign n19826 = n17416 & n19825;
  assign n19827 = ~n17414 & ~n19606;
  assign n19828 = ~n17414 & n19606;
  assign n19829 = ~n19827 & ~n19828;
  assign n19830 = n17473 & n19829;
  assign n19831 = ~n19822 & ~n19826;
  assign n19832 = ~n19830 & n19831;
  assign n19833 = n19818 & n19832;
  assign n19834 = ~n19805 & ~n19810;
  assign n19835 = ~n19812 & n19834;
  assign n19836 = n19833 & n19835;
  assign n19837 = ~n19821 & n19832;
  assign n19838 = ~n19812 & n19837;
  assign n19839 = ~n17360 & n19838;
  assign n19840 = ~n17416 & ~n19825;
  assign n19841 = ~n19830 & n19840;
  assign n19842 = ~n19812 & n19841;
  assign n19843 = ~n19839 & ~n19842;
  assign n19844 = ~n17473 & ~n19829;
  assign n19845 = ~n19812 & n19844;
  assign n19846 = n17549 & n19611;
  assign n19847 = ~n19815 & n19832;
  assign n19848 = ~n19812 & n19847;
  assign n19849 = ~n17299 & n19848;
  assign n19850 = ~n19845 & ~n19846;
  assign n19851 = ~n19849 & n19850;
  assign n19852 = ~n19617 & ~n19836;
  assign n19853 = n19843 & n19852;
  assign n19854 = n19851 & n19853;
  assign n19855 = n15709 & n19854;
  assign n19856 = n15715 & ~n19854;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = ~n19083 & n19857;
  assign n19859 = ~n19531 & n19858;
  assign n19860 = ~n19598 & ~n19605;
  assign n19861 = n19859 & n19860;
  assign n3620 = n19535 & ~n19861;
  assign n19863 = n15505 & ~n17681;
  assign n19864 = ~n15639 & n19863;
  assign n19865 = n15627 & n15641;
  assign n19866 = ~n15706 & ~n19087;
  assign n19867 = ~n17564 & n19866;
  assign n19868 = ~n19865 & n19867;
  assign n19869 = ~n15711 & n19868;
  assign n19870 = ~n15639 & ~n19869;
  assign n19871 = ~n15618 & n15642;
  assign n19872 = ~n15627 & n15691;
  assign n19873 = n15504 & ~n19872;
  assign n19874 = ~n19092 & n19873;
  assign n19875 = ~n19870 & ~n19871;
  assign n19876 = n19874 & n19875;
  assign n19877 = P3_STATE_REG & ~n19876;
  assign n19878 = ~n19864 & ~n19877;
  assign n19879 = ~n16548 & ~n19878;
  assign n19880 = n15639 & n19863;
  assign n19881 = n15505 & n17671;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~n16625 & ~n19882;
  assign n19884 = n15505 & n15645;
  assign n19885 = n15618 & ~n15693;
  assign n19886 = ~n16618 & n19885;
  assign n19887 = n15618 & ~n15767;
  assign n19888 = ~n16491 & n19887;
  assign n19889 = ~n15618 & ~n16548;
  assign n19890 = ~n19886 & ~n19888;
  assign n19891 = ~n19889 & n19890;
  assign n19892 = n19884 & ~n19891;
  assign n19893 = ~n18502 & ~n19892;
  assign n19894 = ~n15557 & n15624;
  assign n19895 = ~n15627 & n19894;
  assign n19896 = n15627 & n15634;
  assign n19897 = ~n19895 & ~n19896;
  assign n19898 = ~n17665 & n19897;
  assign n19899 = ~n16302 & n19898;
  assign n19900 = n16302 & ~n19898;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = ~n16230 & ~n19901;
  assign n19903 = ~n16432 & n19898;
  assign n19904 = n16432 & ~n19898;
  assign n19905 = ~n19903 & ~n19904;
  assign n19906 = n16353 & n19905;
  assign n19907 = ~n16498 & n19898;
  assign n19908 = n16498 & ~n19898;
  assign n19909 = ~n19907 & ~n19908;
  assign n19910 = n16425 & n19909;
  assign n19911 = ~n19906 & ~n19910;
  assign n19912 = ~n16360 & n19898;
  assign n19913 = n16360 & ~n19898;
  assign n19914 = ~n19912 & ~n19913;
  assign n19915 = n16295 & n19914;
  assign n19916 = n19911 & ~n19915;
  assign n19917 = n19902 & n19916;
  assign n19918 = ~n16425 & ~n19909;
  assign n19919 = ~n16353 & ~n19905;
  assign n19920 = ~n19918 & ~n19919;
  assign n19921 = ~n16295 & ~n19914;
  assign n19922 = n19911 & n19921;
  assign n19923 = n19920 & ~n19922;
  assign n19924 = ~n19910 & ~n19923;
  assign n19925 = ~n19917 & ~n19924;
  assign n19926 = ~n16562 & n19898;
  assign n19927 = n16562 & ~n19898;
  assign n19928 = ~n19926 & ~n19927;
  assign n19929 = n16491 & n19928;
  assign n19930 = ~n19925 & ~n19929;
  assign n19931 = ~n16491 & ~n19928;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = n16230 & n19901;
  assign n19934 = n19916 & ~n19933;
  assign n19935 = ~n19929 & n19934;
  assign n19936 = ~n16111 & n19898;
  assign n19937 = n16111 & ~n19898;
  assign n19938 = ~n19936 & ~n19937;
  assign n19939 = ~n16044 & n19898;
  assign n19940 = n16044 & ~n19898;
  assign n19941 = ~n19939 & ~n19940;
  assign n19942 = ~n15978 & ~n19941;
  assign n19943 = n16037 & ~n19942;
  assign n19944 = ~n19938 & ~n19943;
  assign n19945 = ~n16037 & n19942;
  assign n19946 = ~n15985 & n19898;
  assign n19947 = n15985 & ~n19898;
  assign n19948 = ~n19946 & ~n19947;
  assign n19949 = ~n15912 & ~n19948;
  assign n19950 = n15978 & n19941;
  assign n19951 = n16037 & n19938;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = n19949 & n19952;
  assign n19954 = ~n19944 & ~n19945;
  assign n19955 = ~n19953 & n19954;
  assign n19956 = ~n16175 & n19898;
  assign n19957 = n16175 & ~n19898;
  assign n19958 = ~n19956 & ~n19957;
  assign n19959 = n16104 & n19958;
  assign n19960 = ~n19955 & ~n19959;
  assign n19961 = ~n16104 & ~n19958;
  assign n19962 = ~n19960 & ~n19961;
  assign n19963 = n15912 & n19948;
  assign n19964 = n19952 & ~n19963;
  assign n19965 = ~n19959 & n19964;
  assign n19966 = ~n15800 & n19898;
  assign n19967 = n15800 & ~n19898;
  assign n19968 = ~n19966 & ~n19967;
  assign n19969 = ~n15739 & ~n19968;
  assign n19970 = ~n15793 & n19969;
  assign n19971 = ~n15859 & n19898;
  assign n19972 = n15859 & ~n19898;
  assign n19973 = ~n19971 & ~n19972;
  assign n19974 = n15793 & ~n19969;
  assign n19975 = ~n19973 & ~n19974;
  assign n19976 = ~n19970 & ~n19975;
  assign n19977 = n15739 & n19968;
  assign n19978 = n15793 & n19973;
  assign n19979 = ~n19977 & ~n19978;
  assign n19980 = ~n15662 & n19898;
  assign n19981 = n15662 & ~n19898;
  assign n19982 = ~n19980 & ~n19981;
  assign n19983 = ~n19898 & ~n19982;
  assign n19984 = ~n15746 & n19898;
  assign n19985 = n15746 & ~n19898;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = n15701 & n19986;
  assign n19988 = n19983 & ~n19987;
  assign n19989 = ~n15701 & ~n19986;
  assign n19990 = n19898 & n19982;
  assign n19991 = ~n15685 & ~n19990;
  assign n19992 = ~n19987 & n19991;
  assign n19993 = ~n19988 & ~n19989;
  assign n19994 = ~n19992 & n19993;
  assign n19995 = n19979 & ~n19994;
  assign n19996 = n19976 & ~n19995;
  assign n19997 = ~n15852 & ~n19996;
  assign n19998 = ~n15919 & n19898;
  assign n19999 = n15919 & ~n19898;
  assign n20000 = ~n19998 & ~n19999;
  assign n20001 = ~n19996 & ~n20000;
  assign n20002 = ~n15852 & ~n20000;
  assign n20003 = ~n19997 & ~n20001;
  assign n20004 = ~n20002 & n20003;
  assign n20005 = n19965 & ~n20004;
  assign n20006 = n19962 & ~n20005;
  assign n20007 = ~n16168 & ~n20006;
  assign n20008 = ~n16237 & n19898;
  assign n20009 = n16237 & ~n19898;
  assign n20010 = ~n20008 & ~n20009;
  assign n20011 = ~n20006 & ~n20010;
  assign n20012 = ~n16168 & ~n20010;
  assign n20013 = ~n20007 & ~n20011;
  assign n20014 = ~n20012 & n20013;
  assign n20015 = n19935 & ~n20014;
  assign n20016 = n19932 & ~n20015;
  assign n20017 = ~n16625 & n19898;
  assign n20018 = n16625 & ~n19898;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = n16555 & ~n20019;
  assign n20021 = ~n16555 & n20019;
  assign n20022 = ~n20020 & ~n20021;
  assign n20023 = n20016 & ~n20022;
  assign n20024 = ~n20016 & n20022;
  assign n20025 = ~n20023 & ~n20024;
  assign n20026 = n15618 & n15642;
  assign n20027 = n15639 & ~n19869;
  assign n20028 = ~n20026 & ~n20027;
  assign n20029 = n15505 & ~n20028;
  assign n20030 = ~n20025 & n20029;
  assign n20031 = ~n19879 & ~n19883;
  assign n20032 = n19893 & n20031;
  assign n3625 = n20030 | ~n20032;
  assign n20034 = ~n15639 & ~n17681;
  assign n20035 = n19876 & ~n20034;
  assign n20036 = P3_STATE_REG & ~n20035;
  assign n20037 = ~n17233 & n20036;
  assign n20038 = P3_REG3_REG_26_ & ~P3_STATE_REG;
  assign n20039 = ~n17297 & n19885;
  assign n20040 = ~n17177 & n19887;
  assign n20041 = ~n15618 & ~n17233;
  assign n20042 = ~n20039 & ~n20040;
  assign n20043 = ~n20041 & n20042;
  assign n20044 = n19884 & ~n20043;
  assign n20045 = ~n20038 & ~n20044;
  assign n20046 = n15639 & ~n17681;
  assign n20047 = ~n17671 & ~n20046;
  assign n20048 = n15505 & ~n20047;
  assign n20049 = n17299 & n20048;
  assign n20050 = n17299 & n19898;
  assign n20051 = ~n17299 & ~n19898;
  assign n20052 = ~n20050 & ~n20051;
  assign n20053 = ~n17240 & ~n20052;
  assign n20054 = n17242 & n19898;
  assign n20055 = ~n17242 & ~n19898;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = n17177 & n20056;
  assign n20058 = ~n17240 & ~n20057;
  assign n20059 = ~n20052 & ~n20057;
  assign n20060 = ~n20058 & ~n20059;
  assign n20061 = ~n20053 & ~n20060;
  assign n20062 = n17179 & n19898;
  assign n20063 = ~n17179 & ~n19898;
  assign n20064 = ~n20062 & ~n20063;
  assign n20065 = n17118 & n20064;
  assign n20066 = n17120 & n19898;
  assign n20067 = ~n17120 & ~n19898;
  assign n20068 = ~n20066 & ~n20067;
  assign n20069 = ~n17057 & ~n20068;
  assign n20070 = n17057 & n20068;
  assign n20071 = n17059 & n19898;
  assign n20072 = ~n17059 & ~n19898;
  assign n20073 = ~n20071 & ~n20072;
  assign n20074 = ~n16998 & ~n20073;
  assign n20075 = n16998 & n20073;
  assign n20076 = n17000 & n19898;
  assign n20077 = ~n17000 & ~n19898;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = n16940 & n20078;
  assign n20080 = ~n16940 & ~n20078;
  assign n20081 = n16942 & n19898;
  assign n20082 = ~n16942 & ~n19898;
  assign n20083 = ~n20081 & ~n20082;
  assign n20084 = ~n16879 & ~n20083;
  assign n20085 = ~n20080 & ~n20084;
  assign n20086 = ~n16883 & n19898;
  assign n20087 = n16883 & ~n19898;
  assign n20088 = ~n20086 & ~n20087;
  assign n20089 = ~n16814 & ~n20088;
  assign n20090 = n16879 & n20083;
  assign n20091 = ~n20079 & ~n20090;
  assign n20092 = n20089 & n20091;
  assign n20093 = n20085 & ~n20092;
  assign n20094 = ~n20079 & ~n20093;
  assign n20095 = n16814 & n20088;
  assign n20096 = n20091 & ~n20095;
  assign n20097 = ~n16821 & n19898;
  assign n20098 = n16821 & ~n19898;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~n16745 & ~n20099;
  assign n20101 = n16745 & n20099;
  assign n20102 = ~n16686 & n19898;
  assign n20103 = n16686 & ~n19898;
  assign n20104 = ~n20102 & ~n20103;
  assign n20105 = ~n16618 & ~n20104;
  assign n20106 = ~n16679 & n20105;
  assign n20107 = ~n16752 & n19898;
  assign n20108 = n16752 & ~n19898;
  assign n20109 = ~n20107 & ~n20108;
  assign n20110 = n16679 & ~n20105;
  assign n20111 = ~n20109 & ~n20110;
  assign n20112 = ~n20106 & ~n20111;
  assign n20113 = n16618 & n20104;
  assign n20114 = n16679 & n20109;
  assign n20115 = ~n20113 & ~n20114;
  assign n20116 = ~n16555 & ~n20019;
  assign n20117 = n16555 & n20019;
  assign n20118 = ~n20016 & ~n20117;
  assign n20119 = ~n20116 & ~n20118;
  assign n20120 = n20115 & ~n20119;
  assign n20121 = n20112 & ~n20120;
  assign n20122 = ~n20101 & ~n20121;
  assign n20123 = ~n20100 & ~n20122;
  assign n20124 = n20096 & ~n20123;
  assign n20125 = ~n20094 & ~n20124;
  assign n20126 = ~n20075 & ~n20125;
  assign n20127 = ~n20074 & ~n20126;
  assign n20128 = ~n20070 & ~n20127;
  assign n20129 = ~n20069 & ~n20128;
  assign n20130 = ~n20065 & ~n20129;
  assign n20131 = n20061 & n20130;
  assign n20132 = ~n17118 & ~n20064;
  assign n20133 = ~n17177 & ~n20056;
  assign n20134 = ~n20132 & ~n20133;
  assign n20135 = n17240 & ~n20052;
  assign n20136 = ~n17240 & n20052;
  assign n20137 = ~n20135 & ~n20136;
  assign n20138 = n20134 & n20137;
  assign n20139 = ~n20130 & n20138;
  assign n20140 = ~n20053 & n20133;
  assign n20141 = ~n20060 & n20140;
  assign n20142 = n20057 & n20137;
  assign n20143 = ~n20053 & n20132;
  assign n20144 = ~n20060 & n20143;
  assign n20145 = ~n20141 & ~n20142;
  assign n20146 = ~n20144 & n20145;
  assign n20147 = ~n20131 & ~n20139;
  assign n20148 = n20146 & n20147;
  assign n20149 = n20029 & n20148;
  assign n20150 = ~n20037 & n20045;
  assign n20151 = ~n20049 & n20150;
  assign n3630 = n20149 | ~n20151;
  assign n20153 = ~n15971 & ~n19878;
  assign n20154 = ~n16044 & ~n19882;
  assign n20155 = ~n16037 & n19885;
  assign n20156 = ~n15912 & n19887;
  assign n20157 = ~n15618 & ~n15971;
  assign n20158 = ~n20155 & ~n20156;
  assign n20159 = ~n20157 & n20158;
  assign n20160 = n19884 & ~n20159;
  assign n20161 = ~n18778 & ~n20160;
  assign n20162 = n15978 & ~n19941;
  assign n20163 = ~n15978 & n19941;
  assign n20164 = ~n20162 & ~n20163;
  assign n20165 = ~n19963 & ~n20004;
  assign n20166 = ~n19949 & ~n20165;
  assign n20167 = ~n20164 & n20166;
  assign n20168 = ~n19942 & ~n19950;
  assign n20169 = ~n20166 & ~n20168;
  assign n20170 = ~n20167 & ~n20169;
  assign n20171 = n20029 & ~n20170;
  assign n20172 = ~n20153 & ~n20154;
  assign n20173 = n20161 & n20172;
  assign n3635 = n20171 | ~n20173;
  assign n20175 = ~n16738 & ~n19878;
  assign n20176 = ~n16821 & ~n19882;
  assign n20177 = ~n16814 & n19885;
  assign n20178 = ~n16679 & n19887;
  assign n20179 = ~n15618 & ~n16738;
  assign n20180 = ~n20177 & ~n20178;
  assign n20181 = ~n20179 & n20180;
  assign n20182 = n19884 & ~n20181;
  assign n20183 = ~n18402 & ~n20182;
  assign n20184 = n16745 & ~n20099;
  assign n20185 = ~n16745 & n20099;
  assign n20186 = ~n20184 & ~n20185;
  assign n20187 = n20121 & ~n20186;
  assign n20188 = ~n20121 & n20186;
  assign n20189 = ~n20187 & ~n20188;
  assign n20190 = n20029 & ~n20189;
  assign n20191 = ~n20175 & ~n20176;
  assign n20192 = n20183 & n20191;
  assign n3640 = n20190 | ~n20192;
  assign n20194 = n15739 & ~n19968;
  assign n20195 = ~n15739 & n19968;
  assign n20196 = ~n20194 & ~n20195;
  assign n20197 = n19994 & ~n20196;
  assign n20198 = ~n19969 & ~n19977;
  assign n20199 = ~n19994 & ~n20198;
  assign n20200 = ~n20197 & ~n20199;
  assign n20201 = n20029 & ~n20200;
  assign n20202 = ~n15800 & ~n19882;
  assign n20203 = ~n20201 & ~n20202;
  assign n20204 = P3_REG3_REG_2_ & ~n19878;
  assign n20205 = ~n15793 & n19885;
  assign n20206 = ~n15701 & n19887;
  assign n20207 = P3_REG3_REG_2_ & ~n15618;
  assign n20208 = ~n20205 & ~n20206;
  assign n20209 = ~n20207 & n20208;
  assign n20210 = n19884 & ~n20209;
  assign n20211 = ~n18914 & ~n20210;
  assign n20212 = n20203 & ~n20204;
  assign n3645 = ~n20211 | ~n20212;
  assign n20214 = ~n16288 & ~n19878;
  assign n20215 = ~n16360 & ~n19882;
  assign n20216 = ~n16353 & n19885;
  assign n20217 = ~n16230 & n19887;
  assign n20218 = ~n15618 & ~n16288;
  assign n20219 = ~n20216 & ~n20217;
  assign n20220 = ~n20218 & n20219;
  assign n20221 = n19884 & ~n20220;
  assign n20222 = ~n18628 & ~n20221;
  assign n20223 = ~n19933 & ~n20014;
  assign n20224 = ~n19902 & ~n20223;
  assign n20225 = n16295 & ~n19914;
  assign n20226 = ~n16295 & n19914;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = n20224 & ~n20227;
  assign n20229 = ~n19915 & ~n19921;
  assign n20230 = ~n20224 & ~n20229;
  assign n20231 = ~n20228 & ~n20230;
  assign n20232 = n20029 & ~n20231;
  assign n20233 = ~n20214 & ~n20215;
  assign n20234 = n20222 & n20233;
  assign n3650 = n20232 | ~n20234;
  assign n20236 = ~n16991 & n20036;
  assign n20237 = P3_REG3_REG_22_ & ~P3_STATE_REG;
  assign n20238 = ~n17057 & n19885;
  assign n20239 = ~n16940 & n19887;
  assign n20240 = ~n15618 & ~n16991;
  assign n20241 = ~n20238 & ~n20239;
  assign n20242 = ~n20240 & n20241;
  assign n20243 = n19884 & ~n20242;
  assign n20244 = ~n20237 & ~n20243;
  assign n20245 = n17059 & n20048;
  assign n20246 = n16998 & ~n20073;
  assign n20247 = ~n16998 & n20073;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = n20125 & ~n20248;
  assign n20250 = ~n20125 & n20248;
  assign n20251 = ~n20249 & ~n20250;
  assign n20252 = n20029 & ~n20251;
  assign n20253 = ~n20236 & n20244;
  assign n20254 = ~n20245 & n20253;
  assign n3655 = n20252 | ~n20254;
  assign n20256 = ~n16418 & ~n19878;
  assign n20257 = ~n16498 & ~n19882;
  assign n20258 = ~n16491 & n19885;
  assign n20259 = ~n16353 & n19887;
  assign n20260 = ~n15618 & ~n16418;
  assign n20261 = ~n20258 & ~n20259;
  assign n20262 = ~n20260 & n20261;
  assign n20263 = n19884 & ~n20262;
  assign n20264 = ~n18562 & ~n20263;
  assign n20265 = n19911 & ~n19918;
  assign n20266 = ~n19915 & ~n20224;
  assign n20267 = ~n19921 & ~n20266;
  assign n20268 = ~n19919 & n20267;
  assign n20269 = n20265 & ~n20268;
  assign n20270 = n16425 & ~n19909;
  assign n20271 = ~n16425 & n19909;
  assign n20272 = ~n20270 & ~n20271;
  assign n20273 = ~n19919 & n20272;
  assign n20274 = ~n19906 & ~n20267;
  assign n20275 = n20273 & ~n20274;
  assign n20276 = ~n20269 & ~n20275;
  assign n20277 = n20029 & n20276;
  assign n20278 = ~n20256 & ~n20257;
  assign n20279 = n20264 & n20278;
  assign n3660 = n20277 | ~n20279;
  assign n20281 = ~n16872 & n20036;
  assign n20282 = P3_REG3_REG_20_ & ~P3_STATE_REG;
  assign n20283 = ~n16940 & n19885;
  assign n20284 = ~n16814 & n19887;
  assign n20285 = ~n15618 & ~n16872;
  assign n20286 = ~n20283 & ~n20284;
  assign n20287 = ~n20285 & n20286;
  assign n20288 = n19884 & ~n20287;
  assign n20289 = ~n20282 & ~n20288;
  assign n20290 = n16942 & n20048;
  assign n20291 = n16879 & ~n20083;
  assign n20292 = ~n16879 & n20083;
  assign n20293 = ~n20291 & ~n20292;
  assign n20294 = ~n20095 & ~n20123;
  assign n20295 = ~n20089 & ~n20294;
  assign n20296 = ~n20293 & n20295;
  assign n20297 = ~n20084 & ~n20090;
  assign n20298 = ~n20295 & ~n20297;
  assign n20299 = ~n20296 & ~n20298;
  assign n20300 = n20029 & ~n20299;
  assign n20301 = ~n20281 & n20289;
  assign n20302 = ~n20290 & n20301;
  assign n3665 = n20300 | ~n20302;
  assign n20304 = ~n15618 & n19884;
  assign n20305 = n19878 & ~n20304;
  assign n20306 = P3_REG3_REG_0_ & ~n20305;
  assign n20307 = ~n19898 & n19982;
  assign n20308 = n19898 & ~n19982;
  assign n20309 = ~n20307 & ~n20308;
  assign n20310 = n15685 & ~n20309;
  assign n20311 = ~n15685 & n20309;
  assign n20312 = ~n20310 & ~n20311;
  assign n20313 = n20029 & ~n20312;
  assign n20314 = ~n15662 & ~n19882;
  assign n20315 = ~n15701 & n19884;
  assign n20316 = n19885 & n20315;
  assign n20317 = ~n20314 & ~n20316;
  assign n20318 = ~n18974 & ~n20313;
  assign n20319 = n20317 & n20318;
  assign n3670 = n20306 | ~n20319;
  assign n20321 = ~n16161 & ~n19878;
  assign n20322 = ~n16237 & ~n19882;
  assign n20323 = ~n16230 & n19885;
  assign n20324 = ~n16104 & n19887;
  assign n20325 = ~n15618 & ~n16161;
  assign n20326 = ~n20323 & ~n20324;
  assign n20327 = ~n20325 & n20326;
  assign n20328 = n19884 & ~n20327;
  assign n20329 = ~n18688 & ~n20328;
  assign n20330 = n16168 & ~n20010;
  assign n20331 = ~n16168 & n20010;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = n20006 & ~n20332;
  assign n20334 = ~n20006 & n20332;
  assign n20335 = ~n20333 & ~n20334;
  assign n20336 = n20029 & ~n20335;
  assign n20337 = ~n20321 & ~n20322;
  assign n20338 = n20329 & n20337;
  assign n3675 = n20336 | ~n20338;
  assign n20340 = n15852 & ~n20000;
  assign n20341 = ~n15852 & n20000;
  assign n20342 = ~n20340 & ~n20341;
  assign n20343 = n19996 & ~n20342;
  assign n20344 = ~n19996 & n20342;
  assign n20345 = ~n20343 & ~n20344;
  assign n20346 = n20029 & ~n20345;
  assign n20347 = ~n15919 & ~n19882;
  assign n20348 = ~n20346 & ~n20347;
  assign n20349 = ~n15845 & ~n19878;
  assign n20350 = ~n15912 & n19885;
  assign n20351 = ~n15793 & n19887;
  assign n20352 = ~n15618 & ~n15845;
  assign n20353 = ~n20350 & ~n20351;
  assign n20354 = ~n20352 & n20353;
  assign n20355 = n19884 & ~n20354;
  assign n20356 = ~n18844 & ~n20355;
  assign n20357 = n20348 & ~n20349;
  assign n3680 = ~n20356 | ~n20357;
  assign n20359 = ~n17111 & n20036;
  assign n20360 = P3_REG3_REG_24_ & ~P3_STATE_REG;
  assign n20361 = ~n17177 & n19885;
  assign n20362 = ~n17057 & n19887;
  assign n20363 = ~n15618 & ~n17111;
  assign n20364 = ~n20361 & ~n20362;
  assign n20365 = ~n20363 & n20364;
  assign n20366 = n19884 & ~n20365;
  assign n20367 = ~n20360 & ~n20366;
  assign n20368 = n17179 & n20048;
  assign n20369 = n17118 & ~n20064;
  assign n20370 = ~n17118 & n20064;
  assign n20371 = ~n20369 & ~n20370;
  assign n20372 = n20129 & ~n20371;
  assign n20373 = ~n20065 & ~n20132;
  assign n20374 = ~n20129 & ~n20373;
  assign n20375 = ~n20372 & ~n20374;
  assign n20376 = n20029 & ~n20375;
  assign n20377 = ~n20359 & n20367;
  assign n20378 = ~n20368 & n20377;
  assign n3685 = n20376 | ~n20378;
  assign n20380 = ~n16672 & ~n19878;
  assign n20381 = ~n16752 & ~n19882;
  assign n20382 = ~n16745 & n19885;
  assign n20383 = ~n16618 & n19887;
  assign n20384 = ~n15618 & ~n16672;
  assign n20385 = ~n20382 & ~n20383;
  assign n20386 = ~n20384 & n20385;
  assign n20387 = n19884 & ~n20386;
  assign n20388 = ~n18432 & ~n20387;
  assign n20389 = ~n16679 & ~n20109;
  assign n20390 = n20115 & ~n20389;
  assign n20391 = ~n20105 & n20119;
  assign n20392 = n20390 & ~n20391;
  assign n20393 = n16679 & ~n20109;
  assign n20394 = ~n16679 & n20109;
  assign n20395 = ~n20393 & ~n20394;
  assign n20396 = ~n20105 & n20395;
  assign n20397 = ~n20113 & ~n20119;
  assign n20398 = n20396 & ~n20397;
  assign n20399 = ~n20392 & ~n20398;
  assign n20400 = n20029 & n20399;
  assign n20401 = ~n20380 & ~n20381;
  assign n20402 = n20388 & n20401;
  assign n3690 = n20400 | ~n20402;
  assign n20404 = ~n15905 & ~n19878;
  assign n20405 = ~n15985 & ~n19882;
  assign n20406 = ~n15978 & n19885;
  assign n20407 = ~n15852 & n19887;
  assign n20408 = ~n15618 & ~n15905;
  assign n20409 = ~n20406 & ~n20407;
  assign n20410 = ~n20408 & n20409;
  assign n20411 = n19884 & ~n20410;
  assign n20412 = ~n18815 & ~n20411;
  assign n20413 = n15912 & ~n19948;
  assign n20414 = ~n15912 & n19948;
  assign n20415 = ~n20413 & ~n20414;
  assign n20416 = n20004 & ~n20415;
  assign n20417 = ~n20004 & n20415;
  assign n20418 = ~n20416 & ~n20417;
  assign n20419 = n20029 & ~n20418;
  assign n20420 = ~n20404 & ~n20405;
  assign n20421 = n20412 & n20420;
  assign n3695 = n20419 | ~n20421;
  assign n20423 = ~n16611 & ~n19878;
  assign n20424 = ~n16686 & ~n19882;
  assign n20425 = ~n16679 & n19885;
  assign n20426 = ~n16555 & n19887;
  assign n20427 = ~n15618 & ~n16611;
  assign n20428 = ~n20425 & ~n20426;
  assign n20429 = ~n20427 & n20428;
  assign n20430 = n19884 & ~n20429;
  assign n20431 = ~n18468 & ~n20430;
  assign n20432 = n16618 & ~n20104;
  assign n20433 = ~n16618 & n20104;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = n20119 & ~n20434;
  assign n20436 = ~n20105 & ~n20113;
  assign n20437 = ~n20119 & ~n20436;
  assign n20438 = ~n20435 & ~n20437;
  assign n20439 = n20029 & ~n20438;
  assign n20440 = ~n20423 & ~n20424;
  assign n20441 = n20431 & n20440;
  assign n3700 = n20439 | ~n20441;
  assign n20443 = ~n17170 & n20036;
  assign n20444 = P3_REG3_REG_25_ & ~P3_STATE_REG;
  assign n20445 = ~n17240 & n19885;
  assign n20446 = ~n17118 & n19887;
  assign n20447 = ~n15618 & ~n17170;
  assign n20448 = ~n20445 & ~n20446;
  assign n20449 = ~n20447 & n20448;
  assign n20450 = n19884 & ~n20449;
  assign n20451 = ~n20444 & ~n20450;
  assign n20452 = n17242 & n20048;
  assign n20453 = ~n20130 & ~n20132;
  assign n20454 = n17177 & ~n20056;
  assign n20455 = ~n17177 & n20056;
  assign n20456 = ~n20454 & ~n20455;
  assign n20457 = n20453 & ~n20456;
  assign n20458 = ~n20057 & ~n20133;
  assign n20459 = ~n20453 & ~n20458;
  assign n20460 = ~n20457 & ~n20459;
  assign n20461 = n20029 & ~n20460;
  assign n20462 = ~n20443 & n20451;
  assign n20463 = ~n20452 & n20462;
  assign n3705 = n20461 | ~n20463;
  assign n20465 = ~n16346 & ~n19878;
  assign n20466 = ~n16432 & ~n19882;
  assign n20467 = ~n16425 & n19885;
  assign n20468 = ~n16295 & n19887;
  assign n20469 = ~n15618 & ~n16346;
  assign n20470 = ~n20467 & ~n20468;
  assign n20471 = ~n20469 & n20470;
  assign n20472 = n19884 & ~n20471;
  assign n20473 = ~n18592 & ~n20472;
  assign n20474 = n16353 & ~n19905;
  assign n20475 = ~n16353 & n19905;
  assign n20476 = ~n20474 & ~n20475;
  assign n20477 = n20267 & ~n20476;
  assign n20478 = ~n19906 & ~n19919;
  assign n20479 = ~n20267 & ~n20478;
  assign n20480 = ~n20477 & ~n20479;
  assign n20481 = n20029 & ~n20480;
  assign n20482 = ~n20465 & ~n20466;
  assign n20483 = n20473 & n20482;
  assign n3710 = n20481 | ~n20483;
  assign n20485 = ~n16933 & n20036;
  assign n20486 = P3_REG3_REG_21_ & ~P3_STATE_REG;
  assign n20487 = ~n16998 & n19885;
  assign n20488 = ~n16879 & n19887;
  assign n20489 = ~n15618 & ~n16933;
  assign n20490 = ~n20487 & ~n20488;
  assign n20491 = ~n20489 & n20490;
  assign n20492 = n19884 & ~n20491;
  assign n20493 = ~n20486 & ~n20492;
  assign n20494 = n17000 & n20048;
  assign n20495 = ~n20080 & n20091;
  assign n20496 = ~n20084 & n20295;
  assign n20497 = n20495 & ~n20496;
  assign n20498 = n16940 & ~n20078;
  assign n20499 = ~n16940 & n20078;
  assign n20500 = ~n20498 & ~n20499;
  assign n20501 = ~n20084 & n20500;
  assign n20502 = ~n20090 & ~n20295;
  assign n20503 = n20501 & ~n20502;
  assign n20504 = ~n20497 & ~n20503;
  assign n20505 = n20029 & n20504;
  assign n20506 = ~n20485 & n20493;
  assign n20507 = ~n20494 & n20506;
  assign n3715 = n20505 | ~n20507;
  assign n20509 = ~n19983 & ~n19991;
  assign n20510 = n15701 & ~n19986;
  assign n20511 = ~n15701 & n19986;
  assign n20512 = ~n20510 & ~n20511;
  assign n20513 = n20509 & ~n20512;
  assign n20514 = ~n20509 & n20512;
  assign n20515 = ~n20513 & ~n20514;
  assign n20516 = n20029 & ~n20515;
  assign n20517 = ~n15746 & ~n19882;
  assign n20518 = ~n20516 & ~n20517;
  assign n20519 = P3_REG3_REG_1_ & ~n19878;
  assign n20520 = ~n15739 & n19885;
  assign n20521 = ~n15685 & n19887;
  assign n20522 = P3_REG3_REG_1_ & ~n15618;
  assign n20523 = ~n20520 & ~n20521;
  assign n20524 = ~n20522 & n20523;
  assign n20525 = n19884 & ~n20524;
  assign n20526 = ~n18950 & ~n20525;
  assign n20527 = n20518 & ~n20519;
  assign n3720 = ~n20526 | ~n20527;
  assign n20529 = ~n16097 & ~n19878;
  assign n20530 = ~n16175 & ~n19882;
  assign n20531 = ~n16168 & n19885;
  assign n20532 = ~n16037 & n19887;
  assign n20533 = ~n15618 & ~n16097;
  assign n20534 = ~n20531 & ~n20532;
  assign n20535 = ~n20533 & n20534;
  assign n20536 = n19884 & ~n20535;
  assign n20537 = ~n18723 & ~n20536;
  assign n20538 = n19964 & ~n20004;
  assign n20539 = n19955 & ~n20538;
  assign n20540 = n16104 & ~n19958;
  assign n20541 = ~n16104 & n19958;
  assign n20542 = ~n20540 & ~n20541;
  assign n20543 = n20539 & ~n20542;
  assign n20544 = ~n20539 & n20542;
  assign n20545 = ~n20543 & ~n20544;
  assign n20546 = n20029 & ~n20545;
  assign n20547 = ~n20529 & ~n20530;
  assign n20548 = n20537 & n20547;
  assign n3725 = n20546 | ~n20548;
  assign n20550 = ~n17351 & n20036;
  assign n20551 = P3_REG3_REG_28_ & ~P3_STATE_REG;
  assign n20552 = ~n17414 & n19885;
  assign n20553 = ~n17297 & n19887;
  assign n20554 = ~n15618 & ~n17351;
  assign n20555 = ~n20552 & ~n20553;
  assign n20556 = ~n20554 & n20555;
  assign n20557 = n19884 & ~n20556;
  assign n20558 = ~n20551 & ~n20557;
  assign n20559 = n17416 & n20048;
  assign n20560 = n17360 & n19898;
  assign n20561 = ~n17360 & ~n19898;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = n17297 & n20562;
  assign n20564 = ~n20053 & n20134;
  assign n20565 = ~n20563 & ~n20564;
  assign n20566 = ~n20053 & ~n20059;
  assign n20567 = ~n20058 & n20566;
  assign n20568 = n20565 & ~n20567;
  assign n20569 = ~n17297 & ~n20562;
  assign n20570 = ~n20568 & ~n20569;
  assign n20571 = n20058 & ~n20065;
  assign n20572 = ~n20057 & ~n20065;
  assign n20573 = ~n20052 & n20572;
  assign n20574 = ~n20571 & ~n20573;
  assign n20575 = ~n20563 & ~n20574;
  assign n20576 = ~n20129 & n20575;
  assign n20577 = ~n17358 & n19898;
  assign n20578 = n17358 & ~n19898;
  assign n20579 = ~n20577 & ~n20578;
  assign n20580 = ~n17416 & ~n20579;
  assign n20581 = n17416 & n20579;
  assign n20582 = ~n20580 & ~n20581;
  assign n20583 = n20570 & ~n20576;
  assign n20584 = ~n20582 & n20583;
  assign n20585 = ~n20564 & ~n20567;
  assign n20586 = ~n20569 & ~n20585;
  assign n20587 = ~n20129 & ~n20574;
  assign n20588 = n20586 & ~n20587;
  assign n20589 = ~n20563 & ~n20588;
  assign n20590 = n20582 & n20589;
  assign n20591 = ~n20584 & ~n20590;
  assign n20592 = n20029 & ~n20591;
  assign n20593 = ~n20550 & n20558;
  assign n20594 = ~n20559 & n20593;
  assign n3730 = n20592 | ~n20594;
  assign n20596 = ~n16807 & ~n19878;
  assign n20597 = ~n16879 & n19885;
  assign n20598 = ~n16745 & n19887;
  assign n20599 = ~n15618 & ~n16807;
  assign n20600 = ~n20597 & ~n20598;
  assign n20601 = ~n20599 & n20600;
  assign n20602 = n19884 & ~n20601;
  assign n20603 = ~n18369 & ~n20602;
  assign n20604 = ~n16883 & ~n19882;
  assign n20605 = n16814 & ~n20088;
  assign n20606 = ~n16814 & n20088;
  assign n20607 = ~n20605 & ~n20606;
  assign n20608 = n20123 & ~n20607;
  assign n20609 = ~n20089 & ~n20095;
  assign n20610 = ~n20123 & ~n20609;
  assign n20611 = ~n20608 & ~n20610;
  assign n20612 = n20029 & ~n20611;
  assign n20613 = ~n20596 & n20603;
  assign n20614 = ~n20604 & n20613;
  assign n3735 = n20612 | ~n20614;
  assign n20616 = ~n15793 & ~n19973;
  assign n20617 = n19979 & ~n20616;
  assign n20618 = ~n19969 & n19994;
  assign n20619 = n20617 & ~n20618;
  assign n20620 = n15793 & ~n19973;
  assign n20621 = ~n15793 & n19973;
  assign n20622 = ~n20620 & ~n20621;
  assign n20623 = ~n19969 & n20622;
  assign n20624 = ~n19977 & ~n19994;
  assign n20625 = n20623 & ~n20624;
  assign n20626 = ~n20619 & ~n20625;
  assign n20627 = n20029 & n20626;
  assign n20628 = ~n15859 & ~n19882;
  assign n20629 = ~n20627 & ~n20628;
  assign n20630 = ~P3_REG3_REG_3_ & ~n19878;
  assign n20631 = ~n15852 & n19885;
  assign n20632 = ~n15739 & n19887;
  assign n20633 = ~P3_REG3_REG_3_ & ~n15618;
  assign n20634 = ~n20631 & ~n20632;
  assign n20635 = ~n20633 & n20634;
  assign n20636 = n19884 & ~n20635;
  assign n20637 = ~n18874 & ~n20636;
  assign n20638 = n20629 & ~n20630;
  assign n3740 = ~n20637 | ~n20638;
  assign n20640 = ~n16223 & ~n19878;
  assign n20641 = ~n16302 & ~n19882;
  assign n20642 = ~n16295 & n19885;
  assign n20643 = ~n16168 & n19887;
  assign n20644 = ~n15618 & ~n16223;
  assign n20645 = ~n20642 & ~n20643;
  assign n20646 = ~n20644 & n20645;
  assign n20647 = n19884 & ~n20646;
  assign n20648 = ~n18658 & ~n20647;
  assign n20649 = n16230 & ~n19901;
  assign n20650 = ~n16230 & n19901;
  assign n20651 = ~n20649 & ~n20650;
  assign n20652 = n20014 & ~n20651;
  assign n20653 = ~n20014 & n20651;
  assign n20654 = ~n20652 & ~n20653;
  assign n20655 = n20029 & ~n20654;
  assign n20656 = ~n20640 & ~n20641;
  assign n20657 = n20648 & n20656;
  assign n3745 = n20655 | ~n20657;
  assign n20659 = ~n17050 & n20036;
  assign n20660 = P3_REG3_REG_23_ & ~P3_STATE_REG;
  assign n20661 = ~n17118 & n19885;
  assign n20662 = ~n16998 & n19887;
  assign n20663 = ~n15618 & ~n17050;
  assign n20664 = ~n20661 & ~n20662;
  assign n20665 = ~n20663 & n20664;
  assign n20666 = n19884 & ~n20665;
  assign n20667 = ~n20660 & ~n20666;
  assign n20668 = n17120 & n20048;
  assign n20669 = n17057 & ~n20068;
  assign n20670 = ~n17057 & n20068;
  assign n20671 = ~n20669 & ~n20670;
  assign n20672 = n20127 & ~n20671;
  assign n20673 = ~n20127 & n20671;
  assign n20674 = ~n20672 & ~n20673;
  assign n20675 = n20029 & ~n20674;
  assign n20676 = ~n20659 & n20667;
  assign n20677 = ~n20668 & n20676;
  assign n3750 = n20675 | ~n20677;
  assign n20679 = ~n16484 & ~n19878;
  assign n20680 = ~n16562 & ~n19882;
  assign n20681 = ~n16555 & n19885;
  assign n20682 = ~n16425 & n19887;
  assign n20683 = ~n15618 & ~n16484;
  assign n20684 = ~n20681 & ~n20682;
  assign n20685 = ~n20683 & n20684;
  assign n20686 = n19884 & ~n20685;
  assign n20687 = ~n18532 & ~n20686;
  assign n20688 = n19934 & ~n20014;
  assign n20689 = n19925 & ~n20688;
  assign n20690 = n16491 & ~n19928;
  assign n20691 = ~n16491 & n19928;
  assign n20692 = ~n20690 & ~n20691;
  assign n20693 = n20689 & ~n20692;
  assign n20694 = ~n20689 & n20692;
  assign n20695 = ~n20693 & ~n20694;
  assign n20696 = n20029 & ~n20695;
  assign n20697 = ~n20679 & ~n20680;
  assign n20698 = n20687 & n20697;
  assign n3755 = n20696 | ~n20698;
  assign n20700 = ~n17293 & n20036;
  assign n20701 = P3_REG3_REG_27_ & ~P3_STATE_REG;
  assign n20702 = ~n17358 & n19885;
  assign n20703 = ~n17240 & n19887;
  assign n20704 = ~n15618 & ~n17293;
  assign n20705 = ~n20702 & ~n20703;
  assign n20706 = ~n20704 & n20705;
  assign n20707 = n19884 & ~n20706;
  assign n20708 = ~n20701 & ~n20707;
  assign n20709 = n17360 & n20048;
  assign n20710 = ~n20585 & ~n20587;
  assign n20711 = n17297 & ~n20562;
  assign n20712 = ~n17297 & n20562;
  assign n20713 = ~n20711 & ~n20712;
  assign n20714 = n20710 & ~n20713;
  assign n20715 = ~n20710 & n20713;
  assign n20716 = ~n20714 & ~n20715;
  assign n20717 = n20029 & ~n20716;
  assign n20718 = ~n20700 & n20708;
  assign n20719 = ~n20709 & n20718;
  assign n3760 = n20717 | ~n20719;
  assign n20721 = ~n16030 & ~n19878;
  assign n20722 = ~n16111 & ~n19882;
  assign n20723 = ~n16104 & n19885;
  assign n20724 = ~n15978 & n19887;
  assign n20725 = ~n15618 & ~n16030;
  assign n20726 = ~n20723 & ~n20724;
  assign n20727 = ~n20725 & n20726;
  assign n20728 = n19884 & ~n20727;
  assign n20729 = ~n18753 & ~n20728;
  assign n20730 = ~n16037 & ~n19938;
  assign n20731 = n19952 & ~n20730;
  assign n20732 = ~n19942 & n20166;
  assign n20733 = n20731 & ~n20732;
  assign n20734 = n16037 & ~n19938;
  assign n20735 = ~n16037 & n19938;
  assign n20736 = ~n20734 & ~n20735;
  assign n20737 = ~n19942 & n20736;
  assign n20738 = ~n19950 & ~n20166;
  assign n20739 = n20737 & ~n20738;
  assign n20740 = ~n20733 & ~n20739;
  assign n20741 = n20029 & n20740;
  assign n20742 = ~n20721 & ~n20722;
  assign n20743 = n20729 & n20742;
  assign n3765 = n20741 | ~n20743;
  assign n20745 = P3_STATE_REG & ~n18020;
  assign n20746 = n15504 & n18021;
  assign n3775 = ~n20745 | n20746;
  assign n1320 = ~P1_STATE_REG;
  assign n2545 = ~P2_STATE_REG;
  assign n3770 = ~P3_STATE_REG;
  always @ (posedge clock) begin
    P1_IR_REG_0_ <= n110;
    P1_IR_REG_1_ <= n115;
    P1_IR_REG_2_ <= n120;
    P1_IR_REG_3_ <= n125;
    P1_IR_REG_4_ <= n130;
    P1_IR_REG_5_ <= n135;
    P1_IR_REG_6_ <= n140;
    P1_IR_REG_7_ <= n145;
    P1_IR_REG_8_ <= n150;
    P1_IR_REG_9_ <= n155;
    P1_IR_REG_10_ <= n160;
    P1_IR_REG_11_ <= n165;
    P1_IR_REG_12_ <= n170;
    P1_IR_REG_13_ <= n175;
    P1_IR_REG_14_ <= n180;
    P1_IR_REG_15_ <= n185;
    P1_IR_REG_16_ <= n190;
    P1_IR_REG_17_ <= n195;
    P1_IR_REG_18_ <= n200;
    P1_IR_REG_19_ <= n205;
    P1_IR_REG_20_ <= n210;
    P1_IR_REG_21_ <= n215;
    P1_IR_REG_22_ <= n220;
    P1_IR_REG_23_ <= n225;
    P1_IR_REG_24_ <= n230;
    P1_IR_REG_25_ <= n235;
    P1_IR_REG_26_ <= n240;
    P1_IR_REG_27_ <= n245;
    P1_IR_REG_28_ <= n250;
    P1_IR_REG_29_ <= n255;
    P1_IR_REG_30_ <= n260;
    P1_IR_REG_31_ <= n265;
    P1_D_REG_0_ <= n270;
    P1_D_REG_1_ <= n275;
    P1_D_REG_2_ <= n280;
    P1_D_REG_3_ <= n285;
    P1_D_REG_4_ <= n290;
    P1_D_REG_5_ <= n295;
    P1_D_REG_6_ <= n300;
    P1_D_REG_7_ <= n305;
    P1_D_REG_8_ <= n310;
    P1_D_REG_9_ <= n315;
    P1_D_REG_10_ <= n320;
    P1_D_REG_11_ <= n325;
    P1_D_REG_12_ <= n330;
    P1_D_REG_13_ <= n335;
    P1_D_REG_14_ <= n340;
    P1_D_REG_15_ <= n345;
    P1_D_REG_16_ <= n350;
    P1_D_REG_17_ <= n355;
    P1_D_REG_18_ <= n360;
    P1_D_REG_19_ <= n365;
    P1_D_REG_20_ <= n370;
    P1_D_REG_21_ <= n375;
    P1_D_REG_22_ <= n380;
    P1_D_REG_23_ <= n385;
    P1_D_REG_24_ <= n390;
    P1_D_REG_25_ <= n395;
    P1_D_REG_26_ <= n400;
    P1_D_REG_27_ <= n405;
    P1_D_REG_28_ <= n410;
    P1_D_REG_29_ <= n415;
    P1_D_REG_30_ <= n420;
    P1_D_REG_31_ <= n425;
    P1_REG0_REG_0_ <= n430;
    P1_REG0_REG_1_ <= n435;
    P1_REG0_REG_2_ <= n440;
    P1_REG0_REG_3_ <= n445;
    P1_REG0_REG_4_ <= n450;
    P1_REG0_REG_5_ <= n455;
    P1_REG0_REG_6_ <= n460;
    P1_REG0_REG_7_ <= n465;
    P1_REG0_REG_8_ <= n470;
    P1_REG0_REG_9_ <= n475;
    P1_REG0_REG_10_ <= n480;
    P1_REG0_REG_11_ <= n485;
    P1_REG0_REG_12_ <= n490;
    P1_REG0_REG_13_ <= n495;
    P1_REG0_REG_14_ <= n500;
    P1_REG0_REG_15_ <= n505;
    P1_REG0_REG_16_ <= n510;
    P1_REG0_REG_17_ <= n515;
    P1_REG0_REG_18_ <= n520;
    P1_REG0_REG_19_ <= n525;
    P1_REG0_REG_20_ <= n530;
    P1_REG0_REG_21_ <= n535;
    P1_REG0_REG_22_ <= n540;
    P1_REG0_REG_23_ <= n545;
    P1_REG0_REG_24_ <= n550;
    P1_REG0_REG_25_ <= n555;
    P1_REG0_REG_26_ <= n560;
    P1_REG0_REG_27_ <= n565;
    P1_REG0_REG_28_ <= n570;
    P1_REG0_REG_29_ <= n575;
    P1_REG0_REG_30_ <= n580;
    P1_REG0_REG_31_ <= n585;
    P1_REG1_REG_0_ <= n590;
    P1_REG1_REG_1_ <= n595;
    P1_REG1_REG_2_ <= n600;
    P1_REG1_REG_3_ <= n605;
    P1_REG1_REG_4_ <= n610;
    P1_REG1_REG_5_ <= n615;
    P1_REG1_REG_6_ <= n620;
    P1_REG1_REG_7_ <= n625;
    P1_REG1_REG_8_ <= n630;
    P1_REG1_REG_9_ <= n635;
    P1_REG1_REG_10_ <= n640;
    P1_REG1_REG_11_ <= n645;
    P1_REG1_REG_12_ <= n650;
    P1_REG1_REG_13_ <= n655;
    P1_REG1_REG_14_ <= n660;
    P1_REG1_REG_15_ <= n665;
    P1_REG1_REG_16_ <= n670;
    P1_REG1_REG_17_ <= n675;
    P1_REG1_REG_18_ <= n680;
    P1_REG1_REG_19_ <= n685;
    P1_REG1_REG_20_ <= n690;
    P1_REG1_REG_21_ <= n695;
    P1_REG1_REG_22_ <= n700;
    P1_REG1_REG_23_ <= n705;
    P1_REG1_REG_24_ <= n710;
    P1_REG1_REG_25_ <= n715;
    P1_REG1_REG_26_ <= n720;
    P1_REG1_REG_27_ <= n725;
    P1_REG1_REG_28_ <= n730;
    P1_REG1_REG_29_ <= n735;
    P1_REG1_REG_30_ <= n740;
    P1_REG1_REG_31_ <= n745;
    P1_REG2_REG_0_ <= n750;
    P1_REG2_REG_1_ <= n755;
    P1_REG2_REG_2_ <= n760;
    P1_REG2_REG_3_ <= n765;
    P1_REG2_REG_4_ <= n770;
    P1_REG2_REG_5_ <= n775;
    P1_REG2_REG_6_ <= n780;
    P1_REG2_REG_7_ <= n785;
    P1_REG2_REG_8_ <= n790;
    P1_REG2_REG_9_ <= n795;
    P1_REG2_REG_10_ <= n800;
    P1_REG2_REG_11_ <= n805;
    P1_REG2_REG_12_ <= n810;
    P1_REG2_REG_13_ <= n815;
    P1_REG2_REG_14_ <= n820;
    P1_REG2_REG_15_ <= n825;
    P1_REG2_REG_16_ <= n830;
    P1_REG2_REG_17_ <= n835;
    P1_REG2_REG_18_ <= n840;
    P1_REG2_REG_19_ <= n845;
    P1_REG2_REG_20_ <= n850;
    P1_REG2_REG_21_ <= n855;
    P1_REG2_REG_22_ <= n860;
    P1_REG2_REG_23_ <= n865;
    P1_REG2_REG_24_ <= n870;
    P1_REG2_REG_25_ <= n875;
    P1_REG2_REG_26_ <= n880;
    P1_REG2_REG_27_ <= n885;
    P1_REG2_REG_28_ <= n890;
    P1_REG2_REG_29_ <= n895;
    P1_REG2_REG_30_ <= n900;
    P1_REG2_REG_31_ <= n905;
    P1_ADDR_REG_19_ <= n910;
    P1_ADDR_REG_18_ <= n915;
    P1_ADDR_REG_17_ <= n920;
    P1_ADDR_REG_16_ <= n925;
    P1_ADDR_REG_15_ <= n930;
    P1_ADDR_REG_14_ <= n935;
    P1_ADDR_REG_13_ <= n940;
    P1_ADDR_REG_12_ <= n945;
    P1_ADDR_REG_11_ <= n950;
    P1_ADDR_REG_10_ <= n955;
    P1_ADDR_REG_9_ <= n960;
    P1_ADDR_REG_8_ <= n965;
    P1_ADDR_REG_7_ <= n970;
    P1_ADDR_REG_6_ <= n975;
    P1_ADDR_REG_5_ <= n980;
    P1_ADDR_REG_4_ <= n985;
    P1_ADDR_REG_3_ <= n990;
    P1_ADDR_REG_2_ <= n995;
    P1_ADDR_REG_1_ <= n1000;
    P1_ADDR_REG_0_ <= n1005;
    P1_DATAO_REG_0_ <= n1010;
    P1_DATAO_REG_1_ <= n1015;
    P1_DATAO_REG_2_ <= n1020;
    P1_DATAO_REG_3_ <= n1025;
    P1_DATAO_REG_4_ <= n1030;
    P1_DATAO_REG_5_ <= n1035;
    P1_DATAO_REG_6_ <= n1040;
    P1_DATAO_REG_7_ <= n1045;
    P1_DATAO_REG_8_ <= n1050;
    P1_DATAO_REG_9_ <= n1055;
    P1_DATAO_REG_10_ <= n1060;
    P1_DATAO_REG_11_ <= n1065;
    P1_DATAO_REG_12_ <= n1070;
    P1_DATAO_REG_13_ <= n1075;
    P1_DATAO_REG_14_ <= n1080;
    P1_DATAO_REG_15_ <= n1085;
    P1_DATAO_REG_16_ <= n1090;
    P1_DATAO_REG_17_ <= n1095;
    P1_DATAO_REG_18_ <= n1100;
    P1_DATAO_REG_19_ <= n1105;
    P1_DATAO_REG_20_ <= n1110;
    P1_DATAO_REG_21_ <= n1115;
    P1_DATAO_REG_22_ <= n1120;
    P1_DATAO_REG_23_ <= n1125;
    P1_DATAO_REG_24_ <= n1130;
    P1_DATAO_REG_25_ <= n1135;
    P1_DATAO_REG_26_ <= n1140;
    P1_DATAO_REG_27_ <= n1145;
    P1_DATAO_REG_28_ <= n1150;
    P1_DATAO_REG_29_ <= n1155;
    P1_DATAO_REG_30_ <= n1160;
    P1_DATAO_REG_31_ <= n1165;
    P1_B_REG <= n1170;
    P1_REG3_REG_15_ <= n1175;
    P1_REG3_REG_26_ <= n1180;
    P1_REG3_REG_6_ <= n1185;
    P1_REG3_REG_18_ <= n1190;
    P1_REG3_REG_2_ <= n1195;
    P1_REG3_REG_11_ <= n1200;
    P1_REG3_REG_22_ <= n1205;
    P1_REG3_REG_13_ <= n1210;
    P1_REG3_REG_20_ <= n1215;
    P1_REG3_REG_0_ <= n1220;
    P1_REG3_REG_9_ <= n1225;
    P1_REG3_REG_4_ <= n1230;
    P1_REG3_REG_24_ <= n1235;
    P1_REG3_REG_17_ <= n1240;
    P1_REG3_REG_5_ <= n1245;
    P1_REG3_REG_16_ <= n1250;
    P1_REG3_REG_25_ <= n1255;
    P1_REG3_REG_12_ <= n1260;
    P1_REG3_REG_21_ <= n1265;
    P1_REG3_REG_1_ <= n1270;
    P1_REG3_REG_8_ <= n1275;
    P1_REG3_REG_28_ <= n1280;
    P1_REG3_REG_19_ <= n1285;
    P1_REG3_REG_3_ <= n1290;
    P1_REG3_REG_10_ <= n1295;
    P1_REG3_REG_23_ <= n1300;
    P1_REG3_REG_14_ <= n1305;
    P1_REG3_REG_27_ <= n1310;
    P1_REG3_REG_7_ <= n1315;
    P1_STATE_REG <= n1320;
    P1_RD_REG <= n1325;
    P1_WR_REG <= n1330;
    P2_IR_REG_0_ <= n1335;
    P2_IR_REG_1_ <= n1340;
    P2_IR_REG_2_ <= n1345;
    P2_IR_REG_3_ <= n1350;
    P2_IR_REG_4_ <= n1355;
    P2_IR_REG_5_ <= n1360;
    P2_IR_REG_6_ <= n1365;
    P2_IR_REG_7_ <= n1370;
    P2_IR_REG_8_ <= n1375;
    P2_IR_REG_9_ <= n1380;
    P2_IR_REG_10_ <= n1385;
    P2_IR_REG_11_ <= n1390;
    P2_IR_REG_12_ <= n1395;
    P2_IR_REG_13_ <= n1400;
    P2_IR_REG_14_ <= n1405;
    P2_IR_REG_15_ <= n1410;
    P2_IR_REG_16_ <= n1415;
    P2_IR_REG_17_ <= n1420;
    P2_IR_REG_18_ <= n1425;
    P2_IR_REG_19_ <= n1430;
    P2_IR_REG_20_ <= n1435;
    P2_IR_REG_21_ <= n1440;
    P2_IR_REG_22_ <= n1445;
    P2_IR_REG_23_ <= n1450;
    P2_IR_REG_24_ <= n1455;
    P2_IR_REG_25_ <= n1460;
    P2_IR_REG_26_ <= n1465;
    P2_IR_REG_27_ <= n1470;
    P2_IR_REG_28_ <= n1475;
    P2_IR_REG_29_ <= n1480;
    P2_IR_REG_30_ <= n1485;
    P2_IR_REG_31_ <= n1490;
    P2_D_REG_0_ <= n1495;
    P2_D_REG_1_ <= n1500;
    P2_D_REG_2_ <= n1505;
    P2_D_REG_3_ <= n1510;
    P2_D_REG_4_ <= n1515;
    P2_D_REG_5_ <= n1520;
    P2_D_REG_6_ <= n1525;
    P2_D_REG_7_ <= n1530;
    P2_D_REG_8_ <= n1535;
    P2_D_REG_9_ <= n1540;
    P2_D_REG_10_ <= n1545;
    P2_D_REG_11_ <= n1550;
    P2_D_REG_12_ <= n1555;
    P2_D_REG_13_ <= n1560;
    P2_D_REG_14_ <= n1565;
    P2_D_REG_15_ <= n1570;
    P2_D_REG_16_ <= n1575;
    P2_D_REG_17_ <= n1580;
    P2_D_REG_18_ <= n1585;
    P2_D_REG_19_ <= n1590;
    P2_D_REG_20_ <= n1595;
    P2_D_REG_21_ <= n1600;
    P2_D_REG_22_ <= n1605;
    P2_D_REG_23_ <= n1610;
    P2_D_REG_24_ <= n1615;
    P2_D_REG_25_ <= n1620;
    P2_D_REG_26_ <= n1625;
    P2_D_REG_27_ <= n1630;
    P2_D_REG_28_ <= n1635;
    P2_D_REG_29_ <= n1640;
    P2_D_REG_30_ <= n1645;
    P2_D_REG_31_ <= n1650;
    P2_REG0_REG_0_ <= n1655;
    P2_REG0_REG_1_ <= n1660;
    P2_REG0_REG_2_ <= n1665;
    P2_REG0_REG_3_ <= n1670;
    P2_REG0_REG_4_ <= n1675;
    P2_REG0_REG_5_ <= n1680;
    P2_REG0_REG_6_ <= n1685;
    P2_REG0_REG_7_ <= n1690;
    P2_REG0_REG_8_ <= n1695;
    P2_REG0_REG_9_ <= n1700;
    P2_REG0_REG_10_ <= n1705;
    P2_REG0_REG_11_ <= n1710;
    P2_REG0_REG_12_ <= n1715;
    P2_REG0_REG_13_ <= n1720;
    P2_REG0_REG_14_ <= n1725;
    P2_REG0_REG_15_ <= n1730;
    P2_REG0_REG_16_ <= n1735;
    P2_REG0_REG_17_ <= n1740;
    P2_REG0_REG_18_ <= n1745;
    P2_REG0_REG_19_ <= n1750;
    P2_REG0_REG_20_ <= n1755;
    P2_REG0_REG_21_ <= n1760;
    P2_REG0_REG_22_ <= n1765;
    P2_REG0_REG_23_ <= n1770;
    P2_REG0_REG_24_ <= n1775;
    P2_REG0_REG_25_ <= n1780;
    P2_REG0_REG_26_ <= n1785;
    P2_REG0_REG_27_ <= n1790;
    P2_REG0_REG_28_ <= n1795;
    P2_REG0_REG_29_ <= n1800;
    P2_REG0_REG_30_ <= n1805;
    P2_REG0_REG_31_ <= n1810;
    P2_REG1_REG_0_ <= n1815;
    P2_REG1_REG_1_ <= n1820;
    P2_REG1_REG_2_ <= n1825;
    P2_REG1_REG_3_ <= n1830;
    P2_REG1_REG_4_ <= n1835;
    P2_REG1_REG_5_ <= n1840;
    P2_REG1_REG_6_ <= n1845;
    P2_REG1_REG_7_ <= n1850;
    P2_REG1_REG_8_ <= n1855;
    P2_REG1_REG_9_ <= n1860;
    P2_REG1_REG_10_ <= n1865;
    P2_REG1_REG_11_ <= n1870;
    P2_REG1_REG_12_ <= n1875;
    P2_REG1_REG_13_ <= n1880;
    P2_REG1_REG_14_ <= n1885;
    P2_REG1_REG_15_ <= n1890;
    P2_REG1_REG_16_ <= n1895;
    P2_REG1_REG_17_ <= n1900;
    P2_REG1_REG_18_ <= n1905;
    P2_REG1_REG_19_ <= n1910;
    P2_REG1_REG_20_ <= n1915;
    P2_REG1_REG_21_ <= n1920;
    P2_REG1_REG_22_ <= n1925;
    P2_REG1_REG_23_ <= n1930;
    P2_REG1_REG_24_ <= n1935;
    P2_REG1_REG_25_ <= n1940;
    P2_REG1_REG_26_ <= n1945;
    P2_REG1_REG_27_ <= n1950;
    P2_REG1_REG_28_ <= n1955;
    P2_REG1_REG_29_ <= n1960;
    P2_REG1_REG_30_ <= n1965;
    P2_REG1_REG_31_ <= n1970;
    P2_REG2_REG_0_ <= n1975;
    P2_REG2_REG_1_ <= n1980;
    P2_REG2_REG_2_ <= n1985;
    P2_REG2_REG_3_ <= n1990;
    P2_REG2_REG_4_ <= n1995;
    P2_REG2_REG_5_ <= n2000;
    P2_REG2_REG_6_ <= n2005;
    P2_REG2_REG_7_ <= n2010;
    P2_REG2_REG_8_ <= n2015;
    P2_REG2_REG_9_ <= n2020;
    P2_REG2_REG_10_ <= n2025;
    P2_REG2_REG_11_ <= n2030;
    P2_REG2_REG_12_ <= n2035;
    P2_REG2_REG_13_ <= n2040;
    P2_REG2_REG_14_ <= n2045;
    P2_REG2_REG_15_ <= n2050;
    P2_REG2_REG_16_ <= n2055;
    P2_REG2_REG_17_ <= n2060;
    P2_REG2_REG_18_ <= n2065;
    P2_REG2_REG_19_ <= n2070;
    P2_REG2_REG_20_ <= n2075;
    P2_REG2_REG_21_ <= n2080;
    P2_REG2_REG_22_ <= n2085;
    P2_REG2_REG_23_ <= n2090;
    P2_REG2_REG_24_ <= n2095;
    P2_REG2_REG_25_ <= n2100;
    P2_REG2_REG_26_ <= n2105;
    P2_REG2_REG_27_ <= n2110;
    P2_REG2_REG_28_ <= n2115;
    P2_REG2_REG_29_ <= n2120;
    P2_REG2_REG_30_ <= n2125;
    P2_REG2_REG_31_ <= n2130;
    P2_ADDR_REG_19_ <= n2135;
    P2_ADDR_REG_18_ <= n2140;
    P2_ADDR_REG_17_ <= n2145;
    P2_ADDR_REG_16_ <= n2150;
    P2_ADDR_REG_15_ <= n2155;
    P2_ADDR_REG_14_ <= n2160;
    P2_ADDR_REG_13_ <= n2165;
    P2_ADDR_REG_12_ <= n2170;
    P2_ADDR_REG_11_ <= n2175;
    P2_ADDR_REG_10_ <= n2180;
    P2_ADDR_REG_9_ <= n2185;
    P2_ADDR_REG_8_ <= n2190;
    P2_ADDR_REG_7_ <= n2195;
    P2_ADDR_REG_6_ <= n2200;
    P2_ADDR_REG_5_ <= n2205;
    P2_ADDR_REG_4_ <= n2210;
    P2_ADDR_REG_3_ <= n2215;
    P2_ADDR_REG_2_ <= n2220;
    P2_ADDR_REG_1_ <= n2225;
    P2_ADDR_REG_0_ <= n2230;
    P2_DATAO_REG_0_ <= n2235;
    P2_DATAO_REG_1_ <= n2240;
    P2_DATAO_REG_2_ <= n2245;
    P2_DATAO_REG_3_ <= n2250;
    P2_DATAO_REG_4_ <= n2255;
    P2_DATAO_REG_5_ <= n2260;
    P2_DATAO_REG_6_ <= n2265;
    P2_DATAO_REG_7_ <= n2270;
    P2_DATAO_REG_8_ <= n2275;
    P2_DATAO_REG_9_ <= n2280;
    P2_DATAO_REG_10_ <= n2285;
    P2_DATAO_REG_11_ <= n2290;
    P2_DATAO_REG_12_ <= n2295;
    P2_DATAO_REG_13_ <= n2300;
    P2_DATAO_REG_14_ <= n2305;
    P2_DATAO_REG_15_ <= n2310;
    P2_DATAO_REG_16_ <= n2315;
    P2_DATAO_REG_17_ <= n2320;
    P2_DATAO_REG_18_ <= n2325;
    P2_DATAO_REG_19_ <= n2330;
    P2_DATAO_REG_20_ <= n2335;
    P2_DATAO_REG_21_ <= n2340;
    P2_DATAO_REG_22_ <= n2345;
    P2_DATAO_REG_23_ <= n2350;
    P2_DATAO_REG_24_ <= n2355;
    P2_DATAO_REG_25_ <= n2360;
    P2_DATAO_REG_26_ <= n2365;
    P2_DATAO_REG_27_ <= n2370;
    P2_DATAO_REG_28_ <= n2375;
    P2_DATAO_REG_29_ <= n2380;
    P2_DATAO_REG_30_ <= n2385;
    P2_DATAO_REG_31_ <= n2390;
    P2_B_REG <= n2395;
    P2_REG3_REG_15_ <= n2400;
    P2_REG3_REG_26_ <= n2405;
    P2_REG3_REG_6_ <= n2410;
    P2_REG3_REG_18_ <= n2415;
    P2_REG3_REG_2_ <= n2420;
    P2_REG3_REG_11_ <= n2425;
    P2_REG3_REG_22_ <= n2430;
    P2_REG3_REG_13_ <= n2435;
    P2_REG3_REG_20_ <= n2440;
    P2_REG3_REG_0_ <= n2445;
    P2_REG3_REG_9_ <= n2450;
    P2_REG3_REG_4_ <= n2455;
    P2_REG3_REG_24_ <= n2460;
    P2_REG3_REG_17_ <= n2465;
    P2_REG3_REG_5_ <= n2470;
    P2_REG3_REG_16_ <= n2475;
    P2_REG3_REG_25_ <= n2480;
    P2_REG3_REG_12_ <= n2485;
    P2_REG3_REG_21_ <= n2490;
    P2_REG3_REG_1_ <= n2495;
    P2_REG3_REG_8_ <= n2500;
    P2_REG3_REG_28_ <= n2505;
    P2_REG3_REG_19_ <= n2510;
    P2_REG3_REG_3_ <= n2515;
    P2_REG3_REG_10_ <= n2520;
    P2_REG3_REG_23_ <= n2525;
    P2_REG3_REG_14_ <= n2530;
    P2_REG3_REG_27_ <= n2535;
    P2_REG3_REG_7_ <= n2540;
    P2_STATE_REG <= n2545;
    P2_RD_REG <= n2550;
    P2_WR_REG <= n2555;
    P3_IR_REG_0_ <= n2560;
    P3_IR_REG_1_ <= n2565;
    P3_IR_REG_2_ <= n2570;
    P3_IR_REG_3_ <= n2575;
    P3_IR_REG_4_ <= n2580;
    P3_IR_REG_5_ <= n2585;
    P3_IR_REG_6_ <= n2590;
    P3_IR_REG_7_ <= n2595;
    P3_IR_REG_8_ <= n2600;
    P3_IR_REG_9_ <= n2605;
    P3_IR_REG_10_ <= n2610;
    P3_IR_REG_11_ <= n2615;
    P3_IR_REG_12_ <= n2620;
    P3_IR_REG_13_ <= n2625;
    P3_IR_REG_14_ <= n2630;
    P3_IR_REG_15_ <= n2635;
    P3_IR_REG_16_ <= n2640;
    P3_IR_REG_17_ <= n2645;
    P3_IR_REG_18_ <= n2650;
    P3_IR_REG_19_ <= n2655;
    P3_IR_REG_20_ <= n2660;
    P3_IR_REG_21_ <= n2665;
    P3_IR_REG_22_ <= n2670;
    P3_IR_REG_23_ <= n2675;
    P3_IR_REG_24_ <= n2680;
    P3_IR_REG_25_ <= n2685;
    P3_IR_REG_26_ <= n2690;
    P3_IR_REG_27_ <= n2695;
    P3_IR_REG_28_ <= n2700;
    P3_IR_REG_29_ <= n2705;
    P3_IR_REG_30_ <= n2710;
    P3_IR_REG_31_ <= n2715;
    P3_D_REG_0_ <= n2720;
    P3_D_REG_1_ <= n2725;
    P3_D_REG_2_ <= n2730;
    P3_D_REG_3_ <= n2735;
    P3_D_REG_4_ <= n2740;
    P3_D_REG_5_ <= n2745;
    P3_D_REG_6_ <= n2750;
    P3_D_REG_7_ <= n2755;
    P3_D_REG_8_ <= n2760;
    P3_D_REG_9_ <= n2765;
    P3_D_REG_10_ <= n2770;
    P3_D_REG_11_ <= n2775;
    P3_D_REG_12_ <= n2780;
    P3_D_REG_13_ <= n2785;
    P3_D_REG_14_ <= n2790;
    P3_D_REG_15_ <= n2795;
    P3_D_REG_16_ <= n2800;
    P3_D_REG_17_ <= n2805;
    P3_D_REG_18_ <= n2810;
    P3_D_REG_19_ <= n2815;
    P3_D_REG_20_ <= n2820;
    P3_D_REG_21_ <= n2825;
    P3_D_REG_22_ <= n2830;
    P3_D_REG_23_ <= n2835;
    P3_D_REG_24_ <= n2840;
    P3_D_REG_25_ <= n2845;
    P3_D_REG_26_ <= n2850;
    P3_D_REG_27_ <= n2855;
    P3_D_REG_28_ <= n2860;
    P3_D_REG_29_ <= n2865;
    P3_D_REG_30_ <= n2870;
    P3_D_REG_31_ <= n2875;
    P3_REG0_REG_0_ <= n2880;
    P3_REG0_REG_1_ <= n2885;
    P3_REG0_REG_2_ <= n2890;
    P3_REG0_REG_3_ <= n2895;
    P3_REG0_REG_4_ <= n2900;
    P3_REG0_REG_5_ <= n2905;
    P3_REG0_REG_6_ <= n2910;
    P3_REG0_REG_7_ <= n2915;
    P3_REG0_REG_8_ <= n2920;
    P3_REG0_REG_9_ <= n2925;
    P3_REG0_REG_10_ <= n2930;
    P3_REG0_REG_11_ <= n2935;
    P3_REG0_REG_12_ <= n2940;
    P3_REG0_REG_13_ <= n2945;
    P3_REG0_REG_14_ <= n2950;
    P3_REG0_REG_15_ <= n2955;
    P3_REG0_REG_16_ <= n2960;
    P3_REG0_REG_17_ <= n2965;
    P3_REG0_REG_18_ <= n2970;
    P3_REG0_REG_19_ <= n2975;
    P3_REG0_REG_20_ <= n2980;
    P3_REG0_REG_21_ <= n2985;
    P3_REG0_REG_22_ <= n2990;
    P3_REG0_REG_23_ <= n2995;
    P3_REG0_REG_24_ <= n3000;
    P3_REG0_REG_25_ <= n3005;
    P3_REG0_REG_26_ <= n3010;
    P3_REG0_REG_27_ <= n3015;
    P3_REG0_REG_28_ <= n3020;
    P3_REG0_REG_29_ <= n3025;
    P3_REG0_REG_30_ <= n3030;
    P3_REG0_REG_31_ <= n3035;
    P3_REG1_REG_0_ <= n3040;
    P3_REG1_REG_1_ <= n3045;
    P3_REG1_REG_2_ <= n3050;
    P3_REG1_REG_3_ <= n3055;
    P3_REG1_REG_4_ <= n3060;
    P3_REG1_REG_5_ <= n3065;
    P3_REG1_REG_6_ <= n3070;
    P3_REG1_REG_7_ <= n3075;
    P3_REG1_REG_8_ <= n3080;
    P3_REG1_REG_9_ <= n3085;
    P3_REG1_REG_10_ <= n3090;
    P3_REG1_REG_11_ <= n3095;
    P3_REG1_REG_12_ <= n3100;
    P3_REG1_REG_13_ <= n3105;
    P3_REG1_REG_14_ <= n3110;
    P3_REG1_REG_15_ <= n3115;
    P3_REG1_REG_16_ <= n3120;
    P3_REG1_REG_17_ <= n3125;
    P3_REG1_REG_18_ <= n3130;
    P3_REG1_REG_19_ <= n3135;
    P3_REG1_REG_20_ <= n3140;
    P3_REG1_REG_21_ <= n3145;
    P3_REG1_REG_22_ <= n3150;
    P3_REG1_REG_23_ <= n3155;
    P3_REG1_REG_24_ <= n3160;
    P3_REG1_REG_25_ <= n3165;
    P3_REG1_REG_26_ <= n3170;
    P3_REG1_REG_27_ <= n3175;
    P3_REG1_REG_28_ <= n3180;
    P3_REG1_REG_29_ <= n3185;
    P3_REG1_REG_30_ <= n3190;
    P3_REG1_REG_31_ <= n3195;
    P3_REG2_REG_0_ <= n3200;
    P3_REG2_REG_1_ <= n3205;
    P3_REG2_REG_2_ <= n3210;
    P3_REG2_REG_3_ <= n3215;
    P3_REG2_REG_4_ <= n3220;
    P3_REG2_REG_5_ <= n3225;
    P3_REG2_REG_6_ <= n3230;
    P3_REG2_REG_7_ <= n3235;
    P3_REG2_REG_8_ <= n3240;
    P3_REG2_REG_9_ <= n3245;
    P3_REG2_REG_10_ <= n3250;
    P3_REG2_REG_11_ <= n3255;
    P3_REG2_REG_12_ <= n3260;
    P3_REG2_REG_13_ <= n3265;
    P3_REG2_REG_14_ <= n3270;
    P3_REG2_REG_15_ <= n3275;
    P3_REG2_REG_16_ <= n3280;
    P3_REG2_REG_17_ <= n3285;
    P3_REG2_REG_18_ <= n3290;
    P3_REG2_REG_19_ <= n3295;
    P3_REG2_REG_20_ <= n3300;
    P3_REG2_REG_21_ <= n3305;
    P3_REG2_REG_22_ <= n3310;
    P3_REG2_REG_23_ <= n3315;
    P3_REG2_REG_24_ <= n3320;
    P3_REG2_REG_25_ <= n3325;
    P3_REG2_REG_26_ <= n3330;
    P3_REG2_REG_27_ <= n3335;
    P3_REG2_REG_28_ <= n3340;
    P3_REG2_REG_29_ <= n3345;
    P3_REG2_REG_30_ <= n3350;
    P3_REG2_REG_31_ <= n3355;
    P3_ADDR_REG_19_ <= n3360;
    P3_ADDR_REG_18_ <= n3365;
    P3_ADDR_REG_17_ <= n3370;
    P3_ADDR_REG_16_ <= n3375;
    P3_ADDR_REG_15_ <= n3380;
    P3_ADDR_REG_14_ <= n3385;
    P3_ADDR_REG_13_ <= n3390;
    P3_ADDR_REG_12_ <= n3395;
    P3_ADDR_REG_11_ <= n3400;
    P3_ADDR_REG_10_ <= n3405;
    P3_ADDR_REG_9_ <= n3410;
    P3_ADDR_REG_8_ <= n3415;
    P3_ADDR_REG_7_ <= n3420;
    P3_ADDR_REG_6_ <= n3425;
    P3_ADDR_REG_5_ <= n3430;
    P3_ADDR_REG_4_ <= n3435;
    P3_ADDR_REG_3_ <= n3440;
    P3_ADDR_REG_2_ <= n3445;
    P3_ADDR_REG_1_ <= n3450;
    P3_ADDR_REG_0_ <= n3455;
    P3_DATAO_REG_0_ <= n3460;
    P3_DATAO_REG_1_ <= n3465;
    P3_DATAO_REG_2_ <= n3470;
    P3_DATAO_REG_3_ <= n3475;
    P3_DATAO_REG_4_ <= n3480;
    P3_DATAO_REG_5_ <= n3485;
    P3_DATAO_REG_6_ <= n3490;
    P3_DATAO_REG_7_ <= n3495;
    P3_DATAO_REG_8_ <= n3500;
    P3_DATAO_REG_9_ <= n3505;
    P3_DATAO_REG_10_ <= n3510;
    P3_DATAO_REG_11_ <= n3515;
    P3_DATAO_REG_12_ <= n3520;
    P3_DATAO_REG_13_ <= n3525;
    P3_DATAO_REG_14_ <= n3530;
    P3_DATAO_REG_15_ <= n3535;
    P3_DATAO_REG_16_ <= n3540;
    P3_DATAO_REG_17_ <= n3545;
    P3_DATAO_REG_18_ <= n3550;
    P3_DATAO_REG_19_ <= n3555;
    P3_DATAO_REG_20_ <= n3560;
    P3_DATAO_REG_21_ <= n3565;
    P3_DATAO_REG_22_ <= n3570;
    P3_DATAO_REG_23_ <= n3575;
    P3_DATAO_REG_24_ <= n3580;
    P3_DATAO_REG_25_ <= n3585;
    P3_DATAO_REG_26_ <= n3590;
    P3_DATAO_REG_27_ <= n3595;
    P3_DATAO_REG_28_ <= n3600;
    P3_DATAO_REG_29_ <= n3605;
    P3_DATAO_REG_30_ <= n3610;
    P3_DATAO_REG_31_ <= n3615;
    P3_B_REG <= n3620;
    P3_REG3_REG_15_ <= n3625;
    P3_REG3_REG_26_ <= n3630;
    P3_REG3_REG_6_ <= n3635;
    P3_REG3_REG_18_ <= n3640;
    P3_REG3_REG_2_ <= n3645;
    P3_REG3_REG_11_ <= n3650;
    P3_REG3_REG_22_ <= n3655;
    P3_REG3_REG_13_ <= n3660;
    P3_REG3_REG_20_ <= n3665;
    P3_REG3_REG_0_ <= n3670;
    P3_REG3_REG_9_ <= n3675;
    P3_REG3_REG_4_ <= n3680;
    P3_REG3_REG_24_ <= n3685;
    P3_REG3_REG_17_ <= n3690;
    P3_REG3_REG_5_ <= n3695;
    P3_REG3_REG_16_ <= n3700;
    P3_REG3_REG_25_ <= n3705;
    P3_REG3_REG_12_ <= n3710;
    P3_REG3_REG_21_ <= n3715;
    P3_REG3_REG_1_ <= n3720;
    P3_REG3_REG_8_ <= n3725;
    P3_REG3_REG_28_ <= n3730;
    P3_REG3_REG_19_ <= n3735;
    P3_REG3_REG_3_ <= n3740;
    P3_REG3_REG_10_ <= n3745;
    P3_REG3_REG_23_ <= n3750;
    P3_REG3_REG_14_ <= n3755;
    P3_REG3_REG_27_ <= n3760;
    P3_REG3_REG_7_ <= n3765;
    P3_STATE_REG <= n3770;
    P3_RD_REG <= n3775;
    P3_WR_REG <= n3780;
  end
endmodule


