module top ( 
    \1 , 8, 13, 17, 26, 29, 36, 42, 51, 55, 59, 68, 72, 73, 74, 75, 80, 85,
    86, 87, 88, 89, 90, 91, 96, 101, 106, 111, 116, 121, 126, 130, 135,
    138, 143, 146, 149, 152, 153, 156, 159, 165, 171, 177, 183, 189, 195,
    201, 207, 210, 219, 228, 237, 246, 255, 259, 260, 261, 267, 268,
    388, 389, 390, 391, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449,
    450, 767, 768, 850, 863, 864, 865, 866, 874, 878, 879, 880  );
  input  \1 , 8, 13, 17, 26, 29, 36, 42, 51, 55, 59, 68, 72, 73, 74, 75,
    80, 85, 86, 87, 88, 89, 90, 91, 96, 101, 106, 111, 116, 121, 126, 130,
    135, 138, 143, 146, 149, 152, 153, 156, 159, 165, 171, 177, 183, 189,
    195, 201, 207, 210, 219, 228, 237, 246, 255, 259, 260, 261, 267, 268;
  output 388, 389, 390, 391, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449,
    450, 767, 768, 850, 863, 864, 865, 866, 874, 878, 879, 880;
  wire n87, n89, n93, n94, n96, n97, n98, n100, n102, n105, n109, n110, n112,
    n113, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412;
  assign n87 = 29 & 75;
  assign 388 = 42 & n87;
  assign n89 = 29 & 36;
  assign 389 = 80 & n89;
  assign 390 = 42 & n89;
  assign 391 = 85 & 86;
  assign n93 = \1  & 8;
  assign n94 = 13 & n93;
  assign 418 = 17 & n94;
  assign n96 = \1  & 26;
  assign n97 = 13 & n96;
  assign n98 = 17 & n97;
  assign 419 = 390 | ~n98;
  assign n100 = 59 & 75;
  assign 420 = ~80 | ~n100;
  assign n102 = 36 & 59;
  assign 421 = ~80 | ~n102;
  assign 422 = ~42 | ~n102;
  assign n105 = ~87 & ~88;
  assign 423 = 90 & ~n105;
  assign 446 = ~390 | ~n98;
  assign 447 = 51 & n96;
  assign n109 = 55 & n94;
  assign n110 = 29 & 68;
  assign 448 = n109 & n110;
  assign n112 = 59 & 68;
  assign n113 = 74 & n112;
  assign 449 = n109 & n113;
  assign 450 = 89 & ~n105;
  assign n116 = 91 & 96;
  assign n117 = ~91 & ~96;
  assign n118 = ~n116 & ~n117;
  assign n119 = 101 & 106;
  assign n120 = ~101 & ~106;
  assign n121 = ~n119 & ~n120;
  assign n122 = ~n118 & ~n121;
  assign n123 = n118 & n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = 130 & n124;
  assign n126 = ~130 & ~n124;
  assign n127 = ~n125 & ~n126;
  assign n128 = 111 & 116;
  assign n129 = ~111 & ~116;
  assign n130 = ~n128 & ~n129;
  assign n131 = 121 & 126;
  assign n132 = ~121 & ~126;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n130 & ~n133;
  assign n135 = n130 & n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = 135 & n136;
  assign n138 = ~135 & ~n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~n127 & ~n139;
  assign n141 = n127 & n139;
  assign 767 = ~n140 & ~n141;
  assign n143 = 159 & 165;
  assign n144 = ~159 & ~165;
  assign n145 = ~n143 & ~n144;
  assign n146 = 171 & 177;
  assign n147 = ~171 & ~177;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = n145 & n148;
  assign n151 = ~n149 & ~n150;
  assign n152 = 130 & n151;
  assign n153 = ~130 & ~n151;
  assign n154 = ~n152 & ~n153;
  assign n155 = 183 & 189;
  assign n156 = ~183 & ~189;
  assign n157 = ~n155 & ~n156;
  assign n158 = 195 & 201;
  assign n159 = ~195 & ~201;
  assign n160 = ~n158 & ~n159;
  assign n161 = ~n157 & ~n160;
  assign n162 = n157 & n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = 207 & n163;
  assign n165 = ~207 & ~n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = ~n154 & ~n166;
  assign n168 = n154 & n166;
  assign 768 = ~n167 & ~n168;
  assign n170 = 121 & 210;
  assign n171 = 80 & n87;
  assign n172 = 447 & n171;
  assign n173 = 55 & n172;
  assign n174 = ~268 & n173;
  assign n175 = 59 & 156;
  assign n176 = 447 & ~n175;
  assign n177 = 17 & n176;
  assign n178 = \1  & ~n177;
  assign n179 = 153 & ~n178;
  assign n180 = ~17 & ~42;
  assign n181 = 17 & 42;
  assign n182 = ~n180 & ~n181;
  assign n183 = 59 & n182;
  assign n184 = 156 & n183;
  assign n185 = 447 & n184;
  assign n186 = 51 & n93;
  assign n187 = 17 & n186;
  assign n188 = 42 & n100;
  assign n189 = n187 & ~n188;
  assign n190 = ~n185 & ~n189;
  assign n191 = 126 & ~n190;
  assign n192 = ~n179 & ~n191;
  assign n193 = ~n174 & n192;
  assign n194 = ~201 & n193;
  assign n195 = 201 & ~n193;
  assign n196 = ~n194 & ~n195;
  assign n197 = ~261 & ~n196;
  assign n198 = 261 & n196;
  assign n199 = ~n197 & ~n198;
  assign n200 = 219 & n199;
  assign n201 = ~n170 & ~n200;
  assign n202 = 228 & n196;
  assign n203 = 237 & n195;
  assign n204 = ~n202 & ~n203;
  assign n205 = 255 & 267;
  assign n206 = 246 & ~n193;
  assign n207 = ~n205 & ~n206;
  assign n208 = 42 & 59;
  assign n209 = 68 & n208;
  assign n210 = 72 & n209;
  assign n211 = n109 & n210;
  assign n212 = 73 & n211;
  assign n213 = 201 & n212;
  assign n214 = n201 & n204;
  assign n215 = n207 & n214;
  assign 850 = n213 | ~n215;
  assign n217 = 106 & 210;
  assign n218 = 143 & ~n178;
  assign n219 = 111 & ~n190;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~n174 & n220;
  assign n222 = ~183 & n221;
  assign n223 = 183 & ~n221;
  assign n224 = ~n222 & ~n223;
  assign n225 = 146 & ~n178;
  assign n226 = 116 & ~n190;
  assign n227 = ~n225 & ~n226;
  assign n228 = ~n174 & n227;
  assign n229 = 189 & ~n228;
  assign n230 = ~189 & n228;
  assign n231 = 149 & ~n178;
  assign n232 = 121 & ~n190;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n174 & n233;
  assign n235 = 195 & ~n234;
  assign n236 = ~n230 & n235;
  assign n237 = ~195 & n234;
  assign n238 = ~n230 & ~n237;
  assign n239 = n195 & n238;
  assign n240 = ~n194 & n238;
  assign n241 = 261 & n240;
  assign n242 = ~n229 & ~n236;
  assign n243 = ~n239 & n242;
  assign n244 = ~n241 & n243;
  assign n245 = ~n224 & n244;
  assign n246 = n224 & ~n244;
  assign n247 = ~n245 & ~n246;
  assign n248 = 219 & n247;
  assign n249 = ~n217 & ~n248;
  assign n250 = 228 & n224;
  assign n251 = 237 & n223;
  assign n252 = ~n250 & ~n251;
  assign n253 = 246 & ~n221;
  assign n254 = 183 & n212;
  assign n255 = ~n253 & ~n254;
  assign n256 = n249 & n252;
  assign 863 = ~n255 | ~n256;
  assign n258 = 111 & 210;
  assign n259 = ~n229 & ~n230;
  assign n260 = n195 & ~n237;
  assign n261 = ~n194 & ~n237;
  assign n262 = 261 & n261;
  assign n263 = ~n235 & ~n260;
  assign n264 = ~n262 & n263;
  assign n265 = ~n259 & n264;
  assign n266 = n259 & ~n264;
  assign n267 = ~n265 & ~n266;
  assign n268 = 219 & n267;
  assign n269 = ~n258 & ~n268;
  assign n270 = 228 & n259;
  assign n271 = 237 & n229;
  assign n272 = ~n270 & ~n271;
  assign n273 = 255 & 259;
  assign n274 = 246 & ~n228;
  assign n275 = ~n273 & ~n274;
  assign n276 = 189 & n212;
  assign n277 = n269 & n272;
  assign n278 = n275 & n277;
  assign 864 = n276 | ~n278;
  assign n280 = 116 & 210;
  assign n281 = ~n235 & ~n237;
  assign n282 = 261 & ~n194;
  assign n283 = ~n195 & ~n282;
  assign n284 = ~n281 & n283;
  assign n285 = n281 & ~n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = 219 & n286;
  assign n288 = ~n280 & ~n287;
  assign n289 = 228 & n281;
  assign n290 = 237 & n235;
  assign n291 = ~n289 & ~n290;
  assign n292 = 255 & 260;
  assign n293 = 246 & ~n234;
  assign n294 = ~n292 & ~n293;
  assign n295 = 195 & n212;
  assign n296 = n288 & n291;
  assign n297 = n294 & n296;
  assign 865 = n295 | ~n297;
  assign n299 = 8 & 138;
  assign n300 = 91 & ~n190;
  assign n301 = ~n299 & ~n300;
  assign n302 = 55 & n176;
  assign n303 = 143 & n302;
  assign n304 = 17 & 447;
  assign n305 = n171 & n304;
  assign n306 = ~268 & n305;
  assign n307 = ~n303 & ~n306;
  assign n308 = n301 & n307;
  assign n309 = 159 & ~n308;
  assign n310 = 51 & 138;
  assign n311 = 96 & ~n190;
  assign n312 = ~n310 & ~n311;
  assign n313 = 146 & n302;
  assign n314 = ~n306 & ~n313;
  assign n315 = n312 & n314;
  assign n316 = 165 & ~n315;
  assign n317 = ~165 & n315;
  assign n318 = 17 & 138;
  assign n319 = 101 & ~n190;
  assign n320 = ~n318 & ~n319;
  assign n321 = 149 & n302;
  assign n322 = ~n306 & ~n321;
  assign n323 = n320 & n322;
  assign n324 = 171 & ~n323;
  assign n325 = ~n317 & n324;
  assign n326 = ~171 & n323;
  assign n327 = 138 & 152;
  assign n328 = 106 & ~n190;
  assign n329 = ~n327 & ~n328;
  assign n330 = 153 & n302;
  assign n331 = ~n306 & ~n330;
  assign n332 = n329 & n331;
  assign n333 = 177 & ~n332;
  assign n334 = ~n317 & ~n326;
  assign n335 = n333 & n334;
  assign n336 = ~177 & n332;
  assign n337 = ~n222 & ~n244;
  assign n338 = ~n223 & ~n337;
  assign n339 = n334 & ~n336;
  assign n340 = ~n338 & n339;
  assign n341 = ~n316 & ~n325;
  assign n342 = ~n335 & n341;
  assign n343 = ~n340 & n342;
  assign n344 = ~159 & n308;
  assign n345 = ~n343 & ~n344;
  assign 866 = n309 | n345;
  assign n347 = 101 & 210;
  assign n348 = ~n333 & ~n336;
  assign n349 = n338 & ~n348;
  assign n350 = ~n338 & n348;
  assign n351 = ~n349 & ~n350;
  assign n352 = 219 & n351;
  assign n353 = ~n347 & ~n352;
  assign n354 = 228 & n348;
  assign n355 = 237 & n333;
  assign n356 = ~n354 & ~n355;
  assign n357 = 246 & ~n332;
  assign n358 = 177 & n212;
  assign n359 = ~n357 & ~n358;
  assign n360 = n353 & n356;
  assign 874 = ~n359 | ~n360;
  assign n362 = 210 & 268;
  assign n363 = ~n309 & ~n344;
  assign n364 = n343 & ~n363;
  assign n365 = ~n343 & n363;
  assign n366 = ~n364 & ~n365;
  assign n367 = 219 & n366;
  assign n368 = ~n362 & ~n367;
  assign n369 = 228 & n363;
  assign n370 = 237 & n309;
  assign n371 = ~n369 & ~n370;
  assign n372 = 246 & ~n308;
  assign n373 = 159 & n212;
  assign n374 = ~n372 & ~n373;
  assign n375 = n368 & n371;
  assign 878 = ~n374 | ~n375;
  assign n377 = 91 & 210;
  assign n378 = ~n316 & ~n317;
  assign n379 = ~n326 & n333;
  assign n380 = ~n326 & ~n336;
  assign n381 = ~n338 & n380;
  assign n382 = ~n324 & ~n379;
  assign n383 = ~n381 & n382;
  assign n384 = ~n378 & n383;
  assign n385 = n378 & ~n383;
  assign n386 = ~n384 & ~n385;
  assign n387 = 219 & n386;
  assign n388 = ~n377 & ~n387;
  assign n389 = 228 & n378;
  assign n390 = 237 & n316;
  assign n391 = ~n389 & ~n390;
  assign n392 = 246 & ~n315;
  assign n393 = 165 & n212;
  assign n394 = ~n392 & ~n393;
  assign n395 = n388 & n391;
  assign 879 = ~n394 | ~n395;
  assign n397 = 96 & 210;
  assign n398 = ~n324 & ~n326;
  assign n399 = ~n336 & ~n338;
  assign n400 = ~n333 & ~n399;
  assign n401 = ~n398 & n400;
  assign n402 = n398 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = 219 & n403;
  assign n405 = ~n397 & ~n404;
  assign n406 = 228 & n398;
  assign n407 = 237 & n324;
  assign n408 = ~n406 & ~n407;
  assign n409 = 246 & ~n323;
  assign n410 = 171 & n212;
  assign n411 = ~n409 & ~n410;
  assign n412 = n405 & n408;
  assign 880 = ~n411 | ~n412;
endmodule


