// Benchmark "top" written by ABC on Mon Nov 27 16:55:46 2023

module top ( 
    \1 , \8 , \15 , \22 , \29 , \36 , \43 , \50 , \57 , \64 , \71 , \78 ,
    \85 , \92 , \99 , \106 , \113 , \120 , \127 , \134 , \141 , \148 ,
    \155 , \162 , \169 , \176 , \183 , \190 , \197 , \204 , \211 , \218 ,
    \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ,
    \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
    \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
    \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
    \1351 , \1352 , \1353 , \1354 , \1355   );
  input  \1 , \8 , \15 , \22 , \29 , \36 , \43 , \50 , \57 , \64 , \71 ,
    \78 , \85 , \92 , \99 , \106 , \113 , \120 , \127 , \134 , \141 ,
    \148 , \155 , \162 , \169 , \176 , \183 , \190 , \197 , \204 , \211 ,
    \218 , \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ;
  output \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
    \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
    \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 ,
    \1350 , \1351 , \1352 , \1353 , \1354 , \1355 ;
  wire new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n326, new_n327, new_n328, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n336, new_n337, new_n338, new_n340,
    new_n341, new_n342, new_n344, new_n345, new_n346, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n354, new_n355, new_n356, new_n358,
    new_n359, new_n360, new_n362, new_n363, new_n364, new_n366, new_n367,
    new_n368, new_n369, new_n371, new_n372, new_n373, new_n375, new_n376,
    new_n377, new_n379, new_n380, new_n381, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n390, new_n391, new_n392, new_n394,
    new_n395, new_n396, new_n398, new_n399, new_n400, new_n402, new_n403,
    new_n404, new_n405, new_n407, new_n408, new_n409, new_n411, new_n412,
    new_n413, new_n415, new_n416, new_n417, new_n419, new_n420, new_n421,
    new_n422, new_n424, new_n425, new_n426, new_n428, new_n429, new_n430,
    new_n432, new_n433, new_n434, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n442, new_n443, new_n444, new_n446, new_n447, new_n448,
    new_n450, new_n451, new_n452;
  assign new_n74 = ~\113  & ~\120 ;
  assign new_n75 = \113  & \120 ;
  assign new_n76 = ~new_n74 & ~new_n75;
  assign new_n77 = \127  & ~\134 ;
  assign new_n78 = ~\127  & \134 ;
  assign new_n79 = ~new_n77 & ~new_n78;
  assign new_n80 = new_n76 & new_n79;
  assign new_n81 = ~new_n76 & ~new_n79;
  assign new_n82 = ~new_n80 & ~new_n81;
  assign new_n83 = \225  & \233 ;
  assign new_n84 = \29  & ~new_n83;
  assign new_n85 = ~\29  & new_n83;
  assign new_n86 = ~new_n84 & ~new_n85;
  assign new_n87 = ~new_n82 & new_n86;
  assign new_n88 = new_n82 & ~new_n86;
  assign new_n89 = ~new_n87 & ~new_n88;
  assign new_n90 = ~\141  & ~\148 ;
  assign new_n91 = \141  & \148 ;
  assign new_n92 = ~new_n90 & ~new_n91;
  assign new_n93 = \155  & ~\162 ;
  assign new_n94 = ~\155  & \162 ;
  assign new_n95 = ~new_n93 & ~new_n94;
  assign new_n96 = new_n92 & new_n95;
  assign new_n97 = ~new_n92 & ~new_n95;
  assign new_n98 = ~new_n96 & ~new_n97;
  assign new_n99 = ~\1  & ~\85 ;
  assign new_n100 = \1  & \85 ;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = \57  & new_n101;
  assign new_n103 = ~\57  & ~new_n101;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = ~new_n98 & new_n104;
  assign new_n106 = new_n98 & ~new_n104;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = new_n89 & new_n107;
  assign new_n109 = ~new_n89 & ~new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = \230  & \233 ;
  assign new_n112 = \176  & ~new_n111;
  assign new_n113 = ~\176  & new_n111;
  assign new_n114 = ~new_n112 & ~new_n113;
  assign new_n115 = ~\85  & ~\92 ;
  assign new_n116 = \85  & \92 ;
  assign new_n117 = ~new_n115 & ~new_n116;
  assign new_n118 = \99  & ~\106 ;
  assign new_n119 = ~\99  & \106 ;
  assign new_n120 = ~new_n118 & ~new_n119;
  assign new_n121 = new_n117 & new_n120;
  assign new_n122 = ~new_n117 & ~new_n120;
  assign new_n123 = ~new_n121 & ~new_n122;
  assign new_n124 = new_n114 & ~new_n123;
  assign new_n125 = ~new_n114 & new_n123;
  assign new_n126 = ~new_n124 & ~new_n125;
  assign new_n127 = ~\120  & ~\148 ;
  assign new_n128 = \120  & \148 ;
  assign new_n129 = ~new_n127 & ~new_n128;
  assign new_n130 = \204  & new_n129;
  assign new_n131 = ~\204  & ~new_n129;
  assign new_n132 = ~new_n130 & ~new_n131;
  assign new_n133 = ~\57  & ~\64 ;
  assign new_n134 = \57  & \64 ;
  assign new_n135 = ~new_n133 & ~new_n134;
  assign new_n136 = \71  & ~\78 ;
  assign new_n137 = ~\71  & \78 ;
  assign new_n138 = ~new_n136 & ~new_n137;
  assign new_n139 = new_n135 & new_n138;
  assign new_n140 = ~new_n135 & ~new_n138;
  assign new_n141 = ~new_n139 & ~new_n140;
  assign new_n142 = new_n132 & ~new_n141;
  assign new_n143 = ~new_n132 & new_n141;
  assign new_n144 = ~new_n142 & ~new_n143;
  assign new_n145 = new_n126 & new_n144;
  assign new_n146 = ~new_n126 & ~new_n144;
  assign new_n147 = ~new_n145 & ~new_n146;
  assign new_n148 = \232  & \233 ;
  assign new_n149 = \190  & ~new_n148;
  assign new_n150 = ~\190  & new_n148;
  assign new_n151 = ~new_n149 & ~new_n150;
  assign new_n152 = ~new_n123 & new_n151;
  assign new_n153 = new_n123 & ~new_n151;
  assign new_n154 = ~new_n152 & ~new_n153;
  assign new_n155 = ~\134  & ~\162 ;
  assign new_n156 = \134  & \162 ;
  assign new_n157 = ~new_n155 & ~new_n156;
  assign new_n158 = \218  & new_n157;
  assign new_n159 = ~\218  & ~new_n157;
  assign new_n160 = ~new_n158 & ~new_n159;
  assign new_n161 = ~\29  & ~\36 ;
  assign new_n162 = \29  & \36 ;
  assign new_n163 = ~new_n161 & ~new_n162;
  assign new_n164 = \43  & ~\50 ;
  assign new_n165 = ~\43  & \50 ;
  assign new_n166 = ~new_n164 & ~new_n165;
  assign new_n167 = new_n163 & new_n166;
  assign new_n168 = ~new_n163 & ~new_n166;
  assign new_n169 = ~new_n167 & ~new_n168;
  assign new_n170 = new_n160 & ~new_n169;
  assign new_n171 = ~new_n160 & new_n169;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = new_n154 & new_n172;
  assign new_n174 = ~new_n154 & ~new_n172;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176 = new_n147 & new_n175;
  assign new_n177 = ~\197  & ~\204 ;
  assign new_n178 = \197  & \204 ;
  assign new_n179 = ~new_n177 & ~new_n178;
  assign new_n180 = \211  & ~\218 ;
  assign new_n181 = ~\211  & \218 ;
  assign new_n182 = ~new_n180 & ~new_n181;
  assign new_n183 = new_n179 & new_n182;
  assign new_n184 = ~new_n179 & ~new_n182;
  assign new_n185 = ~new_n183 & ~new_n184;
  assign new_n186 = \226  & \233 ;
  assign new_n187 = \64  & ~new_n186;
  assign new_n188 = ~\64  & new_n186;
  assign new_n189 = ~new_n187 & ~new_n188;
  assign new_n190 = new_n185 & ~new_n189;
  assign new_n191 = ~new_n185 & new_n189;
  assign new_n192 = ~new_n190 & ~new_n191;
  assign new_n193 = ~\169  & ~\176 ;
  assign new_n194 = \169  & \176 ;
  assign new_n195 = ~new_n193 & ~new_n194;
  assign new_n196 = \183  & ~\190 ;
  assign new_n197 = ~\183  & \190 ;
  assign new_n198 = ~new_n196 & ~new_n197;
  assign new_n199 = new_n195 & new_n198;
  assign new_n200 = ~new_n195 & ~new_n198;
  assign new_n201 = ~new_n199 & ~new_n200;
  assign new_n202 = ~\8  & ~\36 ;
  assign new_n203 = \8  & \36 ;
  assign new_n204 = ~new_n202 & ~new_n203;
  assign new_n205 = \92  & ~new_n204;
  assign new_n206 = ~\92  & new_n204;
  assign new_n207 = ~new_n205 & ~new_n206;
  assign new_n208 = new_n201 & ~new_n207;
  assign new_n209 = ~new_n201 & new_n207;
  assign new_n210 = ~new_n208 & ~new_n209;
  assign new_n211 = new_n192 & new_n210;
  assign new_n212 = ~new_n192 & ~new_n210;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = \227  & \233 ;
  assign new_n215 = \71  & ~new_n214;
  assign new_n216 = ~\71  & new_n214;
  assign new_n217 = ~new_n215 & ~new_n216;
  assign new_n218 = new_n82 & ~new_n217;
  assign new_n219 = ~new_n82 & new_n217;
  assign new_n220 = ~new_n218 & ~new_n219;
  assign new_n221 = ~\15  & ~\43 ;
  assign new_n222 = \15  & \43 ;
  assign new_n223 = ~new_n221 & ~new_n222;
  assign new_n224 = \99  & ~new_n223;
  assign new_n225 = ~\99  & new_n223;
  assign new_n226 = ~new_n224 & ~new_n225;
  assign new_n227 = new_n201 & ~new_n226;
  assign new_n228 = ~new_n201 & new_n226;
  assign new_n229 = ~new_n227 & ~new_n228;
  assign new_n230 = new_n220 & new_n229;
  assign new_n231 = ~new_n220 & ~new_n229;
  assign new_n232 = ~new_n230 & ~new_n231;
  assign new_n233 = ~new_n213 & ~new_n232;
  assign new_n234 = \228  & \233 ;
  assign new_n235 = \78  & ~new_n234;
  assign new_n236 = ~\78  & new_n234;
  assign new_n237 = ~new_n235 & ~new_n236;
  assign new_n238 = new_n98 & ~new_n237;
  assign new_n239 = ~new_n98 & new_n237;
  assign new_n240 = ~new_n238 & ~new_n239;
  assign new_n241 = ~\22  & ~\50 ;
  assign new_n242 = \22  & \50 ;
  assign new_n243 = ~new_n241 & ~new_n242;
  assign new_n244 = \106  & ~new_n243;
  assign new_n245 = ~\106  & new_n243;
  assign new_n246 = ~new_n244 & ~new_n245;
  assign new_n247 = new_n185 & ~new_n246;
  assign new_n248 = ~new_n185 & new_n246;
  assign new_n249 = ~new_n247 & ~new_n248;
  assign new_n250 = new_n240 & new_n249;
  assign new_n251 = ~new_n240 & ~new_n249;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253 = ~new_n233 & new_n252;
  assign new_n254 = new_n233 & ~new_n252;
  assign new_n255 = new_n213 & new_n232;
  assign new_n256 = new_n110 & ~new_n255;
  assign new_n257 = ~new_n254 & ~new_n256;
  assign new_n258 = ~new_n253 & ~new_n257;
  assign new_n259 = \231  & \233 ;
  assign new_n260 = \183  & ~new_n259;
  assign new_n261 = ~\183  & new_n259;
  assign new_n262 = ~new_n260 & ~new_n261;
  assign new_n263 = new_n141 & ~new_n262;
  assign new_n264 = ~new_n141 & new_n262;
  assign new_n265 = ~new_n263 & ~new_n264;
  assign new_n266 = ~\1  & ~\8 ;
  assign new_n267 = \1  & \8 ;
  assign new_n268 = ~new_n266 & ~new_n267;
  assign new_n269 = \15  & ~\22 ;
  assign new_n270 = ~\15  & \22 ;
  assign new_n271 = ~new_n269 & ~new_n270;
  assign new_n272 = new_n268 & new_n271;
  assign new_n273 = ~new_n268 & ~new_n271;
  assign new_n274 = ~new_n272 & ~new_n273;
  assign new_n275 = ~\127  & ~\155 ;
  assign new_n276 = \127  & \155 ;
  assign new_n277 = ~new_n275 & ~new_n276;
  assign new_n278 = \211  & ~new_n277;
  assign new_n279 = ~\211  & new_n277;
  assign new_n280 = ~new_n278 & ~new_n279;
  assign new_n281 = new_n274 & ~new_n280;
  assign new_n282 = ~new_n274 & new_n280;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = new_n265 & new_n283;
  assign new_n285 = ~new_n265 & ~new_n283;
  assign new_n286 = ~new_n284 & ~new_n285;
  assign new_n287 = ~new_n176 & new_n286;
  assign new_n288 = new_n176 & ~new_n286;
  assign new_n289 = ~new_n147 & ~new_n175;
  assign new_n290 = \229  & \233 ;
  assign new_n291 = \169  & ~new_n290;
  assign new_n292 = ~\169  & new_n290;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294 = new_n169 & ~new_n293;
  assign new_n295 = ~new_n169 & new_n293;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = ~\113  & ~\141 ;
  assign new_n298 = \113  & \141 ;
  assign new_n299 = ~new_n297 & ~new_n298;
  assign new_n300 = \197  & ~new_n299;
  assign new_n301 = ~\197  & new_n299;
  assign new_n302 = ~new_n300 & ~new_n301;
  assign new_n303 = new_n274 & ~new_n302;
  assign new_n304 = ~new_n274 & new_n302;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = new_n296 & new_n305;
  assign new_n307 = ~new_n296 & ~new_n305;
  assign new_n308 = ~new_n306 & ~new_n307;
  assign new_n309 = ~new_n289 & ~new_n308;
  assign new_n310 = ~new_n288 & ~new_n309;
  assign new_n311 = ~new_n287 & ~new_n310;
  assign new_n312 = new_n258 & ~new_n311;
  assign new_n313 = new_n176 & new_n312;
  assign new_n314 = ~new_n110 & new_n313;
  assign new_n315 = \1  & ~new_n314;
  assign new_n316 = ~\1  & new_n314;
  assign \1324  = new_n315 | new_n316;
  assign new_n318 = new_n213 & new_n313;
  assign new_n319 = \8  & ~new_n318;
  assign new_n320 = ~\8  & new_n318;
  assign \1325  = new_n319 | new_n320;
  assign new_n322 = new_n232 & new_n313;
  assign new_n323 = \15  & ~new_n322;
  assign new_n324 = ~\15  & new_n322;
  assign \1326  = new_n323 | new_n324;
  assign new_n326 = new_n252 & new_n313;
  assign new_n327 = \22  & ~new_n326;
  assign new_n328 = ~\22  & new_n326;
  assign \1327  = new_n327 | new_n328;
  assign new_n330 = ~new_n286 & new_n312;
  assign new_n331 = new_n147 & new_n330;
  assign new_n332 = ~new_n110 & new_n331;
  assign new_n333 = \29  & ~new_n332;
  assign new_n334 = ~\29  & new_n332;
  assign \1328  = new_n333 | new_n334;
  assign new_n336 = new_n213 & new_n331;
  assign new_n337 = \36  & ~new_n336;
  assign new_n338 = ~\36  & new_n336;
  assign \1329  = new_n337 | new_n338;
  assign new_n340 = new_n232 & new_n331;
  assign new_n341 = \43  & ~new_n340;
  assign new_n342 = ~\43  & new_n340;
  assign \1330  = new_n341 | new_n342;
  assign new_n344 = new_n252 & new_n331;
  assign new_n345 = \50  & ~new_n344;
  assign new_n346 = ~\50  & new_n344;
  assign \1331  = new_n345 | new_n346;
  assign new_n348 = new_n175 & ~new_n308;
  assign new_n349 = new_n312 & new_n348;
  assign new_n350 = ~new_n110 & new_n349;
  assign new_n351 = \57  & ~new_n350;
  assign new_n352 = ~\57  & new_n350;
  assign \1332  = new_n351 | new_n352;
  assign new_n354 = new_n213 & new_n349;
  assign new_n355 = \64  & ~new_n354;
  assign new_n356 = ~\64  & new_n354;
  assign \1333  = new_n355 | new_n356;
  assign new_n358 = new_n232 & new_n349;
  assign new_n359 = ~\71  & ~new_n358;
  assign new_n360 = \71  & new_n358;
  assign \1334  = ~new_n359 & ~new_n360;
  assign new_n362 = new_n252 & new_n349;
  assign new_n363 = ~\78  & ~new_n362;
  assign new_n364 = \78  & new_n362;
  assign \1335  = ~new_n363 & ~new_n364;
  assign new_n366 = ~new_n308 & new_n330;
  assign new_n367 = ~new_n110 & new_n366;
  assign new_n368 = \85  & ~new_n367;
  assign new_n369 = ~\85  & new_n367;
  assign \1336  = new_n368 | new_n369;
  assign new_n371 = new_n213 & new_n366;
  assign new_n372 = \92  & ~new_n371;
  assign new_n373 = ~\92  & new_n371;
  assign \1337  = new_n372 | new_n373;
  assign new_n375 = new_n232 & new_n366;
  assign new_n376 = \99  & ~new_n375;
  assign new_n377 = ~\99  & new_n375;
  assign \1338  = new_n376 | new_n377;
  assign new_n379 = new_n252 & new_n366;
  assign new_n380 = \106  & ~new_n379;
  assign new_n381 = ~\106  & new_n379;
  assign \1339  = new_n380 | new_n381;
  assign new_n383 = ~new_n258 & new_n311;
  assign new_n384 = ~new_n252 & new_n383;
  assign new_n385 = ~new_n213 & new_n384;
  assign new_n386 = new_n308 & new_n385;
  assign new_n387 = ~\113  & ~new_n386;
  assign new_n388 = \113  & new_n386;
  assign \1340  = ~new_n387 & ~new_n388;
  assign new_n390 = ~new_n147 & new_n385;
  assign new_n391 = \120  & new_n390;
  assign new_n392 = ~\120  & ~new_n390;
  assign \1341  = ~new_n391 & ~new_n392;
  assign new_n394 = new_n286 & new_n385;
  assign new_n395 = ~\127  & ~new_n394;
  assign new_n396 = \127  & new_n394;
  assign \1342  = ~new_n395 & ~new_n396;
  assign new_n398 = ~new_n175 & new_n385;
  assign new_n399 = \134  & new_n398;
  assign new_n400 = ~\134  & ~new_n398;
  assign \1343  = ~new_n399 & ~new_n400;
  assign new_n402 = new_n233 & new_n383;
  assign new_n403 = new_n308 & new_n402;
  assign new_n404 = ~\141  & ~new_n403;
  assign new_n405 = \141  & new_n403;
  assign \1344  = ~new_n404 & ~new_n405;
  assign new_n407 = ~new_n147 & new_n402;
  assign new_n408 = \148  & ~new_n407;
  assign new_n409 = ~\148  & new_n407;
  assign \1345  = new_n408 | new_n409;
  assign new_n411 = new_n286 & new_n402;
  assign new_n412 = \155  & ~new_n411;
  assign new_n413 = ~\155  & new_n411;
  assign \1346  = new_n412 | new_n413;
  assign new_n415 = ~new_n175 & new_n402;
  assign new_n416 = \162  & ~new_n415;
  assign new_n417 = ~\162  & new_n415;
  assign \1347  = new_n416 | new_n417;
  assign new_n419 = new_n110 & new_n384;
  assign new_n420 = new_n308 & new_n419;
  assign new_n421 = ~\169  & ~new_n420;
  assign new_n422 = \169  & new_n420;
  assign \1348  = ~new_n421 & ~new_n422;
  assign new_n424 = ~new_n147 & new_n419;
  assign new_n425 = \176  & ~new_n424;
  assign new_n426 = ~\176  & new_n424;
  assign \1349  = new_n425 | new_n426;
  assign new_n428 = new_n286 & new_n419;
  assign new_n429 = ~\183  & ~new_n428;
  assign new_n430 = \183  & new_n428;
  assign \1350  = ~new_n429 & ~new_n430;
  assign new_n432 = ~new_n175 & new_n419;
  assign new_n433 = \190  & ~new_n432;
  assign new_n434 = ~\190  & new_n432;
  assign \1351  = new_n433 | new_n434;
  assign new_n436 = new_n110 & ~new_n232;
  assign new_n437 = new_n383 & new_n436;
  assign new_n438 = new_n308 & new_n437;
  assign new_n439 = \197  & ~new_n438;
  assign new_n440 = ~\197  & new_n438;
  assign \1352  = new_n439 | new_n440;
  assign new_n442 = ~new_n147 & new_n437;
  assign new_n443 = \204  & ~new_n442;
  assign new_n444 = ~\204  & new_n442;
  assign \1353  = new_n443 | new_n444;
  assign new_n446 = new_n286 & new_n437;
  assign new_n447 = \211  & ~new_n446;
  assign new_n448 = ~\211  & new_n446;
  assign \1354  = new_n447 | new_n448;
  assign new_n450 = ~new_n175 & new_n437;
  assign new_n451 = \218  & new_n450;
  assign new_n452 = ~\218  & ~new_n450;
  assign \1355  = ~new_n451 & ~new_n452;
endmodule


