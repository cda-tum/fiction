module c1355 ( 
    \1 , 8, 15, 22, 29, 36, 43, 50, 57, 64, 71, 78, 85, 92, 99, 106, 113,
    120, 127, 134, 141, 148, 155, 162, 169, 176, 183, 190, 197, 204, 211,
    218, 225, 226, 227, 228, 229, 230, 231, 232, 233,
    1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335,
    1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347,
    1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355  );
  input  \1 , 8, 15, 22, 29, 36, 43, 50, 57, 64, 71, 78, 85, 92, 99, 106,
    113, 120, 127, 134, 141, 148, 155, 162, 169, 176, 183, 190, 197, 204,
    211, 218, 225, 226, 227, 228, 229, 230, 231, 232, 233;
  output 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334,
    1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346,
    1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355;
  wire n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n393, n394, n395, n396, n398, n399, n400, n401, n403, n404,
    n405, n406, n408, n409, n410, n411, n412, n413, n414, n416, n417, n418,
    n419, n421, n422, n423, n424, n426, n427, n428, n429, n431, n432, n433,
    n434, n435, n436, n437, n438, n440, n441, n442, n443, n445, n446, n447,
    n448, n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461,
    n463, n464, n465, n466, n468, n469, n470, n471, n473, n474, n475, n476,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n496, n497, n498, n499, n501, n502, n503,
    n504, n506, n507, n508, n509, n511, n512, n513, n514, n515, n516, n518,
    n519, n520, n521, n523, n524, n525, n526, n528, n529, n530, n531, n533,
    n534, n535, n536, n537, n538, n539, n541, n542, n543, n544, n546, n547,
    n548, n549, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561,
    n563, n564, n565, n566, n568, n569, n570, n571, n573, n574, n575, n576;
  assign n74 = \1  & 29;
  assign n75 = \1  & ~n74;
  assign n76 = 29 & ~n74;
  assign n77 = ~n75 & ~n76;
  assign n78 = 57 & 85;
  assign n79 = 57 & ~n78;
  assign n80 = 85 & ~n78;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~n77 & ~n81;
  assign n83 = ~n77 & ~n82;
  assign n84 = ~n81 & ~n82;
  assign n85 = ~n83 & ~n84;
  assign n86 = 225 & 233;
  assign n87 = 113 & 120;
  assign n88 = 113 & ~n87;
  assign n89 = 120 & ~n87;
  assign n90 = ~n88 & ~n89;
  assign n91 = 127 & 134;
  assign n92 = 127 & ~n91;
  assign n93 = 134 & ~n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = ~n90 & ~n94;
  assign n96 = ~n90 & ~n95;
  assign n97 = ~n94 & ~n95;
  assign n98 = ~n96 & ~n97;
  assign n99 = 141 & 148;
  assign n100 = 141 & ~n99;
  assign n101 = 148 & ~n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = 155 & 162;
  assign n104 = 155 & ~n103;
  assign n105 = 162 & ~n103;
  assign n106 = ~n104 & ~n105;
  assign n107 = ~n102 & ~n106;
  assign n108 = ~n102 & ~n107;
  assign n109 = ~n106 & ~n107;
  assign n110 = ~n108 & ~n109;
  assign n111 = ~n98 & ~n110;
  assign n112 = ~n98 & ~n111;
  assign n113 = ~n110 & ~n111;
  assign n114 = ~n112 & ~n113;
  assign n115 = n86 & ~n114;
  assign n116 = n86 & ~n115;
  assign n117 = ~n114 & ~n115;
  assign n118 = ~n116 & ~n117;
  assign n119 = ~n85 & ~n118;
  assign n120 = ~n85 & ~n119;
  assign n121 = ~n118 & ~n119;
  assign n122 = ~n120 & ~n121;
  assign n123 = 113 & 141;
  assign n124 = 113 & ~n123;
  assign n125 = 141 & ~n123;
  assign n126 = ~n124 & ~n125;
  assign n127 = 169 & 197;
  assign n128 = 169 & ~n127;
  assign n129 = 197 & ~n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = ~n126 & ~n130;
  assign n132 = ~n126 & ~n131;
  assign n133 = ~n130 & ~n131;
  assign n134 = ~n132 & ~n133;
  assign n135 = 229 & 233;
  assign n136 = \1  & 8;
  assign n137 = \1  & ~n136;
  assign n138 = 8 & ~n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = 15 & 22;
  assign n141 = 15 & ~n140;
  assign n142 = 22 & ~n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = ~n139 & ~n143;
  assign n145 = ~n139 & ~n144;
  assign n146 = ~n143 & ~n144;
  assign n147 = ~n145 & ~n146;
  assign n148 = 29 & 36;
  assign n149 = 29 & ~n148;
  assign n150 = 36 & ~n148;
  assign n151 = ~n149 & ~n150;
  assign n152 = 43 & 50;
  assign n153 = 43 & ~n152;
  assign n154 = 50 & ~n152;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n151 & ~n155;
  assign n157 = ~n151 & ~n156;
  assign n158 = ~n155 & ~n156;
  assign n159 = ~n157 & ~n158;
  assign n160 = ~n147 & ~n159;
  assign n161 = ~n147 & ~n160;
  assign n162 = ~n159 & ~n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = n135 & ~n163;
  assign n165 = n135 & ~n164;
  assign n166 = ~n163 & ~n164;
  assign n167 = ~n165 & ~n166;
  assign n168 = ~n134 & ~n167;
  assign n169 = ~n134 & ~n168;
  assign n170 = ~n167 & ~n168;
  assign n171 = ~n169 & ~n170;
  assign n172 = 120 & 148;
  assign n173 = 120 & ~n172;
  assign n174 = 148 & ~n172;
  assign n175 = ~n173 & ~n174;
  assign n176 = 176 & 204;
  assign n177 = 176 & ~n176;
  assign n178 = 204 & ~n176;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~n175 & ~n180;
  assign n182 = ~n179 & ~n180;
  assign n183 = ~n181 & ~n182;
  assign n184 = 230 & 233;
  assign n185 = 57 & 64;
  assign n186 = 57 & ~n185;
  assign n187 = 64 & ~n185;
  assign n188 = ~n186 & ~n187;
  assign n189 = 71 & 78;
  assign n190 = 71 & ~n189;
  assign n191 = 78 & ~n189;
  assign n192 = ~n190 & ~n191;
  assign n193 = ~n188 & ~n192;
  assign n194 = ~n188 & ~n193;
  assign n195 = ~n192 & ~n193;
  assign n196 = ~n194 & ~n195;
  assign n197 = 85 & 92;
  assign n198 = 85 & ~n197;
  assign n199 = 92 & ~n197;
  assign n200 = ~n198 & ~n199;
  assign n201 = 99 & 106;
  assign n202 = 99 & ~n201;
  assign n203 = 106 & ~n201;
  assign n204 = ~n202 & ~n203;
  assign n205 = ~n200 & ~n204;
  assign n206 = ~n200 & ~n205;
  assign n207 = ~n204 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n196 & ~n208;
  assign n210 = ~n196 & ~n209;
  assign n211 = ~n208 & ~n209;
  assign n212 = ~n210 & ~n211;
  assign n213 = n184 & ~n212;
  assign n214 = n184 & ~n213;
  assign n215 = ~n212 & ~n213;
  assign n216 = ~n214 & ~n215;
  assign n217 = ~n183 & ~n216;
  assign n218 = ~n183 & ~n217;
  assign n219 = ~n216 & ~n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = 127 & 155;
  assign n222 = 127 & ~n221;
  assign n223 = 155 & ~n221;
  assign n224 = ~n222 & ~n223;
  assign n225 = 183 & 211;
  assign n226 = 183 & ~n225;
  assign n227 = 211 & ~n225;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n224 & ~n228;
  assign n230 = ~n224 & ~n229;
  assign n231 = ~n228 & ~n229;
  assign n232 = ~n230 & ~n231;
  assign n233 = 231 & 233;
  assign n234 = ~n147 & ~n196;
  assign n235 = ~n147 & ~n234;
  assign n236 = ~n196 & ~n234;
  assign n237 = ~n235 & ~n236;
  assign n238 = n233 & ~n237;
  assign n239 = n233 & ~n238;
  assign n240 = ~n237 & ~n238;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~n232 & ~n241;
  assign n243 = ~n232 & ~n242;
  assign n244 = ~n241 & ~n242;
  assign n245 = ~n243 & ~n244;
  assign n246 = 134 & 162;
  assign n247 = 134 & ~n246;
  assign n248 = 162 & ~n246;
  assign n249 = ~n247 & ~n248;
  assign n250 = 190 & 218;
  assign n251 = 190 & ~n250;
  assign n252 = 218 & ~n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n249 & ~n253;
  assign n255 = ~n249 & ~n254;
  assign n256 = ~n253 & ~n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = 232 & 233;
  assign n259 = ~n159 & ~n208;
  assign n260 = ~n159 & ~n259;
  assign n261 = ~n208 & ~n259;
  assign n262 = ~n260 & ~n261;
  assign n263 = n258 & ~n262;
  assign n264 = n258 & ~n263;
  assign n265 = ~n262 & ~n263;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~n257 & ~n266;
  assign n268 = ~n257 & ~n267;
  assign n269 = ~n266 & ~n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = 8 & 36;
  assign n272 = 8 & ~n271;
  assign n273 = 36 & ~n271;
  assign n274 = ~n272 & ~n273;
  assign n275 = 64 & 92;
  assign n276 = 64 & ~n275;
  assign n277 = 92 & ~n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~n274 & ~n278;
  assign n280 = ~n274 & ~n279;
  assign n281 = ~n278 & ~n279;
  assign n282 = ~n280 & ~n281;
  assign n283 = 226 & 233;
  assign n284 = 169 & 176;
  assign n285 = 169 & ~n284;
  assign n286 = 176 & ~n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = 183 & 190;
  assign n289 = 183 & ~n288;
  assign n290 = 190 & ~n288;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n287 & ~n291;
  assign n293 = ~n287 & ~n292;
  assign n294 = ~n291 & ~n292;
  assign n295 = ~n293 & ~n294;
  assign n296 = 197 & 204;
  assign n297 = 197 & ~n296;
  assign n298 = 204 & ~n296;
  assign n299 = ~n297 & ~n298;
  assign n300 = 211 & 218;
  assign n301 = 211 & ~n300;
  assign n302 = 218 & ~n300;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n299 & ~n303;
  assign n305 = ~n299 & ~n304;
  assign n306 = ~n303 & ~n304;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~n295 & ~n307;
  assign n309 = ~n295 & ~n308;
  assign n310 = ~n307 & ~n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = n283 & ~n311;
  assign n313 = n283 & ~n312;
  assign n314 = ~n311 & ~n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = ~n282 & ~n315;
  assign n317 = ~n282 & ~n316;
  assign n318 = ~n315 & ~n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = 15 & 43;
  assign n321 = 15 & ~n320;
  assign n322 = 43 & ~n320;
  assign n323 = ~n321 & ~n322;
  assign n324 = 71 & 99;
  assign n325 = 71 & ~n324;
  assign n326 = 99 & ~n324;
  assign n327 = ~n325 & ~n326;
  assign n328 = ~n323 & ~n327;
  assign n329 = ~n323 & ~n328;
  assign n330 = ~n327 & ~n328;
  assign n331 = ~n329 & ~n330;
  assign n332 = 227 & 233;
  assign n333 = ~n98 & ~n295;
  assign n334 = ~n98 & ~n333;
  assign n335 = ~n295 & ~n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = n332 & ~n336;
  assign n338 = n332 & ~n337;
  assign n339 = ~n336 & ~n337;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~n331 & ~n340;
  assign n342 = ~n331 & ~n341;
  assign n343 = ~n340 & ~n341;
  assign n344 = ~n342 & ~n343;
  assign n345 = 22 & 50;
  assign n346 = 22 & ~n345;
  assign n347 = 50 & ~n345;
  assign n348 = ~n346 & ~n347;
  assign n349 = 78 & 106;
  assign n350 = 78 & ~n349;
  assign n351 = 106 & ~n349;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~n348 & ~n352;
  assign n354 = ~n348 & ~n353;
  assign n355 = ~n352 & ~n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = 228 & 233;
  assign n358 = ~n110 & ~n307;
  assign n359 = ~n110 & ~n358;
  assign n360 = ~n307 & ~n358;
  assign n361 = ~n359 & ~n360;
  assign n362 = n357 & ~n361;
  assign n363 = n357 & ~n362;
  assign n364 = ~n361 & ~n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n356 & ~n365;
  assign n367 = ~n356 & ~n366;
  assign n368 = ~n365 & ~n366;
  assign n369 = ~n367 & ~n368;
  assign n370 = n122 & n319;
  assign n371 = n344 & n370;
  assign n372 = ~n369 & n371;
  assign n373 = ~n344 & n370;
  assign n374 = n369 & n373;
  assign n375 = n122 & ~n319;
  assign n376 = n344 & n375;
  assign n377 = n369 & n376;
  assign n378 = ~n122 & n319;
  assign n379 = n344 & n378;
  assign n380 = n369 & n379;
  assign n381 = ~n372 & ~n374;
  assign n382 = ~n377 & n381;
  assign n383 = ~n380 & n382;
  assign n384 = ~n171 & n220;
  assign n385 = ~n245 & n384;
  assign n386 = n270 & n385;
  assign n387 = ~n383 & n386;
  assign n388 = ~n122 & n387;
  assign n389 = \1  & n388;
  assign n390 = \1  & ~n389;
  assign n391 = n388 & ~n389;
  assign 1324 = n390 | n391;
  assign n393 = ~n319 & n387;
  assign n394 = 8 & n393;
  assign n395 = 8 & ~n394;
  assign n396 = n393 & ~n394;
  assign 1325 = n395 | n396;
  assign n398 = ~n344 & n387;
  assign n399 = 15 & n398;
  assign n400 = 15 & ~n399;
  assign n401 = n398 & ~n399;
  assign 1326 = n400 | n401;
  assign n403 = ~n369 & n387;
  assign n404 = 22 & n403;
  assign n405 = 22 & ~n404;
  assign n406 = n403 & ~n404;
  assign 1327 = n405 | n406;
  assign n408 = n245 & n384;
  assign n409 = ~n270 & n408;
  assign n410 = ~n383 & n409;
  assign n411 = ~n122 & n410;
  assign n412 = 29 & n411;
  assign n413 = 29 & ~n412;
  assign n414 = n411 & ~n412;
  assign 1328 = n413 | n414;
  assign n416 = ~n319 & n410;
  assign n417 = 36 & n416;
  assign n418 = 36 & ~n417;
  assign n419 = n416 & ~n417;
  assign 1329 = n418 | n419;
  assign n421 = ~n344 & n410;
  assign n422 = 43 & n421;
  assign n423 = 43 & ~n422;
  assign n424 = n421 & ~n422;
  assign 1330 = n423 | n424;
  assign n426 = ~n369 & n410;
  assign n427 = 50 & n426;
  assign n428 = 50 & ~n427;
  assign n429 = n426 & ~n427;
  assign 1331 = n428 | n429;
  assign n431 = n171 & ~n220;
  assign n432 = ~n245 & n431;
  assign n433 = n270 & n432;
  assign n434 = ~n383 & n433;
  assign n435 = ~n122 & n434;
  assign n436 = 57 & n435;
  assign n437 = 57 & ~n436;
  assign n438 = n435 & ~n436;
  assign 1332 = n437 | n438;
  assign n440 = ~n319 & n434;
  assign n441 = 64 & n440;
  assign n442 = 64 & ~n441;
  assign n443 = n440 & ~n441;
  assign 1333 = n442 | n443;
  assign n445 = ~n344 & n434;
  assign n446 = 71 & n445;
  assign n447 = 71 & ~n446;
  assign n448 = n445 & ~n446;
  assign 1334 = n447 | n448;
  assign n450 = ~n369 & n434;
  assign n451 = 78 & n450;
  assign n452 = 78 & ~n451;
  assign n453 = n450 & ~n451;
  assign 1335 = n452 | n453;
  assign n455 = n245 & n431;
  assign n456 = ~n270 & n455;
  assign n457 = ~n383 & n456;
  assign n458 = ~n122 & n457;
  assign n459 = 85 & n458;
  assign n460 = 85 & ~n459;
  assign n461 = n458 & ~n459;
  assign 1336 = n460 | n461;
  assign n463 = ~n319 & n457;
  assign n464 = 92 & n463;
  assign n465 = 92 & ~n464;
  assign n466 = n463 & ~n464;
  assign 1337 = n465 | n466;
  assign n468 = ~n344 & n457;
  assign n469 = 99 & n468;
  assign n470 = 99 & ~n469;
  assign n471 = n468 & ~n469;
  assign 1338 = n470 | n471;
  assign n473 = ~n369 & n457;
  assign n474 = 106 & n473;
  assign n475 = 106 & ~n474;
  assign n476 = n473 & ~n474;
  assign 1339 = n475 | n476;
  assign n478 = n171 & n220;
  assign n479 = n245 & n478;
  assign n480 = ~n270 & n479;
  assign n481 = ~n245 & n478;
  assign n482 = n270 & n481;
  assign n483 = n270 & n455;
  assign n484 = n270 & n408;
  assign n485 = ~n480 & ~n482;
  assign n486 = ~n483 & n485;
  assign n487 = ~n484 & n486;
  assign n488 = ~n344 & n378;
  assign n489 = n369 & n488;
  assign n490 = ~n487 & n489;
  assign n491 = ~n171 & n490;
  assign n492 = 113 & n491;
  assign n493 = 113 & ~n492;
  assign n494 = n491 & ~n492;
  assign 1340 = n493 | n494;
  assign n496 = ~n220 & n490;
  assign n497 = 120 & n496;
  assign n498 = 120 & ~n497;
  assign n499 = n496 & ~n497;
  assign 1341 = n498 | n499;
  assign n501 = ~n245 & n490;
  assign n502 = 127 & n501;
  assign n503 = 127 & ~n502;
  assign n504 = n501 & ~n502;
  assign 1342 = n503 | n504;
  assign n506 = ~n270 & n490;
  assign n507 = 134 & n506;
  assign n508 = 134 & ~n507;
  assign n509 = n506 & ~n507;
  assign 1343 = n508 | n509;
  assign n511 = ~n369 & n379;
  assign n512 = ~n487 & n511;
  assign n513 = ~n171 & n512;
  assign n514 = 141 & n513;
  assign n515 = 141 & ~n514;
  assign n516 = n513 & ~n514;
  assign 1344 = n515 | n516;
  assign n518 = ~n220 & n512;
  assign n519 = 148 & n518;
  assign n520 = 148 & ~n519;
  assign n521 = n518 & ~n519;
  assign 1345 = n520 | n521;
  assign n523 = ~n245 & n512;
  assign n524 = 155 & n523;
  assign n525 = 155 & ~n524;
  assign n526 = n523 & ~n524;
  assign 1346 = n525 | n526;
  assign n528 = ~n270 & n512;
  assign n529 = 162 & n528;
  assign n530 = 162 & ~n529;
  assign n531 = n528 & ~n529;
  assign 1347 = n530 | n531;
  assign n533 = ~n344 & n375;
  assign n534 = n369 & n533;
  assign n535 = ~n487 & n534;
  assign n536 = ~n171 & n535;
  assign n537 = 169 & n536;
  assign n538 = 169 & ~n537;
  assign n539 = n536 & ~n537;
  assign 1348 = n538 | n539;
  assign n541 = ~n220 & n535;
  assign n542 = 176 & n541;
  assign n543 = 176 & ~n542;
  assign n544 = n541 & ~n542;
  assign 1349 = n543 | n544;
  assign n546 = ~n245 & n535;
  assign n547 = 183 & n546;
  assign n548 = 183 & ~n547;
  assign n549 = n546 & ~n547;
  assign 1350 = n548 | n549;
  assign n551 = ~n270 & n535;
  assign n552 = 190 & n551;
  assign n553 = 190 & ~n552;
  assign n554 = n551 & ~n552;
  assign 1351 = n553 | n554;
  assign n556 = ~n369 & n376;
  assign n557 = ~n487 & n556;
  assign n558 = ~n171 & n557;
  assign n559 = 197 & n558;
  assign n560 = 197 & ~n559;
  assign n561 = n558 & ~n559;
  assign 1352 = n560 | n561;
  assign n563 = ~n220 & n557;
  assign n564 = 204 & n563;
  assign n565 = 204 & ~n564;
  assign n566 = n563 & ~n564;
  assign 1353 = n565 | n566;
  assign n568 = ~n245 & n557;
  assign n569 = 211 & n568;
  assign n570 = 211 & ~n569;
  assign n571 = n568 & ~n569;
  assign 1354 = n570 | n571;
  assign n573 = ~n270 & n557;
  assign n574 = 218 & n573;
  assign n575 = 218 & ~n574;
  assign n576 = n573 & ~n574;
  assign 1355 = n575 | n576;
endmodule


