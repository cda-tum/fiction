// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_, i_77_,
    i_62_, i_40_, i_120_, i_72_, i_67_, i_121_, i_71_, i_68_, i_122_,
    i_74_, i_65_, i_30_, i_123_, i_73_, i_66_, i_124_, i_94_, i_81_,
    i_125_, i_93_, i_82_, i_20_, i_126_, i_92_, i_83_, i_69_, i_9_, i_127_,
    i_91_, i_84_, i_128_, i_98_, i_85_, i_10_, i_7_, i_129_, i_97_, i_86_,
    i_79_, i_8_, i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_, i_14_,
    i_3_, i_39_, i_28_, i_13_, i_4_, i_119_, i_108_, i_25_, i_12_, i_1_,
    i_118_, i_109_, i_26_, i_11_, i_2_, i_117_, i_106_, i_90_, i_49_,
    i_23_, i_18_, i_116_, i_107_, i_24_, i_17_, i_0_, i_115_, i_104_,
    i_21_, i_16_, i_114_, i_105_, i_80_, i_59_, i_22_, i_15_, i_113_,
    i_102_, i_58_, i_45_, i_32_, i_112_, i_103_, i_57_, i_46_, i_31_,
    i_111_, i_100_, i_70_, i_56_, i_47_, i_34_, i_110_, i_101_, i_55_,
    i_48_, i_33_, i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_,
    i_52_, i_43_, i_38_, i_29_, i_51_, i_44_, i_37_,
    o_0_  );
  input  i_89_, i_76_, i_63_, i_50_, i_75_, i_64_, i_78_, i_61_, i_99_,
    i_77_, i_62_, i_40_, i_120_, i_72_, i_67_, i_121_, i_71_, i_68_,
    i_122_, i_74_, i_65_, i_30_, i_123_, i_73_, i_66_, i_124_, i_94_,
    i_81_, i_125_, i_93_, i_82_, i_20_, i_126_, i_92_, i_83_, i_69_, i_9_,
    i_127_, i_91_, i_84_, i_128_, i_98_, i_85_, i_10_, i_7_, i_129_, i_97_,
    i_86_, i_79_, i_8_, i_96_, i_87_, i_5_, i_95_, i_88_, i_6_, i_27_,
    i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_119_, i_108_, i_25_, i_12_,
    i_1_, i_118_, i_109_, i_26_, i_11_, i_2_, i_117_, i_106_, i_90_, i_49_,
    i_23_, i_18_, i_116_, i_107_, i_24_, i_17_, i_0_, i_115_, i_104_,
    i_21_, i_16_, i_114_, i_105_, i_80_, i_59_, i_22_, i_15_, i_113_,
    i_102_, i_58_, i_45_, i_32_, i_112_, i_103_, i_57_, i_46_, i_31_,
    i_111_, i_100_, i_70_, i_56_, i_47_, i_34_, i_110_, i_101_, i_55_,
    i_48_, i_33_, i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_,
    i_52_, i_43_, i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_0_;
  wire new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259;
  assign new_n132 = i_105_ & i_41_;
  assign new_n133 = i_106_ & i_42_;
  assign new_n134 = i_40_ & i_104_;
  assign new_n135 = ~new_n132 & ~new_n133;
  assign new_n136 = ~new_n134 & new_n135;
  assign new_n137 = i_108_ & i_44_;
  assign new_n138 = i_109_ & i_45_;
  assign new_n139 = i_107_ & i_43_;
  assign new_n140 = ~new_n137 & ~new_n138;
  assign new_n141 = ~new_n139 & new_n140;
  assign new_n142 = i_102_ & i_38_;
  assign new_n143 = i_39_ & i_103_;
  assign new_n144 = i_101_ & i_37_;
  assign new_n145 = ~new_n142 & ~new_n143;
  assign new_n146 = ~new_n144 & new_n145;
  assign new_n147 = new_n136 & new_n141;
  assign new_n148 = new_n146 & new_n147;
  assign new_n149 = i_50_ & i_114_;
  assign new_n150 = i_115_ & i_51_;
  assign new_n151 = i_49_ & i_113_;
  assign new_n152 = ~new_n149 & ~new_n150;
  assign new_n153 = ~new_n151 & new_n152;
  assign new_n154 = i_117_ & i_53_;
  assign new_n155 = i_118_ & i_54_;
  assign new_n156 = i_116_ & i_52_;
  assign new_n157 = ~new_n154 & ~new_n155;
  assign new_n158 = ~new_n156 & new_n157;
  assign new_n159 = i_111_ & i_47_;
  assign new_n160 = i_112_ & i_48_;
  assign new_n161 = i_46_ & i_110_;
  assign new_n162 = ~new_n159 & ~new_n160;
  assign new_n163 = ~new_n161 & new_n162;
  assign new_n164 = new_n153 & new_n158;
  assign new_n165 = new_n163 & new_n164;
  assign new_n166 = i_96_ & i_32_;
  assign new_n167 = i_97_ & i_33_;
  assign new_n168 = i_95_ & i_31_;
  assign new_n169 = ~new_n166 & ~new_n167;
  assign new_n170 = ~new_n168 & new_n169;
  assign new_n171 = i_99_ & i_35_;
  assign new_n172 = i_100_ & i_36_;
  assign new_n173 = i_98_ & i_34_;
  assign new_n174 = ~new_n171 & ~new_n172;
  assign new_n175 = ~new_n173 & new_n174;
  assign new_n176 = i_93_ & i_29_;
  assign new_n177 = i_30_ & i_94_;
  assign new_n178 = i_92_ & i_28_;
  assign new_n179 = ~new_n176 & ~new_n177;
  assign new_n180 = ~new_n178 & new_n179;
  assign new_n181 = new_n170 & new_n175;
  assign new_n182 = new_n180 & new_n181;
  assign new_n183 = new_n148 & new_n165;
  assign new_n184 = new_n182 & new_n183;
  assign new_n185 = i_129_ & i_0_;
  assign new_n186 = i_64_ & i_128_;
  assign new_n187 = ~new_n185 & ~new_n186;
  assign new_n188 = i_123_ & i_59_;
  assign new_n189 = i_124_ & i_60_;
  assign new_n190 = i_122_ & i_58_;
  assign new_n191 = ~new_n188 & ~new_n189;
  assign new_n192 = ~new_n190 & new_n191;
  assign new_n193 = i_62_ & i_126_;
  assign new_n194 = i_63_ & i_127_;
  assign new_n195 = i_61_ & i_125_;
  assign new_n196 = ~new_n193 & ~new_n194;
  assign new_n197 = ~new_n195 & new_n196;
  assign new_n198 = i_120_ & i_56_;
  assign new_n199 = i_121_ & i_57_;
  assign new_n200 = i_119_ & i_55_;
  assign new_n201 = ~new_n198 & ~new_n199;
  assign new_n202 = ~new_n200 & new_n201;
  assign new_n203 = new_n192 & new_n197;
  assign new_n204 = new_n202 & new_n203;
  assign new_n205 = new_n187 & new_n204;
  assign new_n206 = i_78_ & i_14_;
  assign new_n207 = i_79_ & i_15_;
  assign new_n208 = i_77_ & i_13_;
  assign new_n209 = ~new_n206 & ~new_n207;
  assign new_n210 = ~new_n208 & new_n209;
  assign new_n211 = i_81_ & i_17_;
  assign new_n212 = i_82_ & i_18_;
  assign new_n213 = i_16_ & i_80_;
  assign new_n214 = ~new_n211 & ~new_n212;
  assign new_n215 = ~new_n213 & new_n214;
  assign new_n216 = i_75_ & i_11_;
  assign new_n217 = i_76_ & i_12_;
  assign new_n218 = i_74_ & i_10_;
  assign new_n219 = ~new_n216 & ~new_n217;
  assign new_n220 = ~new_n218 & new_n219;
  assign new_n221 = new_n210 & new_n215;
  assign new_n222 = new_n220 & new_n221;
  assign new_n223 = i_87_ & i_23_;
  assign new_n224 = i_88_ & i_24_;
  assign new_n225 = i_86_ & i_22_;
  assign new_n226 = ~new_n223 & ~new_n224;
  assign new_n227 = ~new_n225 & new_n226;
  assign new_n228 = i_26_ & i_90_;
  assign new_n229 = i_91_ & i_27_;
  assign new_n230 = i_89_ & i_25_;
  assign new_n231 = ~new_n228 & ~new_n229;
  assign new_n232 = ~new_n230 & new_n231;
  assign new_n233 = i_20_ & i_84_;
  assign new_n234 = i_85_ & i_21_;
  assign new_n235 = i_83_ & i_19_;
  assign new_n236 = ~new_n233 & ~new_n234;
  assign new_n237 = ~new_n235 & new_n236;
  assign new_n238 = new_n227 & new_n232;
  assign new_n239 = new_n237 & new_n238;
  assign new_n240 = i_69_ & i_5_;
  assign new_n241 = i_6_ & i_70_;
  assign new_n242 = i_68_ & i_4_;
  assign new_n243 = ~new_n240 & ~new_n241;
  assign new_n244 = ~new_n242 & new_n243;
  assign new_n245 = i_72_ & i_8_;
  assign new_n246 = i_73_ & i_9_;
  assign new_n247 = i_71_ & i_7_;
  assign new_n248 = ~new_n245 & ~new_n246;
  assign new_n249 = ~new_n247 & new_n248;
  assign new_n250 = i_66_ & i_2_;
  assign new_n251 = i_67_ & i_3_;
  assign new_n252 = i_65_ & i_1_;
  assign new_n253 = ~new_n250 & ~new_n251;
  assign new_n254 = ~new_n252 & new_n253;
  assign new_n255 = new_n244 & new_n249;
  assign new_n256 = new_n254 & new_n255;
  assign new_n257 = new_n222 & new_n239;
  assign new_n258 = new_n256 & new_n257;
  assign new_n259 = new_n184 & new_n205;
  assign o_0_ = ~new_n258 | ~new_n259;
endmodule


