// Benchmark "top" written by ABC on Mon Nov 27 16:53:14 2023

module top ( 
    \1 , \18 , \35 , \52 , \69 , \86 , \103 , \120 , \137 , \154 , \171 ,
    \188 , \205 , \222 , \239 , \256 , \273 , \290 , \307 , \324 , \341 ,
    \358 , \375 , \392 , \409 , \426 , \443 , \460 , \477 , \494 , \511 ,
    \528 ,
    \545 , \1581 , \1901 , \2223 , \2548 , \2877 , \3211 , \3552 , \3895 ,
    \4241 , \4591 , \4946 , \5308 , \5672 , \5971 , \6123 , \6150 , \6160 ,
    \6170 , \6180 , \6190 , \6200 , \6210 , \6220 , \6230 , \6240 , \6250 ,
    \6260 , \6270 , \6280 , \6287 , \6288   );
  input  \1 , \18 , \35 , \52 , \69 , \86 , \103 , \120 , \137 , \154 ,
    \171 , \188 , \205 , \222 , \239 , \256 , \273 , \290 , \307 , \324 ,
    \341 , \358 , \375 , \392 , \409 , \426 , \443 , \460 , \477 , \494 ,
    \511 , \528 ;
  output \545 , \1581 , \1901 , \2223 , \2548 , \2877 , \3211 , \3552 ,
    \3895 , \4241 , \4591 , \4946 , \5308 , \5672 , \5971 , \6123 , \6150 ,
    \6160 , \6170 , \6180 , \6190 , \6200 , \6210 , \6220 , \6230 , \6240 ,
    \6250 , \6260 , \6270 , \6280 , \6287 , \6288 ;
  wire new_n66, new_n67, new_n68, new_n69, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n94, new_n95, new_n96, new_n97, new_n98,
    new_n99, new_n100, new_n101, new_n102, new_n103, new_n104, new_n105,
    new_n106, new_n107, new_n108, new_n109, new_n110, new_n111, new_n112,
    new_n113, new_n114, new_n115, new_n116, new_n117, new_n118, new_n119,
    new_n120, new_n122, new_n123, new_n124, new_n125, new_n126, new_n127,
    new_n128, new_n129, new_n130, new_n131, new_n132, new_n133, new_n134,
    new_n135, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1830, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1837, new_n1838, new_n1839, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1979, new_n1980, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2123, new_n2124, new_n2125, new_n2126, new_n2127, new_n2128,
    new_n2129, new_n2130, new_n2131, new_n2132, new_n2133, new_n2134,
    new_n2135, new_n2136, new_n2137, new_n2138, new_n2139, new_n2140,
    new_n2141, new_n2142, new_n2143, new_n2144, new_n2145, new_n2146,
    new_n2147, new_n2148, new_n2149, new_n2150, new_n2151, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2160, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165,
    new_n2166, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171,
    new_n2172, new_n2173, new_n2174, new_n2175, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187;
  assign \545  = \1  & \273 ;
  assign new_n66 = \1  & \290 ;
  assign new_n67 = \18  & \273 ;
  assign new_n68 = ~new_n66 & new_n67;
  assign new_n69 = new_n66 & ~new_n67;
  assign \1581  = new_n68 | new_n69;
  assign new_n71 = \273  & \307 ;
  assign new_n72 = ~\35  & new_n71;
  assign new_n73 = ~\273  & \307 ;
  assign new_n74 = ~\290  & new_n73;
  assign new_n75 = \273  & ~\307 ;
  assign new_n76 = \35  & new_n75;
  assign new_n77 = ~new_n72 & ~new_n74;
  assign new_n78 = ~new_n76 & new_n77;
  assign new_n79 = \1  & ~new_n78;
  assign new_n80 = \1  & \307 ;
  assign new_n81 = \18  & new_n80;
  assign new_n82 = \18  & \290 ;
  assign new_n83 = ~new_n80 & ~new_n82;
  assign new_n84 = ~\273  & ~new_n81;
  assign new_n85 = ~new_n83 & new_n84;
  assign new_n86 = \35  & \273 ;
  assign new_n87 = ~new_n82 & ~new_n86;
  assign new_n88 = \35  & \290 ;
  assign new_n89 = new_n82 & new_n88;
  assign new_n90 = ~\1  & ~new_n87;
  assign new_n91 = ~new_n89 & new_n90;
  assign new_n92 = ~new_n85 & ~new_n91;
  assign \1901  = new_n79 | ~new_n92;
  assign new_n94 = \1  & \324 ;
  assign new_n95 = \307  & ~new_n87;
  assign new_n96 = \273  & new_n82;
  assign new_n97 = ~new_n88 & new_n96;
  assign new_n98 = ~new_n95 & ~new_n97;
  assign new_n99 = \1  & ~new_n98;
  assign new_n100 = ~\273  & \290 ;
  assign new_n101 = ~\307  & new_n100;
  assign new_n102 = \35  & new_n101;
  assign new_n103 = \52  & new_n75;
  assign new_n104 = ~\273  & new_n88;
  assign new_n105 = \52  & \273 ;
  assign new_n106 = \307  & ~new_n105;
  assign new_n107 = ~new_n104 & new_n106;
  assign new_n108 = ~new_n103 & ~new_n107;
  assign new_n109 = \18  & ~new_n108;
  assign new_n110 = new_n88 & new_n105;
  assign new_n111 = ~new_n88 & ~new_n105;
  assign new_n112 = ~\18  & ~new_n110;
  assign new_n113 = ~new_n111 & new_n112;
  assign new_n114 = ~new_n102 & ~new_n113;
  assign new_n115 = ~new_n109 & new_n114;
  assign new_n116 = ~new_n99 & new_n115;
  assign new_n117 = new_n99 & ~new_n115;
  assign new_n118 = ~new_n116 & ~new_n117;
  assign new_n119 = new_n94 & ~new_n118;
  assign new_n120 = ~new_n94 & new_n118;
  assign \2223  = new_n119 | new_n120;
  assign new_n122 = \324  & ~new_n116;
  assign new_n123 = ~new_n117 & ~new_n122;
  assign new_n124 = \341  & ~new_n123;
  assign new_n125 = ~new_n103 & ~new_n111;
  assign new_n126 = ~new_n102 & new_n125;
  assign new_n127 = \324  & new_n126;
  assign new_n128 = ~\324  & ~new_n126;
  assign new_n129 = \18  & ~new_n128;
  assign new_n130 = ~new_n127 & new_n129;
  assign new_n131 = \52  & new_n101;
  assign new_n132 = \52  & \290 ;
  assign new_n133 = new_n73 & ~new_n132;
  assign new_n134 = \69  & new_n71;
  assign new_n135 = \69  & \273 ;
  assign new_n136 = ~new_n71 & ~new_n135;
  assign new_n137 = ~new_n134 & ~new_n136;
  assign new_n138 = ~new_n133 & ~new_n137;
  assign new_n139 = \35  & ~new_n138;
  assign new_n140 = ~new_n132 & ~new_n135;
  assign new_n141 = new_n132 & new_n135;
  assign new_n142 = ~\35  & ~new_n140;
  assign new_n143 = ~new_n141 & new_n142;
  assign new_n144 = ~new_n131 & ~new_n143;
  assign new_n145 = ~new_n139 & new_n144;
  assign new_n146 = ~new_n130 & new_n145;
  assign new_n147 = new_n130 & ~new_n145;
  assign new_n148 = ~new_n146 & ~new_n147;
  assign new_n149 = \1  & new_n124;
  assign new_n150 = ~\341  & new_n123;
  assign new_n151 = ~\1  & ~new_n117;
  assign new_n152 = ~new_n124 & ~new_n151;
  assign new_n153 = ~new_n150 & new_n152;
  assign new_n154 = ~new_n149 & ~new_n153;
  assign new_n155 = new_n148 & ~new_n154;
  assign new_n156 = ~new_n124 & new_n155;
  assign new_n157 = ~new_n148 & ~new_n153;
  assign \2548  = ~new_n156 & ~new_n157;
  assign new_n159 = ~new_n127 & new_n145;
  assign new_n160 = new_n129 & ~new_n159;
  assign new_n161 = \341  & new_n160;
  assign new_n162 = \18  & \341 ;
  assign new_n163 = ~new_n160 & ~new_n162;
  assign new_n164 = ~new_n161 & ~new_n163;
  assign new_n165 = \290  & \307 ;
  assign new_n166 = \273  & \290 ;
  assign new_n167 = ~\69  & new_n166;
  assign new_n168 = ~new_n165 & ~new_n167;
  assign new_n169 = \52  & ~new_n168;
  assign new_n170 = ~new_n134 & ~new_n169;
  assign new_n171 = ~\324  & new_n170;
  assign new_n172 = \35  & \324 ;
  assign new_n173 = ~new_n170 & new_n172;
  assign new_n174 = \35  & ~new_n171;
  assign new_n175 = ~new_n173 & new_n174;
  assign new_n176 = \69  & \290 ;
  assign new_n177 = \86  & \273 ;
  assign new_n178 = ~new_n176 & ~new_n177;
  assign new_n179 = new_n176 & new_n177;
  assign new_n180 = ~\52  & ~new_n178;
  assign new_n181 = ~new_n179 & new_n180;
  assign new_n182 = \69  & new_n101;
  assign new_n183 = \86  & new_n75;
  assign new_n184 = new_n73 & ~new_n176;
  assign new_n185 = ~\86  & new_n71;
  assign new_n186 = ~new_n183 & ~new_n184;
  assign new_n187 = ~new_n185 & new_n186;
  assign new_n188 = \52  & ~new_n187;
  assign new_n189 = ~new_n181 & ~new_n182;
  assign new_n190 = ~new_n188 & new_n189;
  assign new_n191 = ~new_n175 & new_n190;
  assign new_n192 = new_n175 & ~new_n190;
  assign new_n193 = ~new_n191 & ~new_n192;
  assign new_n194 = ~new_n164 & ~new_n193;
  assign new_n195 = new_n164 & new_n193;
  assign new_n196 = ~new_n194 & ~new_n195;
  assign new_n197 = ~new_n149 & ~new_n155;
  assign new_n198 = \1  & \358 ;
  assign new_n199 = new_n197 & ~new_n198;
  assign new_n200 = ~new_n197 & new_n198;
  assign new_n201 = ~new_n199 & ~new_n200;
  assign new_n202 = new_n196 & new_n201;
  assign new_n203 = ~new_n196 & ~new_n201;
  assign \2877  = ~new_n202 & ~new_n203;
  assign new_n205 = \1  & \375 ;
  assign new_n206 = ~new_n161 & ~new_n195;
  assign new_n207 = ~new_n173 & ~new_n192;
  assign new_n208 = \341  & ~new_n207;
  assign new_n209 = \35  & \341 ;
  assign new_n210 = new_n207 & ~new_n209;
  assign new_n211 = ~new_n208 & ~new_n210;
  assign new_n212 = ~new_n178 & ~new_n183;
  assign new_n213 = ~new_n182 & new_n212;
  assign new_n214 = \86  & new_n101;
  assign new_n215 = \86  & \290 ;
  assign new_n216 = new_n73 & ~new_n215;
  assign new_n217 = ~\103  & \273 ;
  assign new_n218 = \307  & new_n217;
  assign new_n219 = \103  & new_n75;
  assign new_n220 = ~new_n216 & ~new_n218;
  assign new_n221 = ~new_n219 & new_n220;
  assign new_n222 = \69  & ~new_n221;
  assign new_n223 = \103  & \290 ;
  assign new_n224 = new_n177 & new_n223;
  assign new_n225 = \103  & \273 ;
  assign new_n226 = ~new_n215 & ~new_n225;
  assign new_n227 = ~\69  & ~new_n224;
  assign new_n228 = ~new_n226 & new_n227;
  assign new_n229 = ~new_n214 & ~new_n228;
  assign new_n230 = ~new_n222 & new_n229;
  assign new_n231 = new_n213 & ~new_n230;
  assign new_n232 = ~new_n213 & new_n230;
  assign new_n233 = ~new_n231 & ~new_n232;
  assign new_n234 = ~\52  & ~new_n213;
  assign new_n235 = \52  & ~\324 ;
  assign new_n236 = ~new_n234 & ~new_n235;
  assign new_n237 = new_n233 & new_n236;
  assign new_n238 = ~new_n233 & ~new_n236;
  assign new_n239 = ~new_n237 & ~new_n238;
  assign new_n240 = ~new_n211 & new_n239;
  assign new_n241 = new_n211 & ~new_n239;
  assign new_n242 = ~new_n240 & ~new_n241;
  assign new_n243 = \18  & \358 ;
  assign new_n244 = new_n242 & ~new_n243;
  assign new_n245 = ~new_n242 & new_n243;
  assign new_n246 = ~new_n244 & ~new_n245;
  assign new_n247 = new_n206 & new_n246;
  assign new_n248 = ~new_n206 & ~new_n246;
  assign new_n249 = ~new_n247 & ~new_n248;
  assign new_n250 = ~new_n205 & new_n249;
  assign new_n251 = new_n205 & ~new_n249;
  assign new_n252 = ~new_n250 & ~new_n251;
  assign new_n253 = ~new_n200 & ~new_n202;
  assign new_n254 = new_n252 & ~new_n253;
  assign new_n255 = ~new_n252 & new_n253;
  assign \3211  = ~new_n254 & ~new_n255;
  assign new_n257 = \35  & \358 ;
  assign new_n258 = ~new_n210 & ~new_n241;
  assign new_n259 = ~new_n257 & ~new_n258;
  assign new_n260 = new_n257 & new_n258;
  assign new_n261 = ~new_n259 & ~new_n260;
  assign new_n262 = \324  & ~new_n232;
  assign new_n263 = ~new_n231 & ~new_n262;
  assign new_n264 = ~\341  & new_n263;
  assign new_n265 = \52  & ~new_n264;
  assign new_n266 = \341  & ~new_n263;
  assign new_n267 = new_n265 & ~new_n266;
  assign new_n268 = ~new_n219 & ~new_n226;
  assign new_n269 = ~new_n214 & new_n268;
  assign new_n270 = \103  & new_n101;
  assign new_n271 = ~\120  & new_n71;
  assign new_n272 = \120  & new_n75;
  assign new_n273 = ~new_n74 & ~new_n271;
  assign new_n274 = ~new_n272 & new_n273;
  assign new_n275 = \86  & ~new_n274;
  assign new_n276 = \120  & new_n166;
  assign new_n277 = \120  & \273 ;
  assign new_n278 = ~new_n223 & ~new_n277;
  assign new_n279 = ~\86  & ~new_n276;
  assign new_n280 = ~new_n278 & new_n279;
  assign new_n281 = \86  & ~new_n73;
  assign new_n282 = ~\86  & ~new_n277;
  assign new_n283 = ~\103  & ~new_n281;
  assign new_n284 = ~new_n282 & new_n283;
  assign new_n285 = ~new_n270 & ~new_n280;
  assign new_n286 = ~new_n284 & new_n285;
  assign new_n287 = ~new_n275 & new_n286;
  assign new_n288 = ~new_n269 & new_n287;
  assign new_n289 = new_n269 & ~new_n287;
  assign new_n290 = ~new_n288 & ~new_n289;
  assign new_n291 = \69  & ~\324 ;
  assign new_n292 = ~\69  & ~new_n269;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294 = new_n290 & ~new_n293;
  assign new_n295 = ~new_n290 & new_n293;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = new_n267 & new_n296;
  assign new_n298 = ~new_n267 & ~new_n296;
  assign new_n299 = ~new_n297 & ~new_n298;
  assign new_n300 = new_n261 & ~new_n299;
  assign new_n301 = ~new_n261 & new_n299;
  assign new_n302 = ~new_n300 & ~new_n301;
  assign new_n303 = ~new_n244 & ~new_n247;
  assign new_n304 = ~new_n302 & ~new_n303;
  assign new_n305 = new_n302 & new_n303;
  assign new_n306 = ~new_n304 & ~new_n305;
  assign new_n307 = \18  & \375 ;
  assign new_n308 = ~new_n306 & new_n307;
  assign new_n309 = new_n306 & ~new_n307;
  assign new_n310 = ~new_n308 & ~new_n309;
  assign new_n311 = \1  & \392 ;
  assign new_n312 = ~new_n251 & ~new_n254;
  assign new_n313 = ~new_n311 & new_n312;
  assign new_n314 = new_n311 & ~new_n312;
  assign new_n315 = ~new_n313 & ~new_n314;
  assign new_n316 = new_n310 & new_n315;
  assign new_n317 = ~new_n310 & ~new_n315;
  assign \3552  = new_n316 | new_n317;
  assign new_n319 = ~\324  & ~new_n289;
  assign new_n320 = ~new_n288 & ~new_n319;
  assign new_n321 = \341  & new_n320;
  assign new_n322 = ~\341  & ~new_n320;
  assign new_n323 = \69  & ~new_n322;
  assign new_n324 = ~new_n321 & new_n323;
  assign new_n325 = ~new_n272 & ~new_n278;
  assign new_n326 = ~new_n270 & new_n325;
  assign new_n327 = \103  & new_n73;
  assign new_n328 = \137  & new_n217;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = ~\120  & ~new_n329;
  assign new_n331 = \273  & ~\290 ;
  assign new_n332 = ~\103  & new_n331;
  assign new_n333 = ~new_n219 & ~new_n332;
  assign new_n334 = \137  & ~new_n333;
  assign new_n335 = ~\137  & \273 ;
  assign new_n336 = \307  & new_n335;
  assign new_n337 = ~new_n74 & ~new_n336;
  assign new_n338 = \103  & ~new_n337;
  assign new_n339 = \120  & \290 ;
  assign new_n340 = ~new_n225 & new_n339;
  assign new_n341 = new_n329 & new_n340;
  assign new_n342 = ~new_n330 & ~new_n334;
  assign new_n343 = ~new_n338 & ~new_n341;
  assign new_n344 = new_n342 & new_n343;
  assign new_n345 = new_n326 & ~new_n344;
  assign new_n346 = ~new_n326 & new_n344;
  assign new_n347 = ~new_n345 & ~new_n346;
  assign new_n348 = \86  & ~\324 ;
  assign new_n349 = ~\86  & ~new_n326;
  assign new_n350 = ~new_n348 & ~new_n349;
  assign new_n351 = new_n347 & ~new_n350;
  assign new_n352 = ~new_n347 & new_n350;
  assign new_n353 = ~new_n351 & ~new_n352;
  assign new_n354 = ~new_n324 & ~new_n353;
  assign new_n355 = new_n324 & new_n353;
  assign new_n356 = ~new_n354 & ~new_n355;
  assign new_n357 = new_n265 & ~new_n297;
  assign new_n358 = \358  & new_n357;
  assign new_n359 = \52  & \358 ;
  assign new_n360 = ~new_n357 & ~new_n359;
  assign new_n361 = ~new_n358 & ~new_n360;
  assign new_n362 = new_n356 & ~new_n361;
  assign new_n363 = ~new_n356 & new_n361;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = ~new_n260 & ~new_n300;
  assign new_n366 = \35  & \375 ;
  assign new_n367 = new_n365 & ~new_n366;
  assign new_n368 = \375  & ~new_n365;
  assign new_n369 = ~new_n367 & ~new_n368;
  assign new_n370 = ~new_n364 & ~new_n369;
  assign new_n371 = new_n364 & new_n369;
  assign new_n372 = ~new_n370 & ~new_n371;
  assign new_n373 = ~new_n304 & ~new_n309;
  assign new_n374 = ~new_n372 & ~new_n373;
  assign new_n375 = new_n372 & new_n373;
  assign new_n376 = ~new_n374 & ~new_n375;
  assign new_n377 = \18  & \392 ;
  assign new_n378 = ~new_n376 & new_n377;
  assign new_n379 = new_n376 & ~new_n377;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = \1  & \409 ;
  assign new_n382 = ~new_n313 & ~new_n316;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = \409  & new_n382;
  assign new_n385 = ~new_n383 & ~new_n384;
  assign new_n386 = new_n380 & new_n385;
  assign new_n387 = ~new_n380 & ~new_n385;
  assign \3895  = new_n386 | new_n387;
  assign new_n389 = new_n323 & ~new_n355;
  assign new_n390 = \358  & new_n389;
  assign new_n391 = \69  & \358 ;
  assign new_n392 = ~new_n389 & ~new_n391;
  assign new_n393 = ~new_n390 & ~new_n392;
  assign new_n394 = \103  & \324 ;
  assign new_n395 = \137  & new_n101;
  assign new_n396 = \120  & ~\154 ;
  assign new_n397 = new_n71 & new_n396;
  assign new_n398 = \137  & \290 ;
  assign new_n399 = ~\120  & \154 ;
  assign new_n400 = \273  & new_n399;
  assign new_n401 = ~new_n398 & new_n400;
  assign new_n402 = \154  & new_n75;
  assign new_n403 = new_n73 & ~new_n398;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = \120  & ~new_n404;
  assign new_n406 = \154  & \273 ;
  assign new_n407 = ~\120  & new_n398;
  assign new_n408 = ~new_n406 & new_n407;
  assign new_n409 = ~new_n395 & ~new_n397;
  assign new_n410 = ~new_n401 & ~new_n408;
  assign new_n411 = new_n409 & new_n410;
  assign new_n412 = ~new_n405 & new_n411;
  assign new_n413 = \137  & \307 ;
  assign new_n414 = new_n225 & new_n413;
  assign new_n415 = ~\307  & ~new_n335;
  assign new_n416 = \120  & new_n223;
  assign new_n417 = ~new_n415 & new_n416;
  assign new_n418 = ~new_n414 & ~new_n417;
  assign new_n419 = ~new_n412 & ~new_n418;
  assign new_n420 = new_n412 & new_n418;
  assign new_n421 = ~new_n419 & ~new_n420;
  assign new_n422 = new_n394 & ~new_n421;
  assign new_n423 = ~new_n394 & new_n421;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = ~\324  & ~new_n345;
  assign new_n426 = ~new_n346 & ~new_n425;
  assign new_n427 = ~\341  & ~new_n426;
  assign new_n428 = \341  & new_n426;
  assign new_n429 = \86  & ~new_n427;
  assign new_n430 = ~new_n428 & new_n429;
  assign new_n431 = new_n424 & new_n430;
  assign new_n432 = ~new_n424 & ~new_n430;
  assign new_n433 = ~new_n431 & ~new_n432;
  assign new_n434 = ~new_n393 & ~new_n433;
  assign new_n435 = new_n393 & new_n433;
  assign new_n436 = ~new_n434 & ~new_n435;
  assign new_n437 = ~new_n358 & ~new_n363;
  assign new_n438 = \52  & \375 ;
  assign new_n439 = new_n437 & ~new_n438;
  assign new_n440 = \375  & ~new_n437;
  assign new_n441 = ~new_n439 & ~new_n440;
  assign new_n442 = new_n436 & new_n441;
  assign new_n443 = ~new_n436 & ~new_n441;
  assign new_n444 = ~new_n442 & ~new_n443;
  assign new_n445 = \35  & \392 ;
  assign new_n446 = ~new_n368 & ~new_n371;
  assign new_n447 = ~new_n445 & new_n446;
  assign new_n448 = new_n445 & ~new_n446;
  assign new_n449 = ~new_n447 & ~new_n448;
  assign new_n450 = new_n444 & new_n449;
  assign new_n451 = ~new_n444 & ~new_n449;
  assign new_n452 = ~new_n450 & ~new_n451;
  assign new_n453 = \18  & \409 ;
  assign new_n454 = ~new_n374 & ~new_n379;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = \409  & new_n454;
  assign new_n457 = ~new_n455 & ~new_n456;
  assign new_n458 = ~new_n452 & new_n457;
  assign new_n459 = new_n452 & ~new_n457;
  assign new_n460 = ~new_n458 & ~new_n459;
  assign new_n461 = \1  & \426 ;
  assign new_n462 = ~new_n383 & ~new_n386;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = \426  & new_n462;
  assign new_n465 = ~new_n463 & ~new_n464;
  assign new_n466 = new_n460 & new_n465;
  assign new_n467 = ~new_n460 & ~new_n465;
  assign \4241  = ~new_n466 & ~new_n467;
  assign new_n469 = ~new_n447 & ~new_n450;
  assign new_n470 = \409  & new_n469;
  assign new_n471 = \35  & \409 ;
  assign new_n472 = ~new_n469 & ~new_n471;
  assign new_n473 = ~new_n470 & ~new_n472;
  assign new_n474 = \52  & \392 ;
  assign new_n475 = ~new_n439 & ~new_n442;
  assign new_n476 = ~new_n474 & ~new_n475;
  assign new_n477 = new_n474 & new_n475;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = \120  & \324 ;
  assign new_n480 = \154  & new_n101;
  assign new_n481 = ~\171  & new_n71;
  assign new_n482 = \154  & \290 ;
  assign new_n483 = new_n73 & ~new_n482;
  assign new_n484 = \171  & new_n75;
  assign new_n485 = ~new_n481 & ~new_n483;
  assign new_n486 = ~new_n484 & new_n485;
  assign new_n487 = \137  & ~new_n486;
  assign new_n488 = \171  & \273 ;
  assign new_n489 = ~new_n482 & ~new_n488;
  assign new_n490 = new_n482 & new_n488;
  assign new_n491 = ~\137  & ~new_n489;
  assign new_n492 = ~new_n490 & new_n491;
  assign new_n493 = ~new_n480 & ~new_n492;
  assign new_n494 = ~new_n487 & new_n493;
  assign new_n495 = ~new_n398 & ~new_n406;
  assign new_n496 = ~\154  & \273 ;
  assign new_n497 = ~\307  & ~new_n496;
  assign new_n498 = \120  & ~new_n495;
  assign new_n499 = ~new_n497 & new_n498;
  assign new_n500 = ~new_n494 & new_n499;
  assign new_n501 = new_n494 & ~new_n499;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = \324  & ~new_n420;
  assign new_n504 = ~new_n419 & ~new_n503;
  assign new_n505 = \341  & ~new_n504;
  assign new_n506 = ~\341  & new_n504;
  assign new_n507 = \103  & ~new_n506;
  assign new_n508 = ~new_n505 & new_n507;
  assign new_n509 = new_n502 & ~new_n508;
  assign new_n510 = ~new_n502 & new_n508;
  assign new_n511 = ~new_n509 & ~new_n510;
  assign new_n512 = new_n479 & new_n511;
  assign new_n513 = ~new_n479 & ~new_n511;
  assign new_n514 = ~new_n512 & ~new_n513;
  assign new_n515 = new_n424 & ~new_n428;
  assign new_n516 = ~new_n427 & ~new_n515;
  assign new_n517 = ~\358  & ~new_n516;
  assign new_n518 = \86  & \358 ;
  assign new_n519 = new_n516 & new_n518;
  assign new_n520 = \86  & ~new_n517;
  assign new_n521 = ~new_n519 & new_n520;
  assign new_n522 = ~new_n514 & new_n521;
  assign new_n523 = new_n514 & ~new_n521;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = ~new_n392 & ~new_n435;
  assign new_n526 = ~new_n524 & ~new_n525;
  assign new_n527 = new_n524 & new_n525;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign new_n529 = \69  & \375 ;
  assign new_n530 = new_n528 & new_n529;
  assign new_n531 = ~new_n528 & ~new_n529;
  assign new_n532 = ~new_n530 & ~new_n531;
  assign new_n533 = new_n478 & ~new_n532;
  assign new_n534 = ~new_n478 & new_n532;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536 = ~new_n473 & ~new_n535;
  assign new_n537 = new_n473 & new_n535;
  assign new_n538 = ~new_n536 & ~new_n537;
  assign new_n539 = \18  & \426 ;
  assign new_n540 = ~new_n456 & ~new_n458;
  assign new_n541 = ~new_n539 & new_n540;
  assign new_n542 = new_n539 & ~new_n540;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign new_n544 = new_n538 & new_n543;
  assign new_n545 = ~new_n538 & ~new_n543;
  assign new_n546 = ~new_n544 & ~new_n545;
  assign new_n547 = ~new_n464 & ~new_n466;
  assign new_n548 = new_n546 & new_n547;
  assign new_n549 = ~new_n546 & ~new_n547;
  assign new_n550 = ~new_n548 & ~new_n549;
  assign new_n551 = \1  & \443 ;
  assign new_n552 = ~new_n550 & new_n551;
  assign new_n553 = new_n550 & ~new_n551;
  assign \4591  = new_n552 | new_n553;
  assign new_n555 = \35  & \426 ;
  assign new_n556 = ~\324  & ~new_n500;
  assign new_n557 = ~new_n501 & ~new_n556;
  assign new_n558 = \341  & new_n557;
  assign new_n559 = ~\341  & ~new_n557;
  assign new_n560 = \120  & ~new_n559;
  assign new_n561 = ~new_n558 & new_n560;
  assign new_n562 = ~\171  & new_n166;
  assign new_n563 = ~new_n165 & ~new_n562;
  assign new_n564 = \154  & ~new_n563;
  assign new_n565 = \307  & new_n488;
  assign new_n566 = ~new_n564 & ~new_n565;
  assign new_n567 = ~\171  & \188 ;
  assign new_n568 = new_n496 & new_n567;
  assign new_n569 = ~\154  & new_n331;
  assign new_n570 = ~new_n402 & ~new_n569;
  assign new_n571 = \188  & ~new_n570;
  assign new_n572 = \154  & ~new_n101;
  assign new_n573 = ~\188  & \290 ;
  assign new_n574 = ~new_n100 & ~new_n573;
  assign new_n575 = \171  & ~new_n574;
  assign new_n576 = ~new_n572 & new_n575;
  assign new_n577 = ~\188  & new_n71;
  assign new_n578 = ~\171  & new_n73;
  assign new_n579 = ~new_n74 & ~new_n577;
  assign new_n580 = ~new_n578 & new_n579;
  assign new_n581 = \154  & ~new_n580;
  assign new_n582 = ~new_n568 & ~new_n571;
  assign new_n583 = ~new_n576 & new_n582;
  assign new_n584 = ~new_n581 & new_n583;
  assign new_n585 = ~new_n566 & ~new_n584;
  assign new_n586 = new_n566 & new_n584;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = \137  & ~\324 ;
  assign new_n589 = ~\137  & new_n566;
  assign new_n590 = ~new_n588 & ~new_n589;
  assign new_n591 = new_n587 & ~new_n590;
  assign new_n592 = ~new_n587 & new_n590;
  assign new_n593 = ~new_n591 & ~new_n592;
  assign new_n594 = new_n561 & new_n593;
  assign new_n595 = ~new_n561 & ~new_n593;
  assign new_n596 = ~new_n594 & ~new_n595;
  assign new_n597 = ~new_n505 & ~new_n514;
  assign new_n598 = new_n507 & ~new_n597;
  assign new_n599 = \358  & new_n598;
  assign new_n600 = \103  & \358 ;
  assign new_n601 = ~new_n598 & ~new_n600;
  assign new_n602 = ~new_n599 & ~new_n601;
  assign new_n603 = new_n596 & ~new_n602;
  assign new_n604 = ~new_n596 & new_n602;
  assign new_n605 = ~new_n603 & ~new_n604;
  assign new_n606 = ~new_n519 & ~new_n522;
  assign new_n607 = ~new_n605 & new_n606;
  assign new_n608 = new_n605 & ~new_n606;
  assign new_n609 = ~new_n607 & ~new_n608;
  assign new_n610 = \86  & \375 ;
  assign new_n611 = ~new_n609 & new_n610;
  assign new_n612 = new_n609 & ~new_n610;
  assign new_n613 = ~new_n611 & ~new_n612;
  assign new_n614 = \69  & \392 ;
  assign new_n615 = ~new_n527 & ~new_n530;
  assign new_n616 = ~new_n614 & new_n615;
  assign new_n617 = new_n614 & ~new_n615;
  assign new_n618 = ~new_n616 & ~new_n617;
  assign new_n619 = new_n613 & new_n618;
  assign new_n620 = ~new_n613 & ~new_n618;
  assign new_n621 = ~new_n619 & ~new_n620;
  assign new_n622 = ~new_n476 & ~new_n533;
  assign new_n623 = new_n621 & ~new_n622;
  assign new_n624 = ~new_n621 & new_n622;
  assign new_n625 = ~new_n623 & ~new_n624;
  assign new_n626 = \52  & \409 ;
  assign new_n627 = ~new_n625 & new_n626;
  assign new_n628 = new_n625 & ~new_n626;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = ~new_n472 & ~new_n537;
  assign new_n631 = ~new_n629 & new_n630;
  assign new_n632 = new_n629 & ~new_n630;
  assign new_n633 = ~new_n631 & ~new_n632;
  assign new_n634 = new_n555 & new_n633;
  assign new_n635 = ~new_n555 & ~new_n633;
  assign new_n636 = ~new_n634 & ~new_n635;
  assign new_n637 = ~new_n541 & ~new_n544;
  assign new_n638 = \443  & new_n637;
  assign new_n639 = \18  & \443 ;
  assign new_n640 = ~new_n637 & ~new_n639;
  assign new_n641 = ~new_n638 & ~new_n640;
  assign new_n642 = ~new_n636 & new_n641;
  assign new_n643 = new_n636 & ~new_n641;
  assign new_n644 = ~new_n642 & ~new_n643;
  assign new_n645 = ~new_n548 & ~new_n553;
  assign new_n646 = new_n644 & ~new_n645;
  assign new_n647 = ~new_n644 & new_n645;
  assign new_n648 = ~new_n646 & ~new_n647;
  assign new_n649 = \1  & \460 ;
  assign new_n650 = ~new_n648 & new_n649;
  assign new_n651 = new_n648 & ~new_n649;
  assign \4946  = new_n650 | new_n651;
  assign new_n653 = \18  & \460 ;
  assign new_n654 = ~new_n640 & ~new_n642;
  assign new_n655 = ~new_n653 & ~new_n654;
  assign new_n656 = new_n653 & new_n654;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign new_n658 = \52  & \426 ;
  assign new_n659 = ~new_n607 & ~new_n612;
  assign new_n660 = \324  & ~new_n586;
  assign new_n661 = ~new_n585 & ~new_n660;
  assign new_n662 = ~\341  & new_n661;
  assign new_n663 = \137  & ~new_n662;
  assign new_n664 = \341  & ~new_n661;
  assign new_n665 = new_n663 & ~new_n664;
  assign new_n666 = \188  & new_n71;
  assign new_n667 = ~\188  & new_n166;
  assign new_n668 = ~new_n165 & ~new_n667;
  assign new_n669 = \171  & ~new_n668;
  assign new_n670 = ~new_n666 & ~new_n669;
  assign new_n671 = \154  & ~new_n670;
  assign new_n672 = ~new_n331 & ~new_n667;
  assign new_n673 = ~\171  & ~new_n672;
  assign new_n674 = ~new_n484 & ~new_n673;
  assign new_n675 = \205  & ~new_n674;
  assign new_n676 = \188  & new_n165;
  assign new_n677 = new_n73 & ~new_n676;
  assign new_n678 = ~\205  & \273 ;
  assign new_n679 = \307  & new_n678;
  assign new_n680 = ~new_n677 & ~new_n679;
  assign new_n681 = \171  & ~new_n680;
  assign new_n682 = ~\205  & \290 ;
  assign new_n683 = ~new_n100 & ~new_n682;
  assign new_n684 = ~\171  & ~new_n683;
  assign new_n685 = ~new_n101 & ~new_n684;
  assign new_n686 = \188  & ~new_n685;
  assign new_n687 = ~new_n681 & ~new_n686;
  assign new_n688 = ~new_n675 & new_n687;
  assign new_n689 = new_n671 & ~new_n688;
  assign new_n690 = ~new_n671 & new_n688;
  assign new_n691 = ~new_n689 & ~new_n690;
  assign new_n692 = \154  & \324 ;
  assign new_n693 = ~new_n691 & new_n692;
  assign new_n694 = new_n691 & ~new_n692;
  assign new_n695 = ~new_n693 & ~new_n694;
  assign new_n696 = new_n665 & new_n695;
  assign new_n697 = ~new_n665 & ~new_n695;
  assign new_n698 = ~new_n696 & ~new_n697;
  assign new_n699 = new_n560 & ~new_n594;
  assign new_n700 = ~new_n698 & new_n699;
  assign new_n701 = new_n698 & ~new_n699;
  assign new_n702 = ~new_n700 & ~new_n701;
  assign new_n703 = \120  & \358 ;
  assign new_n704 = ~new_n702 & new_n703;
  assign new_n705 = new_n702 & ~new_n703;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = ~new_n599 & ~new_n604;
  assign new_n708 = \103  & \375 ;
  assign new_n709 = new_n707 & ~new_n708;
  assign new_n710 = \375  & ~new_n707;
  assign new_n711 = ~new_n709 & ~new_n710;
  assign new_n712 = ~new_n706 & ~new_n711;
  assign new_n713 = new_n706 & new_n711;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = \86  & \392 ;
  assign new_n716 = new_n714 & ~new_n715;
  assign new_n717 = ~new_n714 & new_n715;
  assign new_n718 = ~new_n716 & ~new_n717;
  assign new_n719 = new_n659 & new_n718;
  assign new_n720 = ~new_n659 & ~new_n718;
  assign new_n721 = ~new_n719 & ~new_n720;
  assign new_n722 = \69  & \409 ;
  assign new_n723 = ~new_n616 & ~new_n619;
  assign new_n724 = ~new_n722 & ~new_n723;
  assign new_n725 = \409  & new_n723;
  assign new_n726 = ~new_n724 & ~new_n725;
  assign new_n727 = new_n721 & new_n726;
  assign new_n728 = ~new_n721 & ~new_n726;
  assign new_n729 = ~new_n727 & ~new_n728;
  assign new_n730 = ~new_n623 & ~new_n628;
  assign new_n731 = ~new_n729 & ~new_n730;
  assign new_n732 = new_n729 & new_n730;
  assign new_n733 = ~new_n731 & ~new_n732;
  assign new_n734 = new_n658 & ~new_n733;
  assign new_n735 = ~new_n658 & new_n733;
  assign new_n736 = ~new_n734 & ~new_n735;
  assign new_n737 = ~new_n631 & ~new_n634;
  assign new_n738 = new_n736 & new_n737;
  assign new_n739 = ~new_n736 & ~new_n737;
  assign new_n740 = ~new_n738 & ~new_n739;
  assign new_n741 = \35  & \443 ;
  assign new_n742 = ~new_n740 & new_n741;
  assign new_n743 = new_n740 & ~new_n741;
  assign new_n744 = ~new_n742 & ~new_n743;
  assign new_n745 = ~new_n657 & new_n744;
  assign new_n746 = new_n657 & ~new_n744;
  assign new_n747 = ~new_n745 & ~new_n746;
  assign new_n748 = ~new_n646 & ~new_n651;
  assign new_n749 = ~new_n747 & ~new_n748;
  assign new_n750 = new_n747 & new_n748;
  assign new_n751 = ~new_n749 & ~new_n750;
  assign new_n752 = \1  & \477 ;
  assign new_n753 = ~new_n751 & new_n752;
  assign new_n754 = new_n751 & ~new_n752;
  assign \5308  = new_n753 | new_n754;
  assign new_n756 = \1  & \494 ;
  assign new_n757 = ~new_n749 & ~new_n754;
  assign new_n758 = ~new_n756 & ~new_n757;
  assign new_n759 = \494  & new_n757;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = \324  & ~new_n690;
  assign new_n762 = ~new_n689 & ~new_n761;
  assign new_n763 = ~\341  & new_n762;
  assign new_n764 = \154  & ~new_n763;
  assign new_n765 = \341  & ~new_n762;
  assign new_n766 = new_n764 & ~new_n765;
  assign new_n767 = \188  & ~\205 ;
  assign new_n768 = new_n166 & new_n767;
  assign new_n769 = \205  & new_n71;
  assign new_n770 = ~new_n676 & ~new_n768;
  assign new_n771 = ~new_n769 & new_n770;
  assign new_n772 = \205  & ~\222 ;
  assign new_n773 = new_n573 & new_n772;
  assign new_n774 = \222  & new_n75;
  assign new_n775 = ~new_n74 & ~new_n774;
  assign new_n776 = \188  & ~new_n775;
  assign new_n777 = ~\222  & new_n666;
  assign new_n778 = new_n73 & new_n767;
  assign new_n779 = ~new_n331 & ~new_n678;
  assign new_n780 = ~\188  & \222 ;
  assign new_n781 = ~new_n779 & new_n780;
  assign new_n782 = \205  & new_n100;
  assign new_n783 = ~new_n676 & new_n782;
  assign new_n784 = ~new_n773 & ~new_n778;
  assign new_n785 = ~new_n777 & new_n784;
  assign new_n786 = ~new_n781 & ~new_n783;
  assign new_n787 = new_n785 & new_n786;
  assign new_n788 = ~new_n776 & new_n787;
  assign new_n789 = new_n771 & new_n788;
  assign new_n790 = ~new_n771 & ~new_n788;
  assign new_n791 = ~new_n789 & ~new_n790;
  assign new_n792 = \171  & ~\324 ;
  assign new_n793 = ~\171  & new_n771;
  assign new_n794 = ~new_n792 & ~new_n793;
  assign new_n795 = new_n791 & ~new_n794;
  assign new_n796 = ~new_n791 & new_n794;
  assign new_n797 = ~new_n795 & ~new_n796;
  assign new_n798 = new_n766 & new_n797;
  assign new_n799 = ~new_n766 & ~new_n797;
  assign new_n800 = ~new_n798 & ~new_n799;
  assign new_n801 = new_n663 & ~new_n696;
  assign new_n802 = \358  & new_n801;
  assign new_n803 = \137  & \358 ;
  assign new_n804 = ~new_n801 & ~new_n803;
  assign new_n805 = ~new_n802 & ~new_n804;
  assign new_n806 = new_n800 & ~new_n805;
  assign new_n807 = ~new_n800 & new_n805;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = ~new_n701 & ~new_n705;
  assign new_n810 = ~new_n808 & ~new_n809;
  assign new_n811 = new_n808 & new_n809;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = \120  & \375 ;
  assign new_n814 = ~new_n812 & new_n813;
  assign new_n815 = new_n812 & ~new_n813;
  assign new_n816 = ~new_n814 & ~new_n815;
  assign new_n817 = \103  & \392 ;
  assign new_n818 = ~new_n709 & ~new_n713;
  assign new_n819 = ~new_n817 & ~new_n818;
  assign new_n820 = new_n817 & new_n818;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = new_n816 & new_n821;
  assign new_n823 = ~new_n816 & ~new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = ~new_n717 & ~new_n719;
  assign new_n826 = new_n824 & new_n825;
  assign new_n827 = ~new_n824 & ~new_n825;
  assign new_n828 = ~new_n826 & ~new_n827;
  assign new_n829 = \86  & \409 ;
  assign new_n830 = ~new_n828 & new_n829;
  assign new_n831 = new_n828 & ~new_n829;
  assign new_n832 = ~new_n830 & ~new_n831;
  assign new_n833 = \69  & \426 ;
  assign new_n834 = new_n832 & ~new_n833;
  assign new_n835 = ~new_n832 & new_n833;
  assign new_n836 = ~new_n834 & ~new_n835;
  assign new_n837 = ~new_n725 & ~new_n727;
  assign new_n838 = new_n836 & new_n837;
  assign new_n839 = ~new_n836 & ~new_n837;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = \52  & \443 ;
  assign new_n842 = ~new_n732 & ~new_n841;
  assign new_n843 = ~new_n731 & new_n841;
  assign new_n844 = ~new_n735 & new_n843;
  assign new_n845 = ~new_n842 & ~new_n844;
  assign new_n846 = ~\443  & new_n658;
  assign new_n847 = ~new_n731 & new_n846;
  assign new_n848 = ~new_n845 & ~new_n847;
  assign new_n849 = new_n840 & new_n848;
  assign new_n850 = ~new_n840 & ~new_n848;
  assign new_n851 = ~new_n849 & ~new_n850;
  assign new_n852 = ~new_n738 & ~new_n743;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = new_n851 & new_n852;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign new_n856 = \35  & \460 ;
  assign new_n857 = ~new_n855 & new_n856;
  assign new_n858 = new_n855 & ~new_n856;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = ~new_n656 & ~new_n746;
  assign new_n861 = new_n859 & new_n860;
  assign new_n862 = ~new_n859 & ~new_n860;
  assign new_n863 = ~new_n861 & ~new_n862;
  assign new_n864 = \18  & \477 ;
  assign new_n865 = new_n863 & new_n864;
  assign new_n866 = ~new_n863 & ~new_n864;
  assign new_n867 = ~new_n865 & ~new_n866;
  assign new_n868 = ~new_n760 & new_n867;
  assign new_n869 = new_n760 & ~new_n867;
  assign \5672  = new_n868 | new_n869;
  assign new_n871 = \35  & \477 ;
  assign new_n872 = \52  & \460 ;
  assign new_n873 = ~new_n844 & ~new_n850;
  assign new_n874 = ~new_n872 & new_n873;
  assign new_n875 = new_n872 & ~new_n873;
  assign new_n876 = ~new_n874 & ~new_n875;
  assign new_n877 = \120  & \392 ;
  assign new_n878 = ~new_n810 & ~new_n815;
  assign new_n879 = ~new_n877 & ~new_n878;
  assign new_n880 = new_n877 & new_n878;
  assign new_n881 = ~new_n879 & ~new_n880;
  assign new_n882 = \188  & \324 ;
  assign new_n883 = \205  & new_n165;
  assign new_n884 = \222  & new_n71;
  assign new_n885 = new_n166 & new_n772;
  assign new_n886 = ~new_n883 & ~new_n884;
  assign new_n887 = ~new_n885 & new_n886;
  assign new_n888 = \188  & ~new_n887;
  assign new_n889 = new_n73 & new_n772;
  assign new_n890 = \205  & new_n75;
  assign new_n891 = \222  & \290 ;
  assign new_n892 = new_n678 & ~new_n891;
  assign new_n893 = ~new_n890 & ~new_n892;
  assign new_n894 = \239  & ~new_n893;
  assign new_n895 = ~\239  & new_n71;
  assign new_n896 = ~new_n74 & ~new_n895;
  assign new_n897 = \205  & ~new_n896;
  assign new_n898 = ~\205  & ~\239 ;
  assign new_n899 = new_n891 & new_n898;
  assign new_n900 = \222  & new_n100;
  assign new_n901 = ~new_n883 & new_n900;
  assign new_n902 = ~new_n889 & ~new_n899;
  assign new_n903 = ~new_n901 & new_n902;
  assign new_n904 = ~new_n894 & new_n903;
  assign new_n905 = ~new_n897 & new_n904;
  assign new_n906 = new_n888 & ~new_n905;
  assign new_n907 = ~new_n888 & new_n905;
  assign new_n908 = ~new_n906 & ~new_n907;
  assign new_n909 = new_n882 & ~new_n908;
  assign new_n910 = ~new_n882 & new_n908;
  assign new_n911 = ~new_n909 & ~new_n910;
  assign new_n912 = \324  & ~new_n789;
  assign new_n913 = ~new_n790 & ~new_n912;
  assign new_n914 = \171  & ~new_n913;
  assign new_n915 = \341  & new_n914;
  assign new_n916 = ~\341  & new_n913;
  assign new_n917 = \171  & ~new_n916;
  assign new_n918 = ~new_n915 & new_n917;
  assign new_n919 = new_n911 & new_n918;
  assign new_n920 = ~new_n911 & ~new_n918;
  assign new_n921 = ~new_n919 & ~new_n920;
  assign new_n922 = new_n764 & ~new_n798;
  assign new_n923 = ~\358  & ~new_n922;
  assign new_n924 = \358  & new_n922;
  assign new_n925 = \154  & ~new_n923;
  assign new_n926 = ~new_n924 & new_n925;
  assign new_n927 = ~new_n921 & ~new_n926;
  assign new_n928 = new_n921 & new_n926;
  assign new_n929 = ~new_n927 & ~new_n928;
  assign new_n930 = ~new_n802 & ~new_n807;
  assign new_n931 = \137  & \375 ;
  assign new_n932 = new_n930 & ~new_n931;
  assign new_n933 = \375  & ~new_n930;
  assign new_n934 = ~new_n932 & ~new_n933;
  assign new_n935 = new_n929 & new_n934;
  assign new_n936 = ~new_n929 & ~new_n934;
  assign new_n937 = ~new_n935 & ~new_n936;
  assign new_n938 = ~new_n881 & new_n937;
  assign new_n939 = new_n881 & ~new_n937;
  assign new_n940 = ~new_n938 & ~new_n939;
  assign new_n941 = ~new_n819 & ~new_n822;
  assign new_n942 = ~new_n940 & ~new_n941;
  assign new_n943 = new_n940 & new_n941;
  assign new_n944 = ~new_n942 & ~new_n943;
  assign new_n945 = \103  & \409 ;
  assign new_n946 = ~new_n944 & new_n945;
  assign new_n947 = new_n944 & ~new_n945;
  assign new_n948 = ~new_n946 & ~new_n947;
  assign new_n949 = ~new_n826 & ~new_n831;
  assign new_n950 = new_n948 & ~new_n949;
  assign new_n951 = ~new_n948 & new_n949;
  assign new_n952 = ~new_n950 & ~new_n951;
  assign new_n953 = \86  & \426 ;
  assign new_n954 = ~new_n952 & new_n953;
  assign new_n955 = new_n952 & ~new_n953;
  assign new_n956 = ~new_n954 & ~new_n955;
  assign new_n957 = \69  & \443 ;
  assign new_n958 = ~new_n834 & ~new_n838;
  assign new_n959 = ~new_n957 & ~new_n958;
  assign new_n960 = new_n957 & new_n958;
  assign new_n961 = ~new_n959 & ~new_n960;
  assign new_n962 = new_n956 & new_n961;
  assign new_n963 = ~new_n956 & ~new_n961;
  assign new_n964 = ~new_n962 & ~new_n963;
  assign new_n965 = ~new_n876 & ~new_n964;
  assign new_n966 = new_n876 & new_n964;
  assign new_n967 = ~new_n965 & ~new_n966;
  assign new_n968 = ~new_n853 & ~new_n858;
  assign new_n969 = new_n967 & ~new_n968;
  assign new_n970 = ~new_n967 & new_n968;
  assign new_n971 = ~new_n969 & ~new_n970;
  assign new_n972 = new_n871 & ~new_n971;
  assign new_n973 = ~new_n871 & new_n971;
  assign new_n974 = ~new_n972 & ~new_n973;
  assign new_n975 = ~new_n862 & ~new_n865;
  assign new_n976 = new_n974 & new_n975;
  assign new_n977 = ~new_n974 & ~new_n975;
  assign new_n978 = ~new_n976 & ~new_n977;
  assign new_n979 = \18  & \494 ;
  assign new_n980 = ~new_n978 & new_n979;
  assign new_n981 = new_n978 & ~new_n979;
  assign new_n982 = ~new_n980 & ~new_n981;
  assign new_n983 = ~new_n758 & ~new_n869;
  assign new_n984 = new_n982 & ~new_n983;
  assign new_n985 = ~new_n982 & new_n983;
  assign new_n986 = ~new_n984 & ~new_n985;
  assign new_n987 = \1  & \511 ;
  assign new_n988 = new_n986 & new_n987;
  assign new_n989 = ~new_n986 & ~new_n987;
  assign \5971  = ~new_n988 & ~new_n989;
  assign new_n991 = \1  & \528 ;
  assign new_n992 = ~new_n985 & ~new_n988;
  assign new_n993 = ~new_n991 & new_n992;
  assign new_n994 = new_n991 & ~new_n992;
  assign new_n995 = ~new_n993 & ~new_n994;
  assign new_n996 = ~new_n874 & ~new_n966;
  assign new_n997 = \69  & \460 ;
  assign new_n998 = ~new_n959 & ~new_n962;
  assign new_n999 = ~new_n997 & ~new_n998;
  assign new_n1000 = new_n997 & new_n998;
  assign new_n1001 = ~new_n999 & ~new_n1000;
  assign new_n1002 = \86  & \443 ;
  assign new_n1003 = \205  & \324 ;
  assign new_n1004 = \239  & new_n769;
  assign new_n1005 = ~\307  & ~new_n166;
  assign new_n1006 = ~\239  & ~\307 ;
  assign new_n1007 = ~new_n165 & ~new_n1006;
  assign new_n1008 = ~new_n1005 & new_n1007;
  assign new_n1009 = \205  & \222 ;
  assign new_n1010 = ~new_n1005 & new_n1009;
  assign new_n1011 = ~new_n1008 & new_n1010;
  assign new_n1012 = ~new_n1004 & ~new_n1011;
  assign new_n1013 = ~new_n1003 & new_n1012;
  assign new_n1014 = \324  & ~new_n1012;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = \239  & new_n101;
  assign new_n1017 = ~\256  & new_n71;
  assign new_n1018 = \256  & new_n75;
  assign new_n1019 = ~new_n74 & ~new_n1017;
  assign new_n1020 = ~new_n1018 & new_n1019;
  assign new_n1021 = \222  & ~new_n1020;
  assign new_n1022 = \256  & new_n166;
  assign new_n1023 = \256  & \273 ;
  assign new_n1024 = \239  & \290 ;
  assign new_n1025 = ~new_n1023 & ~new_n1024;
  assign new_n1026 = ~\222  & ~new_n1022;
  assign new_n1027 = ~new_n1025 & new_n1026;
  assign new_n1028 = \222  & ~new_n73;
  assign new_n1029 = ~\222  & ~new_n1023;
  assign new_n1030 = ~\239  & ~new_n1028;
  assign new_n1031 = ~new_n1029 & new_n1030;
  assign new_n1032 = ~new_n1016 & ~new_n1027;
  assign new_n1033 = ~new_n1031 & new_n1032;
  assign new_n1034 = ~new_n1021 & new_n1033;
  assign new_n1035 = ~new_n1015 & new_n1034;
  assign new_n1036 = new_n1015 & ~new_n1034;
  assign new_n1037 = ~new_n1035 & ~new_n1036;
  assign new_n1038 = \324  & ~new_n907;
  assign new_n1039 = ~new_n906 & ~new_n1038;
  assign new_n1040 = \341  & ~new_n1039;
  assign new_n1041 = ~\341  & new_n1039;
  assign new_n1042 = \188  & ~new_n1041;
  assign new_n1043 = ~new_n1040 & new_n1042;
  assign new_n1044 = new_n1037 & ~new_n1043;
  assign new_n1045 = ~new_n1037 & new_n1043;
  assign new_n1046 = ~new_n1044 & ~new_n1045;
  assign new_n1047 = ~\341  & ~new_n914;
  assign new_n1048 = ~new_n911 & ~new_n1047;
  assign new_n1049 = ~new_n915 & ~new_n1048;
  assign new_n1050 = \358  & ~new_n1049;
  assign new_n1051 = ~\358  & new_n1049;
  assign new_n1052 = \171  & ~new_n1051;
  assign new_n1053 = ~new_n1050 & new_n1052;
  assign new_n1054 = new_n1046 & new_n1053;
  assign new_n1055 = ~new_n1046 & ~new_n1053;
  assign new_n1056 = ~new_n1054 & ~new_n1055;
  assign new_n1057 = \154  & \375 ;
  assign new_n1058 = ~new_n921 & ~new_n923;
  assign new_n1059 = ~new_n924 & ~new_n1058;
  assign new_n1060 = ~new_n1057 & new_n1059;
  assign new_n1061 = new_n1057 & ~new_n1059;
  assign new_n1062 = \154  & ~new_n1060;
  assign new_n1063 = ~new_n1061 & new_n1062;
  assign new_n1064 = ~new_n1056 & new_n1063;
  assign new_n1065 = new_n1056 & ~new_n1063;
  assign new_n1066 = ~new_n1064 & ~new_n1065;
  assign new_n1067 = ~new_n932 & ~new_n935;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n1066 & new_n1067;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = \137  & \392 ;
  assign new_n1072 = ~new_n1070 & new_n1071;
  assign new_n1073 = new_n1070 & ~new_n1071;
  assign new_n1074 = ~new_n1072 & ~new_n1073;
  assign new_n1075 = ~new_n880 & ~new_n939;
  assign new_n1076 = new_n1074 & new_n1075;
  assign new_n1077 = ~new_n1074 & ~new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = \120  & \409 ;
  assign new_n1080 = ~new_n1078 & new_n1079;
  assign new_n1081 = new_n1078 & ~new_n1079;
  assign new_n1082 = ~new_n1080 & ~new_n1081;
  assign new_n1083 = ~new_n942 & ~new_n947;
  assign new_n1084 = \103  & \426 ;
  assign new_n1085 = ~new_n1083 & ~new_n1084;
  assign new_n1086 = \426  & new_n1083;
  assign new_n1087 = ~new_n1085 & ~new_n1086;
  assign new_n1088 = new_n1082 & new_n1087;
  assign new_n1089 = ~new_n1082 & ~new_n1087;
  assign new_n1090 = ~new_n1088 & ~new_n1089;
  assign new_n1091 = ~new_n950 & ~new_n955;
  assign new_n1092 = ~new_n1090 & new_n1091;
  assign new_n1093 = new_n1090 & ~new_n1091;
  assign new_n1094 = ~new_n1092 & ~new_n1093;
  assign new_n1095 = new_n1002 & new_n1094;
  assign new_n1096 = ~new_n1002 & ~new_n1094;
  assign new_n1097 = ~new_n1095 & ~new_n1096;
  assign new_n1098 = ~new_n1001 & new_n1097;
  assign new_n1099 = new_n1001 & ~new_n1097;
  assign new_n1100 = ~new_n1098 & ~new_n1099;
  assign new_n1101 = \52  & \477 ;
  assign new_n1102 = new_n1100 & ~new_n1101;
  assign new_n1103 = ~new_n1100 & new_n1101;
  assign new_n1104 = ~new_n1102 & ~new_n1103;
  assign new_n1105 = new_n996 & new_n1104;
  assign new_n1106 = ~new_n996 & ~new_n1104;
  assign new_n1107 = ~new_n1105 & ~new_n1106;
  assign new_n1108 = \35  & \494 ;
  assign new_n1109 = ~new_n969 & ~new_n973;
  assign new_n1110 = ~new_n1108 & ~new_n1109;
  assign new_n1111 = \494  & new_n1109;
  assign new_n1112 = ~new_n1110 & ~new_n1111;
  assign new_n1113 = new_n1107 & new_n1112;
  assign new_n1114 = ~new_n1107 & ~new_n1112;
  assign new_n1115 = ~new_n1113 & ~new_n1114;
  assign new_n1116 = ~new_n976 & ~new_n981;
  assign new_n1117 = ~\511  & new_n1116;
  assign new_n1118 = \18  & \511 ;
  assign new_n1119 = ~new_n1116 & new_n1118;
  assign new_n1120 = ~new_n1117 & ~new_n1119;
  assign new_n1121 = new_n1115 & ~new_n1120;
  assign new_n1122 = ~new_n1115 & new_n1120;
  assign new_n1123 = ~new_n1121 & ~new_n1122;
  assign new_n1124 = new_n995 & new_n1123;
  assign new_n1125 = ~new_n995 & ~new_n1123;
  assign \6123  = ~new_n1124 & ~new_n1125;
  assign new_n1127 = ~new_n994 & ~new_n1124;
  assign new_n1128 = \69  & \477 ;
  assign new_n1129 = ~new_n1061 & ~new_n1064;
  assign new_n1130 = \392  & ~new_n1129;
  assign new_n1131 = \154  & \392 ;
  assign new_n1132 = new_n1129 & ~new_n1131;
  assign new_n1133 = ~new_n1130 & ~new_n1132;
  assign new_n1134 = new_n1052 & ~new_n1054;
  assign new_n1135 = \171  & \375 ;
  assign new_n1136 = ~new_n1018 & ~new_n1025;
  assign new_n1137 = ~new_n1016 & new_n1136;
  assign new_n1138 = \324  & new_n1137;
  assign new_n1139 = ~\324  & ~new_n1137;
  assign new_n1140 = \222  & ~new_n1138;
  assign new_n1141 = ~new_n1139 & new_n1140;
  assign new_n1142 = \239  & \307 ;
  assign new_n1143 = \256  & \290 ;
  assign new_n1144 = new_n1142 & ~new_n1143;
  assign new_n1145 = \256  & new_n101;
  assign new_n1146 = \239  & ~new_n71;
  assign new_n1147 = new_n1143 & ~new_n1146;
  assign new_n1148 = ~new_n1144 & ~new_n1145;
  assign new_n1149 = ~new_n1147 & new_n1148;
  assign new_n1150 = ~new_n1141 & new_n1149;
  assign new_n1151 = new_n1141 & ~new_n1149;
  assign new_n1152 = ~new_n1150 & ~new_n1151;
  assign new_n1153 = ~new_n1012 & ~new_n1034;
  assign new_n1154 = \205  & \341 ;
  assign new_n1155 = ~new_n1153 & ~new_n1154;
  assign new_n1156 = ~new_n1014 & ~new_n1036;
  assign new_n1157 = \341  & ~new_n1156;
  assign new_n1158 = ~new_n1155 & ~new_n1157;
  assign new_n1159 = \205  & ~new_n1034;
  assign new_n1160 = new_n1012 & ~new_n1159;
  assign new_n1161 = \324  & ~\341 ;
  assign new_n1162 = ~new_n1160 & new_n1161;
  assign new_n1163 = ~new_n1158 & ~new_n1162;
  assign new_n1164 = new_n1152 & new_n1163;
  assign new_n1165 = ~new_n1152 & ~new_n1163;
  assign new_n1166 = ~new_n1164 & ~new_n1165;
  assign new_n1167 = new_n1042 & ~new_n1045;
  assign new_n1168 = new_n1166 & ~new_n1167;
  assign new_n1169 = ~new_n1166 & new_n1167;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = \188  & \358 ;
  assign new_n1172 = new_n1170 & ~new_n1171;
  assign new_n1173 = ~new_n1170 & new_n1171;
  assign new_n1174 = ~new_n1172 & ~new_n1173;
  assign new_n1175 = new_n1135 & new_n1174;
  assign new_n1176 = ~new_n1135 & ~new_n1174;
  assign new_n1177 = ~new_n1175 & ~new_n1176;
  assign new_n1178 = new_n1134 & ~new_n1177;
  assign new_n1179 = ~new_n1134 & new_n1177;
  assign new_n1180 = ~new_n1178 & ~new_n1179;
  assign new_n1181 = ~new_n1133 & ~new_n1180;
  assign new_n1182 = new_n1133 & new_n1180;
  assign new_n1183 = ~new_n1181 & ~new_n1182;
  assign new_n1184 = ~new_n1068 & ~new_n1073;
  assign new_n1185 = ~new_n1183 & ~new_n1184;
  assign new_n1186 = new_n1183 & new_n1184;
  assign new_n1187 = ~new_n1185 & ~new_n1186;
  assign new_n1188 = \137  & \409 ;
  assign new_n1189 = ~new_n1187 & new_n1188;
  assign new_n1190 = new_n1187 & ~new_n1188;
  assign new_n1191 = ~new_n1189 & ~new_n1190;
  assign new_n1192 = \120  & \426 ;
  assign new_n1193 = ~new_n1076 & ~new_n1081;
  assign new_n1194 = ~new_n1192 & ~new_n1193;
  assign new_n1195 = \426  & new_n1193;
  assign new_n1196 = ~new_n1194 & ~new_n1195;
  assign new_n1197 = new_n1191 & ~new_n1196;
  assign new_n1198 = ~new_n1191 & new_n1196;
  assign new_n1199 = ~new_n1197 & ~new_n1198;
  assign new_n1200 = \103  & \443 ;
  assign new_n1201 = ~new_n1085 & ~new_n1088;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign new_n1203 = \443  & new_n1201;
  assign new_n1204 = ~new_n1202 & ~new_n1203;
  assign new_n1205 = new_n1199 & new_n1204;
  assign new_n1206 = ~new_n1199 & ~new_n1204;
  assign new_n1207 = ~new_n1205 & ~new_n1206;
  assign new_n1208 = ~new_n1092 & ~new_n1095;
  assign new_n1209 = new_n1207 & ~new_n1208;
  assign new_n1210 = ~new_n1207 & new_n1208;
  assign new_n1211 = ~new_n1209 & ~new_n1210;
  assign new_n1212 = \86  & \460 ;
  assign new_n1213 = ~new_n1211 & new_n1212;
  assign new_n1214 = new_n1211 & ~new_n1212;
  assign new_n1215 = ~new_n1213 & ~new_n1214;
  assign new_n1216 = ~new_n999 & ~new_n1099;
  assign new_n1217 = ~new_n1215 & new_n1216;
  assign new_n1218 = new_n1215 & ~new_n1216;
  assign new_n1219 = ~new_n1217 & ~new_n1218;
  assign new_n1220 = new_n1128 & new_n1219;
  assign new_n1221 = ~new_n1128 & ~new_n1219;
  assign new_n1222 = ~new_n1220 & ~new_n1221;
  assign new_n1223 = ~new_n1103 & ~new_n1105;
  assign new_n1224 = new_n1222 & ~new_n1223;
  assign new_n1225 = ~new_n1222 & new_n1223;
  assign new_n1226 = ~new_n1224 & ~new_n1225;
  assign new_n1227 = \52  & \494 ;
  assign new_n1228 = ~new_n1226 & new_n1227;
  assign new_n1229 = new_n1226 & ~new_n1227;
  assign new_n1230 = ~new_n1228 & ~new_n1229;
  assign new_n1231 = ~new_n1111 & ~new_n1113;
  assign new_n1232 = new_n1230 & new_n1231;
  assign new_n1233 = ~new_n1230 & ~new_n1231;
  assign new_n1234 = ~new_n1232 & ~new_n1233;
  assign new_n1235 = \35  & \511 ;
  assign new_n1236 = ~new_n1234 & new_n1235;
  assign new_n1237 = new_n1234 & ~new_n1235;
  assign new_n1238 = ~new_n1236 & ~new_n1237;
  assign new_n1239 = ~\511  & ~new_n1115;
  assign new_n1240 = new_n1116 & ~new_n1239;
  assign new_n1241 = \511  & new_n1115;
  assign new_n1242 = ~\528  & ~new_n1241;
  assign new_n1243 = \18  & ~new_n1242;
  assign new_n1244 = ~new_n1240 & ~new_n1243;
  assign new_n1245 = \18  & new_n1240;
  assign new_n1246 = ~new_n1116 & new_n1241;
  assign new_n1247 = ~new_n1245 & ~new_n1246;
  assign new_n1248 = \528  & ~new_n1247;
  assign new_n1249 = ~new_n1244 & ~new_n1248;
  assign new_n1250 = new_n1238 & new_n1249;
  assign new_n1251 = ~new_n1238 & ~new_n1249;
  assign new_n1252 = ~new_n1250 & ~new_n1251;
  assign new_n1253 = ~new_n1127 & ~new_n1252;
  assign new_n1254 = new_n1127 & new_n1252;
  assign \6150  = ~new_n1253 & ~new_n1254;
  assign new_n1256 = \35  & \528 ;
  assign new_n1257 = ~new_n1138 & new_n1149;
  assign new_n1258 = ~new_n1139 & ~new_n1257;
  assign new_n1259 = ~\341  & ~new_n1258;
  assign new_n1260 = \341  & new_n1258;
  assign new_n1261 = \222  & ~new_n1259;
  assign new_n1262 = ~new_n1260 & new_n1261;
  assign new_n1263 = \256  & ~\324 ;
  assign new_n1264 = new_n1008 & new_n1263;
  assign new_n1265 = \239  & \256 ;
  assign new_n1266 = \324  & new_n1265;
  assign new_n1267 = ~new_n1005 & new_n1266;
  assign new_n1268 = \239  & ~new_n1267;
  assign new_n1269 = \324  & new_n1268;
  assign new_n1270 = ~\239  & \256 ;
  assign new_n1271 = \324  & new_n1143;
  assign new_n1272 = ~new_n1270 & ~new_n1271;
  assign new_n1273 = \307  & ~new_n1272;
  assign new_n1274 = ~new_n1264 & ~new_n1273;
  assign new_n1275 = ~new_n1269 & new_n1274;
  assign new_n1276 = ~new_n1262 & new_n1275;
  assign new_n1277 = new_n1262 & ~new_n1275;
  assign new_n1278 = ~new_n1276 & ~new_n1277;
  assign new_n1279 = ~new_n1154 & new_n1156;
  assign new_n1280 = ~new_n1165 & ~new_n1279;
  assign new_n1281 = ~new_n1278 & ~new_n1280;
  assign new_n1282 = new_n1278 & new_n1280;
  assign new_n1283 = ~new_n1281 & ~new_n1282;
  assign new_n1284 = \205  & \358 ;
  assign new_n1285 = ~new_n1283 & new_n1284;
  assign new_n1286 = new_n1283 & ~new_n1284;
  assign new_n1287 = ~new_n1285 & ~new_n1286;
  assign new_n1288 = ~new_n1168 & ~new_n1172;
  assign new_n1289 = \188  & \375 ;
  assign new_n1290 = ~new_n1288 & ~new_n1289;
  assign new_n1291 = \375  & new_n1288;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = new_n1287 & new_n1292;
  assign new_n1294 = ~new_n1287 & ~new_n1292;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = \171  & \392 ;
  assign new_n1297 = new_n1295 & ~new_n1296;
  assign new_n1298 = ~new_n1295 & new_n1296;
  assign new_n1299 = ~new_n1297 & ~new_n1298;
  assign new_n1300 = new_n1135 & ~new_n1174;
  assign new_n1301 = ~new_n1178 & ~new_n1300;
  assign new_n1302 = new_n1299 & new_n1301;
  assign new_n1303 = ~new_n1299 & ~new_n1301;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = ~new_n1130 & ~new_n1182;
  assign new_n1306 = \409  & ~new_n1305;
  assign new_n1307 = \154  & \409 ;
  assign new_n1308 = new_n1305 & ~new_n1307;
  assign new_n1309 = ~new_n1306 & ~new_n1308;
  assign new_n1310 = ~new_n1304 & new_n1309;
  assign new_n1311 = new_n1304 & ~new_n1309;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = ~new_n1185 & ~new_n1190;
  assign new_n1314 = new_n1312 & new_n1313;
  assign new_n1315 = ~new_n1312 & ~new_n1313;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = \137  & \426 ;
  assign new_n1318 = ~new_n1316 & new_n1317;
  assign new_n1319 = new_n1316 & ~new_n1317;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = ~new_n1195 & ~new_n1198;
  assign new_n1322 = \120  & \443 ;
  assign new_n1323 = new_n1321 & ~new_n1322;
  assign new_n1324 = ~new_n1321 & new_n1322;
  assign new_n1325 = ~new_n1323 & ~new_n1324;
  assign new_n1326 = new_n1320 & new_n1325;
  assign new_n1327 = ~new_n1320 & ~new_n1325;
  assign new_n1328 = ~new_n1326 & ~new_n1327;
  assign new_n1329 = ~new_n1203 & ~new_n1205;
  assign new_n1330 = new_n1328 & new_n1329;
  assign new_n1331 = ~new_n1328 & ~new_n1329;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = \103  & \460 ;
  assign new_n1334 = ~new_n1332 & new_n1333;
  assign new_n1335 = new_n1332 & ~new_n1333;
  assign new_n1336 = ~new_n1334 & ~new_n1335;
  assign new_n1337 = ~new_n1210 & ~new_n1214;
  assign new_n1338 = new_n1336 & ~new_n1337;
  assign new_n1339 = ~new_n1336 & new_n1337;
  assign new_n1340 = ~new_n1338 & ~new_n1339;
  assign new_n1341 = \86  & \477 ;
  assign new_n1342 = ~new_n1340 & new_n1341;
  assign new_n1343 = new_n1340 & ~new_n1341;
  assign new_n1344 = ~new_n1342 & ~new_n1343;
  assign new_n1345 = \69  & \494 ;
  assign new_n1346 = ~new_n1217 & ~new_n1220;
  assign new_n1347 = ~new_n1345 & new_n1346;
  assign new_n1348 = new_n1345 & ~new_n1346;
  assign new_n1349 = ~new_n1347 & ~new_n1348;
  assign new_n1350 = new_n1344 & new_n1349;
  assign new_n1351 = ~new_n1344 & ~new_n1349;
  assign new_n1352 = ~new_n1350 & ~new_n1351;
  assign new_n1353 = ~new_n1225 & ~new_n1229;
  assign new_n1354 = new_n1352 & ~new_n1353;
  assign new_n1355 = ~new_n1352 & new_n1353;
  assign new_n1356 = ~new_n1354 & ~new_n1355;
  assign new_n1357 = \52  & \511 ;
  assign new_n1358 = ~new_n1356 & new_n1357;
  assign new_n1359 = new_n1356 & ~new_n1357;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = ~new_n1232 & ~new_n1237;
  assign new_n1362 = ~new_n1360 & new_n1361;
  assign new_n1363 = new_n1360 & ~new_n1361;
  assign new_n1364 = ~new_n1362 & ~new_n1363;
  assign new_n1365 = new_n1256 & new_n1364;
  assign new_n1366 = ~new_n1256 & ~new_n1364;
  assign new_n1367 = ~new_n1365 & ~new_n1366;
  assign new_n1368 = ~new_n1244 & ~new_n1250;
  assign new_n1369 = ~new_n1367 & ~new_n1368;
  assign new_n1370 = new_n1367 & new_n1368;
  assign new_n1371 = ~new_n1369 & ~new_n1370;
  assign new_n1372 = new_n1253 & ~new_n1371;
  assign new_n1373 = ~new_n1253 & new_n1371;
  assign \6160  = new_n1372 | new_n1373;
  assign new_n1375 = \52  & \528 ;
  assign new_n1376 = ~new_n1354 & ~new_n1359;
  assign new_n1377 = ~new_n1375 & ~new_n1376;
  assign new_n1378 = new_n1375 & new_n1376;
  assign new_n1379 = ~new_n1377 & ~new_n1378;
  assign new_n1380 = \103  & \477 ;
  assign new_n1381 = \205  & \375 ;
  assign new_n1382 = \222  & new_n1260;
  assign new_n1383 = ~new_n1277 & ~new_n1382;
  assign new_n1384 = \358  & ~new_n1383;
  assign new_n1385 = \222  & \358 ;
  assign new_n1386 = new_n1383 & ~new_n1385;
  assign new_n1387 = ~new_n1384 & ~new_n1386;
  assign new_n1388 = \256  & \324 ;
  assign new_n1389 = new_n1142 & new_n1143;
  assign new_n1390 = ~new_n1267 & ~new_n1389;
  assign new_n1391 = \341  & ~new_n1390;
  assign new_n1392 = \239  & \341 ;
  assign new_n1393 = new_n1390 & ~new_n1392;
  assign new_n1394 = ~new_n1391 & ~new_n1393;
  assign new_n1395 = new_n1388 & ~new_n1394;
  assign new_n1396 = ~new_n1388 & new_n1394;
  assign new_n1397 = ~new_n1395 & ~new_n1396;
  assign new_n1398 = ~new_n1387 & ~new_n1397;
  assign new_n1399 = new_n1387 & new_n1397;
  assign new_n1400 = ~new_n1398 & ~new_n1399;
  assign new_n1401 = ~new_n1281 & ~new_n1286;
  assign new_n1402 = ~new_n1400 & new_n1401;
  assign new_n1403 = new_n1400 & ~new_n1401;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = new_n1381 & new_n1404;
  assign new_n1406 = ~new_n1381 & ~new_n1404;
  assign new_n1407 = ~new_n1405 & ~new_n1406;
  assign new_n1408 = \188  & \392 ;
  assign new_n1409 = ~new_n1290 & ~new_n1293;
  assign new_n1410 = ~new_n1408 & ~new_n1409;
  assign new_n1411 = \392  & new_n1409;
  assign new_n1412 = ~new_n1410 & ~new_n1411;
  assign new_n1413 = new_n1407 & new_n1412;
  assign new_n1414 = ~new_n1407 & ~new_n1412;
  assign new_n1415 = ~new_n1413 & ~new_n1414;
  assign new_n1416 = ~new_n1297 & ~new_n1302;
  assign new_n1417 = ~new_n1415 & ~new_n1416;
  assign new_n1418 = new_n1415 & new_n1416;
  assign new_n1419 = ~new_n1417 & ~new_n1418;
  assign new_n1420 = \171  & \409 ;
  assign new_n1421 = ~new_n1419 & new_n1420;
  assign new_n1422 = new_n1419 & ~new_n1420;
  assign new_n1423 = ~new_n1421 & ~new_n1422;
  assign new_n1424 = \154  & \426 ;
  assign new_n1425 = new_n1423 & ~new_n1424;
  assign new_n1426 = ~new_n1423 & new_n1424;
  assign new_n1427 = ~new_n1425 & ~new_n1426;
  assign new_n1428 = ~new_n1306 & ~new_n1310;
  assign new_n1429 = new_n1427 & new_n1428;
  assign new_n1430 = ~new_n1427 & ~new_n1428;
  assign new_n1431 = ~new_n1429 & ~new_n1430;
  assign new_n1432 = ~new_n1315 & ~new_n1319;
  assign new_n1433 = new_n1431 & ~new_n1432;
  assign new_n1434 = ~new_n1431 & new_n1432;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = \137  & \443 ;
  assign new_n1437 = ~new_n1435 & new_n1436;
  assign new_n1438 = new_n1435 & ~new_n1436;
  assign new_n1439 = ~new_n1437 & ~new_n1438;
  assign new_n1440 = \120  & \460 ;
  assign new_n1441 = ~new_n1323 & ~new_n1326;
  assign new_n1442 = ~new_n1440 & ~new_n1441;
  assign new_n1443 = \460  & new_n1441;
  assign new_n1444 = ~new_n1442 & ~new_n1443;
  assign new_n1445 = ~new_n1439 & ~new_n1444;
  assign new_n1446 = new_n1439 & new_n1444;
  assign new_n1447 = ~new_n1445 & ~new_n1446;
  assign new_n1448 = ~new_n1330 & ~new_n1335;
  assign new_n1449 = new_n1447 & ~new_n1448;
  assign new_n1450 = ~new_n1447 & new_n1448;
  assign new_n1451 = ~new_n1449 & ~new_n1450;
  assign new_n1452 = new_n1380 & ~new_n1451;
  assign new_n1453 = ~new_n1380 & new_n1451;
  assign new_n1454 = ~new_n1452 & ~new_n1453;
  assign new_n1455 = ~new_n1338 & ~new_n1343;
  assign new_n1456 = \86  & \494 ;
  assign new_n1457 = ~new_n1455 & ~new_n1456;
  assign new_n1458 = \494  & new_n1455;
  assign new_n1459 = ~new_n1457 & ~new_n1458;
  assign new_n1460 = new_n1454 & new_n1459;
  assign new_n1461 = ~new_n1454 & ~new_n1459;
  assign new_n1462 = ~new_n1460 & ~new_n1461;
  assign new_n1463 = ~new_n1347 & ~new_n1350;
  assign new_n1464 = \69  & \511 ;
  assign new_n1465 = ~new_n1463 & ~new_n1464;
  assign new_n1466 = \511  & new_n1463;
  assign new_n1467 = ~new_n1465 & ~new_n1466;
  assign new_n1468 = new_n1462 & new_n1467;
  assign new_n1469 = ~new_n1462 & ~new_n1467;
  assign new_n1470 = ~new_n1468 & ~new_n1469;
  assign new_n1471 = ~new_n1379 & new_n1470;
  assign new_n1472 = new_n1379 & ~new_n1470;
  assign new_n1473 = ~new_n1471 & ~new_n1472;
  assign new_n1474 = ~new_n1362 & ~new_n1365;
  assign new_n1475 = new_n1473 & ~new_n1474;
  assign new_n1476 = ~new_n1473 & new_n1474;
  assign new_n1477 = ~new_n1475 & ~new_n1476;
  assign new_n1478 = ~new_n1369 & ~new_n1373;
  assign new_n1479 = new_n1477 & new_n1478;
  assign new_n1480 = ~new_n1477 & ~new_n1478;
  assign \6170  = ~new_n1479 & ~new_n1480;
  assign new_n1482 = \86  & \511 ;
  assign new_n1483 = ~new_n1457 & ~new_n1460;
  assign new_n1484 = ~new_n1482 & ~new_n1483;
  assign new_n1485 = new_n1482 & new_n1483;
  assign new_n1486 = ~new_n1484 & ~new_n1485;
  assign new_n1487 = ~new_n1433 & ~new_n1438;
  assign new_n1488 = ~new_n1386 & ~new_n1399;
  assign new_n1489 = \256  & \341 ;
  assign new_n1490 = ~new_n1268 & ~new_n1392;
  assign new_n1491 = \358  & ~new_n1490;
  assign new_n1492 = ~\358  & new_n1266;
  assign new_n1493 = ~new_n1489 & ~new_n1492;
  assign new_n1494 = ~new_n1491 & new_n1493;
  assign new_n1495 = \256  & \358 ;
  assign new_n1496 = ~new_n1388 & ~new_n1495;
  assign new_n1497 = new_n1392 & ~new_n1496;
  assign new_n1498 = ~new_n1390 & new_n1397;
  assign new_n1499 = ~new_n1497 & ~new_n1498;
  assign new_n1500 = \358  & ~new_n1499;
  assign new_n1501 = ~\341  & ~\358 ;
  assign new_n1502 = ~new_n1499 & ~new_n1501;
  assign new_n1503 = ~new_n1495 & ~new_n1502;
  assign new_n1504 = ~new_n1500 & ~new_n1503;
  assign new_n1505 = new_n1392 & new_n1504;
  assign new_n1506 = ~\324  & new_n1497;
  assign new_n1507 = ~new_n1501 & ~new_n1506;
  assign new_n1508 = new_n1390 & ~new_n1507;
  assign new_n1509 = ~new_n1494 & ~new_n1508;
  assign new_n1510 = ~new_n1505 & new_n1509;
  assign new_n1511 = new_n1488 & new_n1510;
  assign new_n1512 = ~new_n1488 & ~new_n1510;
  assign new_n1513 = ~new_n1511 & ~new_n1512;
  assign new_n1514 = \222  & \375 ;
  assign new_n1515 = ~new_n1513 & new_n1514;
  assign new_n1516 = new_n1513 & ~new_n1514;
  assign new_n1517 = ~new_n1515 & ~new_n1516;
  assign new_n1518 = \205  & \392 ;
  assign new_n1519 = new_n1517 & ~new_n1518;
  assign new_n1520 = ~new_n1517 & new_n1518;
  assign new_n1521 = ~new_n1519 & ~new_n1520;
  assign new_n1522 = ~new_n1402 & ~new_n1405;
  assign new_n1523 = new_n1521 & new_n1522;
  assign new_n1524 = ~new_n1521 & ~new_n1522;
  assign new_n1525 = ~new_n1523 & ~new_n1524;
  assign new_n1526 = ~new_n1411 & ~new_n1413;
  assign new_n1527 = \188  & \409 ;
  assign new_n1528 = new_n1526 & ~new_n1527;
  assign new_n1529 = ~new_n1526 & new_n1527;
  assign new_n1530 = ~new_n1528 & ~new_n1529;
  assign new_n1531 = new_n1525 & new_n1530;
  assign new_n1532 = ~new_n1525 & ~new_n1530;
  assign new_n1533 = ~new_n1531 & ~new_n1532;
  assign new_n1534 = ~new_n1417 & ~new_n1422;
  assign new_n1535 = new_n1533 & ~new_n1534;
  assign new_n1536 = ~new_n1533 & new_n1534;
  assign new_n1537 = ~new_n1535 & ~new_n1536;
  assign new_n1538 = \171  & \426 ;
  assign new_n1539 = ~new_n1537 & new_n1538;
  assign new_n1540 = new_n1537 & ~new_n1538;
  assign new_n1541 = ~new_n1539 & ~new_n1540;
  assign new_n1542 = ~new_n1425 & ~new_n1429;
  assign new_n1543 = \154  & \443 ;
  assign new_n1544 = ~new_n1542 & ~new_n1543;
  assign new_n1545 = \443  & new_n1542;
  assign new_n1546 = ~new_n1544 & ~new_n1545;
  assign new_n1547 = new_n1541 & new_n1546;
  assign new_n1548 = ~new_n1541 & ~new_n1546;
  assign new_n1549 = ~new_n1547 & ~new_n1548;
  assign new_n1550 = \137  & \460 ;
  assign new_n1551 = new_n1549 & ~new_n1550;
  assign new_n1552 = ~new_n1549 & new_n1550;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = new_n1487 & new_n1553;
  assign new_n1555 = ~new_n1487 & ~new_n1553;
  assign new_n1556 = ~new_n1554 & ~new_n1555;
  assign new_n1557 = ~new_n1442 & ~new_n1446;
  assign new_n1558 = ~new_n1556 & ~new_n1557;
  assign new_n1559 = new_n1556 & new_n1557;
  assign new_n1560 = ~new_n1558 & ~new_n1559;
  assign new_n1561 = \120  & \477 ;
  assign new_n1562 = ~new_n1560 & new_n1561;
  assign new_n1563 = new_n1560 & ~new_n1561;
  assign new_n1564 = ~new_n1562 & ~new_n1563;
  assign new_n1565 = ~new_n1449 & ~new_n1453;
  assign new_n1566 = \494  & new_n1565;
  assign new_n1567 = \103  & \494 ;
  assign new_n1568 = ~new_n1565 & ~new_n1567;
  assign new_n1569 = ~new_n1566 & ~new_n1568;
  assign new_n1570 = new_n1564 & ~new_n1569;
  assign new_n1571 = ~new_n1564 & new_n1569;
  assign new_n1572 = ~new_n1570 & ~new_n1571;
  assign new_n1573 = ~new_n1486 & new_n1572;
  assign new_n1574 = new_n1486 & ~new_n1572;
  assign new_n1575 = ~new_n1573 & ~new_n1574;
  assign new_n1576 = ~new_n1465 & ~new_n1468;
  assign new_n1577 = ~new_n1575 & new_n1576;
  assign new_n1578 = new_n1575 & ~new_n1576;
  assign new_n1579 = ~new_n1577 & ~new_n1578;
  assign new_n1580 = \69  & \528 ;
  assign new_n1581 = ~new_n1579 & new_n1580;
  assign new_n1582 = new_n1579 & ~new_n1580;
  assign new_n1583 = ~new_n1581 & ~new_n1582;
  assign new_n1584 = ~new_n1378 & ~new_n1472;
  assign new_n1585 = ~new_n1583 & ~new_n1584;
  assign new_n1586 = new_n1583 & new_n1584;
  assign new_n1587 = ~new_n1585 & ~new_n1586;
  assign new_n1588 = ~new_n1475 & ~new_n1479;
  assign new_n1589 = new_n1587 & new_n1588;
  assign new_n1590 = ~new_n1587 & ~new_n1588;
  assign \6180  = new_n1589 | new_n1590;
  assign new_n1592 = \86  & \528 ;
  assign new_n1593 = ~new_n1558 & ~new_n1563;
  assign new_n1594 = \494  & new_n1593;
  assign new_n1595 = \120  & \494 ;
  assign new_n1596 = ~new_n1593 & ~new_n1595;
  assign new_n1597 = ~new_n1594 & ~new_n1596;
  assign new_n1598 = \137  & \477 ;
  assign new_n1599 = ~new_n1552 & ~new_n1554;
  assign new_n1600 = ~new_n1598 & new_n1599;
  assign new_n1601 = new_n1598 & ~new_n1599;
  assign new_n1602 = ~new_n1600 & ~new_n1601;
  assign new_n1603 = \205  & \409 ;
  assign new_n1604 = ~new_n1519 & ~new_n1523;
  assign new_n1605 = ~new_n1603 & ~new_n1604;
  assign new_n1606 = new_n1603 & new_n1604;
  assign new_n1607 = ~new_n1605 & ~new_n1606;
  assign new_n1608 = ~new_n1512 & ~new_n1516;
  assign new_n1609 = \239  & \375 ;
  assign new_n1610 = ~new_n1504 & new_n1609;
  assign new_n1611 = new_n1504 & ~new_n1609;
  assign new_n1612 = ~new_n1610 & ~new_n1611;
  assign new_n1613 = new_n1608 & ~new_n1612;
  assign new_n1614 = ~new_n1608 & new_n1612;
  assign new_n1615 = ~new_n1613 & ~new_n1614;
  assign new_n1616 = \222  & \392 ;
  assign new_n1617 = ~new_n1615 & new_n1616;
  assign new_n1618 = new_n1615 & ~new_n1616;
  assign new_n1619 = ~new_n1617 & ~new_n1618;
  assign new_n1620 = ~new_n1607 & new_n1619;
  assign new_n1621 = new_n1607 & ~new_n1619;
  assign new_n1622 = ~new_n1620 & ~new_n1621;
  assign new_n1623 = ~new_n1528 & ~new_n1531;
  assign new_n1624 = new_n1622 & new_n1623;
  assign new_n1625 = ~new_n1622 & ~new_n1623;
  assign new_n1626 = ~new_n1624 & ~new_n1625;
  assign new_n1627 = \188  & \426 ;
  assign new_n1628 = ~new_n1626 & new_n1627;
  assign new_n1629 = new_n1626 & ~new_n1627;
  assign new_n1630 = ~new_n1628 & ~new_n1629;
  assign new_n1631 = ~new_n1535 & ~new_n1540;
  assign new_n1632 = ~new_n1630 & new_n1631;
  assign new_n1633 = new_n1630 & ~new_n1631;
  assign new_n1634 = ~new_n1632 & ~new_n1633;
  assign new_n1635 = \171  & \443 ;
  assign new_n1636 = ~new_n1634 & new_n1635;
  assign new_n1637 = new_n1634 & ~new_n1635;
  assign new_n1638 = ~new_n1636 & ~new_n1637;
  assign new_n1639 = ~new_n1544 & ~new_n1547;
  assign new_n1640 = \154  & \460 ;
  assign new_n1641 = ~new_n1639 & ~new_n1640;
  assign new_n1642 = new_n1639 & new_n1640;
  assign new_n1643 = ~new_n1641 & ~new_n1642;
  assign new_n1644 = ~new_n1638 & ~new_n1643;
  assign new_n1645 = new_n1638 & new_n1643;
  assign new_n1646 = ~new_n1644 & ~new_n1645;
  assign new_n1647 = new_n1602 & ~new_n1646;
  assign new_n1648 = ~new_n1602 & new_n1646;
  assign new_n1649 = ~new_n1647 & ~new_n1648;
  assign new_n1650 = ~new_n1597 & ~new_n1649;
  assign new_n1651 = new_n1597 & new_n1649;
  assign new_n1652 = ~new_n1650 & ~new_n1651;
  assign new_n1653 = ~new_n1566 & ~new_n1571;
  assign new_n1654 = ~new_n1652 & new_n1653;
  assign new_n1655 = new_n1652 & ~new_n1653;
  assign new_n1656 = ~new_n1654 & ~new_n1655;
  assign new_n1657 = \103  & \511 ;
  assign new_n1658 = ~new_n1656 & new_n1657;
  assign new_n1659 = new_n1656 & ~new_n1657;
  assign new_n1660 = ~new_n1658 & ~new_n1659;
  assign new_n1661 = ~new_n1484 & ~new_n1574;
  assign new_n1662 = ~new_n1660 & new_n1661;
  assign new_n1663 = new_n1660 & ~new_n1661;
  assign new_n1664 = ~new_n1662 & ~new_n1663;
  assign new_n1665 = new_n1592 & new_n1664;
  assign new_n1666 = ~new_n1592 & ~new_n1664;
  assign new_n1667 = ~new_n1665 & ~new_n1666;
  assign new_n1668 = ~new_n1578 & ~new_n1582;
  assign new_n1669 = ~new_n1667 & ~new_n1668;
  assign new_n1670 = new_n1667 & new_n1668;
  assign new_n1671 = ~new_n1669 & ~new_n1670;
  assign new_n1672 = ~new_n1586 & ~new_n1589;
  assign new_n1673 = new_n1671 & new_n1672;
  assign new_n1674 = ~new_n1671 & ~new_n1672;
  assign \6190  = ~new_n1673 & ~new_n1674;
  assign new_n1676 = \154  & \477 ;
  assign new_n1677 = \256  & \392 ;
  assign new_n1678 = ~new_n1500 & ~new_n1609;
  assign new_n1679 = new_n1677 & ~new_n1678;
  assign new_n1680 = \239  & ~new_n1679;
  assign new_n1681 = ~\375  & ~new_n1680;
  assign new_n1682 = ~\358  & ~\375 ;
  assign new_n1683 = \256  & ~new_n1682;
  assign new_n1684 = ~\239  & ~\256 ;
  assign new_n1685 = \392  & ~new_n1684;
  assign new_n1686 = ~new_n1683 & ~new_n1685;
  assign new_n1687 = \358  & ~\392 ;
  assign new_n1688 = ~\358  & \375 ;
  assign new_n1689 = new_n1677 & new_n1688;
  assign new_n1690 = ~new_n1687 & ~new_n1689;
  assign new_n1691 = \239  & ~new_n1690;
  assign new_n1692 = ~new_n1502 & new_n1691;
  assign new_n1693 = \375  & ~new_n1677;
  assign new_n1694 = new_n1502 & new_n1693;
  assign new_n1695 = ~new_n1686 & ~new_n1692;
  assign new_n1696 = ~new_n1694 & new_n1695;
  assign new_n1697 = ~new_n1681 & new_n1696;
  assign new_n1698 = \222  & \409 ;
  assign new_n1699 = new_n1697 & new_n1698;
  assign new_n1700 = ~new_n1697 & ~new_n1698;
  assign new_n1701 = ~new_n1699 & ~new_n1700;
  assign new_n1702 = ~new_n1614 & ~new_n1618;
  assign new_n1703 = new_n1701 & new_n1702;
  assign new_n1704 = ~new_n1701 & ~new_n1702;
  assign new_n1705 = ~new_n1703 & ~new_n1704;
  assign new_n1706 = ~new_n1606 & ~new_n1621;
  assign new_n1707 = ~new_n1705 & new_n1706;
  assign new_n1708 = new_n1705 & ~new_n1706;
  assign new_n1709 = ~new_n1707 & ~new_n1708;
  assign new_n1710 = \205  & \426 ;
  assign new_n1711 = ~new_n1709 & new_n1710;
  assign new_n1712 = new_n1709 & ~new_n1710;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = \188  & \443 ;
  assign new_n1715 = new_n1713 & ~new_n1714;
  assign new_n1716 = ~new_n1713 & new_n1714;
  assign new_n1717 = ~new_n1715 & ~new_n1716;
  assign new_n1718 = ~new_n1625 & ~new_n1629;
  assign new_n1719 = new_n1717 & ~new_n1718;
  assign new_n1720 = ~new_n1717 & new_n1718;
  assign new_n1721 = ~new_n1719 & ~new_n1720;
  assign new_n1722 = ~new_n1633 & ~new_n1637;
  assign new_n1723 = \460  & new_n1722;
  assign new_n1724 = \171  & \460 ;
  assign new_n1725 = ~new_n1722 & ~new_n1724;
  assign new_n1726 = ~new_n1723 & ~new_n1725;
  assign new_n1727 = ~new_n1721 & new_n1726;
  assign new_n1728 = new_n1721 & ~new_n1726;
  assign new_n1729 = ~new_n1727 & ~new_n1728;
  assign new_n1730 = ~new_n1641 & ~new_n1645;
  assign new_n1731 = ~new_n1729 & ~new_n1730;
  assign new_n1732 = new_n1729 & new_n1730;
  assign new_n1733 = ~new_n1731 & ~new_n1732;
  assign new_n1734 = new_n1676 & ~new_n1733;
  assign new_n1735 = ~new_n1676 & new_n1733;
  assign new_n1736 = ~new_n1734 & ~new_n1735;
  assign new_n1737 = ~new_n1601 & ~new_n1647;
  assign new_n1738 = new_n1736 & new_n1737;
  assign new_n1739 = ~new_n1736 & ~new_n1737;
  assign new_n1740 = ~new_n1738 & ~new_n1739;
  assign new_n1741 = \137  & \494 ;
  assign new_n1742 = ~new_n1740 & new_n1741;
  assign new_n1743 = new_n1740 & ~new_n1741;
  assign new_n1744 = ~new_n1742 & ~new_n1743;
  assign new_n1745 = \120  & \511 ;
  assign new_n1746 = ~new_n1594 & ~new_n1651;
  assign new_n1747 = ~new_n1745 & new_n1746;
  assign new_n1748 = \511  & ~new_n1746;
  assign new_n1749 = ~new_n1747 & ~new_n1748;
  assign new_n1750 = new_n1744 & new_n1749;
  assign new_n1751 = ~new_n1744 & ~new_n1749;
  assign new_n1752 = ~new_n1750 & ~new_n1751;
  assign new_n1753 = ~new_n1654 & ~new_n1659;
  assign new_n1754 = ~new_n1752 & new_n1753;
  assign new_n1755 = new_n1752 & ~new_n1753;
  assign new_n1756 = ~new_n1754 & ~new_n1755;
  assign new_n1757 = \103  & \528 ;
  assign new_n1758 = ~new_n1756 & new_n1757;
  assign new_n1759 = new_n1756 & ~new_n1757;
  assign new_n1760 = ~new_n1758 & ~new_n1759;
  assign new_n1761 = ~new_n1662 & ~new_n1665;
  assign new_n1762 = new_n1760 & new_n1761;
  assign new_n1763 = ~new_n1760 & ~new_n1761;
  assign new_n1764 = ~new_n1762 & ~new_n1763;
  assign new_n1765 = ~new_n1670 & ~new_n1673;
  assign new_n1766 = ~new_n1764 & new_n1765;
  assign new_n1767 = new_n1764 & ~new_n1765;
  assign \6200  = ~new_n1766 & ~new_n1767;
  assign new_n1769 = ~new_n1755 & ~new_n1759;
  assign new_n1770 = ~new_n1747 & ~new_n1750;
  assign new_n1771 = ~new_n1731 & ~new_n1735;
  assign new_n1772 = \205  & \443 ;
  assign new_n1773 = ~new_n1707 & ~new_n1712;
  assign new_n1774 = ~new_n1699 & ~new_n1703;
  assign new_n1775 = \222  & \426 ;
  assign new_n1776 = ~new_n1503 & new_n1609;
  assign new_n1777 = ~new_n1677 & ~new_n1776;
  assign new_n1778 = ~new_n1679 & ~new_n1777;
  assign new_n1779 = \239  & \409 ;
  assign new_n1780 = new_n1778 & ~new_n1779;
  assign new_n1781 = ~new_n1778 & new_n1779;
  assign new_n1782 = ~new_n1780 & ~new_n1781;
  assign new_n1783 = new_n1775 & new_n1782;
  assign new_n1784 = ~new_n1775 & ~new_n1782;
  assign new_n1785 = ~new_n1783 & ~new_n1784;
  assign new_n1786 = new_n1774 & ~new_n1785;
  assign new_n1787 = ~new_n1774 & new_n1785;
  assign new_n1788 = ~new_n1786 & ~new_n1787;
  assign new_n1789 = new_n1773 & ~new_n1788;
  assign new_n1790 = ~new_n1773 & new_n1788;
  assign new_n1791 = ~new_n1789 & ~new_n1790;
  assign new_n1792 = new_n1772 & new_n1791;
  assign new_n1793 = ~new_n1772 & ~new_n1791;
  assign new_n1794 = ~new_n1792 & ~new_n1793;
  assign new_n1795 = ~new_n1715 & ~new_n1719;
  assign new_n1796 = ~new_n1794 & ~new_n1795;
  assign new_n1797 = new_n1794 & new_n1795;
  assign new_n1798 = ~new_n1796 & ~new_n1797;
  assign new_n1799 = \188  & \460 ;
  assign new_n1800 = ~new_n1798 & new_n1799;
  assign new_n1801 = new_n1798 & ~new_n1799;
  assign new_n1802 = ~new_n1800 & ~new_n1801;
  assign new_n1803 = \171  & \477 ;
  assign new_n1804 = ~new_n1723 & ~new_n1727;
  assign new_n1805 = ~new_n1803 & new_n1804;
  assign new_n1806 = new_n1803 & ~new_n1804;
  assign new_n1807 = ~new_n1805 & ~new_n1806;
  assign new_n1808 = new_n1802 & new_n1807;
  assign new_n1809 = ~new_n1802 & ~new_n1807;
  assign new_n1810 = ~new_n1808 & ~new_n1809;
  assign new_n1811 = ~new_n1771 & new_n1810;
  assign new_n1812 = new_n1771 & ~new_n1810;
  assign new_n1813 = ~new_n1811 & ~new_n1812;
  assign new_n1814 = \154  & \494 ;
  assign new_n1815 = ~new_n1813 & new_n1814;
  assign new_n1816 = new_n1813 & ~new_n1814;
  assign new_n1817 = ~new_n1815 & ~new_n1816;
  assign new_n1818 = ~new_n1738 & ~new_n1743;
  assign new_n1819 = \137  & \511 ;
  assign new_n1820 = ~new_n1818 & ~new_n1819;
  assign new_n1821 = \511  & new_n1818;
  assign new_n1822 = ~new_n1820 & ~new_n1821;
  assign new_n1823 = new_n1817 & new_n1822;
  assign new_n1824 = ~new_n1817 & ~new_n1822;
  assign new_n1825 = ~new_n1823 & ~new_n1824;
  assign new_n1826 = \120  & \528 ;
  assign new_n1827 = new_n1825 & ~new_n1826;
  assign new_n1828 = ~new_n1825 & new_n1826;
  assign new_n1829 = ~new_n1827 & ~new_n1828;
  assign new_n1830 = new_n1770 & new_n1829;
  assign new_n1831 = ~new_n1770 & ~new_n1829;
  assign new_n1832 = ~new_n1830 & ~new_n1831;
  assign new_n1833 = new_n1769 & new_n1832;
  assign new_n1834 = ~new_n1769 & ~new_n1832;
  assign new_n1835 = ~new_n1833 & ~new_n1834;
  assign new_n1836 = ~new_n1762 & ~new_n1765;
  assign new_n1837 = ~new_n1763 & ~new_n1836;
  assign new_n1838 = new_n1835 & new_n1837;
  assign new_n1839 = ~new_n1835 & ~new_n1837;
  assign \6210  = new_n1838 | new_n1839;
  assign new_n1841 = ~new_n1775 & new_n1782;
  assign new_n1842 = ~new_n1786 & ~new_n1841;
  assign new_n1843 = \443  & new_n1842;
  assign new_n1844 = \222  & \443 ;
  assign new_n1845 = ~new_n1842 & ~new_n1844;
  assign new_n1846 = ~new_n1843 & ~new_n1845;
  assign new_n1847 = \256  & \426 ;
  assign new_n1848 = \409  & ~new_n1777;
  assign new_n1849 = new_n1847 & new_n1848;
  assign new_n1850 = \239  & \426 ;
  assign new_n1851 = ~\409  & ~new_n1850;
  assign new_n1852 = new_n1679 & new_n1851;
  assign new_n1853 = ~\256  & ~new_n1850;
  assign new_n1854 = \409  & ~\426 ;
  assign new_n1855 = \256  & ~new_n1854;
  assign new_n1856 = ~new_n1853 & ~new_n1855;
  assign new_n1857 = new_n1777 & new_n1856;
  assign new_n1858 = \409  & ~new_n1270;
  assign new_n1859 = ~new_n1851 & ~new_n1858;
  assign new_n1860 = ~new_n1679 & new_n1859;
  assign new_n1861 = ~new_n1852 & ~new_n1860;
  assign new_n1862 = ~new_n1857 & new_n1861;
  assign new_n1863 = ~new_n1849 & new_n1862;
  assign new_n1864 = ~new_n1846 & new_n1863;
  assign new_n1865 = new_n1846 & ~new_n1863;
  assign new_n1866 = ~new_n1864 & ~new_n1865;
  assign new_n1867 = ~new_n1789 & ~new_n1792;
  assign new_n1868 = ~new_n1866 & new_n1867;
  assign new_n1869 = new_n1866 & ~new_n1867;
  assign new_n1870 = ~new_n1868 & ~new_n1869;
  assign new_n1871 = \205  & \460 ;
  assign new_n1872 = ~new_n1870 & new_n1871;
  assign new_n1873 = new_n1870 & ~new_n1871;
  assign new_n1874 = ~new_n1872 & ~new_n1873;
  assign new_n1875 = ~new_n1796 & ~new_n1801;
  assign new_n1876 = \477  & new_n1875;
  assign new_n1877 = \188  & \477 ;
  assign new_n1878 = ~new_n1875 & ~new_n1877;
  assign new_n1879 = ~new_n1876 & ~new_n1878;
  assign new_n1880 = new_n1874 & ~new_n1879;
  assign new_n1881 = ~new_n1874 & new_n1879;
  assign new_n1882 = ~new_n1880 & ~new_n1881;
  assign new_n1883 = ~new_n1805 & ~new_n1808;
  assign new_n1884 = \494  & new_n1883;
  assign new_n1885 = \171  & \494 ;
  assign new_n1886 = ~new_n1883 & ~new_n1885;
  assign new_n1887 = ~new_n1884 & ~new_n1886;
  assign new_n1888 = new_n1882 & ~new_n1887;
  assign new_n1889 = ~new_n1882 & new_n1887;
  assign new_n1890 = ~new_n1888 & ~new_n1889;
  assign new_n1891 = ~new_n1811 & ~new_n1816;
  assign new_n1892 = new_n1890 & ~new_n1891;
  assign new_n1893 = ~new_n1890 & new_n1891;
  assign new_n1894 = ~new_n1892 & ~new_n1893;
  assign new_n1895 = \154  & \511 ;
  assign new_n1896 = ~new_n1894 & new_n1895;
  assign new_n1897 = new_n1894 & ~new_n1895;
  assign new_n1898 = ~new_n1896 & ~new_n1897;
  assign new_n1899 = \137  & \528 ;
  assign new_n1900 = new_n1898 & ~new_n1899;
  assign new_n1901 = ~new_n1898 & new_n1899;
  assign new_n1902 = ~new_n1900 & ~new_n1901;
  assign new_n1903 = ~new_n1820 & ~new_n1823;
  assign new_n1904 = new_n1902 & ~new_n1903;
  assign new_n1905 = ~new_n1902 & new_n1903;
  assign new_n1906 = ~new_n1904 & ~new_n1905;
  assign new_n1907 = ~new_n1828 & ~new_n1830;
  assign new_n1908 = ~new_n1906 & ~new_n1907;
  assign new_n1909 = new_n1906 & new_n1907;
  assign new_n1910 = ~new_n1908 & ~new_n1909;
  assign new_n1911 = ~new_n1834 & ~new_n1838;
  assign new_n1912 = new_n1910 & ~new_n1911;
  assign new_n1913 = ~new_n1910 & new_n1911;
  assign \6220  = new_n1912 | new_n1913;
  assign new_n1915 = \154  & \528 ;
  assign new_n1916 = ~new_n1892 & ~new_n1897;
  assign new_n1917 = ~new_n1915 & ~new_n1916;
  assign new_n1918 = new_n1915 & new_n1916;
  assign new_n1919 = ~new_n1917 & ~new_n1918;
  assign new_n1920 = ~new_n1886 & ~new_n1889;
  assign new_n1921 = \222  & \460 ;
  assign new_n1922 = \239  & new_n1848;
  assign new_n1923 = ~new_n1679 & ~new_n1922;
  assign new_n1924 = new_n1854 & ~new_n1923;
  assign new_n1925 = new_n1847 & new_n1923;
  assign new_n1926 = ~new_n1924 & ~new_n1925;
  assign new_n1927 = \239  & \443 ;
  assign new_n1928 = new_n1926 & new_n1927;
  assign new_n1929 = ~\239  & ~new_n1926;
  assign new_n1930 = ~\443  & new_n1924;
  assign new_n1931 = ~\409  & ~\443 ;
  assign new_n1932 = \409  & \443 ;
  assign new_n1933 = ~new_n1931 & ~new_n1932;
  assign new_n1934 = new_n1925 & ~new_n1933;
  assign new_n1935 = ~new_n1930 & ~new_n1934;
  assign new_n1936 = ~new_n1928 & new_n1935;
  assign new_n1937 = ~new_n1929 & new_n1936;
  assign new_n1938 = ~new_n1921 & new_n1937;
  assign new_n1939 = new_n1921 & ~new_n1937;
  assign new_n1940 = ~new_n1938 & ~new_n1939;
  assign new_n1941 = ~new_n1843 & ~new_n1865;
  assign new_n1942 = new_n1940 & ~new_n1941;
  assign new_n1943 = ~new_n1940 & new_n1941;
  assign new_n1944 = ~new_n1942 & ~new_n1943;
  assign new_n1945 = ~new_n1868 & ~new_n1873;
  assign new_n1946 = ~new_n1944 & ~new_n1945;
  assign new_n1947 = new_n1944 & new_n1945;
  assign new_n1948 = ~new_n1946 & ~new_n1947;
  assign new_n1949 = \205  & \477 ;
  assign new_n1950 = ~new_n1948 & new_n1949;
  assign new_n1951 = new_n1948 & ~new_n1949;
  assign new_n1952 = ~new_n1950 & ~new_n1951;
  assign new_n1953 = ~new_n1876 & ~new_n1881;
  assign new_n1954 = ~new_n1952 & ~new_n1953;
  assign new_n1955 = new_n1952 & new_n1953;
  assign new_n1956 = ~new_n1954 & ~new_n1955;
  assign new_n1957 = \188  & \494 ;
  assign new_n1958 = new_n1956 & new_n1957;
  assign new_n1959 = ~new_n1956 & ~new_n1957;
  assign new_n1960 = ~new_n1958 & ~new_n1959;
  assign new_n1961 = new_n1920 & new_n1960;
  assign new_n1962 = ~new_n1920 & ~new_n1960;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = \171  & \511 ;
  assign new_n1965 = ~new_n1963 & new_n1964;
  assign new_n1966 = new_n1963 & ~new_n1964;
  assign new_n1967 = ~new_n1965 & ~new_n1966;
  assign new_n1968 = ~new_n1919 & new_n1967;
  assign new_n1969 = new_n1919 & ~new_n1967;
  assign new_n1970 = ~new_n1968 & ~new_n1969;
  assign new_n1971 = ~new_n1900 & ~new_n1904;
  assign new_n1972 = ~new_n1970 & ~new_n1971;
  assign new_n1973 = new_n1970 & new_n1971;
  assign new_n1974 = ~new_n1972 & ~new_n1973;
  assign new_n1975 = ~new_n1909 & ~new_n1912;
  assign new_n1976 = ~new_n1974 & new_n1975;
  assign new_n1977 = new_n1974 & ~new_n1975;
  assign \6230  = new_n1976 | new_n1977;
  assign new_n1979 = \171  & \528 ;
  assign new_n1980 = ~new_n1962 & ~new_n1966;
  assign new_n1981 = ~new_n1979 & ~new_n1980;
  assign new_n1982 = \528  & new_n1980;
  assign new_n1983 = ~new_n1981 & ~new_n1982;
  assign new_n1984 = ~new_n1946 & ~new_n1951;
  assign new_n1985 = \494  & new_n1984;
  assign new_n1986 = \205  & \494 ;
  assign new_n1987 = ~new_n1984 & ~new_n1986;
  assign new_n1988 = ~new_n1985 & ~new_n1987;
  assign new_n1989 = \222  & \477 ;
  assign new_n1990 = ~new_n1939 & ~new_n1942;
  assign new_n1991 = \239  & \460 ;
  assign new_n1992 = \443  & new_n1779;
  assign new_n1993 = ~\426  & ~new_n1992;
  assign new_n1994 = ~new_n1923 & ~new_n1993;
  assign new_n1995 = new_n1265 & new_n1850;
  assign new_n1996 = ~new_n1931 & new_n1995;
  assign new_n1997 = ~new_n1994 & ~new_n1996;
  assign new_n1998 = ~new_n1991 & new_n1997;
  assign new_n1999 = new_n1991 & ~new_n1997;
  assign new_n2000 = ~new_n1998 & ~new_n1999;
  assign new_n2001 = \256  & \443 ;
  assign new_n2002 = ~new_n2000 & new_n2001;
  assign new_n2003 = new_n2000 & ~new_n2001;
  assign new_n2004 = ~new_n2002 & ~new_n2003;
  assign new_n2005 = new_n1990 & new_n2004;
  assign new_n2006 = ~new_n1990 & ~new_n2004;
  assign new_n2007 = ~new_n2005 & ~new_n2006;
  assign new_n2008 = new_n1989 & new_n2007;
  assign new_n2009 = ~new_n1989 & ~new_n2007;
  assign new_n2010 = ~new_n2008 & ~new_n2009;
  assign new_n2011 = ~new_n1988 & new_n2010;
  assign new_n2012 = new_n1988 & ~new_n2010;
  assign new_n2013 = ~new_n2011 & ~new_n2012;
  assign new_n2014 = \188  & \511 ;
  assign new_n2015 = ~new_n1954 & ~new_n1958;
  assign new_n2016 = ~new_n2014 & new_n2015;
  assign new_n2017 = new_n2014 & ~new_n2015;
  assign new_n2018 = ~new_n2016 & ~new_n2017;
  assign new_n2019 = new_n2013 & new_n2018;
  assign new_n2020 = ~new_n2013 & ~new_n2018;
  assign new_n2021 = ~new_n2019 & ~new_n2020;
  assign new_n2022 = new_n1983 & ~new_n2021;
  assign new_n2023 = ~new_n1983 & new_n2021;
  assign new_n2024 = ~new_n2022 & ~new_n2023;
  assign new_n2025 = ~new_n1918 & ~new_n1969;
  assign new_n2026 = new_n2024 & ~new_n2025;
  assign new_n2027 = ~new_n2024 & new_n2025;
  assign new_n2028 = ~new_n2026 & ~new_n2027;
  assign new_n2029 = ~new_n1973 & ~new_n1975;
  assign new_n2030 = ~new_n1972 & ~new_n2029;
  assign new_n2031 = new_n2028 & new_n2030;
  assign new_n2032 = ~new_n2028 & ~new_n2030;
  assign \6240  = ~new_n2031 & ~new_n2032;
  assign new_n2034 = ~new_n2026 & ~new_n2030;
  assign new_n2035 = ~new_n2027 & ~new_n2034;
  assign new_n2036 = \188  & \528 ;
  assign new_n2037 = ~new_n2016 & ~new_n2019;
  assign new_n2038 = ~new_n2036 & ~new_n2037;
  assign new_n2039 = new_n2036 & new_n2037;
  assign new_n2040 = ~new_n2038 & ~new_n2039;
  assign new_n2041 = ~new_n1987 & ~new_n2012;
  assign new_n2042 = \222  & \494 ;
  assign new_n2043 = ~new_n1989 & ~new_n2006;
  assign new_n2044 = ~new_n2005 & ~new_n2043;
  assign new_n2045 = \256  & \460 ;
  assign new_n2046 = ~new_n1998 & ~new_n2003;
  assign new_n2047 = \239  & \477 ;
  assign new_n2048 = new_n2046 & ~new_n2047;
  assign new_n2049 = ~new_n2046 & new_n2047;
  assign new_n2050 = ~new_n2048 & ~new_n2049;
  assign new_n2051 = new_n2045 & new_n2050;
  assign new_n2052 = ~new_n2045 & ~new_n2050;
  assign new_n2053 = ~new_n2051 & ~new_n2052;
  assign new_n2054 = new_n2044 & ~new_n2053;
  assign new_n2055 = ~new_n2044 & new_n2053;
  assign new_n2056 = ~new_n2054 & ~new_n2055;
  assign new_n2057 = new_n2042 & ~new_n2056;
  assign new_n2058 = ~new_n2042 & new_n2056;
  assign new_n2059 = ~new_n2057 & ~new_n2058;
  assign new_n2060 = new_n2041 & ~new_n2059;
  assign new_n2061 = ~new_n2041 & new_n2059;
  assign new_n2062 = ~new_n2060 & ~new_n2061;
  assign new_n2063 = \205  & \511 ;
  assign new_n2064 = ~new_n2062 & new_n2063;
  assign new_n2065 = new_n2062 & ~new_n2063;
  assign new_n2066 = ~new_n2064 & ~new_n2065;
  assign new_n2067 = ~new_n2040 & new_n2066;
  assign new_n2068 = new_n2040 & ~new_n2066;
  assign new_n2069 = ~new_n2067 & ~new_n2068;
  assign new_n2070 = ~new_n1982 & ~new_n2022;
  assign new_n2071 = ~new_n2069 & new_n2070;
  assign new_n2072 = new_n2069 & ~new_n2070;
  assign new_n2073 = ~new_n2071 & ~new_n2072;
  assign new_n2074 = new_n2035 & ~new_n2073;
  assign new_n2075 = ~new_n2035 & new_n2073;
  assign \6250  = new_n2074 | new_n2075;
  assign new_n2077 = \256  & new_n2047;
  assign new_n2078 = ~\494  & new_n2077;
  assign new_n2079 = ~\239  & \460 ;
  assign new_n2080 = ~\477  & ~new_n2045;
  assign new_n2081 = \256  & \477 ;
  assign new_n2082 = \494  & ~new_n2081;
  assign new_n2083 = ~new_n2080 & new_n2082;
  assign new_n2084 = ~new_n2078 & ~new_n2079;
  assign new_n2085 = ~new_n2083 & new_n2084;
  assign new_n2086 = new_n2046 & new_n2085;
  assign new_n2087 = ~\460  & \494 ;
  assign new_n2088 = new_n2077 & new_n2087;
  assign new_n2089 = \256  & ~new_n1991;
  assign new_n2090 = ~\494  & ~new_n2089;
  assign new_n2091 = ~new_n2088 & ~new_n2090;
  assign new_n2092 = ~new_n2046 & new_n2091;
  assign new_n2093 = ~new_n2086 & ~new_n2092;
  assign new_n2094 = ~\494  & new_n2080;
  assign new_n2095 = \239  & ~new_n2094;
  assign new_n2096 = ~new_n2081 & ~new_n2095;
  assign new_n2097 = ~new_n2093 & ~new_n2096;
  assign new_n2098 = ~new_n2055 & ~new_n2058;
  assign new_n2099 = new_n2097 & new_n2098;
  assign new_n2100 = ~new_n2097 & ~new_n2098;
  assign new_n2101 = ~new_n2099 & ~new_n2100;
  assign new_n2102 = \222  & \511 ;
  assign new_n2103 = ~new_n2101 & new_n2102;
  assign new_n2104 = new_n2101 & ~new_n2102;
  assign new_n2105 = ~new_n2103 & ~new_n2104;
  assign new_n2106 = ~new_n2061 & ~new_n2065;
  assign new_n2107 = new_n2105 & ~new_n2106;
  assign new_n2108 = ~new_n2105 & new_n2106;
  assign new_n2109 = ~new_n2107 & ~new_n2108;
  assign new_n2110 = \205  & \528 ;
  assign new_n2111 = ~new_n2109 & new_n2110;
  assign new_n2112 = new_n2109 & ~new_n2110;
  assign new_n2113 = ~new_n2111 & ~new_n2112;
  assign new_n2114 = ~new_n2039 & ~new_n2068;
  assign new_n2115 = new_n2113 & new_n2114;
  assign new_n2116 = ~new_n2113 & ~new_n2114;
  assign new_n2117 = ~new_n2115 & ~new_n2116;
  assign new_n2118 = ~new_n2035 & ~new_n2072;
  assign new_n2119 = ~new_n2071 & ~new_n2118;
  assign new_n2120 = new_n2117 & ~new_n2119;
  assign new_n2121 = ~new_n2117 & new_n2119;
  assign \6260  = new_n2120 | new_n2121;
  assign new_n2123 = \222  & \528 ;
  assign new_n2124 = ~new_n2100 & ~new_n2104;
  assign new_n2125 = ~new_n2123 & ~new_n2124;
  assign new_n2126 = new_n2123 & new_n2124;
  assign new_n2127 = ~new_n2125 & ~new_n2126;
  assign new_n2128 = \239  & \511 ;
  assign new_n2129 = ~\460  & ~\477 ;
  assign new_n2130 = new_n2046 & ~new_n2129;
  assign new_n2131 = ~new_n2077 & ~new_n2130;
  assign new_n2132 = \494  & ~new_n2131;
  assign new_n2133 = ~\460  & ~new_n2046;
  assign new_n2134 = new_n2047 & ~new_n2133;
  assign new_n2135 = ~\494  & ~new_n2134;
  assign new_n2136 = \256  & ~new_n2135;
  assign new_n2137 = ~new_n2132 & new_n2136;
  assign new_n2138 = new_n2128 & ~new_n2137;
  assign new_n2139 = ~new_n2128 & new_n2137;
  assign new_n2140 = ~new_n2138 & ~new_n2139;
  assign new_n2141 = ~new_n2127 & new_n2140;
  assign new_n2142 = new_n2127 & ~new_n2140;
  assign new_n2143 = ~new_n2141 & ~new_n2142;
  assign new_n2144 = ~new_n2107 & ~new_n2112;
  assign new_n2145 = ~new_n2143 & ~new_n2144;
  assign new_n2146 = new_n2143 & new_n2144;
  assign new_n2147 = ~new_n2145 & ~new_n2146;
  assign new_n2148 = ~new_n2115 & new_n2119;
  assign new_n2149 = ~new_n2116 & ~new_n2148;
  assign new_n2150 = new_n2147 & ~new_n2149;
  assign new_n2151 = ~new_n2147 & new_n2149;
  assign \6270  = ~new_n2150 & ~new_n2151;
  assign new_n2153 = ~new_n2126 & ~new_n2142;
  assign new_n2154 = ~\528  & new_n2128;
  assign new_n2155 = ~new_n2135 & new_n2154;
  assign new_n2156 = \256  & \528 ;
  assign new_n2157 = new_n2128 & new_n2156;
  assign new_n2158 = ~\256  & ~\528 ;
  assign new_n2159 = ~new_n2157 & ~new_n2158;
  assign new_n2160 = new_n2135 & ~new_n2159;
  assign new_n2161 = \256  & \511 ;
  assign new_n2162 = ~\239  & ~new_n2161;
  assign new_n2163 = \528  & ~new_n2132;
  assign new_n2164 = ~\528  & new_n2132;
  assign new_n2165 = ~\511  & ~new_n2163;
  assign new_n2166 = ~new_n2164 & new_n2165;
  assign new_n2167 = ~new_n2155 & ~new_n2162;
  assign new_n2168 = ~new_n2160 & new_n2167;
  assign new_n2169 = ~new_n2166 & new_n2168;
  assign new_n2170 = new_n2153 & ~new_n2169;
  assign new_n2171 = ~new_n2153 & new_n2169;
  assign new_n2172 = ~new_n2170 & ~new_n2171;
  assign new_n2173 = ~new_n2146 & ~new_n2150;
  assign new_n2174 = ~new_n2172 & new_n2173;
  assign new_n2175 = new_n2172 & ~new_n2173;
  assign \6280  = ~new_n2174 & ~new_n2175;
  assign new_n2177 = ~\511  & new_n2132;
  assign new_n2178 = ~new_n2128 & ~new_n2177;
  assign new_n2179 = ~new_n2171 & new_n2173;
  assign new_n2180 = ~new_n2170 & ~new_n2179;
  assign new_n2181 = new_n2178 & ~new_n2180;
  assign \6287  = new_n2156 & ~new_n2181;
  assign new_n2183 = new_n2156 & new_n2178;
  assign new_n2184 = new_n2136 & new_n2154;
  assign new_n2185 = ~new_n2183 & ~new_n2184;
  assign new_n2186 = new_n2180 & new_n2185;
  assign new_n2187 = ~new_n2180 & ~new_n2185;
  assign \6288  = new_n2186 | new_n2187;
endmodule


