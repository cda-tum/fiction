// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_, pv118_3_,
    pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_, pv40_14_,
    pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_, pv88_2_,
    pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_, pv88_3_,
    pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_, pv88_13_,
    pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_, pv88_14_,
    pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_, pv100_3_,
    pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_, pv121_3_,
    pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_, pv100_6_,
    pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_, pv28_2_,
    pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_, pv76_10_,
    pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_, pv124_2_,
    pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_, pv52_5_,
    pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_, pv100_9_,
    pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_, pv16_1_,
    pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_, pv106_2_,
    pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_, pv88_1_,
    pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_, pv64_14_,
    pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_, pv115_2_,
    pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_  );
  input  pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_,
    pv118_3_, pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_,
    pv40_14_, pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_,
    pv88_2_, pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_,
    pv88_3_, pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_,
    pv88_13_, pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_,
    pv88_14_, pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_,
    pv100_3_, pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_,
    pv121_3_, pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_,
    pv100_6_, pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_,
    pv28_2_, pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_,
    pv76_10_, pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_,
    pv124_2_, pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_,
    pv52_5_, pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_,
    pv100_9_, pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_,
    pv16_1_, pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_,
    pv106_2_, pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_,
    pv88_1_, pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_,
    pv64_14_, pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_,
    pv115_2_;
  output pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_;
  wire new_n200, new_n201, new_n202, new_n203, new_n205, new_n207, new_n209,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n220, new_n221, new_n222, new_n223, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n234,
    new_n235, new_n236, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n287, new_n289, new_n291,
    new_n292, new_n293, new_n294, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n304, new_n306, new_n308, new_n310,
    new_n311, new_n312, new_n314, new_n315, new_n316, new_n317, new_n319,
    new_n320, new_n321, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n341, new_n342, new_n343,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n354, new_n355, new_n356, new_n357, new_n359, new_n361,
    new_n363, new_n364, new_n365, new_n367, new_n368, new_n369, new_n370,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n380, new_n382, new_n383, new_n384, new_n386, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n396, new_n397,
    new_n398, new_n400, new_n402, new_n403, new_n404, new_n405, new_n407,
    new_n408, new_n409, new_n410, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n420, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n430, new_n431, new_n432,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n443, new_n444, new_n445, new_n446, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n472, new_n474, new_n475,
    new_n476, new_n478, new_n480, new_n482, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n517, new_n519, new_n521,
    new_n523, new_n524, new_n525, new_n526, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534;
  assign new_n200 = pv132_3_ & pv132_2_;
  assign new_n201 = pv133_0_ & new_n200;
  assign new_n202 = pv128_3_ & pv132_2_;
  assign new_n203 = ~pv128_2_ & ~new_n201;
  assign pv183_0_ = new_n202 | ~new_n203;
  assign new_n205 = pv112_3_ & pv183_0_;
  assign pv167_12_ = pv109_3_ | new_n205;
  assign new_n207 = pv52_11_ & pv167_12_;
  assign pv167_11_ = pv40_11_ | new_n207;
  assign new_n209 = pv133_0_ & pv124_3_;
  assign pv199_12_ = pv121_3_ | new_n209;
  assign new_n211 = pv100_10_ & pv100_11_;
  assign new_n212 = pv100_9_ & new_n211;
  assign new_n213 = pv199_12_ & new_n212;
  assign new_n214 = pv88_10_ & pv100_9_;
  assign new_n215 = pv88_11_ & pv100_9_;
  assign new_n216 = pv100_10_ & new_n215;
  assign new_n217 = ~pv88_9_ & ~new_n213;
  assign new_n218 = ~new_n214 & ~new_n216;
  assign pv199_9_ = ~new_n217 | ~new_n218;
  assign new_n220 = pv124_2_ & pv124_3_;
  assign new_n221 = pv133_0_ & new_n220;
  assign new_n222 = pv121_3_ & pv124_2_;
  assign new_n223 = ~pv121_2_ & ~new_n221;
  assign pv199_8_ = new_n222 | ~new_n223;
  assign new_n225 = pv52_14_ & pv52_15_;
  assign new_n226 = pv52_13_ & new_n225;
  assign new_n227 = pv183_0_ & new_n226;
  assign new_n228 = pv40_14_ & pv52_13_;
  assign new_n229 = pv40_15_ & pv52_13_;
  assign new_n230 = pv52_14_ & new_n229;
  assign new_n231 = ~pv40_13_ & ~new_n227;
  assign new_n232 = ~new_n228 & ~new_n230;
  assign pv167_13_ = ~new_n231 | ~new_n232;
  assign new_n234 = pv183_0_ & new_n225;
  assign new_n235 = pv40_15_ & pv52_14_;
  assign new_n236 = ~pv40_14_ & ~new_n234;
  assign pv167_14_ = new_n235 | ~new_n236;
  assign new_n238 = pv132_1_ & new_n200;
  assign new_n239 = pv133_0_ & new_n238;
  assign new_n240 = pv128_2_ & pv132_1_;
  assign new_n241 = pv128_3_ & pv132_1_;
  assign new_n242 = pv132_2_ & new_n241;
  assign new_n243 = ~pv128_1_ & ~new_n239;
  assign new_n244 = ~new_n240 & ~new_n242;
  assign pv167_0_ = ~new_n243 | ~new_n244;
  assign new_n246 = pv106_2_ & pv106_3_;
  assign new_n247 = pv106_1_ & new_n246;
  assign new_n248 = pv167_0_ & new_n247;
  assign new_n249 = pv103_2_ & pv106_1_;
  assign new_n250 = pv103_3_ & pv106_1_;
  assign new_n251 = pv106_2_ & new_n250;
  assign new_n252 = ~pv103_1_ & ~new_n248;
  assign new_n253 = ~new_n249 & ~new_n251;
  assign pv151_4_ = ~new_n252 | ~new_n253;
  assign new_n255 = pv28_2_ & pv28_3_;
  assign new_n256 = pv28_1_ & new_n255;
  assign new_n257 = pv151_4_ & new_n256;
  assign new_n258 = pv28_1_ & pv16_2_;
  assign new_n259 = pv28_1_ & pv16_3_;
  assign new_n260 = pv28_2_ & new_n259;
  assign new_n261 = ~pv16_1_ & ~new_n257;
  assign new_n262 = ~new_n258 & ~new_n260;
  assign pv151_1_ = ~new_n261 | ~new_n262;
  assign new_n264 = pv100_6_ & pv100_7_;
  assign new_n265 = pv100_5_ & new_n264;
  assign new_n266 = pv199_8_ & new_n265;
  assign new_n267 = pv88_6_ & pv100_5_;
  assign new_n268 = pv88_7_ & pv100_5_;
  assign new_n269 = pv100_6_ & new_n268;
  assign new_n270 = ~pv88_5_ & ~new_n266;
  assign new_n271 = ~new_n267 & ~new_n269;
  assign pv199_5_ = ~new_n270 | ~new_n271;
  assign new_n273 = pv128_2_ & pv132_0_;
  assign new_n274 = pv132_1_ & new_n273;
  assign new_n275 = pv132_3_ & pv132_1_;
  assign new_n276 = pv132_2_ & new_n275;
  assign new_n277 = pv132_0_ & new_n276;
  assign new_n278 = pv133_0_ & new_n277;
  assign new_n279 = pv128_1_ & pv132_0_;
  assign new_n280 = pv132_0_ & pv132_1_;
  assign new_n281 = pv128_3_ & new_n280;
  assign new_n282 = pv132_2_ & new_n281;
  assign new_n283 = ~new_n274 & ~new_n278;
  assign new_n284 = ~new_n279 & new_n283;
  assign new_n285 = ~pv128_0_ & ~new_n282;
  assign pv151_0_ = ~new_n284 | ~new_n285;
  assign new_n287 = pv132_3_ & pv133_0_;
  assign pv199_0_ = pv128_3_ | new_n287;
  assign new_n289 = pv118_3_ & pv199_0_;
  assign pv183_12_ = pv115_3_ | new_n289;
  assign new_n291 = pv76_10_ & pv76_11_;
  assign new_n292 = pv183_12_ & new_n291;
  assign new_n293 = pv76_10_ & pv64_11_;
  assign new_n294 = ~pv64_10_ & ~new_n292;
  assign pv183_10_ = new_n293 | ~new_n294;
  assign new_n296 = pv124_1_ & new_n220;
  assign new_n297 = pv133_0_ & new_n296;
  assign new_n298 = pv121_2_ & pv124_1_;
  assign new_n299 = pv121_3_ & pv124_1_;
  assign new_n300 = pv124_2_ & new_n299;
  assign new_n301 = ~pv121_1_ & ~new_n297;
  assign new_n302 = ~new_n298 & ~new_n300;
  assign pv199_4_ = ~new_n301 | ~new_n302;
  assign new_n304 = pv28_3_ & pv151_4_;
  assign pv151_3_ = pv16_3_ | new_n304;
  assign new_n306 = pv76_11_ & pv183_12_;
  assign pv183_11_ = pv64_11_ | new_n306;
  assign new_n308 = pv100_7_ & pv199_8_;
  assign pv199_7_ = pv88_7_ | new_n308;
  assign new_n310 = pv151_4_ & new_n255;
  assign new_n311 = pv28_2_ & pv16_3_;
  assign new_n312 = ~pv16_2_ & ~new_n310;
  assign pv151_2_ = new_n311 | ~new_n312;
  assign new_n314 = pv52_10_ & pv52_11_;
  assign new_n315 = pv167_12_ & new_n314;
  assign new_n316 = pv52_10_ & pv40_11_;
  assign new_n317 = ~pv40_10_ & ~new_n315;
  assign pv167_10_ = new_n316 | ~new_n317;
  assign new_n319 = pv199_8_ & new_n264;
  assign new_n320 = pv88_7_ & pv100_6_;
  assign new_n321 = ~pv88_6_ & ~new_n319;
  assign pv199_6_ = new_n320 | ~new_n321;
  assign new_n323 = pv112_2_ & pv112_3_;
  assign new_n324 = pv112_1_ & new_n323;
  assign new_n325 = pv183_0_ & new_n324;
  assign new_n326 = pv109_2_ & pv112_1_;
  assign new_n327 = pv109_3_ & pv112_1_;
  assign new_n328 = pv112_2_ & new_n327;
  assign new_n329 = ~pv109_1_ & ~new_n325;
  assign new_n330 = ~new_n326 & ~new_n328;
  assign pv167_4_ = ~new_n329 | ~new_n330;
  assign new_n332 = pv100_3_ & pv100_2_;
  assign new_n333 = pv100_1_ & new_n332;
  assign new_n334 = pv199_4_ & new_n333;
  assign new_n335 = pv88_2_ & pv100_1_;
  assign new_n336 = pv88_3_ & pv100_1_;
  assign new_n337 = pv100_2_ & new_n336;
  assign new_n338 = ~pv88_1_ & ~new_n334;
  assign new_n339 = ~new_n335 & ~new_n337;
  assign pv199_1_ = ~new_n338 | ~new_n339;
  assign new_n341 = pv183_0_ & new_n323;
  assign new_n342 = pv109_3_ & pv112_2_;
  assign new_n343 = ~pv109_2_ & ~new_n341;
  assign pv167_8_ = new_n342 | ~new_n343;
  assign new_n345 = pv52_7_ & pv52_6_;
  assign new_n346 = pv52_5_ & new_n345;
  assign new_n347 = pv167_8_ & new_n346;
  assign new_n348 = pv52_5_ & pv40_6_;
  assign new_n349 = pv52_5_ & pv40_7_;
  assign new_n350 = pv52_6_ & new_n349;
  assign new_n351 = ~pv40_5_ & ~new_n347;
  assign new_n352 = ~new_n348 & ~new_n350;
  assign pv167_5_ = ~new_n351 | ~new_n352;
  assign new_n354 = pv52_3_ & pv52_2_;
  assign new_n355 = pv167_4_ & new_n354;
  assign new_n356 = pv52_2_ & pv40_3_;
  assign new_n357 = ~pv40_2_ & ~new_n355;
  assign pv167_2_ = new_n356 | ~new_n357;
  assign new_n359 = pv100_3_ & pv199_4_;
  assign pv199_3_ = pv88_3_ | new_n359;
  assign new_n361 = pv52_3_ & pv167_4_;
  assign pv167_3_ = pv40_3_ | new_n361;
  assign new_n363 = pv199_4_ & new_n332;
  assign new_n364 = pv88_3_ & pv100_2_;
  assign new_n365 = ~pv88_2_ & ~new_n363;
  assign pv199_2_ = new_n364 | ~new_n365;
  assign new_n367 = pv100_14_ & pv100_15_;
  assign new_n368 = pv133_0_ & new_n367;
  assign new_n369 = pv88_15_ & pv100_14_;
  assign new_n370 = ~pv88_14_ & ~new_n368;
  assign pv199_14_ = new_n369 | ~new_n370;
  assign new_n372 = pv52_9_ & new_n314;
  assign new_n373 = pv167_12_ & new_n372;
  assign new_n374 = pv40_10_ & pv52_9_;
  assign new_n375 = pv40_11_ & pv52_9_;
  assign new_n376 = pv52_10_ & new_n375;
  assign new_n377 = ~pv40_9_ & ~new_n373;
  assign new_n378 = ~new_n374 & ~new_n376;
  assign pv167_9_ = ~new_n377 | ~new_n378;
  assign new_n380 = pv100_15_ & pv133_0_;
  assign pv199_15_ = pv88_15_ | new_n380;
  assign new_n382 = pv167_8_ & new_n345;
  assign new_n383 = pv52_6_ & pv40_7_;
  assign new_n384 = ~pv40_6_ & ~new_n382;
  assign pv167_6_ = new_n383 | ~new_n384;
  assign new_n386 = pv52_7_ & pv167_8_;
  assign pv167_7_ = pv40_7_ | new_n386;
  assign new_n388 = pv100_13_ & new_n367;
  assign new_n389 = pv133_0_ & new_n388;
  assign new_n390 = pv100_13_ & pv88_14_;
  assign new_n391 = pv88_15_ & pv100_13_;
  assign new_n392 = pv100_14_ & new_n391;
  assign new_n393 = ~pv88_13_ & ~new_n389;
  assign new_n394 = ~new_n390 & ~new_n392;
  assign pv199_13_ = ~new_n393 | ~new_n394;
  assign new_n396 = pv199_12_ & new_n211;
  assign new_n397 = pv88_11_ & pv100_10_;
  assign new_n398 = ~pv88_10_ & ~new_n396;
  assign pv199_10_ = new_n397 | ~new_n398;
  assign new_n400 = pv100_11_ & pv199_12_;
  assign pv199_11_ = pv88_11_ | new_n400;
  assign new_n402 = pv118_3_ & pv118_2_;
  assign new_n403 = pv199_0_ & new_n402;
  assign new_n404 = pv118_2_ & pv115_3_;
  assign new_n405 = ~pv115_2_ & ~new_n403;
  assign pv183_8_ = new_n404 | ~new_n405;
  assign new_n407 = pv76_7_ & pv76_6_;
  assign new_n408 = pv183_8_ & new_n407;
  assign new_n409 = pv64_7_ & pv76_6_;
  assign new_n410 = ~pv64_6_ & ~new_n408;
  assign pv183_6_ = new_n409 | ~new_n410;
  assign new_n412 = pv52_1_ & new_n354;
  assign new_n413 = pv167_4_ & new_n412;
  assign new_n414 = pv52_1_ & pv40_2_;
  assign new_n415 = pv52_1_ & pv40_3_;
  assign new_n416 = pv52_2_ & new_n415;
  assign new_n417 = ~pv40_1_ & ~new_n413;
  assign new_n418 = ~new_n414 & ~new_n416;
  assign pv167_1_ = ~new_n417 | ~new_n418;
  assign new_n420 = pv76_7_ & pv183_8_;
  assign pv183_7_ = pv64_7_ | new_n420;
  assign new_n422 = pv76_9_ & new_n291;
  assign new_n423 = pv183_12_ & new_n422;
  assign new_n424 = pv64_10_ & pv76_9_;
  assign new_n425 = pv64_11_ & pv76_9_;
  assign new_n426 = pv76_10_ & new_n425;
  assign new_n427 = ~pv64_9_ & ~new_n423;
  assign new_n428 = ~new_n424 & ~new_n426;
  assign pv183_9_ = ~new_n427 | ~new_n428;
  assign new_n430 = pv167_0_ & new_n246;
  assign new_n431 = pv103_3_ & pv106_2_;
  assign new_n432 = ~pv103_2_ & ~new_n430;
  assign pv151_8_ = new_n431 | ~new_n432;
  assign new_n434 = pv28_6_ & pv28_7_;
  assign new_n435 = pv28_5_ & new_n434;
  assign new_n436 = pv151_8_ & new_n435;
  assign new_n437 = pv16_6_ & pv28_5_;
  assign new_n438 = pv16_7_ & pv28_5_;
  assign new_n439 = pv28_6_ & new_n438;
  assign new_n440 = ~pv16_5_ & ~new_n436;
  assign new_n441 = ~new_n437 & ~new_n439;
  assign pv151_5_ = ~new_n440 | ~new_n441;
  assign new_n443 = pv28_15_ & pv28_14_;
  assign new_n444 = pv167_0_ & new_n443;
  assign new_n445 = pv16_15_ & pv28_14_;
  assign new_n446 = ~pv16_14_ & ~new_n444;
  assign pv151_14_ = new_n445 | ~new_n446;
  assign new_n448 = pv118_1_ & new_n402;
  assign new_n449 = pv199_0_ & new_n448;
  assign new_n450 = pv118_1_ & pv115_2_;
  assign new_n451 = pv118_1_ & pv115_3_;
  assign new_n452 = pv118_2_ & new_n451;
  assign new_n453 = ~pv115_1_ & ~new_n449;
  assign new_n454 = ~new_n450 & ~new_n452;
  assign pv183_4_ = ~new_n453 | ~new_n454;
  assign new_n456 = pv76_3_ & pv76_2_;
  assign new_n457 = pv183_4_ & new_n456;
  assign new_n458 = pv76_2_ & pv64_3_;
  assign new_n459 = ~pv64_2_ & ~new_n457;
  assign pv183_2_ = new_n458 | ~new_n459;
  assign new_n461 = pv76_14_ & pv76_15_;
  assign new_n462 = pv76_13_ & new_n461;
  assign new_n463 = pv199_0_ & new_n462;
  assign new_n464 = pv76_13_ & pv64_14_;
  assign new_n465 = pv64_15_ & pv76_13_;
  assign new_n466 = pv76_14_ & new_n465;
  assign new_n467 = ~pv64_13_ & ~new_n463;
  assign new_n468 = ~new_n464 & ~new_n466;
  assign pv183_13_ = ~new_n467 | ~new_n468;
  assign new_n470 = pv28_15_ & pv167_0_;
  assign pv151_15_ = pv16_15_ | new_n470;
  assign new_n472 = pv76_3_ & pv183_4_;
  assign pv183_3_ = pv64_3_ | new_n472;
  assign new_n474 = pv199_0_ & new_n461;
  assign new_n475 = pv76_14_ & pv64_15_;
  assign new_n476 = ~pv64_14_ & ~new_n474;
  assign pv183_14_ = new_n475 | ~new_n476;
  assign new_n478 = pv28_7_ & pv151_8_;
  assign pv151_7_ = pv16_7_ | new_n478;
  assign new_n480 = pv106_3_ & pv167_0_;
  assign pv151_12_ = pv103_3_ | new_n480;
  assign new_n482 = pv76_15_ & pv199_0_;
  assign pv183_15_ = pv64_15_ | new_n482;
  assign new_n484 = pv151_8_ & new_n434;
  assign new_n485 = pv16_7_ & pv28_6_;
  assign new_n486 = ~pv16_6_ & ~new_n484;
  assign pv151_6_ = new_n485 | ~new_n486;
  assign new_n488 = pv28_13_ & new_n443;
  assign new_n489 = pv167_0_ & new_n488;
  assign new_n490 = pv16_14_ & pv28_13_;
  assign new_n491 = pv16_15_ & pv28_13_;
  assign new_n492 = pv28_14_ & new_n491;
  assign new_n493 = ~pv16_13_ & ~new_n489;
  assign new_n494 = ~new_n490 & ~new_n492;
  assign pv151_13_ = ~new_n493 | ~new_n494;
  assign new_n496 = pv76_5_ & new_n407;
  assign new_n497 = pv183_8_ & new_n496;
  assign new_n498 = pv64_6_ & pv76_5_;
  assign new_n499 = pv64_7_ & pv76_5_;
  assign new_n500 = pv76_6_ & new_n499;
  assign new_n501 = ~pv64_5_ & ~new_n497;
  assign new_n502 = ~new_n498 & ~new_n500;
  assign pv183_5_ = ~new_n501 | ~new_n502;
  assign new_n504 = pv28_10_ & pv28_11_;
  assign new_n505 = pv28_9_ & new_n504;
  assign new_n506 = pv151_12_ & new_n505;
  assign new_n507 = pv28_9_ & pv16_10_;
  assign new_n508 = pv28_9_ & pv16_11_;
  assign new_n509 = pv28_10_ & new_n508;
  assign new_n510 = ~pv16_9_ & ~new_n506;
  assign new_n511 = ~new_n507 & ~new_n509;
  assign pv151_9_ = ~new_n510 | ~new_n511;
  assign new_n513 = pv151_12_ & new_n504;
  assign new_n514 = pv28_10_ & pv16_11_;
  assign new_n515 = ~pv16_10_ & ~new_n513;
  assign pv151_10_ = new_n514 | ~new_n515;
  assign new_n517 = pv52_15_ & pv183_0_;
  assign pv167_15_ = pv40_15_ | new_n517;
  assign new_n519 = pv28_11_ & pv151_12_;
  assign pv151_11_ = pv16_11_ | new_n519;
  assign new_n521 = pv4_1_ & pv151_0_;
  assign pv135_1_ = pv2_1_ | new_n521;
  assign new_n523 = pv4_0_ & pv4_1_;
  assign new_n524 = pv151_0_ & new_n523;
  assign new_n525 = pv2_1_ & pv4_0_;
  assign new_n526 = ~pv2_0_ & ~new_n524;
  assign pv135_0_ = new_n525 | ~new_n526;
  assign new_n528 = pv76_1_ & new_n456;
  assign new_n529 = pv183_4_ & new_n528;
  assign new_n530 = pv76_1_ & pv64_2_;
  assign new_n531 = pv76_1_ & pv64_3_;
  assign new_n532 = pv76_2_ & new_n531;
  assign new_n533 = ~pv64_1_ & ~new_n529;
  assign new_n534 = ~new_n530 & ~new_n532;
  assign pv183_1_ = ~new_n533 | ~new_n534;
endmodule


