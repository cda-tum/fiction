// Benchmark "top" written by ABC on Mon Nov 27 17:02:17 2023

module top ( 
    a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15,
    a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29,
    a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43,
    a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57,
    a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71,
    a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85,
    a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99,
    a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111,
    a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123,
    a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4, shift5,
    shift6,
    result0, result1, result2, result3, result4, result5, result6, result7,
    result8, result9, result10, result11, result12, result13, result14,
    result15, result16, result17, result18, result19, result20, result21,
    result22, result23, result24, result25, result26, result27, result28,
    result29, result30, result31, result32, result33, result34, result35,
    result36, result37, result38, result39, result40, result41, result42,
    result43, result44, result45, result46, result47, result48, result49,
    result50, result51, result52, result53, result54, result55, result56,
    result57, result58, result59, result60, result61, result62, result63,
    result64, result65, result66, result67, result68, result69, result70,
    result71, result72, result73, result74, result75, result76, result77,
    result78, result79, result80, result81, result82, result83, result84,
    result85, result86, result87, result88, result89, result90, result91,
    result92, result93, result94, result95, result96, result97, result98,
    result99, result100, result101, result102, result103, result104,
    result105, result106, result107, result108, result109, result110,
    result111, result112, result113, result114, result115, result116,
    result117, result118, result119, result120, result121, result122,
    result123, result124, result125, result126, result127  );
  input  a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14,
    a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28,
    a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42,
    a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56,
    a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70,
    a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84,
    a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98,
    a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110,
    a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122,
    a123, a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4,
    shift5, shift6;
  output result0, result1, result2, result3, result4, result5, result6,
    result7, result8, result9, result10, result11, result12, result13,
    result14, result15, result16, result17, result18, result19, result20,
    result21, result22, result23, result24, result25, result26, result27,
    result28, result29, result30, result31, result32, result33, result34,
    result35, result36, result37, result38, result39, result40, result41,
    result42, result43, result44, result45, result46, result47, result48,
    result49, result50, result51, result52, result53, result54, result55,
    result56, result57, result58, result59, result60, result61, result62,
    result63, result64, result65, result66, result67, result68, result69,
    result70, result71, result72, result73, result74, result75, result76,
    result77, result78, result79, result80, result81, result82, result83,
    result84, result85, result86, result87, result88, result89, result90,
    result91, result92, result93, result94, result95, result96, result97,
    result98, result99, result100, result101, result102, result103,
    result104, result105, result106, result107, result108, result109,
    result110, result111, result112, result113, result114, result115,
    result116, result117, result118, result119, result120, result121,
    result122, result123, result124, result125, result126, result127;
  wire new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2194,
    new_n2195, new_n2196, new_n2197, new_n2198, new_n2199, new_n2200,
    new_n2201, new_n2202, new_n2203, new_n2204, new_n2205, new_n2206,
    new_n2207, new_n2208, new_n2209, new_n2210, new_n2211, new_n2212,
    new_n2213, new_n2214, new_n2215, new_n2216, new_n2217, new_n2218,
    new_n2219, new_n2220, new_n2221, new_n2222, new_n2223, new_n2224,
    new_n2225, new_n2226, new_n2227, new_n2228, new_n2229, new_n2230,
    new_n2231, new_n2232, new_n2233, new_n2234, new_n2235, new_n2236,
    new_n2237, new_n2238, new_n2239, new_n2240, new_n2241, new_n2242,
    new_n2243, new_n2244, new_n2245, new_n2246, new_n2247, new_n2248,
    new_n2249, new_n2250, new_n2251, new_n2252, new_n2253, new_n2254,
    new_n2255, new_n2256, new_n2257, new_n2258, new_n2259, new_n2260,
    new_n2261, new_n2262, new_n2263, new_n2264, new_n2265, new_n2267,
    new_n2268, new_n2269, new_n2270, new_n2271, new_n2272, new_n2273,
    new_n2274, new_n2275, new_n2276, new_n2277, new_n2278, new_n2279,
    new_n2280, new_n2281, new_n2282, new_n2283, new_n2284, new_n2285,
    new_n2286, new_n2287, new_n2288, new_n2289, new_n2290, new_n2291,
    new_n2292, new_n2293, new_n2294, new_n2295, new_n2296, new_n2297,
    new_n2298, new_n2299, new_n2300, new_n2301, new_n2302, new_n2303,
    new_n2304, new_n2305, new_n2306, new_n2307, new_n2308, new_n2309,
    new_n2310, new_n2311, new_n2312, new_n2313, new_n2314, new_n2315,
    new_n2316, new_n2317, new_n2318, new_n2319, new_n2320, new_n2321,
    new_n2322, new_n2323, new_n2324, new_n2325, new_n2326, new_n2327,
    new_n2328, new_n2329, new_n2330, new_n2331, new_n2332, new_n2333,
    new_n2334, new_n2335, new_n2336, new_n2337, new_n2338, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2408, new_n2409, new_n2410,
    new_n2411, new_n2412, new_n2413, new_n2414, new_n2415, new_n2416,
    new_n2417, new_n2418, new_n2419, new_n2420, new_n2421, new_n2422,
    new_n2423, new_n2425, new_n2426, new_n2427, new_n2428, new_n2429,
    new_n2430, new_n2431, new_n2432, new_n2433, new_n2434, new_n2435,
    new_n2436, new_n2437, new_n2438, new_n2439, new_n2440, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2510, new_n2511, new_n2512,
    new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518,
    new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2527, new_n2528, new_n2529, new_n2530, new_n2531,
    new_n2532, new_n2533, new_n2534, new_n2535, new_n2536, new_n2537,
    new_n2538, new_n2539, new_n2540, new_n2541, new_n2542, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2561, new_n2562, new_n2563,
    new_n2564, new_n2565, new_n2566, new_n2567, new_n2568, new_n2569,
    new_n2570, new_n2571, new_n2572, new_n2573, new_n2574, new_n2575,
    new_n2576, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2646,
    new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658,
    new_n2659, new_n2660, new_n2661, new_n2663, new_n2664, new_n2665,
    new_n2666, new_n2667, new_n2668, new_n2669, new_n2670, new_n2671,
    new_n2672, new_n2673, new_n2674, new_n2675, new_n2676, new_n2677,
    new_n2678, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2765, new_n2766, new_n2767,
    new_n2768, new_n2769, new_n2770, new_n2771, new_n2772, new_n2773,
    new_n2774, new_n2775, new_n2776, new_n2777, new_n2778, new_n2779,
    new_n2780, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2867, new_n2868, new_n2869,
    new_n2870, new_n2871, new_n2872, new_n2873, new_n2874, new_n2875,
    new_n2876, new_n2877, new_n2878, new_n2879, new_n2880, new_n2881,
    new_n2882, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2901,
    new_n2902, new_n2903, new_n2904, new_n2905, new_n2906, new_n2907,
    new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913,
    new_n2914, new_n2915, new_n2916, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2969, new_n2970, new_n2971,
    new_n2972, new_n2973, new_n2974, new_n2975, new_n2976, new_n2977,
    new_n2978, new_n2979, new_n2980, new_n2981, new_n2982, new_n2983,
    new_n2984, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3003,
    new_n3004, new_n3005, new_n3006, new_n3007, new_n3008, new_n3009,
    new_n3010, new_n3011, new_n3012, new_n3013, new_n3014, new_n3015,
    new_n3016, new_n3017, new_n3018, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3037, new_n3038, new_n3039, new_n3040, new_n3041,
    new_n3042, new_n3043, new_n3044, new_n3045, new_n3046, new_n3047,
    new_n3048, new_n3049, new_n3050, new_n3051, new_n3052, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3071, new_n3072, new_n3073,
    new_n3074, new_n3075, new_n3076, new_n3077, new_n3078, new_n3079,
    new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085,
    new_n3086, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3105,
    new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111,
    new_n3112, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117,
    new_n3118, new_n3119, new_n3120, new_n3122, new_n3123, new_n3124,
    new_n3125, new_n3126, new_n3127, new_n3128, new_n3129, new_n3130,
    new_n3131, new_n3132, new_n3133, new_n3134, new_n3135, new_n3136,
    new_n3137, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3156,
    new_n3157, new_n3159, new_n3160, new_n3162, new_n3163, new_n3165,
    new_n3166, new_n3168, new_n3169, new_n3171, new_n3172, new_n3174,
    new_n3175, new_n3177, new_n3178, new_n3180, new_n3181, new_n3183,
    new_n3184, new_n3186, new_n3187, new_n3189, new_n3190, new_n3192,
    new_n3193, new_n3195, new_n3196, new_n3198, new_n3199, new_n3201,
    new_n3202, new_n3204, new_n3205, new_n3207, new_n3208, new_n3210,
    new_n3211, new_n3213, new_n3214, new_n3216, new_n3217, new_n3219,
    new_n3220, new_n3222, new_n3223, new_n3225, new_n3226, new_n3228,
    new_n3229, new_n3231, new_n3232, new_n3234, new_n3235, new_n3237,
    new_n3238, new_n3240, new_n3241, new_n3243, new_n3244, new_n3246,
    new_n3247, new_n3249, new_n3250, new_n3252, new_n3253, new_n3255,
    new_n3256, new_n3258, new_n3259, new_n3261, new_n3262, new_n3264,
    new_n3265, new_n3267, new_n3268, new_n3270, new_n3271, new_n3273,
    new_n3274, new_n3276, new_n3277, new_n3279, new_n3280, new_n3282,
    new_n3283, new_n3285, new_n3286, new_n3288, new_n3289, new_n3291,
    new_n3292, new_n3294, new_n3295, new_n3297, new_n3298, new_n3300,
    new_n3301, new_n3303, new_n3304, new_n3306, new_n3307, new_n3309,
    new_n3310, new_n3312, new_n3313, new_n3315, new_n3316, new_n3318,
    new_n3319, new_n3321, new_n3322, new_n3324, new_n3325, new_n3327,
    new_n3328, new_n3330, new_n3331, new_n3333, new_n3334, new_n3336,
    new_n3337, new_n3339, new_n3340, new_n3342, new_n3343, new_n3345,
    new_n3346;
  assign new_n264 = ~shift4 & shift5;
  assign new_n265 = ~shift2 & shift3;
  assign new_n266 = ~shift0 & shift1;
  assign new_n267 = a86 & new_n266;
  assign new_n268 = shift0 & shift1;
  assign new_n269 = a85 & new_n268;
  assign new_n270 = ~shift0 & ~shift1;
  assign new_n271 = a88 & new_n270;
  assign new_n272 = shift0 & ~shift1;
  assign new_n273 = a87 & new_n272;
  assign new_n274 = ~new_n267 & ~new_n269;
  assign new_n275 = ~new_n271 & ~new_n273;
  assign new_n276 = new_n274 & new_n275;
  assign new_n277 = new_n265 & new_n276;
  assign new_n278 = ~shift2 & ~shift3;
  assign new_n279 = a94 & new_n266;
  assign new_n280 = a93 & new_n268;
  assign new_n281 = a96 & new_n270;
  assign new_n282 = a95 & new_n272;
  assign new_n283 = ~new_n279 & ~new_n280;
  assign new_n284 = ~new_n281 & ~new_n282;
  assign new_n285 = new_n283 & new_n284;
  assign new_n286 = new_n278 & new_n285;
  assign new_n287 = shift2 & shift3;
  assign new_n288 = a82 & new_n266;
  assign new_n289 = a81 & new_n268;
  assign new_n290 = a84 & new_n270;
  assign new_n291 = a83 & new_n272;
  assign new_n292 = ~new_n288 & ~new_n289;
  assign new_n293 = ~new_n290 & ~new_n291;
  assign new_n294 = new_n292 & new_n293;
  assign new_n295 = new_n287 & new_n294;
  assign new_n296 = shift2 & ~shift3;
  assign new_n297 = a90 & new_n266;
  assign new_n298 = a89 & new_n268;
  assign new_n299 = a92 & new_n270;
  assign new_n300 = a91 & new_n272;
  assign new_n301 = ~new_n297 & ~new_n298;
  assign new_n302 = ~new_n299 & ~new_n300;
  assign new_n303 = new_n301 & new_n302;
  assign new_n304 = new_n296 & new_n303;
  assign new_n305 = ~new_n277 & ~new_n286;
  assign new_n306 = ~new_n295 & ~new_n304;
  assign new_n307 = new_n305 & new_n306;
  assign new_n308 = new_n264 & ~new_n307;
  assign new_n309 = ~shift4 & ~shift5;
  assign new_n310 = a118 & new_n266;
  assign new_n311 = a117 & new_n268;
  assign new_n312 = a120 & new_n270;
  assign new_n313 = a119 & new_n272;
  assign new_n314 = ~new_n310 & ~new_n311;
  assign new_n315 = ~new_n312 & ~new_n313;
  assign new_n316 = new_n314 & new_n315;
  assign new_n317 = new_n265 & new_n316;
  assign new_n318 = a125 & new_n268;
  assign new_n319 = a0 & new_n270;
  assign new_n320 = a127 & new_n272;
  assign new_n321 = a126 & new_n266;
  assign new_n322 = ~new_n318 & ~new_n319;
  assign new_n323 = ~new_n320 & ~new_n321;
  assign new_n324 = new_n322 & new_n323;
  assign new_n325 = new_n278 & new_n324;
  assign new_n326 = a114 & new_n266;
  assign new_n327 = a113 & new_n268;
  assign new_n328 = a116 & new_n270;
  assign new_n329 = a115 & new_n272;
  assign new_n330 = ~new_n326 & ~new_n327;
  assign new_n331 = ~new_n328 & ~new_n329;
  assign new_n332 = new_n330 & new_n331;
  assign new_n333 = new_n287 & new_n332;
  assign new_n334 = a122 & new_n266;
  assign new_n335 = a121 & new_n268;
  assign new_n336 = a124 & new_n270;
  assign new_n337 = a123 & new_n272;
  assign new_n338 = ~new_n334 & ~new_n335;
  assign new_n339 = ~new_n336 & ~new_n337;
  assign new_n340 = new_n338 & new_n339;
  assign new_n341 = new_n296 & new_n340;
  assign new_n342 = ~new_n317 & ~new_n325;
  assign new_n343 = ~new_n333 & ~new_n341;
  assign new_n344 = new_n342 & new_n343;
  assign new_n345 = new_n309 & ~new_n344;
  assign new_n346 = shift4 & shift5;
  assign new_n347 = a70 & new_n266;
  assign new_n348 = a69 & new_n268;
  assign new_n349 = a72 & new_n270;
  assign new_n350 = a71 & new_n272;
  assign new_n351 = ~new_n347 & ~new_n348;
  assign new_n352 = ~new_n349 & ~new_n350;
  assign new_n353 = new_n351 & new_n352;
  assign new_n354 = new_n265 & new_n353;
  assign new_n355 = a78 & new_n266;
  assign new_n356 = a77 & new_n268;
  assign new_n357 = a80 & new_n270;
  assign new_n358 = a79 & new_n272;
  assign new_n359 = ~new_n355 & ~new_n356;
  assign new_n360 = ~new_n357 & ~new_n358;
  assign new_n361 = new_n359 & new_n360;
  assign new_n362 = new_n278 & new_n361;
  assign new_n363 = a66 & new_n266;
  assign new_n364 = a65 & new_n268;
  assign new_n365 = a68 & new_n270;
  assign new_n366 = a67 & new_n272;
  assign new_n367 = ~new_n363 & ~new_n364;
  assign new_n368 = ~new_n365 & ~new_n366;
  assign new_n369 = new_n367 & new_n368;
  assign new_n370 = new_n287 & new_n369;
  assign new_n371 = a74 & new_n266;
  assign new_n372 = a73 & new_n268;
  assign new_n373 = a76 & new_n270;
  assign new_n374 = a75 & new_n272;
  assign new_n375 = ~new_n371 & ~new_n372;
  assign new_n376 = ~new_n373 & ~new_n374;
  assign new_n377 = new_n375 & new_n376;
  assign new_n378 = new_n296 & new_n377;
  assign new_n379 = ~new_n354 & ~new_n362;
  assign new_n380 = ~new_n370 & ~new_n378;
  assign new_n381 = new_n379 & new_n380;
  assign new_n382 = new_n346 & ~new_n381;
  assign new_n383 = shift4 & ~shift5;
  assign new_n384 = a102 & new_n266;
  assign new_n385 = a101 & new_n268;
  assign new_n386 = a104 & new_n270;
  assign new_n387 = a103 & new_n272;
  assign new_n388 = ~new_n384 & ~new_n385;
  assign new_n389 = ~new_n386 & ~new_n387;
  assign new_n390 = new_n388 & new_n389;
  assign new_n391 = new_n265 & new_n390;
  assign new_n392 = a110 & new_n266;
  assign new_n393 = a109 & new_n268;
  assign new_n394 = a112 & new_n270;
  assign new_n395 = a111 & new_n272;
  assign new_n396 = ~new_n392 & ~new_n393;
  assign new_n397 = ~new_n394 & ~new_n395;
  assign new_n398 = new_n396 & new_n397;
  assign new_n399 = new_n278 & new_n398;
  assign new_n400 = a98 & new_n266;
  assign new_n401 = a97 & new_n268;
  assign new_n402 = a100 & new_n270;
  assign new_n403 = a99 & new_n272;
  assign new_n404 = ~new_n400 & ~new_n401;
  assign new_n405 = ~new_n402 & ~new_n403;
  assign new_n406 = new_n404 & new_n405;
  assign new_n407 = new_n287 & new_n406;
  assign new_n408 = a106 & new_n266;
  assign new_n409 = a105 & new_n268;
  assign new_n410 = a108 & new_n270;
  assign new_n411 = a107 & new_n272;
  assign new_n412 = ~new_n408 & ~new_n409;
  assign new_n413 = ~new_n410 & ~new_n411;
  assign new_n414 = new_n412 & new_n413;
  assign new_n415 = new_n296 & new_n414;
  assign new_n416 = ~new_n391 & ~new_n399;
  assign new_n417 = ~new_n407 & ~new_n415;
  assign new_n418 = new_n416 & new_n417;
  assign new_n419 = new_n383 & ~new_n418;
  assign new_n420 = ~new_n308 & ~new_n345;
  assign new_n421 = ~new_n382 & ~new_n419;
  assign new_n422 = new_n420 & new_n421;
  assign new_n423 = ~shift6 & ~new_n422;
  assign new_n424 = a22 & new_n266;
  assign new_n425 = a21 & new_n268;
  assign new_n426 = a24 & new_n270;
  assign new_n427 = a23 & new_n272;
  assign new_n428 = ~new_n424 & ~new_n425;
  assign new_n429 = ~new_n426 & ~new_n427;
  assign new_n430 = new_n428 & new_n429;
  assign new_n431 = new_n265 & new_n430;
  assign new_n432 = a30 & new_n266;
  assign new_n433 = a29 & new_n268;
  assign new_n434 = a32 & new_n270;
  assign new_n435 = a31 & new_n272;
  assign new_n436 = ~new_n432 & ~new_n433;
  assign new_n437 = ~new_n434 & ~new_n435;
  assign new_n438 = new_n436 & new_n437;
  assign new_n439 = new_n278 & new_n438;
  assign new_n440 = a18 & new_n266;
  assign new_n441 = a17 & new_n268;
  assign new_n442 = a20 & new_n270;
  assign new_n443 = a19 & new_n272;
  assign new_n444 = ~new_n440 & ~new_n441;
  assign new_n445 = ~new_n442 & ~new_n443;
  assign new_n446 = new_n444 & new_n445;
  assign new_n447 = new_n287 & new_n446;
  assign new_n448 = a26 & new_n266;
  assign new_n449 = a25 & new_n268;
  assign new_n450 = a28 & new_n270;
  assign new_n451 = a27 & new_n272;
  assign new_n452 = ~new_n448 & ~new_n449;
  assign new_n453 = ~new_n450 & ~new_n451;
  assign new_n454 = new_n452 & new_n453;
  assign new_n455 = new_n296 & new_n454;
  assign new_n456 = ~new_n431 & ~new_n439;
  assign new_n457 = ~new_n447 & ~new_n455;
  assign new_n458 = new_n456 & new_n457;
  assign new_n459 = new_n264 & ~new_n458;
  assign new_n460 = a54 & new_n266;
  assign new_n461 = a53 & new_n268;
  assign new_n462 = a56 & new_n270;
  assign new_n463 = a55 & new_n272;
  assign new_n464 = ~new_n460 & ~new_n461;
  assign new_n465 = ~new_n462 & ~new_n463;
  assign new_n466 = new_n464 & new_n465;
  assign new_n467 = new_n265 & new_n466;
  assign new_n468 = a62 & new_n266;
  assign new_n469 = a61 & new_n268;
  assign new_n470 = a64 & new_n270;
  assign new_n471 = a63 & new_n272;
  assign new_n472 = ~new_n468 & ~new_n469;
  assign new_n473 = ~new_n470 & ~new_n471;
  assign new_n474 = new_n472 & new_n473;
  assign new_n475 = new_n278 & new_n474;
  assign new_n476 = a50 & new_n266;
  assign new_n477 = a49 & new_n268;
  assign new_n478 = a52 & new_n270;
  assign new_n479 = a51 & new_n272;
  assign new_n480 = ~new_n476 & ~new_n477;
  assign new_n481 = ~new_n478 & ~new_n479;
  assign new_n482 = new_n480 & new_n481;
  assign new_n483 = new_n287 & new_n482;
  assign new_n484 = a58 & new_n266;
  assign new_n485 = a57 & new_n268;
  assign new_n486 = a60 & new_n270;
  assign new_n487 = a59 & new_n272;
  assign new_n488 = ~new_n484 & ~new_n485;
  assign new_n489 = ~new_n486 & ~new_n487;
  assign new_n490 = new_n488 & new_n489;
  assign new_n491 = new_n296 & new_n490;
  assign new_n492 = ~new_n467 & ~new_n475;
  assign new_n493 = ~new_n483 & ~new_n491;
  assign new_n494 = new_n492 & new_n493;
  assign new_n495 = new_n309 & ~new_n494;
  assign new_n496 = a6 & new_n266;
  assign new_n497 = a5 & new_n268;
  assign new_n498 = a8 & new_n270;
  assign new_n499 = a7 & new_n272;
  assign new_n500 = ~new_n496 & ~new_n497;
  assign new_n501 = ~new_n498 & ~new_n499;
  assign new_n502 = new_n500 & new_n501;
  assign new_n503 = new_n265 & new_n502;
  assign new_n504 = a14 & new_n266;
  assign new_n505 = a13 & new_n268;
  assign new_n506 = a16 & new_n270;
  assign new_n507 = a15 & new_n272;
  assign new_n508 = ~new_n504 & ~new_n505;
  assign new_n509 = ~new_n506 & ~new_n507;
  assign new_n510 = new_n508 & new_n509;
  assign new_n511 = new_n278 & new_n510;
  assign new_n512 = a2 & new_n266;
  assign new_n513 = a1 & new_n268;
  assign new_n514 = a4 & new_n270;
  assign new_n515 = a3 & new_n272;
  assign new_n516 = ~new_n512 & ~new_n513;
  assign new_n517 = ~new_n514 & ~new_n515;
  assign new_n518 = new_n516 & new_n517;
  assign new_n519 = new_n287 & new_n518;
  assign new_n520 = a10 & new_n266;
  assign new_n521 = a9 & new_n268;
  assign new_n522 = a12 & new_n270;
  assign new_n523 = a11 & new_n272;
  assign new_n524 = ~new_n520 & ~new_n521;
  assign new_n525 = ~new_n522 & ~new_n523;
  assign new_n526 = new_n524 & new_n525;
  assign new_n527 = new_n296 & new_n526;
  assign new_n528 = ~new_n503 & ~new_n511;
  assign new_n529 = ~new_n519 & ~new_n527;
  assign new_n530 = new_n528 & new_n529;
  assign new_n531 = new_n346 & ~new_n530;
  assign new_n532 = a38 & new_n266;
  assign new_n533 = a37 & new_n268;
  assign new_n534 = a40 & new_n270;
  assign new_n535 = a39 & new_n272;
  assign new_n536 = ~new_n532 & ~new_n533;
  assign new_n537 = ~new_n534 & ~new_n535;
  assign new_n538 = new_n536 & new_n537;
  assign new_n539 = new_n265 & new_n538;
  assign new_n540 = a46 & new_n266;
  assign new_n541 = a45 & new_n268;
  assign new_n542 = a48 & new_n270;
  assign new_n543 = a47 & new_n272;
  assign new_n544 = ~new_n540 & ~new_n541;
  assign new_n545 = ~new_n542 & ~new_n543;
  assign new_n546 = new_n544 & new_n545;
  assign new_n547 = new_n278 & new_n546;
  assign new_n548 = a34 & new_n266;
  assign new_n549 = a33 & new_n268;
  assign new_n550 = a36 & new_n270;
  assign new_n551 = a35 & new_n272;
  assign new_n552 = ~new_n548 & ~new_n549;
  assign new_n553 = ~new_n550 & ~new_n551;
  assign new_n554 = new_n552 & new_n553;
  assign new_n555 = new_n287 & new_n554;
  assign new_n556 = a42 & new_n266;
  assign new_n557 = a41 & new_n268;
  assign new_n558 = a44 & new_n270;
  assign new_n559 = a43 & new_n272;
  assign new_n560 = ~new_n556 & ~new_n557;
  assign new_n561 = ~new_n558 & ~new_n559;
  assign new_n562 = new_n560 & new_n561;
  assign new_n563 = new_n296 & new_n562;
  assign new_n564 = ~new_n539 & ~new_n547;
  assign new_n565 = ~new_n555 & ~new_n563;
  assign new_n566 = new_n564 & new_n565;
  assign new_n567 = new_n383 & ~new_n566;
  assign new_n568 = ~new_n459 & ~new_n495;
  assign new_n569 = ~new_n531 & ~new_n567;
  assign new_n570 = new_n568 & new_n569;
  assign new_n571 = shift6 & ~new_n570;
  assign result0 = ~new_n423 & ~new_n571;
  assign new_n573 = a87 & new_n266;
  assign new_n574 = a86 & new_n268;
  assign new_n575 = a89 & new_n270;
  assign new_n576 = a88 & new_n272;
  assign new_n577 = ~new_n573 & ~new_n574;
  assign new_n578 = ~new_n575 & ~new_n576;
  assign new_n579 = new_n577 & new_n578;
  assign new_n580 = new_n265 & new_n579;
  assign new_n581 = a95 & new_n266;
  assign new_n582 = a94 & new_n268;
  assign new_n583 = a97 & new_n270;
  assign new_n584 = a96 & new_n272;
  assign new_n585 = ~new_n581 & ~new_n582;
  assign new_n586 = ~new_n583 & ~new_n584;
  assign new_n587 = new_n585 & new_n586;
  assign new_n588 = new_n278 & new_n587;
  assign new_n589 = a83 & new_n266;
  assign new_n590 = a82 & new_n268;
  assign new_n591 = a85 & new_n270;
  assign new_n592 = a84 & new_n272;
  assign new_n593 = ~new_n589 & ~new_n590;
  assign new_n594 = ~new_n591 & ~new_n592;
  assign new_n595 = new_n593 & new_n594;
  assign new_n596 = new_n287 & new_n595;
  assign new_n597 = a91 & new_n266;
  assign new_n598 = a90 & new_n268;
  assign new_n599 = a93 & new_n270;
  assign new_n600 = a92 & new_n272;
  assign new_n601 = ~new_n597 & ~new_n598;
  assign new_n602 = ~new_n599 & ~new_n600;
  assign new_n603 = new_n601 & new_n602;
  assign new_n604 = new_n296 & new_n603;
  assign new_n605 = ~new_n580 & ~new_n588;
  assign new_n606 = ~new_n596 & ~new_n604;
  assign new_n607 = new_n605 & new_n606;
  assign new_n608 = new_n264 & ~new_n607;
  assign new_n609 = a119 & new_n266;
  assign new_n610 = a118 & new_n268;
  assign new_n611 = a121 & new_n270;
  assign new_n612 = a120 & new_n272;
  assign new_n613 = ~new_n609 & ~new_n610;
  assign new_n614 = ~new_n611 & ~new_n612;
  assign new_n615 = new_n613 & new_n614;
  assign new_n616 = new_n265 & new_n615;
  assign new_n617 = a1 & new_n270;
  assign new_n618 = a0 & new_n272;
  assign new_n619 = a127 & new_n266;
  assign new_n620 = a126 & new_n268;
  assign new_n621 = ~new_n617 & ~new_n618;
  assign new_n622 = ~new_n619 & ~new_n620;
  assign new_n623 = new_n621 & new_n622;
  assign new_n624 = new_n278 & new_n623;
  assign new_n625 = a115 & new_n266;
  assign new_n626 = a114 & new_n268;
  assign new_n627 = a117 & new_n270;
  assign new_n628 = a116 & new_n272;
  assign new_n629 = ~new_n625 & ~new_n626;
  assign new_n630 = ~new_n627 & ~new_n628;
  assign new_n631 = new_n629 & new_n630;
  assign new_n632 = new_n287 & new_n631;
  assign new_n633 = a123 & new_n266;
  assign new_n634 = a122 & new_n268;
  assign new_n635 = a125 & new_n270;
  assign new_n636 = a124 & new_n272;
  assign new_n637 = ~new_n633 & ~new_n634;
  assign new_n638 = ~new_n635 & ~new_n636;
  assign new_n639 = new_n637 & new_n638;
  assign new_n640 = new_n296 & new_n639;
  assign new_n641 = ~new_n616 & ~new_n624;
  assign new_n642 = ~new_n632 & ~new_n640;
  assign new_n643 = new_n641 & new_n642;
  assign new_n644 = new_n309 & ~new_n643;
  assign new_n645 = a71 & new_n266;
  assign new_n646 = a70 & new_n268;
  assign new_n647 = a73 & new_n270;
  assign new_n648 = a72 & new_n272;
  assign new_n649 = ~new_n645 & ~new_n646;
  assign new_n650 = ~new_n647 & ~new_n648;
  assign new_n651 = new_n649 & new_n650;
  assign new_n652 = new_n265 & new_n651;
  assign new_n653 = a79 & new_n266;
  assign new_n654 = a78 & new_n268;
  assign new_n655 = a81 & new_n270;
  assign new_n656 = a80 & new_n272;
  assign new_n657 = ~new_n653 & ~new_n654;
  assign new_n658 = ~new_n655 & ~new_n656;
  assign new_n659 = new_n657 & new_n658;
  assign new_n660 = new_n278 & new_n659;
  assign new_n661 = a67 & new_n266;
  assign new_n662 = a66 & new_n268;
  assign new_n663 = a69 & new_n270;
  assign new_n664 = a68 & new_n272;
  assign new_n665 = ~new_n661 & ~new_n662;
  assign new_n666 = ~new_n663 & ~new_n664;
  assign new_n667 = new_n665 & new_n666;
  assign new_n668 = new_n287 & new_n667;
  assign new_n669 = a75 & new_n266;
  assign new_n670 = a74 & new_n268;
  assign new_n671 = a77 & new_n270;
  assign new_n672 = a76 & new_n272;
  assign new_n673 = ~new_n669 & ~new_n670;
  assign new_n674 = ~new_n671 & ~new_n672;
  assign new_n675 = new_n673 & new_n674;
  assign new_n676 = new_n296 & new_n675;
  assign new_n677 = ~new_n652 & ~new_n660;
  assign new_n678 = ~new_n668 & ~new_n676;
  assign new_n679 = new_n677 & new_n678;
  assign new_n680 = new_n346 & ~new_n679;
  assign new_n681 = a103 & new_n266;
  assign new_n682 = a102 & new_n268;
  assign new_n683 = a105 & new_n270;
  assign new_n684 = a104 & new_n272;
  assign new_n685 = ~new_n681 & ~new_n682;
  assign new_n686 = ~new_n683 & ~new_n684;
  assign new_n687 = new_n685 & new_n686;
  assign new_n688 = new_n265 & new_n687;
  assign new_n689 = a111 & new_n266;
  assign new_n690 = a110 & new_n268;
  assign new_n691 = a113 & new_n270;
  assign new_n692 = a112 & new_n272;
  assign new_n693 = ~new_n689 & ~new_n690;
  assign new_n694 = ~new_n691 & ~new_n692;
  assign new_n695 = new_n693 & new_n694;
  assign new_n696 = new_n278 & new_n695;
  assign new_n697 = a99 & new_n266;
  assign new_n698 = a98 & new_n268;
  assign new_n699 = a101 & new_n270;
  assign new_n700 = a100 & new_n272;
  assign new_n701 = ~new_n697 & ~new_n698;
  assign new_n702 = ~new_n699 & ~new_n700;
  assign new_n703 = new_n701 & new_n702;
  assign new_n704 = new_n287 & new_n703;
  assign new_n705 = a107 & new_n266;
  assign new_n706 = a106 & new_n268;
  assign new_n707 = a109 & new_n270;
  assign new_n708 = a108 & new_n272;
  assign new_n709 = ~new_n705 & ~new_n706;
  assign new_n710 = ~new_n707 & ~new_n708;
  assign new_n711 = new_n709 & new_n710;
  assign new_n712 = new_n296 & new_n711;
  assign new_n713 = ~new_n688 & ~new_n696;
  assign new_n714 = ~new_n704 & ~new_n712;
  assign new_n715 = new_n713 & new_n714;
  assign new_n716 = new_n383 & ~new_n715;
  assign new_n717 = ~new_n608 & ~new_n644;
  assign new_n718 = ~new_n680 & ~new_n716;
  assign new_n719 = new_n717 & new_n718;
  assign new_n720 = ~shift6 & ~new_n719;
  assign new_n721 = a23 & new_n266;
  assign new_n722 = a22 & new_n268;
  assign new_n723 = a25 & new_n270;
  assign new_n724 = a24 & new_n272;
  assign new_n725 = ~new_n721 & ~new_n722;
  assign new_n726 = ~new_n723 & ~new_n724;
  assign new_n727 = new_n725 & new_n726;
  assign new_n728 = new_n265 & new_n727;
  assign new_n729 = a31 & new_n266;
  assign new_n730 = a30 & new_n268;
  assign new_n731 = a33 & new_n270;
  assign new_n732 = a32 & new_n272;
  assign new_n733 = ~new_n729 & ~new_n730;
  assign new_n734 = ~new_n731 & ~new_n732;
  assign new_n735 = new_n733 & new_n734;
  assign new_n736 = new_n278 & new_n735;
  assign new_n737 = a19 & new_n266;
  assign new_n738 = a18 & new_n268;
  assign new_n739 = a21 & new_n270;
  assign new_n740 = a20 & new_n272;
  assign new_n741 = ~new_n737 & ~new_n738;
  assign new_n742 = ~new_n739 & ~new_n740;
  assign new_n743 = new_n741 & new_n742;
  assign new_n744 = new_n287 & new_n743;
  assign new_n745 = a27 & new_n266;
  assign new_n746 = a26 & new_n268;
  assign new_n747 = a29 & new_n270;
  assign new_n748 = a28 & new_n272;
  assign new_n749 = ~new_n745 & ~new_n746;
  assign new_n750 = ~new_n747 & ~new_n748;
  assign new_n751 = new_n749 & new_n750;
  assign new_n752 = new_n296 & new_n751;
  assign new_n753 = ~new_n728 & ~new_n736;
  assign new_n754 = ~new_n744 & ~new_n752;
  assign new_n755 = new_n753 & new_n754;
  assign new_n756 = new_n264 & ~new_n755;
  assign new_n757 = a55 & new_n266;
  assign new_n758 = a54 & new_n268;
  assign new_n759 = a57 & new_n270;
  assign new_n760 = a56 & new_n272;
  assign new_n761 = ~new_n757 & ~new_n758;
  assign new_n762 = ~new_n759 & ~new_n760;
  assign new_n763 = new_n761 & new_n762;
  assign new_n764 = new_n265 & new_n763;
  assign new_n765 = a63 & new_n266;
  assign new_n766 = a62 & new_n268;
  assign new_n767 = a65 & new_n270;
  assign new_n768 = a64 & new_n272;
  assign new_n769 = ~new_n765 & ~new_n766;
  assign new_n770 = ~new_n767 & ~new_n768;
  assign new_n771 = new_n769 & new_n770;
  assign new_n772 = new_n278 & new_n771;
  assign new_n773 = a51 & new_n266;
  assign new_n774 = a50 & new_n268;
  assign new_n775 = a53 & new_n270;
  assign new_n776 = a52 & new_n272;
  assign new_n777 = ~new_n773 & ~new_n774;
  assign new_n778 = ~new_n775 & ~new_n776;
  assign new_n779 = new_n777 & new_n778;
  assign new_n780 = new_n287 & new_n779;
  assign new_n781 = a59 & new_n266;
  assign new_n782 = a58 & new_n268;
  assign new_n783 = a61 & new_n270;
  assign new_n784 = a60 & new_n272;
  assign new_n785 = ~new_n781 & ~new_n782;
  assign new_n786 = ~new_n783 & ~new_n784;
  assign new_n787 = new_n785 & new_n786;
  assign new_n788 = new_n296 & new_n787;
  assign new_n789 = ~new_n764 & ~new_n772;
  assign new_n790 = ~new_n780 & ~new_n788;
  assign new_n791 = new_n789 & new_n790;
  assign new_n792 = new_n309 & ~new_n791;
  assign new_n793 = a7 & new_n266;
  assign new_n794 = a6 & new_n268;
  assign new_n795 = a9 & new_n270;
  assign new_n796 = a8 & new_n272;
  assign new_n797 = ~new_n793 & ~new_n794;
  assign new_n798 = ~new_n795 & ~new_n796;
  assign new_n799 = new_n797 & new_n798;
  assign new_n800 = new_n265 & new_n799;
  assign new_n801 = a15 & new_n266;
  assign new_n802 = a14 & new_n268;
  assign new_n803 = a17 & new_n270;
  assign new_n804 = a16 & new_n272;
  assign new_n805 = ~new_n801 & ~new_n802;
  assign new_n806 = ~new_n803 & ~new_n804;
  assign new_n807 = new_n805 & new_n806;
  assign new_n808 = new_n278 & new_n807;
  assign new_n809 = a3 & new_n266;
  assign new_n810 = a2 & new_n268;
  assign new_n811 = a5 & new_n270;
  assign new_n812 = a4 & new_n272;
  assign new_n813 = ~new_n809 & ~new_n810;
  assign new_n814 = ~new_n811 & ~new_n812;
  assign new_n815 = new_n813 & new_n814;
  assign new_n816 = new_n287 & new_n815;
  assign new_n817 = a11 & new_n266;
  assign new_n818 = a10 & new_n268;
  assign new_n819 = a13 & new_n270;
  assign new_n820 = a12 & new_n272;
  assign new_n821 = ~new_n817 & ~new_n818;
  assign new_n822 = ~new_n819 & ~new_n820;
  assign new_n823 = new_n821 & new_n822;
  assign new_n824 = new_n296 & new_n823;
  assign new_n825 = ~new_n800 & ~new_n808;
  assign new_n826 = ~new_n816 & ~new_n824;
  assign new_n827 = new_n825 & new_n826;
  assign new_n828 = new_n346 & ~new_n827;
  assign new_n829 = a39 & new_n266;
  assign new_n830 = a38 & new_n268;
  assign new_n831 = a41 & new_n270;
  assign new_n832 = a40 & new_n272;
  assign new_n833 = ~new_n829 & ~new_n830;
  assign new_n834 = ~new_n831 & ~new_n832;
  assign new_n835 = new_n833 & new_n834;
  assign new_n836 = new_n265 & new_n835;
  assign new_n837 = a47 & new_n266;
  assign new_n838 = a46 & new_n268;
  assign new_n839 = a49 & new_n270;
  assign new_n840 = a48 & new_n272;
  assign new_n841 = ~new_n837 & ~new_n838;
  assign new_n842 = ~new_n839 & ~new_n840;
  assign new_n843 = new_n841 & new_n842;
  assign new_n844 = new_n278 & new_n843;
  assign new_n845 = a35 & new_n266;
  assign new_n846 = a34 & new_n268;
  assign new_n847 = a37 & new_n270;
  assign new_n848 = a36 & new_n272;
  assign new_n849 = ~new_n845 & ~new_n846;
  assign new_n850 = ~new_n847 & ~new_n848;
  assign new_n851 = new_n849 & new_n850;
  assign new_n852 = new_n287 & new_n851;
  assign new_n853 = a43 & new_n266;
  assign new_n854 = a42 & new_n268;
  assign new_n855 = a45 & new_n270;
  assign new_n856 = a44 & new_n272;
  assign new_n857 = ~new_n853 & ~new_n854;
  assign new_n858 = ~new_n855 & ~new_n856;
  assign new_n859 = new_n857 & new_n858;
  assign new_n860 = new_n296 & new_n859;
  assign new_n861 = ~new_n836 & ~new_n844;
  assign new_n862 = ~new_n852 & ~new_n860;
  assign new_n863 = new_n861 & new_n862;
  assign new_n864 = new_n383 & ~new_n863;
  assign new_n865 = ~new_n756 & ~new_n792;
  assign new_n866 = ~new_n828 & ~new_n864;
  assign new_n867 = new_n865 & new_n866;
  assign new_n868 = shift6 & ~new_n867;
  assign result1 = ~new_n720 & ~new_n868;
  assign new_n870 = a88 & new_n266;
  assign new_n871 = a87 & new_n268;
  assign new_n872 = a90 & new_n270;
  assign new_n873 = a89 & new_n272;
  assign new_n874 = ~new_n870 & ~new_n871;
  assign new_n875 = ~new_n872 & ~new_n873;
  assign new_n876 = new_n874 & new_n875;
  assign new_n877 = new_n265 & new_n876;
  assign new_n878 = a96 & new_n266;
  assign new_n879 = a95 & new_n268;
  assign new_n880 = a98 & new_n270;
  assign new_n881 = a97 & new_n272;
  assign new_n882 = ~new_n878 & ~new_n879;
  assign new_n883 = ~new_n880 & ~new_n881;
  assign new_n884 = new_n882 & new_n883;
  assign new_n885 = new_n278 & new_n884;
  assign new_n886 = a84 & new_n266;
  assign new_n887 = a83 & new_n268;
  assign new_n888 = a86 & new_n270;
  assign new_n889 = a85 & new_n272;
  assign new_n890 = ~new_n886 & ~new_n887;
  assign new_n891 = ~new_n888 & ~new_n889;
  assign new_n892 = new_n890 & new_n891;
  assign new_n893 = new_n287 & new_n892;
  assign new_n894 = a92 & new_n266;
  assign new_n895 = a91 & new_n268;
  assign new_n896 = a94 & new_n270;
  assign new_n897 = a93 & new_n272;
  assign new_n898 = ~new_n894 & ~new_n895;
  assign new_n899 = ~new_n896 & ~new_n897;
  assign new_n900 = new_n898 & new_n899;
  assign new_n901 = new_n296 & new_n900;
  assign new_n902 = ~new_n877 & ~new_n885;
  assign new_n903 = ~new_n893 & ~new_n901;
  assign new_n904 = new_n902 & new_n903;
  assign new_n905 = new_n264 & ~new_n904;
  assign new_n906 = a120 & new_n266;
  assign new_n907 = a119 & new_n268;
  assign new_n908 = a122 & new_n270;
  assign new_n909 = a121 & new_n272;
  assign new_n910 = ~new_n906 & ~new_n907;
  assign new_n911 = ~new_n908 & ~new_n909;
  assign new_n912 = new_n910 & new_n911;
  assign new_n913 = new_n265 & new_n912;
  assign new_n914 = a1 & new_n272;
  assign new_n915 = a0 & new_n266;
  assign new_n916 = a127 & new_n268;
  assign new_n917 = a2 & new_n270;
  assign new_n918 = ~new_n914 & ~new_n915;
  assign new_n919 = ~new_n916 & ~new_n917;
  assign new_n920 = new_n918 & new_n919;
  assign new_n921 = new_n278 & new_n920;
  assign new_n922 = a116 & new_n266;
  assign new_n923 = a115 & new_n268;
  assign new_n924 = a118 & new_n270;
  assign new_n925 = a117 & new_n272;
  assign new_n926 = ~new_n922 & ~new_n923;
  assign new_n927 = ~new_n924 & ~new_n925;
  assign new_n928 = new_n926 & new_n927;
  assign new_n929 = new_n287 & new_n928;
  assign new_n930 = a124 & new_n266;
  assign new_n931 = a123 & new_n268;
  assign new_n932 = a126 & new_n270;
  assign new_n933 = a125 & new_n272;
  assign new_n934 = ~new_n930 & ~new_n931;
  assign new_n935 = ~new_n932 & ~new_n933;
  assign new_n936 = new_n934 & new_n935;
  assign new_n937 = new_n296 & new_n936;
  assign new_n938 = ~new_n913 & ~new_n921;
  assign new_n939 = ~new_n929 & ~new_n937;
  assign new_n940 = new_n938 & new_n939;
  assign new_n941 = new_n309 & ~new_n940;
  assign new_n942 = a72 & new_n266;
  assign new_n943 = a71 & new_n268;
  assign new_n944 = a74 & new_n270;
  assign new_n945 = a73 & new_n272;
  assign new_n946 = ~new_n942 & ~new_n943;
  assign new_n947 = ~new_n944 & ~new_n945;
  assign new_n948 = new_n946 & new_n947;
  assign new_n949 = new_n265 & new_n948;
  assign new_n950 = a80 & new_n266;
  assign new_n951 = a79 & new_n268;
  assign new_n952 = a82 & new_n270;
  assign new_n953 = a81 & new_n272;
  assign new_n954 = ~new_n950 & ~new_n951;
  assign new_n955 = ~new_n952 & ~new_n953;
  assign new_n956 = new_n954 & new_n955;
  assign new_n957 = new_n278 & new_n956;
  assign new_n958 = a68 & new_n266;
  assign new_n959 = a67 & new_n268;
  assign new_n960 = a70 & new_n270;
  assign new_n961 = a69 & new_n272;
  assign new_n962 = ~new_n958 & ~new_n959;
  assign new_n963 = ~new_n960 & ~new_n961;
  assign new_n964 = new_n962 & new_n963;
  assign new_n965 = new_n287 & new_n964;
  assign new_n966 = a76 & new_n266;
  assign new_n967 = a75 & new_n268;
  assign new_n968 = a78 & new_n270;
  assign new_n969 = a77 & new_n272;
  assign new_n970 = ~new_n966 & ~new_n967;
  assign new_n971 = ~new_n968 & ~new_n969;
  assign new_n972 = new_n970 & new_n971;
  assign new_n973 = new_n296 & new_n972;
  assign new_n974 = ~new_n949 & ~new_n957;
  assign new_n975 = ~new_n965 & ~new_n973;
  assign new_n976 = new_n974 & new_n975;
  assign new_n977 = new_n346 & ~new_n976;
  assign new_n978 = a104 & new_n266;
  assign new_n979 = a103 & new_n268;
  assign new_n980 = a106 & new_n270;
  assign new_n981 = a105 & new_n272;
  assign new_n982 = ~new_n978 & ~new_n979;
  assign new_n983 = ~new_n980 & ~new_n981;
  assign new_n984 = new_n982 & new_n983;
  assign new_n985 = new_n265 & new_n984;
  assign new_n986 = a112 & new_n266;
  assign new_n987 = a111 & new_n268;
  assign new_n988 = a114 & new_n270;
  assign new_n989 = a113 & new_n272;
  assign new_n990 = ~new_n986 & ~new_n987;
  assign new_n991 = ~new_n988 & ~new_n989;
  assign new_n992 = new_n990 & new_n991;
  assign new_n993 = new_n278 & new_n992;
  assign new_n994 = a100 & new_n266;
  assign new_n995 = a99 & new_n268;
  assign new_n996 = a102 & new_n270;
  assign new_n997 = a101 & new_n272;
  assign new_n998 = ~new_n994 & ~new_n995;
  assign new_n999 = ~new_n996 & ~new_n997;
  assign new_n1000 = new_n998 & new_n999;
  assign new_n1001 = new_n287 & new_n1000;
  assign new_n1002 = a108 & new_n266;
  assign new_n1003 = a107 & new_n268;
  assign new_n1004 = a110 & new_n270;
  assign new_n1005 = a109 & new_n272;
  assign new_n1006 = ~new_n1002 & ~new_n1003;
  assign new_n1007 = ~new_n1004 & ~new_n1005;
  assign new_n1008 = new_n1006 & new_n1007;
  assign new_n1009 = new_n296 & new_n1008;
  assign new_n1010 = ~new_n985 & ~new_n993;
  assign new_n1011 = ~new_n1001 & ~new_n1009;
  assign new_n1012 = new_n1010 & new_n1011;
  assign new_n1013 = new_n383 & ~new_n1012;
  assign new_n1014 = ~new_n905 & ~new_n941;
  assign new_n1015 = ~new_n977 & ~new_n1013;
  assign new_n1016 = new_n1014 & new_n1015;
  assign new_n1017 = ~shift6 & ~new_n1016;
  assign new_n1018 = a24 & new_n266;
  assign new_n1019 = a23 & new_n268;
  assign new_n1020 = a26 & new_n270;
  assign new_n1021 = a25 & new_n272;
  assign new_n1022 = ~new_n1018 & ~new_n1019;
  assign new_n1023 = ~new_n1020 & ~new_n1021;
  assign new_n1024 = new_n1022 & new_n1023;
  assign new_n1025 = new_n265 & new_n1024;
  assign new_n1026 = a32 & new_n266;
  assign new_n1027 = a31 & new_n268;
  assign new_n1028 = a34 & new_n270;
  assign new_n1029 = a33 & new_n272;
  assign new_n1030 = ~new_n1026 & ~new_n1027;
  assign new_n1031 = ~new_n1028 & ~new_n1029;
  assign new_n1032 = new_n1030 & new_n1031;
  assign new_n1033 = new_n278 & new_n1032;
  assign new_n1034 = a20 & new_n266;
  assign new_n1035 = a19 & new_n268;
  assign new_n1036 = a22 & new_n270;
  assign new_n1037 = a21 & new_n272;
  assign new_n1038 = ~new_n1034 & ~new_n1035;
  assign new_n1039 = ~new_n1036 & ~new_n1037;
  assign new_n1040 = new_n1038 & new_n1039;
  assign new_n1041 = new_n287 & new_n1040;
  assign new_n1042 = a28 & new_n266;
  assign new_n1043 = a27 & new_n268;
  assign new_n1044 = a30 & new_n270;
  assign new_n1045 = a29 & new_n272;
  assign new_n1046 = ~new_n1042 & ~new_n1043;
  assign new_n1047 = ~new_n1044 & ~new_n1045;
  assign new_n1048 = new_n1046 & new_n1047;
  assign new_n1049 = new_n296 & new_n1048;
  assign new_n1050 = ~new_n1025 & ~new_n1033;
  assign new_n1051 = ~new_n1041 & ~new_n1049;
  assign new_n1052 = new_n1050 & new_n1051;
  assign new_n1053 = new_n264 & ~new_n1052;
  assign new_n1054 = a56 & new_n266;
  assign new_n1055 = a55 & new_n268;
  assign new_n1056 = a58 & new_n270;
  assign new_n1057 = a57 & new_n272;
  assign new_n1058 = ~new_n1054 & ~new_n1055;
  assign new_n1059 = ~new_n1056 & ~new_n1057;
  assign new_n1060 = new_n1058 & new_n1059;
  assign new_n1061 = new_n265 & new_n1060;
  assign new_n1062 = a64 & new_n266;
  assign new_n1063 = a63 & new_n268;
  assign new_n1064 = a66 & new_n270;
  assign new_n1065 = a65 & new_n272;
  assign new_n1066 = ~new_n1062 & ~new_n1063;
  assign new_n1067 = ~new_n1064 & ~new_n1065;
  assign new_n1068 = new_n1066 & new_n1067;
  assign new_n1069 = new_n278 & new_n1068;
  assign new_n1070 = a52 & new_n266;
  assign new_n1071 = a51 & new_n268;
  assign new_n1072 = a54 & new_n270;
  assign new_n1073 = a53 & new_n272;
  assign new_n1074 = ~new_n1070 & ~new_n1071;
  assign new_n1075 = ~new_n1072 & ~new_n1073;
  assign new_n1076 = new_n1074 & new_n1075;
  assign new_n1077 = new_n287 & new_n1076;
  assign new_n1078 = a60 & new_n266;
  assign new_n1079 = a59 & new_n268;
  assign new_n1080 = a62 & new_n270;
  assign new_n1081 = a61 & new_n272;
  assign new_n1082 = ~new_n1078 & ~new_n1079;
  assign new_n1083 = ~new_n1080 & ~new_n1081;
  assign new_n1084 = new_n1082 & new_n1083;
  assign new_n1085 = new_n296 & new_n1084;
  assign new_n1086 = ~new_n1061 & ~new_n1069;
  assign new_n1087 = ~new_n1077 & ~new_n1085;
  assign new_n1088 = new_n1086 & new_n1087;
  assign new_n1089 = new_n309 & ~new_n1088;
  assign new_n1090 = a8 & new_n266;
  assign new_n1091 = a7 & new_n268;
  assign new_n1092 = a10 & new_n270;
  assign new_n1093 = a9 & new_n272;
  assign new_n1094 = ~new_n1090 & ~new_n1091;
  assign new_n1095 = ~new_n1092 & ~new_n1093;
  assign new_n1096 = new_n1094 & new_n1095;
  assign new_n1097 = new_n265 & new_n1096;
  assign new_n1098 = a16 & new_n266;
  assign new_n1099 = a15 & new_n268;
  assign new_n1100 = a18 & new_n270;
  assign new_n1101 = a17 & new_n272;
  assign new_n1102 = ~new_n1098 & ~new_n1099;
  assign new_n1103 = ~new_n1100 & ~new_n1101;
  assign new_n1104 = new_n1102 & new_n1103;
  assign new_n1105 = new_n278 & new_n1104;
  assign new_n1106 = a4 & new_n266;
  assign new_n1107 = a3 & new_n268;
  assign new_n1108 = a6 & new_n270;
  assign new_n1109 = a5 & new_n272;
  assign new_n1110 = ~new_n1106 & ~new_n1107;
  assign new_n1111 = ~new_n1108 & ~new_n1109;
  assign new_n1112 = new_n1110 & new_n1111;
  assign new_n1113 = new_n287 & new_n1112;
  assign new_n1114 = a12 & new_n266;
  assign new_n1115 = a11 & new_n268;
  assign new_n1116 = a14 & new_n270;
  assign new_n1117 = a13 & new_n272;
  assign new_n1118 = ~new_n1114 & ~new_n1115;
  assign new_n1119 = ~new_n1116 & ~new_n1117;
  assign new_n1120 = new_n1118 & new_n1119;
  assign new_n1121 = new_n296 & new_n1120;
  assign new_n1122 = ~new_n1097 & ~new_n1105;
  assign new_n1123 = ~new_n1113 & ~new_n1121;
  assign new_n1124 = new_n1122 & new_n1123;
  assign new_n1125 = new_n346 & ~new_n1124;
  assign new_n1126 = a40 & new_n266;
  assign new_n1127 = a39 & new_n268;
  assign new_n1128 = a42 & new_n270;
  assign new_n1129 = a41 & new_n272;
  assign new_n1130 = ~new_n1126 & ~new_n1127;
  assign new_n1131 = ~new_n1128 & ~new_n1129;
  assign new_n1132 = new_n1130 & new_n1131;
  assign new_n1133 = new_n265 & new_n1132;
  assign new_n1134 = a48 & new_n266;
  assign new_n1135 = a47 & new_n268;
  assign new_n1136 = a50 & new_n270;
  assign new_n1137 = a49 & new_n272;
  assign new_n1138 = ~new_n1134 & ~new_n1135;
  assign new_n1139 = ~new_n1136 & ~new_n1137;
  assign new_n1140 = new_n1138 & new_n1139;
  assign new_n1141 = new_n278 & new_n1140;
  assign new_n1142 = a36 & new_n266;
  assign new_n1143 = a35 & new_n268;
  assign new_n1144 = a38 & new_n270;
  assign new_n1145 = a37 & new_n272;
  assign new_n1146 = ~new_n1142 & ~new_n1143;
  assign new_n1147 = ~new_n1144 & ~new_n1145;
  assign new_n1148 = new_n1146 & new_n1147;
  assign new_n1149 = new_n287 & new_n1148;
  assign new_n1150 = a44 & new_n266;
  assign new_n1151 = a43 & new_n268;
  assign new_n1152 = a46 & new_n270;
  assign new_n1153 = a45 & new_n272;
  assign new_n1154 = ~new_n1150 & ~new_n1151;
  assign new_n1155 = ~new_n1152 & ~new_n1153;
  assign new_n1156 = new_n1154 & new_n1155;
  assign new_n1157 = new_n296 & new_n1156;
  assign new_n1158 = ~new_n1133 & ~new_n1141;
  assign new_n1159 = ~new_n1149 & ~new_n1157;
  assign new_n1160 = new_n1158 & new_n1159;
  assign new_n1161 = new_n383 & ~new_n1160;
  assign new_n1162 = ~new_n1053 & ~new_n1089;
  assign new_n1163 = ~new_n1125 & ~new_n1161;
  assign new_n1164 = new_n1162 & new_n1163;
  assign new_n1165 = shift6 & ~new_n1164;
  assign result2 = ~new_n1017 & ~new_n1165;
  assign new_n1167 = a89 & new_n266;
  assign new_n1168 = a88 & new_n268;
  assign new_n1169 = a91 & new_n270;
  assign new_n1170 = a90 & new_n272;
  assign new_n1171 = ~new_n1167 & ~new_n1168;
  assign new_n1172 = ~new_n1169 & ~new_n1170;
  assign new_n1173 = new_n1171 & new_n1172;
  assign new_n1174 = new_n265 & new_n1173;
  assign new_n1175 = a97 & new_n266;
  assign new_n1176 = a96 & new_n268;
  assign new_n1177 = a99 & new_n270;
  assign new_n1178 = a98 & new_n272;
  assign new_n1179 = ~new_n1175 & ~new_n1176;
  assign new_n1180 = ~new_n1177 & ~new_n1178;
  assign new_n1181 = new_n1179 & new_n1180;
  assign new_n1182 = new_n278 & new_n1181;
  assign new_n1183 = a85 & new_n266;
  assign new_n1184 = a84 & new_n268;
  assign new_n1185 = a87 & new_n270;
  assign new_n1186 = a86 & new_n272;
  assign new_n1187 = ~new_n1183 & ~new_n1184;
  assign new_n1188 = ~new_n1185 & ~new_n1186;
  assign new_n1189 = new_n1187 & new_n1188;
  assign new_n1190 = new_n287 & new_n1189;
  assign new_n1191 = a93 & new_n266;
  assign new_n1192 = a92 & new_n268;
  assign new_n1193 = a95 & new_n270;
  assign new_n1194 = a94 & new_n272;
  assign new_n1195 = ~new_n1191 & ~new_n1192;
  assign new_n1196 = ~new_n1193 & ~new_n1194;
  assign new_n1197 = new_n1195 & new_n1196;
  assign new_n1198 = new_n296 & new_n1197;
  assign new_n1199 = ~new_n1174 & ~new_n1182;
  assign new_n1200 = ~new_n1190 & ~new_n1198;
  assign new_n1201 = new_n1199 & new_n1200;
  assign new_n1202 = new_n264 & ~new_n1201;
  assign new_n1203 = a121 & new_n266;
  assign new_n1204 = a120 & new_n268;
  assign new_n1205 = a123 & new_n270;
  assign new_n1206 = a122 & new_n272;
  assign new_n1207 = ~new_n1203 & ~new_n1204;
  assign new_n1208 = ~new_n1205 & ~new_n1206;
  assign new_n1209 = new_n1207 & new_n1208;
  assign new_n1210 = new_n265 & new_n1209;
  assign new_n1211 = a1 & new_n266;
  assign new_n1212 = a0 & new_n268;
  assign new_n1213 = a3 & new_n270;
  assign new_n1214 = a2 & new_n272;
  assign new_n1215 = ~new_n1211 & ~new_n1212;
  assign new_n1216 = ~new_n1213 & ~new_n1214;
  assign new_n1217 = new_n1215 & new_n1216;
  assign new_n1218 = new_n278 & new_n1217;
  assign new_n1219 = a117 & new_n266;
  assign new_n1220 = a116 & new_n268;
  assign new_n1221 = a119 & new_n270;
  assign new_n1222 = a118 & new_n272;
  assign new_n1223 = ~new_n1219 & ~new_n1220;
  assign new_n1224 = ~new_n1221 & ~new_n1222;
  assign new_n1225 = new_n1223 & new_n1224;
  assign new_n1226 = new_n287 & new_n1225;
  assign new_n1227 = a125 & new_n266;
  assign new_n1228 = a124 & new_n268;
  assign new_n1229 = a127 & new_n270;
  assign new_n1230 = a126 & new_n272;
  assign new_n1231 = ~new_n1227 & ~new_n1228;
  assign new_n1232 = ~new_n1229 & ~new_n1230;
  assign new_n1233 = new_n1231 & new_n1232;
  assign new_n1234 = new_n296 & new_n1233;
  assign new_n1235 = ~new_n1210 & ~new_n1218;
  assign new_n1236 = ~new_n1226 & ~new_n1234;
  assign new_n1237 = new_n1235 & new_n1236;
  assign new_n1238 = new_n309 & ~new_n1237;
  assign new_n1239 = a73 & new_n266;
  assign new_n1240 = a72 & new_n268;
  assign new_n1241 = a75 & new_n270;
  assign new_n1242 = a74 & new_n272;
  assign new_n1243 = ~new_n1239 & ~new_n1240;
  assign new_n1244 = ~new_n1241 & ~new_n1242;
  assign new_n1245 = new_n1243 & new_n1244;
  assign new_n1246 = new_n265 & new_n1245;
  assign new_n1247 = a81 & new_n266;
  assign new_n1248 = a80 & new_n268;
  assign new_n1249 = a83 & new_n270;
  assign new_n1250 = a82 & new_n272;
  assign new_n1251 = ~new_n1247 & ~new_n1248;
  assign new_n1252 = ~new_n1249 & ~new_n1250;
  assign new_n1253 = new_n1251 & new_n1252;
  assign new_n1254 = new_n278 & new_n1253;
  assign new_n1255 = a69 & new_n266;
  assign new_n1256 = a68 & new_n268;
  assign new_n1257 = a71 & new_n270;
  assign new_n1258 = a70 & new_n272;
  assign new_n1259 = ~new_n1255 & ~new_n1256;
  assign new_n1260 = ~new_n1257 & ~new_n1258;
  assign new_n1261 = new_n1259 & new_n1260;
  assign new_n1262 = new_n287 & new_n1261;
  assign new_n1263 = a77 & new_n266;
  assign new_n1264 = a76 & new_n268;
  assign new_n1265 = a79 & new_n270;
  assign new_n1266 = a78 & new_n272;
  assign new_n1267 = ~new_n1263 & ~new_n1264;
  assign new_n1268 = ~new_n1265 & ~new_n1266;
  assign new_n1269 = new_n1267 & new_n1268;
  assign new_n1270 = new_n296 & new_n1269;
  assign new_n1271 = ~new_n1246 & ~new_n1254;
  assign new_n1272 = ~new_n1262 & ~new_n1270;
  assign new_n1273 = new_n1271 & new_n1272;
  assign new_n1274 = new_n346 & ~new_n1273;
  assign new_n1275 = a105 & new_n266;
  assign new_n1276 = a104 & new_n268;
  assign new_n1277 = a107 & new_n270;
  assign new_n1278 = a106 & new_n272;
  assign new_n1279 = ~new_n1275 & ~new_n1276;
  assign new_n1280 = ~new_n1277 & ~new_n1278;
  assign new_n1281 = new_n1279 & new_n1280;
  assign new_n1282 = new_n265 & new_n1281;
  assign new_n1283 = a113 & new_n266;
  assign new_n1284 = a112 & new_n268;
  assign new_n1285 = a115 & new_n270;
  assign new_n1286 = a114 & new_n272;
  assign new_n1287 = ~new_n1283 & ~new_n1284;
  assign new_n1288 = ~new_n1285 & ~new_n1286;
  assign new_n1289 = new_n1287 & new_n1288;
  assign new_n1290 = new_n278 & new_n1289;
  assign new_n1291 = a101 & new_n266;
  assign new_n1292 = a100 & new_n268;
  assign new_n1293 = a103 & new_n270;
  assign new_n1294 = a102 & new_n272;
  assign new_n1295 = ~new_n1291 & ~new_n1292;
  assign new_n1296 = ~new_n1293 & ~new_n1294;
  assign new_n1297 = new_n1295 & new_n1296;
  assign new_n1298 = new_n287 & new_n1297;
  assign new_n1299 = a109 & new_n266;
  assign new_n1300 = a108 & new_n268;
  assign new_n1301 = a111 & new_n270;
  assign new_n1302 = a110 & new_n272;
  assign new_n1303 = ~new_n1299 & ~new_n1300;
  assign new_n1304 = ~new_n1301 & ~new_n1302;
  assign new_n1305 = new_n1303 & new_n1304;
  assign new_n1306 = new_n296 & new_n1305;
  assign new_n1307 = ~new_n1282 & ~new_n1290;
  assign new_n1308 = ~new_n1298 & ~new_n1306;
  assign new_n1309 = new_n1307 & new_n1308;
  assign new_n1310 = new_n383 & ~new_n1309;
  assign new_n1311 = ~new_n1202 & ~new_n1238;
  assign new_n1312 = ~new_n1274 & ~new_n1310;
  assign new_n1313 = new_n1311 & new_n1312;
  assign new_n1314 = ~shift6 & ~new_n1313;
  assign new_n1315 = a25 & new_n266;
  assign new_n1316 = a24 & new_n268;
  assign new_n1317 = a27 & new_n270;
  assign new_n1318 = a26 & new_n272;
  assign new_n1319 = ~new_n1315 & ~new_n1316;
  assign new_n1320 = ~new_n1317 & ~new_n1318;
  assign new_n1321 = new_n1319 & new_n1320;
  assign new_n1322 = new_n265 & new_n1321;
  assign new_n1323 = a33 & new_n266;
  assign new_n1324 = a32 & new_n268;
  assign new_n1325 = a35 & new_n270;
  assign new_n1326 = a34 & new_n272;
  assign new_n1327 = ~new_n1323 & ~new_n1324;
  assign new_n1328 = ~new_n1325 & ~new_n1326;
  assign new_n1329 = new_n1327 & new_n1328;
  assign new_n1330 = new_n278 & new_n1329;
  assign new_n1331 = a21 & new_n266;
  assign new_n1332 = a20 & new_n268;
  assign new_n1333 = a23 & new_n270;
  assign new_n1334 = a22 & new_n272;
  assign new_n1335 = ~new_n1331 & ~new_n1332;
  assign new_n1336 = ~new_n1333 & ~new_n1334;
  assign new_n1337 = new_n1335 & new_n1336;
  assign new_n1338 = new_n287 & new_n1337;
  assign new_n1339 = a29 & new_n266;
  assign new_n1340 = a28 & new_n268;
  assign new_n1341 = a31 & new_n270;
  assign new_n1342 = a30 & new_n272;
  assign new_n1343 = ~new_n1339 & ~new_n1340;
  assign new_n1344 = ~new_n1341 & ~new_n1342;
  assign new_n1345 = new_n1343 & new_n1344;
  assign new_n1346 = new_n296 & new_n1345;
  assign new_n1347 = ~new_n1322 & ~new_n1330;
  assign new_n1348 = ~new_n1338 & ~new_n1346;
  assign new_n1349 = new_n1347 & new_n1348;
  assign new_n1350 = new_n264 & ~new_n1349;
  assign new_n1351 = a57 & new_n266;
  assign new_n1352 = a56 & new_n268;
  assign new_n1353 = a59 & new_n270;
  assign new_n1354 = a58 & new_n272;
  assign new_n1355 = ~new_n1351 & ~new_n1352;
  assign new_n1356 = ~new_n1353 & ~new_n1354;
  assign new_n1357 = new_n1355 & new_n1356;
  assign new_n1358 = new_n265 & new_n1357;
  assign new_n1359 = a65 & new_n266;
  assign new_n1360 = a64 & new_n268;
  assign new_n1361 = a67 & new_n270;
  assign new_n1362 = a66 & new_n272;
  assign new_n1363 = ~new_n1359 & ~new_n1360;
  assign new_n1364 = ~new_n1361 & ~new_n1362;
  assign new_n1365 = new_n1363 & new_n1364;
  assign new_n1366 = new_n278 & new_n1365;
  assign new_n1367 = a53 & new_n266;
  assign new_n1368 = a52 & new_n268;
  assign new_n1369 = a55 & new_n270;
  assign new_n1370 = a54 & new_n272;
  assign new_n1371 = ~new_n1367 & ~new_n1368;
  assign new_n1372 = ~new_n1369 & ~new_n1370;
  assign new_n1373 = new_n1371 & new_n1372;
  assign new_n1374 = new_n287 & new_n1373;
  assign new_n1375 = a61 & new_n266;
  assign new_n1376 = a60 & new_n268;
  assign new_n1377 = a63 & new_n270;
  assign new_n1378 = a62 & new_n272;
  assign new_n1379 = ~new_n1375 & ~new_n1376;
  assign new_n1380 = ~new_n1377 & ~new_n1378;
  assign new_n1381 = new_n1379 & new_n1380;
  assign new_n1382 = new_n296 & new_n1381;
  assign new_n1383 = ~new_n1358 & ~new_n1366;
  assign new_n1384 = ~new_n1374 & ~new_n1382;
  assign new_n1385 = new_n1383 & new_n1384;
  assign new_n1386 = new_n309 & ~new_n1385;
  assign new_n1387 = a9 & new_n266;
  assign new_n1388 = a8 & new_n268;
  assign new_n1389 = a11 & new_n270;
  assign new_n1390 = a10 & new_n272;
  assign new_n1391 = ~new_n1387 & ~new_n1388;
  assign new_n1392 = ~new_n1389 & ~new_n1390;
  assign new_n1393 = new_n1391 & new_n1392;
  assign new_n1394 = new_n265 & new_n1393;
  assign new_n1395 = a17 & new_n266;
  assign new_n1396 = a16 & new_n268;
  assign new_n1397 = a19 & new_n270;
  assign new_n1398 = a18 & new_n272;
  assign new_n1399 = ~new_n1395 & ~new_n1396;
  assign new_n1400 = ~new_n1397 & ~new_n1398;
  assign new_n1401 = new_n1399 & new_n1400;
  assign new_n1402 = new_n278 & new_n1401;
  assign new_n1403 = a5 & new_n266;
  assign new_n1404 = a4 & new_n268;
  assign new_n1405 = a7 & new_n270;
  assign new_n1406 = a6 & new_n272;
  assign new_n1407 = ~new_n1403 & ~new_n1404;
  assign new_n1408 = ~new_n1405 & ~new_n1406;
  assign new_n1409 = new_n1407 & new_n1408;
  assign new_n1410 = new_n287 & new_n1409;
  assign new_n1411 = a13 & new_n266;
  assign new_n1412 = a12 & new_n268;
  assign new_n1413 = a15 & new_n270;
  assign new_n1414 = a14 & new_n272;
  assign new_n1415 = ~new_n1411 & ~new_n1412;
  assign new_n1416 = ~new_n1413 & ~new_n1414;
  assign new_n1417 = new_n1415 & new_n1416;
  assign new_n1418 = new_n296 & new_n1417;
  assign new_n1419 = ~new_n1394 & ~new_n1402;
  assign new_n1420 = ~new_n1410 & ~new_n1418;
  assign new_n1421 = new_n1419 & new_n1420;
  assign new_n1422 = new_n346 & ~new_n1421;
  assign new_n1423 = a41 & new_n266;
  assign new_n1424 = a40 & new_n268;
  assign new_n1425 = a43 & new_n270;
  assign new_n1426 = a42 & new_n272;
  assign new_n1427 = ~new_n1423 & ~new_n1424;
  assign new_n1428 = ~new_n1425 & ~new_n1426;
  assign new_n1429 = new_n1427 & new_n1428;
  assign new_n1430 = new_n265 & new_n1429;
  assign new_n1431 = a49 & new_n266;
  assign new_n1432 = a48 & new_n268;
  assign new_n1433 = a51 & new_n270;
  assign new_n1434 = a50 & new_n272;
  assign new_n1435 = ~new_n1431 & ~new_n1432;
  assign new_n1436 = ~new_n1433 & ~new_n1434;
  assign new_n1437 = new_n1435 & new_n1436;
  assign new_n1438 = new_n278 & new_n1437;
  assign new_n1439 = a37 & new_n266;
  assign new_n1440 = a36 & new_n268;
  assign new_n1441 = a39 & new_n270;
  assign new_n1442 = a38 & new_n272;
  assign new_n1443 = ~new_n1439 & ~new_n1440;
  assign new_n1444 = ~new_n1441 & ~new_n1442;
  assign new_n1445 = new_n1443 & new_n1444;
  assign new_n1446 = new_n287 & new_n1445;
  assign new_n1447 = a45 & new_n266;
  assign new_n1448 = a44 & new_n268;
  assign new_n1449 = a47 & new_n270;
  assign new_n1450 = a46 & new_n272;
  assign new_n1451 = ~new_n1447 & ~new_n1448;
  assign new_n1452 = ~new_n1449 & ~new_n1450;
  assign new_n1453 = new_n1451 & new_n1452;
  assign new_n1454 = new_n296 & new_n1453;
  assign new_n1455 = ~new_n1430 & ~new_n1438;
  assign new_n1456 = ~new_n1446 & ~new_n1454;
  assign new_n1457 = new_n1455 & new_n1456;
  assign new_n1458 = new_n383 & ~new_n1457;
  assign new_n1459 = ~new_n1350 & ~new_n1386;
  assign new_n1460 = ~new_n1422 & ~new_n1458;
  assign new_n1461 = new_n1459 & new_n1460;
  assign new_n1462 = shift6 & ~new_n1461;
  assign result3 = ~new_n1314 & ~new_n1462;
  assign new_n1464 = new_n265 & new_n303;
  assign new_n1465 = new_n278 & new_n406;
  assign new_n1466 = new_n276 & new_n287;
  assign new_n1467 = new_n285 & new_n296;
  assign new_n1468 = ~new_n1464 & ~new_n1465;
  assign new_n1469 = ~new_n1466 & ~new_n1467;
  assign new_n1470 = new_n1468 & new_n1469;
  assign new_n1471 = new_n264 & ~new_n1470;
  assign new_n1472 = new_n265 & new_n340;
  assign new_n1473 = new_n278 & new_n518;
  assign new_n1474 = new_n287 & new_n316;
  assign new_n1475 = new_n296 & new_n324;
  assign new_n1476 = ~new_n1472 & ~new_n1473;
  assign new_n1477 = ~new_n1474 & ~new_n1475;
  assign new_n1478 = new_n1476 & new_n1477;
  assign new_n1479 = new_n309 & ~new_n1478;
  assign new_n1480 = new_n265 & new_n377;
  assign new_n1481 = new_n278 & new_n294;
  assign new_n1482 = new_n287 & new_n353;
  assign new_n1483 = new_n296 & new_n361;
  assign new_n1484 = ~new_n1480 & ~new_n1481;
  assign new_n1485 = ~new_n1482 & ~new_n1483;
  assign new_n1486 = new_n1484 & new_n1485;
  assign new_n1487 = new_n346 & ~new_n1486;
  assign new_n1488 = new_n265 & new_n414;
  assign new_n1489 = new_n278 & new_n332;
  assign new_n1490 = new_n287 & new_n390;
  assign new_n1491 = new_n296 & new_n398;
  assign new_n1492 = ~new_n1488 & ~new_n1489;
  assign new_n1493 = ~new_n1490 & ~new_n1491;
  assign new_n1494 = new_n1492 & new_n1493;
  assign new_n1495 = new_n383 & ~new_n1494;
  assign new_n1496 = ~new_n1471 & ~new_n1479;
  assign new_n1497 = ~new_n1487 & ~new_n1495;
  assign new_n1498 = new_n1496 & new_n1497;
  assign new_n1499 = ~shift6 & ~new_n1498;
  assign new_n1500 = new_n265 & new_n454;
  assign new_n1501 = new_n278 & new_n554;
  assign new_n1502 = new_n287 & new_n430;
  assign new_n1503 = new_n296 & new_n438;
  assign new_n1504 = ~new_n1500 & ~new_n1501;
  assign new_n1505 = ~new_n1502 & ~new_n1503;
  assign new_n1506 = new_n1504 & new_n1505;
  assign new_n1507 = new_n264 & ~new_n1506;
  assign new_n1508 = new_n265 & new_n490;
  assign new_n1509 = new_n278 & new_n369;
  assign new_n1510 = new_n287 & new_n466;
  assign new_n1511 = new_n296 & new_n474;
  assign new_n1512 = ~new_n1508 & ~new_n1509;
  assign new_n1513 = ~new_n1510 & ~new_n1511;
  assign new_n1514 = new_n1512 & new_n1513;
  assign new_n1515 = new_n309 & ~new_n1514;
  assign new_n1516 = new_n265 & new_n526;
  assign new_n1517 = new_n278 & new_n446;
  assign new_n1518 = new_n287 & new_n502;
  assign new_n1519 = new_n296 & new_n510;
  assign new_n1520 = ~new_n1516 & ~new_n1517;
  assign new_n1521 = ~new_n1518 & ~new_n1519;
  assign new_n1522 = new_n1520 & new_n1521;
  assign new_n1523 = new_n346 & ~new_n1522;
  assign new_n1524 = new_n265 & new_n562;
  assign new_n1525 = new_n278 & new_n482;
  assign new_n1526 = new_n287 & new_n538;
  assign new_n1527 = new_n296 & new_n546;
  assign new_n1528 = ~new_n1524 & ~new_n1525;
  assign new_n1529 = ~new_n1526 & ~new_n1527;
  assign new_n1530 = new_n1528 & new_n1529;
  assign new_n1531 = new_n383 & ~new_n1530;
  assign new_n1532 = ~new_n1507 & ~new_n1515;
  assign new_n1533 = ~new_n1523 & ~new_n1531;
  assign new_n1534 = new_n1532 & new_n1533;
  assign new_n1535 = shift6 & ~new_n1534;
  assign result4 = ~new_n1499 & ~new_n1535;
  assign new_n1537 = new_n265 & new_n603;
  assign new_n1538 = new_n278 & new_n703;
  assign new_n1539 = new_n287 & new_n579;
  assign new_n1540 = new_n296 & new_n587;
  assign new_n1541 = ~new_n1537 & ~new_n1538;
  assign new_n1542 = ~new_n1539 & ~new_n1540;
  assign new_n1543 = new_n1541 & new_n1542;
  assign new_n1544 = new_n264 & ~new_n1543;
  assign new_n1545 = new_n265 & new_n639;
  assign new_n1546 = new_n278 & new_n815;
  assign new_n1547 = new_n287 & new_n615;
  assign new_n1548 = new_n296 & new_n623;
  assign new_n1549 = ~new_n1545 & ~new_n1546;
  assign new_n1550 = ~new_n1547 & ~new_n1548;
  assign new_n1551 = new_n1549 & new_n1550;
  assign new_n1552 = new_n309 & ~new_n1551;
  assign new_n1553 = new_n265 & new_n675;
  assign new_n1554 = new_n278 & new_n595;
  assign new_n1555 = new_n287 & new_n651;
  assign new_n1556 = new_n296 & new_n659;
  assign new_n1557 = ~new_n1553 & ~new_n1554;
  assign new_n1558 = ~new_n1555 & ~new_n1556;
  assign new_n1559 = new_n1557 & new_n1558;
  assign new_n1560 = new_n346 & ~new_n1559;
  assign new_n1561 = new_n265 & new_n711;
  assign new_n1562 = new_n278 & new_n631;
  assign new_n1563 = new_n287 & new_n687;
  assign new_n1564 = new_n296 & new_n695;
  assign new_n1565 = ~new_n1561 & ~new_n1562;
  assign new_n1566 = ~new_n1563 & ~new_n1564;
  assign new_n1567 = new_n1565 & new_n1566;
  assign new_n1568 = new_n383 & ~new_n1567;
  assign new_n1569 = ~new_n1544 & ~new_n1552;
  assign new_n1570 = ~new_n1560 & ~new_n1568;
  assign new_n1571 = new_n1569 & new_n1570;
  assign new_n1572 = ~shift6 & ~new_n1571;
  assign new_n1573 = new_n265 & new_n751;
  assign new_n1574 = new_n278 & new_n851;
  assign new_n1575 = new_n287 & new_n727;
  assign new_n1576 = new_n296 & new_n735;
  assign new_n1577 = ~new_n1573 & ~new_n1574;
  assign new_n1578 = ~new_n1575 & ~new_n1576;
  assign new_n1579 = new_n1577 & new_n1578;
  assign new_n1580 = new_n264 & ~new_n1579;
  assign new_n1581 = new_n265 & new_n787;
  assign new_n1582 = new_n278 & new_n667;
  assign new_n1583 = new_n287 & new_n763;
  assign new_n1584 = new_n296 & new_n771;
  assign new_n1585 = ~new_n1581 & ~new_n1582;
  assign new_n1586 = ~new_n1583 & ~new_n1584;
  assign new_n1587 = new_n1585 & new_n1586;
  assign new_n1588 = new_n309 & ~new_n1587;
  assign new_n1589 = new_n265 & new_n823;
  assign new_n1590 = new_n278 & new_n743;
  assign new_n1591 = new_n287 & new_n799;
  assign new_n1592 = new_n296 & new_n807;
  assign new_n1593 = ~new_n1589 & ~new_n1590;
  assign new_n1594 = ~new_n1591 & ~new_n1592;
  assign new_n1595 = new_n1593 & new_n1594;
  assign new_n1596 = new_n346 & ~new_n1595;
  assign new_n1597 = new_n265 & new_n859;
  assign new_n1598 = new_n278 & new_n779;
  assign new_n1599 = new_n287 & new_n835;
  assign new_n1600 = new_n296 & new_n843;
  assign new_n1601 = ~new_n1597 & ~new_n1598;
  assign new_n1602 = ~new_n1599 & ~new_n1600;
  assign new_n1603 = new_n1601 & new_n1602;
  assign new_n1604 = new_n383 & ~new_n1603;
  assign new_n1605 = ~new_n1580 & ~new_n1588;
  assign new_n1606 = ~new_n1596 & ~new_n1604;
  assign new_n1607 = new_n1605 & new_n1606;
  assign new_n1608 = shift6 & ~new_n1607;
  assign result5 = ~new_n1572 & ~new_n1608;
  assign new_n1610 = new_n265 & new_n900;
  assign new_n1611 = new_n278 & new_n1000;
  assign new_n1612 = new_n287 & new_n876;
  assign new_n1613 = new_n296 & new_n884;
  assign new_n1614 = ~new_n1610 & ~new_n1611;
  assign new_n1615 = ~new_n1612 & ~new_n1613;
  assign new_n1616 = new_n1614 & new_n1615;
  assign new_n1617 = new_n264 & ~new_n1616;
  assign new_n1618 = new_n265 & new_n936;
  assign new_n1619 = new_n278 & new_n1112;
  assign new_n1620 = new_n287 & new_n912;
  assign new_n1621 = new_n296 & new_n920;
  assign new_n1622 = ~new_n1618 & ~new_n1619;
  assign new_n1623 = ~new_n1620 & ~new_n1621;
  assign new_n1624 = new_n1622 & new_n1623;
  assign new_n1625 = new_n309 & ~new_n1624;
  assign new_n1626 = new_n265 & new_n972;
  assign new_n1627 = new_n278 & new_n892;
  assign new_n1628 = new_n287 & new_n948;
  assign new_n1629 = new_n296 & new_n956;
  assign new_n1630 = ~new_n1626 & ~new_n1627;
  assign new_n1631 = ~new_n1628 & ~new_n1629;
  assign new_n1632 = new_n1630 & new_n1631;
  assign new_n1633 = new_n346 & ~new_n1632;
  assign new_n1634 = new_n265 & new_n1008;
  assign new_n1635 = new_n278 & new_n928;
  assign new_n1636 = new_n287 & new_n984;
  assign new_n1637 = new_n296 & new_n992;
  assign new_n1638 = ~new_n1634 & ~new_n1635;
  assign new_n1639 = ~new_n1636 & ~new_n1637;
  assign new_n1640 = new_n1638 & new_n1639;
  assign new_n1641 = new_n383 & ~new_n1640;
  assign new_n1642 = ~new_n1617 & ~new_n1625;
  assign new_n1643 = ~new_n1633 & ~new_n1641;
  assign new_n1644 = new_n1642 & new_n1643;
  assign new_n1645 = ~shift6 & ~new_n1644;
  assign new_n1646 = new_n265 & new_n1048;
  assign new_n1647 = new_n278 & new_n1148;
  assign new_n1648 = new_n287 & new_n1024;
  assign new_n1649 = new_n296 & new_n1032;
  assign new_n1650 = ~new_n1646 & ~new_n1647;
  assign new_n1651 = ~new_n1648 & ~new_n1649;
  assign new_n1652 = new_n1650 & new_n1651;
  assign new_n1653 = new_n264 & ~new_n1652;
  assign new_n1654 = new_n265 & new_n1084;
  assign new_n1655 = new_n278 & new_n964;
  assign new_n1656 = new_n287 & new_n1060;
  assign new_n1657 = new_n296 & new_n1068;
  assign new_n1658 = ~new_n1654 & ~new_n1655;
  assign new_n1659 = ~new_n1656 & ~new_n1657;
  assign new_n1660 = new_n1658 & new_n1659;
  assign new_n1661 = new_n309 & ~new_n1660;
  assign new_n1662 = new_n265 & new_n1120;
  assign new_n1663 = new_n278 & new_n1040;
  assign new_n1664 = new_n287 & new_n1096;
  assign new_n1665 = new_n296 & new_n1104;
  assign new_n1666 = ~new_n1662 & ~new_n1663;
  assign new_n1667 = ~new_n1664 & ~new_n1665;
  assign new_n1668 = new_n1666 & new_n1667;
  assign new_n1669 = new_n346 & ~new_n1668;
  assign new_n1670 = new_n265 & new_n1156;
  assign new_n1671 = new_n278 & new_n1076;
  assign new_n1672 = new_n287 & new_n1132;
  assign new_n1673 = new_n296 & new_n1140;
  assign new_n1674 = ~new_n1670 & ~new_n1671;
  assign new_n1675 = ~new_n1672 & ~new_n1673;
  assign new_n1676 = new_n1674 & new_n1675;
  assign new_n1677 = new_n383 & ~new_n1676;
  assign new_n1678 = ~new_n1653 & ~new_n1661;
  assign new_n1679 = ~new_n1669 & ~new_n1677;
  assign new_n1680 = new_n1678 & new_n1679;
  assign new_n1681 = shift6 & ~new_n1680;
  assign result6 = ~new_n1645 & ~new_n1681;
  assign new_n1683 = new_n265 & new_n1197;
  assign new_n1684 = new_n278 & new_n1297;
  assign new_n1685 = new_n287 & new_n1173;
  assign new_n1686 = new_n296 & new_n1181;
  assign new_n1687 = ~new_n1683 & ~new_n1684;
  assign new_n1688 = ~new_n1685 & ~new_n1686;
  assign new_n1689 = new_n1687 & new_n1688;
  assign new_n1690 = new_n264 & ~new_n1689;
  assign new_n1691 = new_n265 & new_n1233;
  assign new_n1692 = new_n278 & new_n1409;
  assign new_n1693 = new_n287 & new_n1209;
  assign new_n1694 = new_n296 & new_n1217;
  assign new_n1695 = ~new_n1691 & ~new_n1692;
  assign new_n1696 = ~new_n1693 & ~new_n1694;
  assign new_n1697 = new_n1695 & new_n1696;
  assign new_n1698 = new_n309 & ~new_n1697;
  assign new_n1699 = new_n265 & new_n1269;
  assign new_n1700 = new_n278 & new_n1189;
  assign new_n1701 = new_n287 & new_n1245;
  assign new_n1702 = new_n296 & new_n1253;
  assign new_n1703 = ~new_n1699 & ~new_n1700;
  assign new_n1704 = ~new_n1701 & ~new_n1702;
  assign new_n1705 = new_n1703 & new_n1704;
  assign new_n1706 = new_n346 & ~new_n1705;
  assign new_n1707 = new_n265 & new_n1305;
  assign new_n1708 = new_n278 & new_n1225;
  assign new_n1709 = new_n287 & new_n1281;
  assign new_n1710 = new_n296 & new_n1289;
  assign new_n1711 = ~new_n1707 & ~new_n1708;
  assign new_n1712 = ~new_n1709 & ~new_n1710;
  assign new_n1713 = new_n1711 & new_n1712;
  assign new_n1714 = new_n383 & ~new_n1713;
  assign new_n1715 = ~new_n1690 & ~new_n1698;
  assign new_n1716 = ~new_n1706 & ~new_n1714;
  assign new_n1717 = new_n1715 & new_n1716;
  assign new_n1718 = ~shift6 & ~new_n1717;
  assign new_n1719 = new_n265 & new_n1345;
  assign new_n1720 = new_n278 & new_n1445;
  assign new_n1721 = new_n287 & new_n1321;
  assign new_n1722 = new_n296 & new_n1329;
  assign new_n1723 = ~new_n1719 & ~new_n1720;
  assign new_n1724 = ~new_n1721 & ~new_n1722;
  assign new_n1725 = new_n1723 & new_n1724;
  assign new_n1726 = new_n264 & ~new_n1725;
  assign new_n1727 = new_n265 & new_n1381;
  assign new_n1728 = new_n278 & new_n1261;
  assign new_n1729 = new_n287 & new_n1357;
  assign new_n1730 = new_n296 & new_n1365;
  assign new_n1731 = ~new_n1727 & ~new_n1728;
  assign new_n1732 = ~new_n1729 & ~new_n1730;
  assign new_n1733 = new_n1731 & new_n1732;
  assign new_n1734 = new_n309 & ~new_n1733;
  assign new_n1735 = new_n265 & new_n1417;
  assign new_n1736 = new_n278 & new_n1337;
  assign new_n1737 = new_n287 & new_n1393;
  assign new_n1738 = new_n296 & new_n1401;
  assign new_n1739 = ~new_n1735 & ~new_n1736;
  assign new_n1740 = ~new_n1737 & ~new_n1738;
  assign new_n1741 = new_n1739 & new_n1740;
  assign new_n1742 = new_n346 & ~new_n1741;
  assign new_n1743 = new_n265 & new_n1453;
  assign new_n1744 = new_n278 & new_n1373;
  assign new_n1745 = new_n287 & new_n1429;
  assign new_n1746 = new_n296 & new_n1437;
  assign new_n1747 = ~new_n1743 & ~new_n1744;
  assign new_n1748 = ~new_n1745 & ~new_n1746;
  assign new_n1749 = new_n1747 & new_n1748;
  assign new_n1750 = new_n383 & ~new_n1749;
  assign new_n1751 = ~new_n1726 & ~new_n1734;
  assign new_n1752 = ~new_n1742 & ~new_n1750;
  assign new_n1753 = new_n1751 & new_n1752;
  assign new_n1754 = shift6 & ~new_n1753;
  assign result7 = ~new_n1718 & ~new_n1754;
  assign new_n1756 = new_n265 & new_n285;
  assign new_n1757 = new_n278 & new_n390;
  assign new_n1758 = new_n287 & new_n303;
  assign new_n1759 = new_n296 & new_n406;
  assign new_n1760 = ~new_n1756 & ~new_n1757;
  assign new_n1761 = ~new_n1758 & ~new_n1759;
  assign new_n1762 = new_n1760 & new_n1761;
  assign new_n1763 = new_n264 & ~new_n1762;
  assign new_n1764 = new_n265 & new_n324;
  assign new_n1765 = new_n278 & new_n502;
  assign new_n1766 = new_n287 & new_n340;
  assign new_n1767 = new_n296 & new_n518;
  assign new_n1768 = ~new_n1764 & ~new_n1765;
  assign new_n1769 = ~new_n1766 & ~new_n1767;
  assign new_n1770 = new_n1768 & new_n1769;
  assign new_n1771 = new_n309 & ~new_n1770;
  assign new_n1772 = new_n265 & new_n361;
  assign new_n1773 = new_n276 & new_n278;
  assign new_n1774 = new_n287 & new_n377;
  assign new_n1775 = new_n294 & new_n296;
  assign new_n1776 = ~new_n1772 & ~new_n1773;
  assign new_n1777 = ~new_n1774 & ~new_n1775;
  assign new_n1778 = new_n1776 & new_n1777;
  assign new_n1779 = new_n346 & ~new_n1778;
  assign new_n1780 = new_n265 & new_n398;
  assign new_n1781 = new_n278 & new_n316;
  assign new_n1782 = new_n287 & new_n414;
  assign new_n1783 = new_n296 & new_n332;
  assign new_n1784 = ~new_n1780 & ~new_n1781;
  assign new_n1785 = ~new_n1782 & ~new_n1783;
  assign new_n1786 = new_n1784 & new_n1785;
  assign new_n1787 = new_n383 & ~new_n1786;
  assign new_n1788 = ~new_n1763 & ~new_n1771;
  assign new_n1789 = ~new_n1779 & ~new_n1787;
  assign new_n1790 = new_n1788 & new_n1789;
  assign new_n1791 = ~shift6 & ~new_n1790;
  assign new_n1792 = new_n265 & new_n438;
  assign new_n1793 = new_n278 & new_n538;
  assign new_n1794 = new_n287 & new_n454;
  assign new_n1795 = new_n296 & new_n554;
  assign new_n1796 = ~new_n1792 & ~new_n1793;
  assign new_n1797 = ~new_n1794 & ~new_n1795;
  assign new_n1798 = new_n1796 & new_n1797;
  assign new_n1799 = new_n264 & ~new_n1798;
  assign new_n1800 = new_n265 & new_n474;
  assign new_n1801 = new_n278 & new_n353;
  assign new_n1802 = new_n287 & new_n490;
  assign new_n1803 = new_n296 & new_n369;
  assign new_n1804 = ~new_n1800 & ~new_n1801;
  assign new_n1805 = ~new_n1802 & ~new_n1803;
  assign new_n1806 = new_n1804 & new_n1805;
  assign new_n1807 = new_n309 & ~new_n1806;
  assign new_n1808 = new_n265 & new_n510;
  assign new_n1809 = new_n278 & new_n430;
  assign new_n1810 = new_n287 & new_n526;
  assign new_n1811 = new_n296 & new_n446;
  assign new_n1812 = ~new_n1808 & ~new_n1809;
  assign new_n1813 = ~new_n1810 & ~new_n1811;
  assign new_n1814 = new_n1812 & new_n1813;
  assign new_n1815 = new_n346 & ~new_n1814;
  assign new_n1816 = new_n265 & new_n546;
  assign new_n1817 = new_n278 & new_n466;
  assign new_n1818 = new_n287 & new_n562;
  assign new_n1819 = new_n296 & new_n482;
  assign new_n1820 = ~new_n1816 & ~new_n1817;
  assign new_n1821 = ~new_n1818 & ~new_n1819;
  assign new_n1822 = new_n1820 & new_n1821;
  assign new_n1823 = new_n383 & ~new_n1822;
  assign new_n1824 = ~new_n1799 & ~new_n1807;
  assign new_n1825 = ~new_n1815 & ~new_n1823;
  assign new_n1826 = new_n1824 & new_n1825;
  assign new_n1827 = shift6 & ~new_n1826;
  assign result8 = ~new_n1791 & ~new_n1827;
  assign new_n1829 = new_n265 & new_n587;
  assign new_n1830 = new_n278 & new_n687;
  assign new_n1831 = new_n287 & new_n603;
  assign new_n1832 = new_n296 & new_n703;
  assign new_n1833 = ~new_n1829 & ~new_n1830;
  assign new_n1834 = ~new_n1831 & ~new_n1832;
  assign new_n1835 = new_n1833 & new_n1834;
  assign new_n1836 = new_n264 & ~new_n1835;
  assign new_n1837 = new_n265 & new_n623;
  assign new_n1838 = new_n278 & new_n799;
  assign new_n1839 = new_n287 & new_n639;
  assign new_n1840 = new_n296 & new_n815;
  assign new_n1841 = ~new_n1837 & ~new_n1838;
  assign new_n1842 = ~new_n1839 & ~new_n1840;
  assign new_n1843 = new_n1841 & new_n1842;
  assign new_n1844 = new_n309 & ~new_n1843;
  assign new_n1845 = new_n265 & new_n659;
  assign new_n1846 = new_n278 & new_n579;
  assign new_n1847 = new_n287 & new_n675;
  assign new_n1848 = new_n296 & new_n595;
  assign new_n1849 = ~new_n1845 & ~new_n1846;
  assign new_n1850 = ~new_n1847 & ~new_n1848;
  assign new_n1851 = new_n1849 & new_n1850;
  assign new_n1852 = new_n346 & ~new_n1851;
  assign new_n1853 = new_n265 & new_n695;
  assign new_n1854 = new_n278 & new_n615;
  assign new_n1855 = new_n287 & new_n711;
  assign new_n1856 = new_n296 & new_n631;
  assign new_n1857 = ~new_n1853 & ~new_n1854;
  assign new_n1858 = ~new_n1855 & ~new_n1856;
  assign new_n1859 = new_n1857 & new_n1858;
  assign new_n1860 = new_n383 & ~new_n1859;
  assign new_n1861 = ~new_n1836 & ~new_n1844;
  assign new_n1862 = ~new_n1852 & ~new_n1860;
  assign new_n1863 = new_n1861 & new_n1862;
  assign new_n1864 = ~shift6 & ~new_n1863;
  assign new_n1865 = new_n265 & new_n735;
  assign new_n1866 = new_n278 & new_n835;
  assign new_n1867 = new_n287 & new_n751;
  assign new_n1868 = new_n296 & new_n851;
  assign new_n1869 = ~new_n1865 & ~new_n1866;
  assign new_n1870 = ~new_n1867 & ~new_n1868;
  assign new_n1871 = new_n1869 & new_n1870;
  assign new_n1872 = new_n264 & ~new_n1871;
  assign new_n1873 = new_n265 & new_n771;
  assign new_n1874 = new_n278 & new_n651;
  assign new_n1875 = new_n287 & new_n787;
  assign new_n1876 = new_n296 & new_n667;
  assign new_n1877 = ~new_n1873 & ~new_n1874;
  assign new_n1878 = ~new_n1875 & ~new_n1876;
  assign new_n1879 = new_n1877 & new_n1878;
  assign new_n1880 = new_n309 & ~new_n1879;
  assign new_n1881 = new_n265 & new_n807;
  assign new_n1882 = new_n278 & new_n727;
  assign new_n1883 = new_n287 & new_n823;
  assign new_n1884 = new_n296 & new_n743;
  assign new_n1885 = ~new_n1881 & ~new_n1882;
  assign new_n1886 = ~new_n1883 & ~new_n1884;
  assign new_n1887 = new_n1885 & new_n1886;
  assign new_n1888 = new_n346 & ~new_n1887;
  assign new_n1889 = new_n265 & new_n843;
  assign new_n1890 = new_n278 & new_n763;
  assign new_n1891 = new_n287 & new_n859;
  assign new_n1892 = new_n296 & new_n779;
  assign new_n1893 = ~new_n1889 & ~new_n1890;
  assign new_n1894 = ~new_n1891 & ~new_n1892;
  assign new_n1895 = new_n1893 & new_n1894;
  assign new_n1896 = new_n383 & ~new_n1895;
  assign new_n1897 = ~new_n1872 & ~new_n1880;
  assign new_n1898 = ~new_n1888 & ~new_n1896;
  assign new_n1899 = new_n1897 & new_n1898;
  assign new_n1900 = shift6 & ~new_n1899;
  assign result9 = ~new_n1864 & ~new_n1900;
  assign new_n1902 = new_n265 & new_n884;
  assign new_n1903 = new_n278 & new_n984;
  assign new_n1904 = new_n287 & new_n900;
  assign new_n1905 = new_n296 & new_n1000;
  assign new_n1906 = ~new_n1902 & ~new_n1903;
  assign new_n1907 = ~new_n1904 & ~new_n1905;
  assign new_n1908 = new_n1906 & new_n1907;
  assign new_n1909 = new_n264 & ~new_n1908;
  assign new_n1910 = new_n265 & new_n920;
  assign new_n1911 = new_n278 & new_n1096;
  assign new_n1912 = new_n287 & new_n936;
  assign new_n1913 = new_n296 & new_n1112;
  assign new_n1914 = ~new_n1910 & ~new_n1911;
  assign new_n1915 = ~new_n1912 & ~new_n1913;
  assign new_n1916 = new_n1914 & new_n1915;
  assign new_n1917 = new_n309 & ~new_n1916;
  assign new_n1918 = new_n265 & new_n956;
  assign new_n1919 = new_n278 & new_n876;
  assign new_n1920 = new_n287 & new_n972;
  assign new_n1921 = new_n296 & new_n892;
  assign new_n1922 = ~new_n1918 & ~new_n1919;
  assign new_n1923 = ~new_n1920 & ~new_n1921;
  assign new_n1924 = new_n1922 & new_n1923;
  assign new_n1925 = new_n346 & ~new_n1924;
  assign new_n1926 = new_n265 & new_n992;
  assign new_n1927 = new_n278 & new_n912;
  assign new_n1928 = new_n287 & new_n1008;
  assign new_n1929 = new_n296 & new_n928;
  assign new_n1930 = ~new_n1926 & ~new_n1927;
  assign new_n1931 = ~new_n1928 & ~new_n1929;
  assign new_n1932 = new_n1930 & new_n1931;
  assign new_n1933 = new_n383 & ~new_n1932;
  assign new_n1934 = ~new_n1909 & ~new_n1917;
  assign new_n1935 = ~new_n1925 & ~new_n1933;
  assign new_n1936 = new_n1934 & new_n1935;
  assign new_n1937 = ~shift6 & ~new_n1936;
  assign new_n1938 = new_n265 & new_n1032;
  assign new_n1939 = new_n278 & new_n1132;
  assign new_n1940 = new_n287 & new_n1048;
  assign new_n1941 = new_n296 & new_n1148;
  assign new_n1942 = ~new_n1938 & ~new_n1939;
  assign new_n1943 = ~new_n1940 & ~new_n1941;
  assign new_n1944 = new_n1942 & new_n1943;
  assign new_n1945 = new_n264 & ~new_n1944;
  assign new_n1946 = new_n265 & new_n1068;
  assign new_n1947 = new_n278 & new_n948;
  assign new_n1948 = new_n287 & new_n1084;
  assign new_n1949 = new_n296 & new_n964;
  assign new_n1950 = ~new_n1946 & ~new_n1947;
  assign new_n1951 = ~new_n1948 & ~new_n1949;
  assign new_n1952 = new_n1950 & new_n1951;
  assign new_n1953 = new_n309 & ~new_n1952;
  assign new_n1954 = new_n265 & new_n1104;
  assign new_n1955 = new_n278 & new_n1024;
  assign new_n1956 = new_n287 & new_n1120;
  assign new_n1957 = new_n296 & new_n1040;
  assign new_n1958 = ~new_n1954 & ~new_n1955;
  assign new_n1959 = ~new_n1956 & ~new_n1957;
  assign new_n1960 = new_n1958 & new_n1959;
  assign new_n1961 = new_n346 & ~new_n1960;
  assign new_n1962 = new_n265 & new_n1140;
  assign new_n1963 = new_n278 & new_n1060;
  assign new_n1964 = new_n287 & new_n1156;
  assign new_n1965 = new_n296 & new_n1076;
  assign new_n1966 = ~new_n1962 & ~new_n1963;
  assign new_n1967 = ~new_n1964 & ~new_n1965;
  assign new_n1968 = new_n1966 & new_n1967;
  assign new_n1969 = new_n383 & ~new_n1968;
  assign new_n1970 = ~new_n1945 & ~new_n1953;
  assign new_n1971 = ~new_n1961 & ~new_n1969;
  assign new_n1972 = new_n1970 & new_n1971;
  assign new_n1973 = shift6 & ~new_n1972;
  assign result10 = ~new_n1937 & ~new_n1973;
  assign new_n1975 = new_n265 & new_n1181;
  assign new_n1976 = new_n278 & new_n1281;
  assign new_n1977 = new_n287 & new_n1197;
  assign new_n1978 = new_n296 & new_n1297;
  assign new_n1979 = ~new_n1975 & ~new_n1976;
  assign new_n1980 = ~new_n1977 & ~new_n1978;
  assign new_n1981 = new_n1979 & new_n1980;
  assign new_n1982 = new_n264 & ~new_n1981;
  assign new_n1983 = new_n265 & new_n1217;
  assign new_n1984 = new_n278 & new_n1393;
  assign new_n1985 = new_n287 & new_n1233;
  assign new_n1986 = new_n296 & new_n1409;
  assign new_n1987 = ~new_n1983 & ~new_n1984;
  assign new_n1988 = ~new_n1985 & ~new_n1986;
  assign new_n1989 = new_n1987 & new_n1988;
  assign new_n1990 = new_n309 & ~new_n1989;
  assign new_n1991 = new_n265 & new_n1253;
  assign new_n1992 = new_n278 & new_n1173;
  assign new_n1993 = new_n287 & new_n1269;
  assign new_n1994 = new_n296 & new_n1189;
  assign new_n1995 = ~new_n1991 & ~new_n1992;
  assign new_n1996 = ~new_n1993 & ~new_n1994;
  assign new_n1997 = new_n1995 & new_n1996;
  assign new_n1998 = new_n346 & ~new_n1997;
  assign new_n1999 = new_n265 & new_n1289;
  assign new_n2000 = new_n278 & new_n1209;
  assign new_n2001 = new_n287 & new_n1305;
  assign new_n2002 = new_n296 & new_n1225;
  assign new_n2003 = ~new_n1999 & ~new_n2000;
  assign new_n2004 = ~new_n2001 & ~new_n2002;
  assign new_n2005 = new_n2003 & new_n2004;
  assign new_n2006 = new_n383 & ~new_n2005;
  assign new_n2007 = ~new_n1982 & ~new_n1990;
  assign new_n2008 = ~new_n1998 & ~new_n2006;
  assign new_n2009 = new_n2007 & new_n2008;
  assign new_n2010 = ~shift6 & ~new_n2009;
  assign new_n2011 = new_n265 & new_n1329;
  assign new_n2012 = new_n278 & new_n1429;
  assign new_n2013 = new_n287 & new_n1345;
  assign new_n2014 = new_n296 & new_n1445;
  assign new_n2015 = ~new_n2011 & ~new_n2012;
  assign new_n2016 = ~new_n2013 & ~new_n2014;
  assign new_n2017 = new_n2015 & new_n2016;
  assign new_n2018 = new_n264 & ~new_n2017;
  assign new_n2019 = new_n265 & new_n1365;
  assign new_n2020 = new_n278 & new_n1245;
  assign new_n2021 = new_n287 & new_n1381;
  assign new_n2022 = new_n296 & new_n1261;
  assign new_n2023 = ~new_n2019 & ~new_n2020;
  assign new_n2024 = ~new_n2021 & ~new_n2022;
  assign new_n2025 = new_n2023 & new_n2024;
  assign new_n2026 = new_n309 & ~new_n2025;
  assign new_n2027 = new_n265 & new_n1401;
  assign new_n2028 = new_n278 & new_n1321;
  assign new_n2029 = new_n287 & new_n1417;
  assign new_n2030 = new_n296 & new_n1337;
  assign new_n2031 = ~new_n2027 & ~new_n2028;
  assign new_n2032 = ~new_n2029 & ~new_n2030;
  assign new_n2033 = new_n2031 & new_n2032;
  assign new_n2034 = new_n346 & ~new_n2033;
  assign new_n2035 = new_n265 & new_n1437;
  assign new_n2036 = new_n278 & new_n1357;
  assign new_n2037 = new_n287 & new_n1453;
  assign new_n2038 = new_n296 & new_n1373;
  assign new_n2039 = ~new_n2035 & ~new_n2036;
  assign new_n2040 = ~new_n2037 & ~new_n2038;
  assign new_n2041 = new_n2039 & new_n2040;
  assign new_n2042 = new_n383 & ~new_n2041;
  assign new_n2043 = ~new_n2018 & ~new_n2026;
  assign new_n2044 = ~new_n2034 & ~new_n2042;
  assign new_n2045 = new_n2043 & new_n2044;
  assign new_n2046 = shift6 & ~new_n2045;
  assign result11 = ~new_n2010 & ~new_n2046;
  assign new_n2048 = new_n265 & new_n406;
  assign new_n2049 = new_n278 & new_n414;
  assign new_n2050 = new_n285 & new_n287;
  assign new_n2051 = new_n296 & new_n390;
  assign new_n2052 = ~new_n2048 & ~new_n2049;
  assign new_n2053 = ~new_n2050 & ~new_n2051;
  assign new_n2054 = new_n2052 & new_n2053;
  assign new_n2055 = new_n264 & ~new_n2054;
  assign new_n2056 = new_n265 & new_n518;
  assign new_n2057 = new_n278 & new_n526;
  assign new_n2058 = new_n287 & new_n324;
  assign new_n2059 = new_n296 & new_n502;
  assign new_n2060 = ~new_n2056 & ~new_n2057;
  assign new_n2061 = ~new_n2058 & ~new_n2059;
  assign new_n2062 = new_n2060 & new_n2061;
  assign new_n2063 = new_n309 & ~new_n2062;
  assign new_n2064 = new_n265 & new_n294;
  assign new_n2065 = new_n278 & new_n303;
  assign new_n2066 = new_n287 & new_n361;
  assign new_n2067 = new_n276 & new_n296;
  assign new_n2068 = ~new_n2064 & ~new_n2065;
  assign new_n2069 = ~new_n2066 & ~new_n2067;
  assign new_n2070 = new_n2068 & new_n2069;
  assign new_n2071 = new_n346 & ~new_n2070;
  assign new_n2072 = new_n265 & new_n332;
  assign new_n2073 = new_n278 & new_n340;
  assign new_n2074 = new_n287 & new_n398;
  assign new_n2075 = new_n296 & new_n316;
  assign new_n2076 = ~new_n2072 & ~new_n2073;
  assign new_n2077 = ~new_n2074 & ~new_n2075;
  assign new_n2078 = new_n2076 & new_n2077;
  assign new_n2079 = new_n383 & ~new_n2078;
  assign new_n2080 = ~new_n2055 & ~new_n2063;
  assign new_n2081 = ~new_n2071 & ~new_n2079;
  assign new_n2082 = new_n2080 & new_n2081;
  assign new_n2083 = ~shift6 & ~new_n2082;
  assign new_n2084 = new_n265 & new_n554;
  assign new_n2085 = new_n278 & new_n562;
  assign new_n2086 = new_n287 & new_n438;
  assign new_n2087 = new_n296 & new_n538;
  assign new_n2088 = ~new_n2084 & ~new_n2085;
  assign new_n2089 = ~new_n2086 & ~new_n2087;
  assign new_n2090 = new_n2088 & new_n2089;
  assign new_n2091 = new_n264 & ~new_n2090;
  assign new_n2092 = new_n265 & new_n369;
  assign new_n2093 = new_n278 & new_n377;
  assign new_n2094 = new_n287 & new_n474;
  assign new_n2095 = new_n296 & new_n353;
  assign new_n2096 = ~new_n2092 & ~new_n2093;
  assign new_n2097 = ~new_n2094 & ~new_n2095;
  assign new_n2098 = new_n2096 & new_n2097;
  assign new_n2099 = new_n309 & ~new_n2098;
  assign new_n2100 = new_n265 & new_n446;
  assign new_n2101 = new_n278 & new_n454;
  assign new_n2102 = new_n287 & new_n510;
  assign new_n2103 = new_n296 & new_n430;
  assign new_n2104 = ~new_n2100 & ~new_n2101;
  assign new_n2105 = ~new_n2102 & ~new_n2103;
  assign new_n2106 = new_n2104 & new_n2105;
  assign new_n2107 = new_n346 & ~new_n2106;
  assign new_n2108 = new_n265 & new_n482;
  assign new_n2109 = new_n278 & new_n490;
  assign new_n2110 = new_n287 & new_n546;
  assign new_n2111 = new_n296 & new_n466;
  assign new_n2112 = ~new_n2108 & ~new_n2109;
  assign new_n2113 = ~new_n2110 & ~new_n2111;
  assign new_n2114 = new_n2112 & new_n2113;
  assign new_n2115 = new_n383 & ~new_n2114;
  assign new_n2116 = ~new_n2091 & ~new_n2099;
  assign new_n2117 = ~new_n2107 & ~new_n2115;
  assign new_n2118 = new_n2116 & new_n2117;
  assign new_n2119 = shift6 & ~new_n2118;
  assign result12 = ~new_n2083 & ~new_n2119;
  assign new_n2121 = new_n265 & new_n703;
  assign new_n2122 = new_n278 & new_n711;
  assign new_n2123 = new_n287 & new_n587;
  assign new_n2124 = new_n296 & new_n687;
  assign new_n2125 = ~new_n2121 & ~new_n2122;
  assign new_n2126 = ~new_n2123 & ~new_n2124;
  assign new_n2127 = new_n2125 & new_n2126;
  assign new_n2128 = new_n264 & ~new_n2127;
  assign new_n2129 = new_n265 & new_n815;
  assign new_n2130 = new_n278 & new_n823;
  assign new_n2131 = new_n287 & new_n623;
  assign new_n2132 = new_n296 & new_n799;
  assign new_n2133 = ~new_n2129 & ~new_n2130;
  assign new_n2134 = ~new_n2131 & ~new_n2132;
  assign new_n2135 = new_n2133 & new_n2134;
  assign new_n2136 = new_n309 & ~new_n2135;
  assign new_n2137 = new_n265 & new_n595;
  assign new_n2138 = new_n278 & new_n603;
  assign new_n2139 = new_n287 & new_n659;
  assign new_n2140 = new_n296 & new_n579;
  assign new_n2141 = ~new_n2137 & ~new_n2138;
  assign new_n2142 = ~new_n2139 & ~new_n2140;
  assign new_n2143 = new_n2141 & new_n2142;
  assign new_n2144 = new_n346 & ~new_n2143;
  assign new_n2145 = new_n265 & new_n631;
  assign new_n2146 = new_n278 & new_n639;
  assign new_n2147 = new_n287 & new_n695;
  assign new_n2148 = new_n296 & new_n615;
  assign new_n2149 = ~new_n2145 & ~new_n2146;
  assign new_n2150 = ~new_n2147 & ~new_n2148;
  assign new_n2151 = new_n2149 & new_n2150;
  assign new_n2152 = new_n383 & ~new_n2151;
  assign new_n2153 = ~new_n2128 & ~new_n2136;
  assign new_n2154 = ~new_n2144 & ~new_n2152;
  assign new_n2155 = new_n2153 & new_n2154;
  assign new_n2156 = ~shift6 & ~new_n2155;
  assign new_n2157 = new_n265 & new_n851;
  assign new_n2158 = new_n278 & new_n859;
  assign new_n2159 = new_n287 & new_n735;
  assign new_n2160 = new_n296 & new_n835;
  assign new_n2161 = ~new_n2157 & ~new_n2158;
  assign new_n2162 = ~new_n2159 & ~new_n2160;
  assign new_n2163 = new_n2161 & new_n2162;
  assign new_n2164 = new_n264 & ~new_n2163;
  assign new_n2165 = new_n265 & new_n667;
  assign new_n2166 = new_n278 & new_n675;
  assign new_n2167 = new_n287 & new_n771;
  assign new_n2168 = new_n296 & new_n651;
  assign new_n2169 = ~new_n2165 & ~new_n2166;
  assign new_n2170 = ~new_n2167 & ~new_n2168;
  assign new_n2171 = new_n2169 & new_n2170;
  assign new_n2172 = new_n309 & ~new_n2171;
  assign new_n2173 = new_n265 & new_n743;
  assign new_n2174 = new_n278 & new_n751;
  assign new_n2175 = new_n287 & new_n807;
  assign new_n2176 = new_n296 & new_n727;
  assign new_n2177 = ~new_n2173 & ~new_n2174;
  assign new_n2178 = ~new_n2175 & ~new_n2176;
  assign new_n2179 = new_n2177 & new_n2178;
  assign new_n2180 = new_n346 & ~new_n2179;
  assign new_n2181 = new_n265 & new_n779;
  assign new_n2182 = new_n278 & new_n787;
  assign new_n2183 = new_n287 & new_n843;
  assign new_n2184 = new_n296 & new_n763;
  assign new_n2185 = ~new_n2181 & ~new_n2182;
  assign new_n2186 = ~new_n2183 & ~new_n2184;
  assign new_n2187 = new_n2185 & new_n2186;
  assign new_n2188 = new_n383 & ~new_n2187;
  assign new_n2189 = ~new_n2164 & ~new_n2172;
  assign new_n2190 = ~new_n2180 & ~new_n2188;
  assign new_n2191 = new_n2189 & new_n2190;
  assign new_n2192 = shift6 & ~new_n2191;
  assign result13 = ~new_n2156 & ~new_n2192;
  assign new_n2194 = new_n265 & new_n1000;
  assign new_n2195 = new_n278 & new_n1008;
  assign new_n2196 = new_n287 & new_n884;
  assign new_n2197 = new_n296 & new_n984;
  assign new_n2198 = ~new_n2194 & ~new_n2195;
  assign new_n2199 = ~new_n2196 & ~new_n2197;
  assign new_n2200 = new_n2198 & new_n2199;
  assign new_n2201 = new_n264 & ~new_n2200;
  assign new_n2202 = new_n265 & new_n1112;
  assign new_n2203 = new_n278 & new_n1120;
  assign new_n2204 = new_n287 & new_n920;
  assign new_n2205 = new_n296 & new_n1096;
  assign new_n2206 = ~new_n2202 & ~new_n2203;
  assign new_n2207 = ~new_n2204 & ~new_n2205;
  assign new_n2208 = new_n2206 & new_n2207;
  assign new_n2209 = new_n309 & ~new_n2208;
  assign new_n2210 = new_n265 & new_n892;
  assign new_n2211 = new_n278 & new_n900;
  assign new_n2212 = new_n287 & new_n956;
  assign new_n2213 = new_n296 & new_n876;
  assign new_n2214 = ~new_n2210 & ~new_n2211;
  assign new_n2215 = ~new_n2212 & ~new_n2213;
  assign new_n2216 = new_n2214 & new_n2215;
  assign new_n2217 = new_n346 & ~new_n2216;
  assign new_n2218 = new_n265 & new_n928;
  assign new_n2219 = new_n278 & new_n936;
  assign new_n2220 = new_n287 & new_n992;
  assign new_n2221 = new_n296 & new_n912;
  assign new_n2222 = ~new_n2218 & ~new_n2219;
  assign new_n2223 = ~new_n2220 & ~new_n2221;
  assign new_n2224 = new_n2222 & new_n2223;
  assign new_n2225 = new_n383 & ~new_n2224;
  assign new_n2226 = ~new_n2201 & ~new_n2209;
  assign new_n2227 = ~new_n2217 & ~new_n2225;
  assign new_n2228 = new_n2226 & new_n2227;
  assign new_n2229 = ~shift6 & ~new_n2228;
  assign new_n2230 = new_n265 & new_n1148;
  assign new_n2231 = new_n278 & new_n1156;
  assign new_n2232 = new_n287 & new_n1032;
  assign new_n2233 = new_n296 & new_n1132;
  assign new_n2234 = ~new_n2230 & ~new_n2231;
  assign new_n2235 = ~new_n2232 & ~new_n2233;
  assign new_n2236 = new_n2234 & new_n2235;
  assign new_n2237 = new_n264 & ~new_n2236;
  assign new_n2238 = new_n265 & new_n964;
  assign new_n2239 = new_n278 & new_n972;
  assign new_n2240 = new_n287 & new_n1068;
  assign new_n2241 = new_n296 & new_n948;
  assign new_n2242 = ~new_n2238 & ~new_n2239;
  assign new_n2243 = ~new_n2240 & ~new_n2241;
  assign new_n2244 = new_n2242 & new_n2243;
  assign new_n2245 = new_n309 & ~new_n2244;
  assign new_n2246 = new_n265 & new_n1040;
  assign new_n2247 = new_n278 & new_n1048;
  assign new_n2248 = new_n287 & new_n1104;
  assign new_n2249 = new_n296 & new_n1024;
  assign new_n2250 = ~new_n2246 & ~new_n2247;
  assign new_n2251 = ~new_n2248 & ~new_n2249;
  assign new_n2252 = new_n2250 & new_n2251;
  assign new_n2253 = new_n346 & ~new_n2252;
  assign new_n2254 = new_n265 & new_n1076;
  assign new_n2255 = new_n278 & new_n1084;
  assign new_n2256 = new_n287 & new_n1140;
  assign new_n2257 = new_n296 & new_n1060;
  assign new_n2258 = ~new_n2254 & ~new_n2255;
  assign new_n2259 = ~new_n2256 & ~new_n2257;
  assign new_n2260 = new_n2258 & new_n2259;
  assign new_n2261 = new_n383 & ~new_n2260;
  assign new_n2262 = ~new_n2237 & ~new_n2245;
  assign new_n2263 = ~new_n2253 & ~new_n2261;
  assign new_n2264 = new_n2262 & new_n2263;
  assign new_n2265 = shift6 & ~new_n2264;
  assign result14 = ~new_n2229 & ~new_n2265;
  assign new_n2267 = new_n265 & new_n1297;
  assign new_n2268 = new_n278 & new_n1305;
  assign new_n2269 = new_n287 & new_n1181;
  assign new_n2270 = new_n296 & new_n1281;
  assign new_n2271 = ~new_n2267 & ~new_n2268;
  assign new_n2272 = ~new_n2269 & ~new_n2270;
  assign new_n2273 = new_n2271 & new_n2272;
  assign new_n2274 = new_n264 & ~new_n2273;
  assign new_n2275 = new_n265 & new_n1409;
  assign new_n2276 = new_n278 & new_n1417;
  assign new_n2277 = new_n287 & new_n1217;
  assign new_n2278 = new_n296 & new_n1393;
  assign new_n2279 = ~new_n2275 & ~new_n2276;
  assign new_n2280 = ~new_n2277 & ~new_n2278;
  assign new_n2281 = new_n2279 & new_n2280;
  assign new_n2282 = new_n309 & ~new_n2281;
  assign new_n2283 = new_n265 & new_n1189;
  assign new_n2284 = new_n278 & new_n1197;
  assign new_n2285 = new_n287 & new_n1253;
  assign new_n2286 = new_n296 & new_n1173;
  assign new_n2287 = ~new_n2283 & ~new_n2284;
  assign new_n2288 = ~new_n2285 & ~new_n2286;
  assign new_n2289 = new_n2287 & new_n2288;
  assign new_n2290 = new_n346 & ~new_n2289;
  assign new_n2291 = new_n265 & new_n1225;
  assign new_n2292 = new_n278 & new_n1233;
  assign new_n2293 = new_n287 & new_n1289;
  assign new_n2294 = new_n296 & new_n1209;
  assign new_n2295 = ~new_n2291 & ~new_n2292;
  assign new_n2296 = ~new_n2293 & ~new_n2294;
  assign new_n2297 = new_n2295 & new_n2296;
  assign new_n2298 = new_n383 & ~new_n2297;
  assign new_n2299 = ~new_n2274 & ~new_n2282;
  assign new_n2300 = ~new_n2290 & ~new_n2298;
  assign new_n2301 = new_n2299 & new_n2300;
  assign new_n2302 = ~shift6 & ~new_n2301;
  assign new_n2303 = new_n265 & new_n1445;
  assign new_n2304 = new_n278 & new_n1453;
  assign new_n2305 = new_n287 & new_n1329;
  assign new_n2306 = new_n296 & new_n1429;
  assign new_n2307 = ~new_n2303 & ~new_n2304;
  assign new_n2308 = ~new_n2305 & ~new_n2306;
  assign new_n2309 = new_n2307 & new_n2308;
  assign new_n2310 = new_n264 & ~new_n2309;
  assign new_n2311 = new_n265 & new_n1261;
  assign new_n2312 = new_n278 & new_n1269;
  assign new_n2313 = new_n287 & new_n1365;
  assign new_n2314 = new_n296 & new_n1245;
  assign new_n2315 = ~new_n2311 & ~new_n2312;
  assign new_n2316 = ~new_n2313 & ~new_n2314;
  assign new_n2317 = new_n2315 & new_n2316;
  assign new_n2318 = new_n309 & ~new_n2317;
  assign new_n2319 = new_n265 & new_n1337;
  assign new_n2320 = new_n278 & new_n1345;
  assign new_n2321 = new_n287 & new_n1401;
  assign new_n2322 = new_n296 & new_n1321;
  assign new_n2323 = ~new_n2319 & ~new_n2320;
  assign new_n2324 = ~new_n2321 & ~new_n2322;
  assign new_n2325 = new_n2323 & new_n2324;
  assign new_n2326 = new_n346 & ~new_n2325;
  assign new_n2327 = new_n265 & new_n1373;
  assign new_n2328 = new_n278 & new_n1381;
  assign new_n2329 = new_n287 & new_n1437;
  assign new_n2330 = new_n296 & new_n1357;
  assign new_n2331 = ~new_n2327 & ~new_n2328;
  assign new_n2332 = ~new_n2329 & ~new_n2330;
  assign new_n2333 = new_n2331 & new_n2332;
  assign new_n2334 = new_n383 & ~new_n2333;
  assign new_n2335 = ~new_n2310 & ~new_n2318;
  assign new_n2336 = ~new_n2326 & ~new_n2334;
  assign new_n2337 = new_n2335 & new_n2336;
  assign new_n2338 = shift6 & ~new_n2337;
  assign result15 = ~new_n2302 & ~new_n2338;
  assign new_n2340 = new_n264 & ~new_n418;
  assign new_n2341 = new_n309 & ~new_n530;
  assign new_n2342 = ~new_n307 & new_n346;
  assign new_n2343 = ~new_n344 & new_n383;
  assign new_n2344 = ~new_n2340 & ~new_n2341;
  assign new_n2345 = ~new_n2342 & ~new_n2343;
  assign new_n2346 = new_n2344 & new_n2345;
  assign new_n2347 = ~shift6 & ~new_n2346;
  assign new_n2348 = new_n264 & ~new_n566;
  assign new_n2349 = new_n309 & ~new_n381;
  assign new_n2350 = new_n346 & ~new_n458;
  assign new_n2351 = new_n383 & ~new_n494;
  assign new_n2352 = ~new_n2348 & ~new_n2349;
  assign new_n2353 = ~new_n2350 & ~new_n2351;
  assign new_n2354 = new_n2352 & new_n2353;
  assign new_n2355 = shift6 & ~new_n2354;
  assign result16 = ~new_n2347 & ~new_n2355;
  assign new_n2357 = new_n264 & ~new_n715;
  assign new_n2358 = new_n309 & ~new_n827;
  assign new_n2359 = new_n346 & ~new_n607;
  assign new_n2360 = new_n383 & ~new_n643;
  assign new_n2361 = ~new_n2357 & ~new_n2358;
  assign new_n2362 = ~new_n2359 & ~new_n2360;
  assign new_n2363 = new_n2361 & new_n2362;
  assign new_n2364 = ~shift6 & ~new_n2363;
  assign new_n2365 = new_n264 & ~new_n863;
  assign new_n2366 = new_n309 & ~new_n679;
  assign new_n2367 = new_n346 & ~new_n755;
  assign new_n2368 = new_n383 & ~new_n791;
  assign new_n2369 = ~new_n2365 & ~new_n2366;
  assign new_n2370 = ~new_n2367 & ~new_n2368;
  assign new_n2371 = new_n2369 & new_n2370;
  assign new_n2372 = shift6 & ~new_n2371;
  assign result17 = ~new_n2364 & ~new_n2372;
  assign new_n2374 = new_n264 & ~new_n1012;
  assign new_n2375 = new_n309 & ~new_n1124;
  assign new_n2376 = new_n346 & ~new_n904;
  assign new_n2377 = new_n383 & ~new_n940;
  assign new_n2378 = ~new_n2374 & ~new_n2375;
  assign new_n2379 = ~new_n2376 & ~new_n2377;
  assign new_n2380 = new_n2378 & new_n2379;
  assign new_n2381 = ~shift6 & ~new_n2380;
  assign new_n2382 = new_n264 & ~new_n1160;
  assign new_n2383 = new_n309 & ~new_n976;
  assign new_n2384 = new_n346 & ~new_n1052;
  assign new_n2385 = new_n383 & ~new_n1088;
  assign new_n2386 = ~new_n2382 & ~new_n2383;
  assign new_n2387 = ~new_n2384 & ~new_n2385;
  assign new_n2388 = new_n2386 & new_n2387;
  assign new_n2389 = shift6 & ~new_n2388;
  assign result18 = ~new_n2381 & ~new_n2389;
  assign new_n2391 = new_n264 & ~new_n1309;
  assign new_n2392 = new_n309 & ~new_n1421;
  assign new_n2393 = new_n346 & ~new_n1201;
  assign new_n2394 = new_n383 & ~new_n1237;
  assign new_n2395 = ~new_n2391 & ~new_n2392;
  assign new_n2396 = ~new_n2393 & ~new_n2394;
  assign new_n2397 = new_n2395 & new_n2396;
  assign new_n2398 = ~shift6 & ~new_n2397;
  assign new_n2399 = new_n264 & ~new_n1457;
  assign new_n2400 = new_n309 & ~new_n1273;
  assign new_n2401 = new_n346 & ~new_n1349;
  assign new_n2402 = new_n383 & ~new_n1385;
  assign new_n2403 = ~new_n2399 & ~new_n2400;
  assign new_n2404 = ~new_n2401 & ~new_n2402;
  assign new_n2405 = new_n2403 & new_n2404;
  assign new_n2406 = shift6 & ~new_n2405;
  assign result19 = ~new_n2398 & ~new_n2406;
  assign new_n2408 = new_n264 & ~new_n1494;
  assign new_n2409 = new_n309 & ~new_n1522;
  assign new_n2410 = new_n346 & ~new_n1470;
  assign new_n2411 = new_n383 & ~new_n1478;
  assign new_n2412 = ~new_n2408 & ~new_n2409;
  assign new_n2413 = ~new_n2410 & ~new_n2411;
  assign new_n2414 = new_n2412 & new_n2413;
  assign new_n2415 = ~shift6 & ~new_n2414;
  assign new_n2416 = new_n264 & ~new_n1530;
  assign new_n2417 = new_n309 & ~new_n1486;
  assign new_n2418 = new_n346 & ~new_n1506;
  assign new_n2419 = new_n383 & ~new_n1514;
  assign new_n2420 = ~new_n2416 & ~new_n2417;
  assign new_n2421 = ~new_n2418 & ~new_n2419;
  assign new_n2422 = new_n2420 & new_n2421;
  assign new_n2423 = shift6 & ~new_n2422;
  assign result20 = ~new_n2415 & ~new_n2423;
  assign new_n2425 = new_n264 & ~new_n1567;
  assign new_n2426 = new_n309 & ~new_n1595;
  assign new_n2427 = new_n346 & ~new_n1543;
  assign new_n2428 = new_n383 & ~new_n1551;
  assign new_n2429 = ~new_n2425 & ~new_n2426;
  assign new_n2430 = ~new_n2427 & ~new_n2428;
  assign new_n2431 = new_n2429 & new_n2430;
  assign new_n2432 = ~shift6 & ~new_n2431;
  assign new_n2433 = new_n264 & ~new_n1603;
  assign new_n2434 = new_n309 & ~new_n1559;
  assign new_n2435 = new_n346 & ~new_n1579;
  assign new_n2436 = new_n383 & ~new_n1587;
  assign new_n2437 = ~new_n2433 & ~new_n2434;
  assign new_n2438 = ~new_n2435 & ~new_n2436;
  assign new_n2439 = new_n2437 & new_n2438;
  assign new_n2440 = shift6 & ~new_n2439;
  assign result21 = ~new_n2432 & ~new_n2440;
  assign new_n2442 = new_n264 & ~new_n1640;
  assign new_n2443 = new_n309 & ~new_n1668;
  assign new_n2444 = new_n346 & ~new_n1616;
  assign new_n2445 = new_n383 & ~new_n1624;
  assign new_n2446 = ~new_n2442 & ~new_n2443;
  assign new_n2447 = ~new_n2444 & ~new_n2445;
  assign new_n2448 = new_n2446 & new_n2447;
  assign new_n2449 = ~shift6 & ~new_n2448;
  assign new_n2450 = new_n264 & ~new_n1676;
  assign new_n2451 = new_n309 & ~new_n1632;
  assign new_n2452 = new_n346 & ~new_n1652;
  assign new_n2453 = new_n383 & ~new_n1660;
  assign new_n2454 = ~new_n2450 & ~new_n2451;
  assign new_n2455 = ~new_n2452 & ~new_n2453;
  assign new_n2456 = new_n2454 & new_n2455;
  assign new_n2457 = shift6 & ~new_n2456;
  assign result22 = ~new_n2449 & ~new_n2457;
  assign new_n2459 = new_n264 & ~new_n1713;
  assign new_n2460 = new_n309 & ~new_n1741;
  assign new_n2461 = new_n346 & ~new_n1689;
  assign new_n2462 = new_n383 & ~new_n1697;
  assign new_n2463 = ~new_n2459 & ~new_n2460;
  assign new_n2464 = ~new_n2461 & ~new_n2462;
  assign new_n2465 = new_n2463 & new_n2464;
  assign new_n2466 = ~shift6 & ~new_n2465;
  assign new_n2467 = new_n264 & ~new_n1749;
  assign new_n2468 = new_n309 & ~new_n1705;
  assign new_n2469 = new_n346 & ~new_n1725;
  assign new_n2470 = new_n383 & ~new_n1733;
  assign new_n2471 = ~new_n2467 & ~new_n2468;
  assign new_n2472 = ~new_n2469 & ~new_n2470;
  assign new_n2473 = new_n2471 & new_n2472;
  assign new_n2474 = shift6 & ~new_n2473;
  assign result23 = ~new_n2466 & ~new_n2474;
  assign new_n2476 = new_n264 & ~new_n1786;
  assign new_n2477 = new_n309 & ~new_n1814;
  assign new_n2478 = new_n346 & ~new_n1762;
  assign new_n2479 = new_n383 & ~new_n1770;
  assign new_n2480 = ~new_n2476 & ~new_n2477;
  assign new_n2481 = ~new_n2478 & ~new_n2479;
  assign new_n2482 = new_n2480 & new_n2481;
  assign new_n2483 = ~shift6 & ~new_n2482;
  assign new_n2484 = new_n264 & ~new_n1822;
  assign new_n2485 = new_n309 & ~new_n1778;
  assign new_n2486 = new_n346 & ~new_n1798;
  assign new_n2487 = new_n383 & ~new_n1806;
  assign new_n2488 = ~new_n2484 & ~new_n2485;
  assign new_n2489 = ~new_n2486 & ~new_n2487;
  assign new_n2490 = new_n2488 & new_n2489;
  assign new_n2491 = shift6 & ~new_n2490;
  assign result24 = ~new_n2483 & ~new_n2491;
  assign new_n2493 = new_n264 & ~new_n1859;
  assign new_n2494 = new_n309 & ~new_n1887;
  assign new_n2495 = new_n346 & ~new_n1835;
  assign new_n2496 = new_n383 & ~new_n1843;
  assign new_n2497 = ~new_n2493 & ~new_n2494;
  assign new_n2498 = ~new_n2495 & ~new_n2496;
  assign new_n2499 = new_n2497 & new_n2498;
  assign new_n2500 = ~shift6 & ~new_n2499;
  assign new_n2501 = new_n264 & ~new_n1895;
  assign new_n2502 = new_n309 & ~new_n1851;
  assign new_n2503 = new_n346 & ~new_n1871;
  assign new_n2504 = new_n383 & ~new_n1879;
  assign new_n2505 = ~new_n2501 & ~new_n2502;
  assign new_n2506 = ~new_n2503 & ~new_n2504;
  assign new_n2507 = new_n2505 & new_n2506;
  assign new_n2508 = shift6 & ~new_n2507;
  assign result25 = ~new_n2500 & ~new_n2508;
  assign new_n2510 = new_n264 & ~new_n1932;
  assign new_n2511 = new_n309 & ~new_n1960;
  assign new_n2512 = new_n346 & ~new_n1908;
  assign new_n2513 = new_n383 & ~new_n1916;
  assign new_n2514 = ~new_n2510 & ~new_n2511;
  assign new_n2515 = ~new_n2512 & ~new_n2513;
  assign new_n2516 = new_n2514 & new_n2515;
  assign new_n2517 = ~shift6 & ~new_n2516;
  assign new_n2518 = new_n264 & ~new_n1968;
  assign new_n2519 = new_n309 & ~new_n1924;
  assign new_n2520 = new_n346 & ~new_n1944;
  assign new_n2521 = new_n383 & ~new_n1952;
  assign new_n2522 = ~new_n2518 & ~new_n2519;
  assign new_n2523 = ~new_n2520 & ~new_n2521;
  assign new_n2524 = new_n2522 & new_n2523;
  assign new_n2525 = shift6 & ~new_n2524;
  assign result26 = ~new_n2517 & ~new_n2525;
  assign new_n2527 = new_n264 & ~new_n2005;
  assign new_n2528 = new_n309 & ~new_n2033;
  assign new_n2529 = new_n346 & ~new_n1981;
  assign new_n2530 = new_n383 & ~new_n1989;
  assign new_n2531 = ~new_n2527 & ~new_n2528;
  assign new_n2532 = ~new_n2529 & ~new_n2530;
  assign new_n2533 = new_n2531 & new_n2532;
  assign new_n2534 = ~shift6 & ~new_n2533;
  assign new_n2535 = new_n264 & ~new_n2041;
  assign new_n2536 = new_n309 & ~new_n1997;
  assign new_n2537 = new_n346 & ~new_n2017;
  assign new_n2538 = new_n383 & ~new_n2025;
  assign new_n2539 = ~new_n2535 & ~new_n2536;
  assign new_n2540 = ~new_n2537 & ~new_n2538;
  assign new_n2541 = new_n2539 & new_n2540;
  assign new_n2542 = shift6 & ~new_n2541;
  assign result27 = ~new_n2534 & ~new_n2542;
  assign new_n2544 = new_n264 & ~new_n2078;
  assign new_n2545 = new_n309 & ~new_n2106;
  assign new_n2546 = new_n346 & ~new_n2054;
  assign new_n2547 = new_n383 & ~new_n2062;
  assign new_n2548 = ~new_n2544 & ~new_n2545;
  assign new_n2549 = ~new_n2546 & ~new_n2547;
  assign new_n2550 = new_n2548 & new_n2549;
  assign new_n2551 = ~shift6 & ~new_n2550;
  assign new_n2552 = new_n264 & ~new_n2114;
  assign new_n2553 = new_n309 & ~new_n2070;
  assign new_n2554 = new_n346 & ~new_n2090;
  assign new_n2555 = new_n383 & ~new_n2098;
  assign new_n2556 = ~new_n2552 & ~new_n2553;
  assign new_n2557 = ~new_n2554 & ~new_n2555;
  assign new_n2558 = new_n2556 & new_n2557;
  assign new_n2559 = shift6 & ~new_n2558;
  assign result28 = ~new_n2551 & ~new_n2559;
  assign new_n2561 = new_n264 & ~new_n2151;
  assign new_n2562 = new_n309 & ~new_n2179;
  assign new_n2563 = new_n346 & ~new_n2127;
  assign new_n2564 = new_n383 & ~new_n2135;
  assign new_n2565 = ~new_n2561 & ~new_n2562;
  assign new_n2566 = ~new_n2563 & ~new_n2564;
  assign new_n2567 = new_n2565 & new_n2566;
  assign new_n2568 = ~shift6 & ~new_n2567;
  assign new_n2569 = new_n264 & ~new_n2187;
  assign new_n2570 = new_n309 & ~new_n2143;
  assign new_n2571 = new_n346 & ~new_n2163;
  assign new_n2572 = new_n383 & ~new_n2171;
  assign new_n2573 = ~new_n2569 & ~new_n2570;
  assign new_n2574 = ~new_n2571 & ~new_n2572;
  assign new_n2575 = new_n2573 & new_n2574;
  assign new_n2576 = shift6 & ~new_n2575;
  assign result29 = ~new_n2568 & ~new_n2576;
  assign new_n2578 = new_n264 & ~new_n2224;
  assign new_n2579 = new_n309 & ~new_n2252;
  assign new_n2580 = new_n346 & ~new_n2200;
  assign new_n2581 = new_n383 & ~new_n2208;
  assign new_n2582 = ~new_n2578 & ~new_n2579;
  assign new_n2583 = ~new_n2580 & ~new_n2581;
  assign new_n2584 = new_n2582 & new_n2583;
  assign new_n2585 = ~shift6 & ~new_n2584;
  assign new_n2586 = new_n264 & ~new_n2260;
  assign new_n2587 = new_n309 & ~new_n2216;
  assign new_n2588 = new_n346 & ~new_n2236;
  assign new_n2589 = new_n383 & ~new_n2244;
  assign new_n2590 = ~new_n2586 & ~new_n2587;
  assign new_n2591 = ~new_n2588 & ~new_n2589;
  assign new_n2592 = new_n2590 & new_n2591;
  assign new_n2593 = shift6 & ~new_n2592;
  assign result30 = ~new_n2585 & ~new_n2593;
  assign new_n2595 = new_n264 & ~new_n2297;
  assign new_n2596 = new_n309 & ~new_n2325;
  assign new_n2597 = new_n346 & ~new_n2273;
  assign new_n2598 = new_n383 & ~new_n2281;
  assign new_n2599 = ~new_n2595 & ~new_n2596;
  assign new_n2600 = ~new_n2597 & ~new_n2598;
  assign new_n2601 = new_n2599 & new_n2600;
  assign new_n2602 = ~shift6 & ~new_n2601;
  assign new_n2603 = new_n264 & ~new_n2333;
  assign new_n2604 = new_n309 & ~new_n2289;
  assign new_n2605 = new_n346 & ~new_n2309;
  assign new_n2606 = new_n383 & ~new_n2317;
  assign new_n2607 = ~new_n2603 & ~new_n2604;
  assign new_n2608 = ~new_n2605 & ~new_n2606;
  assign new_n2609 = new_n2607 & new_n2608;
  assign new_n2610 = shift6 & ~new_n2609;
  assign result31 = ~new_n2602 & ~new_n2610;
  assign new_n2612 = new_n264 & ~new_n344;
  assign new_n2613 = new_n309 & ~new_n458;
  assign new_n2614 = new_n346 & ~new_n418;
  assign new_n2615 = new_n383 & ~new_n530;
  assign new_n2616 = ~new_n2612 & ~new_n2613;
  assign new_n2617 = ~new_n2614 & ~new_n2615;
  assign new_n2618 = new_n2616 & new_n2617;
  assign new_n2619 = ~shift6 & ~new_n2618;
  assign new_n2620 = new_n264 & ~new_n494;
  assign new_n2621 = ~new_n307 & new_n309;
  assign new_n2622 = new_n346 & ~new_n566;
  assign new_n2623 = ~new_n381 & new_n383;
  assign new_n2624 = ~new_n2620 & ~new_n2621;
  assign new_n2625 = ~new_n2622 & ~new_n2623;
  assign new_n2626 = new_n2624 & new_n2625;
  assign new_n2627 = shift6 & ~new_n2626;
  assign result32 = ~new_n2619 & ~new_n2627;
  assign new_n2629 = new_n264 & ~new_n643;
  assign new_n2630 = new_n309 & ~new_n755;
  assign new_n2631 = new_n346 & ~new_n715;
  assign new_n2632 = new_n383 & ~new_n827;
  assign new_n2633 = ~new_n2629 & ~new_n2630;
  assign new_n2634 = ~new_n2631 & ~new_n2632;
  assign new_n2635 = new_n2633 & new_n2634;
  assign new_n2636 = ~shift6 & ~new_n2635;
  assign new_n2637 = new_n264 & ~new_n791;
  assign new_n2638 = new_n309 & ~new_n607;
  assign new_n2639 = new_n346 & ~new_n863;
  assign new_n2640 = new_n383 & ~new_n679;
  assign new_n2641 = ~new_n2637 & ~new_n2638;
  assign new_n2642 = ~new_n2639 & ~new_n2640;
  assign new_n2643 = new_n2641 & new_n2642;
  assign new_n2644 = shift6 & ~new_n2643;
  assign result33 = ~new_n2636 & ~new_n2644;
  assign new_n2646 = new_n264 & ~new_n940;
  assign new_n2647 = new_n309 & ~new_n1052;
  assign new_n2648 = new_n346 & ~new_n1012;
  assign new_n2649 = new_n383 & ~new_n1124;
  assign new_n2650 = ~new_n2646 & ~new_n2647;
  assign new_n2651 = ~new_n2648 & ~new_n2649;
  assign new_n2652 = new_n2650 & new_n2651;
  assign new_n2653 = ~shift6 & ~new_n2652;
  assign new_n2654 = new_n264 & ~new_n1088;
  assign new_n2655 = new_n309 & ~new_n904;
  assign new_n2656 = new_n346 & ~new_n1160;
  assign new_n2657 = new_n383 & ~new_n976;
  assign new_n2658 = ~new_n2654 & ~new_n2655;
  assign new_n2659 = ~new_n2656 & ~new_n2657;
  assign new_n2660 = new_n2658 & new_n2659;
  assign new_n2661 = shift6 & ~new_n2660;
  assign result34 = ~new_n2653 & ~new_n2661;
  assign new_n2663 = new_n264 & ~new_n1237;
  assign new_n2664 = new_n309 & ~new_n1349;
  assign new_n2665 = new_n346 & ~new_n1309;
  assign new_n2666 = new_n383 & ~new_n1421;
  assign new_n2667 = ~new_n2663 & ~new_n2664;
  assign new_n2668 = ~new_n2665 & ~new_n2666;
  assign new_n2669 = new_n2667 & new_n2668;
  assign new_n2670 = ~shift6 & ~new_n2669;
  assign new_n2671 = new_n264 & ~new_n1385;
  assign new_n2672 = new_n309 & ~new_n1201;
  assign new_n2673 = new_n346 & ~new_n1457;
  assign new_n2674 = new_n383 & ~new_n1273;
  assign new_n2675 = ~new_n2671 & ~new_n2672;
  assign new_n2676 = ~new_n2673 & ~new_n2674;
  assign new_n2677 = new_n2675 & new_n2676;
  assign new_n2678 = shift6 & ~new_n2677;
  assign result35 = ~new_n2670 & ~new_n2678;
  assign new_n2680 = new_n264 & ~new_n1478;
  assign new_n2681 = new_n309 & ~new_n1506;
  assign new_n2682 = new_n346 & ~new_n1494;
  assign new_n2683 = new_n383 & ~new_n1522;
  assign new_n2684 = ~new_n2680 & ~new_n2681;
  assign new_n2685 = ~new_n2682 & ~new_n2683;
  assign new_n2686 = new_n2684 & new_n2685;
  assign new_n2687 = ~shift6 & ~new_n2686;
  assign new_n2688 = new_n264 & ~new_n1514;
  assign new_n2689 = new_n309 & ~new_n1470;
  assign new_n2690 = new_n346 & ~new_n1530;
  assign new_n2691 = new_n383 & ~new_n1486;
  assign new_n2692 = ~new_n2688 & ~new_n2689;
  assign new_n2693 = ~new_n2690 & ~new_n2691;
  assign new_n2694 = new_n2692 & new_n2693;
  assign new_n2695 = shift6 & ~new_n2694;
  assign result36 = ~new_n2687 & ~new_n2695;
  assign new_n2697 = new_n264 & ~new_n1551;
  assign new_n2698 = new_n309 & ~new_n1579;
  assign new_n2699 = new_n346 & ~new_n1567;
  assign new_n2700 = new_n383 & ~new_n1595;
  assign new_n2701 = ~new_n2697 & ~new_n2698;
  assign new_n2702 = ~new_n2699 & ~new_n2700;
  assign new_n2703 = new_n2701 & new_n2702;
  assign new_n2704 = ~shift6 & ~new_n2703;
  assign new_n2705 = new_n264 & ~new_n1587;
  assign new_n2706 = new_n309 & ~new_n1543;
  assign new_n2707 = new_n346 & ~new_n1603;
  assign new_n2708 = new_n383 & ~new_n1559;
  assign new_n2709 = ~new_n2705 & ~new_n2706;
  assign new_n2710 = ~new_n2707 & ~new_n2708;
  assign new_n2711 = new_n2709 & new_n2710;
  assign new_n2712 = shift6 & ~new_n2711;
  assign result37 = ~new_n2704 & ~new_n2712;
  assign new_n2714 = new_n264 & ~new_n1624;
  assign new_n2715 = new_n309 & ~new_n1652;
  assign new_n2716 = new_n346 & ~new_n1640;
  assign new_n2717 = new_n383 & ~new_n1668;
  assign new_n2718 = ~new_n2714 & ~new_n2715;
  assign new_n2719 = ~new_n2716 & ~new_n2717;
  assign new_n2720 = new_n2718 & new_n2719;
  assign new_n2721 = ~shift6 & ~new_n2720;
  assign new_n2722 = new_n264 & ~new_n1660;
  assign new_n2723 = new_n309 & ~new_n1616;
  assign new_n2724 = new_n346 & ~new_n1676;
  assign new_n2725 = new_n383 & ~new_n1632;
  assign new_n2726 = ~new_n2722 & ~new_n2723;
  assign new_n2727 = ~new_n2724 & ~new_n2725;
  assign new_n2728 = new_n2726 & new_n2727;
  assign new_n2729 = shift6 & ~new_n2728;
  assign result38 = ~new_n2721 & ~new_n2729;
  assign new_n2731 = new_n264 & ~new_n1697;
  assign new_n2732 = new_n309 & ~new_n1725;
  assign new_n2733 = new_n346 & ~new_n1713;
  assign new_n2734 = new_n383 & ~new_n1741;
  assign new_n2735 = ~new_n2731 & ~new_n2732;
  assign new_n2736 = ~new_n2733 & ~new_n2734;
  assign new_n2737 = new_n2735 & new_n2736;
  assign new_n2738 = ~shift6 & ~new_n2737;
  assign new_n2739 = new_n264 & ~new_n1733;
  assign new_n2740 = new_n309 & ~new_n1689;
  assign new_n2741 = new_n346 & ~new_n1749;
  assign new_n2742 = new_n383 & ~new_n1705;
  assign new_n2743 = ~new_n2739 & ~new_n2740;
  assign new_n2744 = ~new_n2741 & ~new_n2742;
  assign new_n2745 = new_n2743 & new_n2744;
  assign new_n2746 = shift6 & ~new_n2745;
  assign result39 = ~new_n2738 & ~new_n2746;
  assign new_n2748 = new_n264 & ~new_n1770;
  assign new_n2749 = new_n309 & ~new_n1798;
  assign new_n2750 = new_n346 & ~new_n1786;
  assign new_n2751 = new_n383 & ~new_n1814;
  assign new_n2752 = ~new_n2748 & ~new_n2749;
  assign new_n2753 = ~new_n2750 & ~new_n2751;
  assign new_n2754 = new_n2752 & new_n2753;
  assign new_n2755 = ~shift6 & ~new_n2754;
  assign new_n2756 = new_n264 & ~new_n1806;
  assign new_n2757 = new_n309 & ~new_n1762;
  assign new_n2758 = new_n346 & ~new_n1822;
  assign new_n2759 = new_n383 & ~new_n1778;
  assign new_n2760 = ~new_n2756 & ~new_n2757;
  assign new_n2761 = ~new_n2758 & ~new_n2759;
  assign new_n2762 = new_n2760 & new_n2761;
  assign new_n2763 = shift6 & ~new_n2762;
  assign result40 = ~new_n2755 & ~new_n2763;
  assign new_n2765 = new_n264 & ~new_n1843;
  assign new_n2766 = new_n309 & ~new_n1871;
  assign new_n2767 = new_n346 & ~new_n1859;
  assign new_n2768 = new_n383 & ~new_n1887;
  assign new_n2769 = ~new_n2765 & ~new_n2766;
  assign new_n2770 = ~new_n2767 & ~new_n2768;
  assign new_n2771 = new_n2769 & new_n2770;
  assign new_n2772 = ~shift6 & ~new_n2771;
  assign new_n2773 = new_n264 & ~new_n1879;
  assign new_n2774 = new_n309 & ~new_n1835;
  assign new_n2775 = new_n346 & ~new_n1895;
  assign new_n2776 = new_n383 & ~new_n1851;
  assign new_n2777 = ~new_n2773 & ~new_n2774;
  assign new_n2778 = ~new_n2775 & ~new_n2776;
  assign new_n2779 = new_n2777 & new_n2778;
  assign new_n2780 = shift6 & ~new_n2779;
  assign result41 = ~new_n2772 & ~new_n2780;
  assign new_n2782 = new_n264 & ~new_n1916;
  assign new_n2783 = new_n309 & ~new_n1944;
  assign new_n2784 = new_n346 & ~new_n1932;
  assign new_n2785 = new_n383 & ~new_n1960;
  assign new_n2786 = ~new_n2782 & ~new_n2783;
  assign new_n2787 = ~new_n2784 & ~new_n2785;
  assign new_n2788 = new_n2786 & new_n2787;
  assign new_n2789 = ~shift6 & ~new_n2788;
  assign new_n2790 = new_n264 & ~new_n1952;
  assign new_n2791 = new_n309 & ~new_n1908;
  assign new_n2792 = new_n346 & ~new_n1968;
  assign new_n2793 = new_n383 & ~new_n1924;
  assign new_n2794 = ~new_n2790 & ~new_n2791;
  assign new_n2795 = ~new_n2792 & ~new_n2793;
  assign new_n2796 = new_n2794 & new_n2795;
  assign new_n2797 = shift6 & ~new_n2796;
  assign result42 = ~new_n2789 & ~new_n2797;
  assign new_n2799 = new_n264 & ~new_n1989;
  assign new_n2800 = new_n309 & ~new_n2017;
  assign new_n2801 = new_n346 & ~new_n2005;
  assign new_n2802 = new_n383 & ~new_n2033;
  assign new_n2803 = ~new_n2799 & ~new_n2800;
  assign new_n2804 = ~new_n2801 & ~new_n2802;
  assign new_n2805 = new_n2803 & new_n2804;
  assign new_n2806 = ~shift6 & ~new_n2805;
  assign new_n2807 = new_n264 & ~new_n2025;
  assign new_n2808 = new_n309 & ~new_n1981;
  assign new_n2809 = new_n346 & ~new_n2041;
  assign new_n2810 = new_n383 & ~new_n1997;
  assign new_n2811 = ~new_n2807 & ~new_n2808;
  assign new_n2812 = ~new_n2809 & ~new_n2810;
  assign new_n2813 = new_n2811 & new_n2812;
  assign new_n2814 = shift6 & ~new_n2813;
  assign result43 = ~new_n2806 & ~new_n2814;
  assign new_n2816 = new_n264 & ~new_n2062;
  assign new_n2817 = new_n309 & ~new_n2090;
  assign new_n2818 = new_n346 & ~new_n2078;
  assign new_n2819 = new_n383 & ~new_n2106;
  assign new_n2820 = ~new_n2816 & ~new_n2817;
  assign new_n2821 = ~new_n2818 & ~new_n2819;
  assign new_n2822 = new_n2820 & new_n2821;
  assign new_n2823 = ~shift6 & ~new_n2822;
  assign new_n2824 = new_n264 & ~new_n2098;
  assign new_n2825 = new_n309 & ~new_n2054;
  assign new_n2826 = new_n346 & ~new_n2114;
  assign new_n2827 = new_n383 & ~new_n2070;
  assign new_n2828 = ~new_n2824 & ~new_n2825;
  assign new_n2829 = ~new_n2826 & ~new_n2827;
  assign new_n2830 = new_n2828 & new_n2829;
  assign new_n2831 = shift6 & ~new_n2830;
  assign result44 = ~new_n2823 & ~new_n2831;
  assign new_n2833 = new_n264 & ~new_n2135;
  assign new_n2834 = new_n309 & ~new_n2163;
  assign new_n2835 = new_n346 & ~new_n2151;
  assign new_n2836 = new_n383 & ~new_n2179;
  assign new_n2837 = ~new_n2833 & ~new_n2834;
  assign new_n2838 = ~new_n2835 & ~new_n2836;
  assign new_n2839 = new_n2837 & new_n2838;
  assign new_n2840 = ~shift6 & ~new_n2839;
  assign new_n2841 = new_n264 & ~new_n2171;
  assign new_n2842 = new_n309 & ~new_n2127;
  assign new_n2843 = new_n346 & ~new_n2187;
  assign new_n2844 = new_n383 & ~new_n2143;
  assign new_n2845 = ~new_n2841 & ~new_n2842;
  assign new_n2846 = ~new_n2843 & ~new_n2844;
  assign new_n2847 = new_n2845 & new_n2846;
  assign new_n2848 = shift6 & ~new_n2847;
  assign result45 = ~new_n2840 & ~new_n2848;
  assign new_n2850 = new_n264 & ~new_n2208;
  assign new_n2851 = new_n309 & ~new_n2236;
  assign new_n2852 = new_n346 & ~new_n2224;
  assign new_n2853 = new_n383 & ~new_n2252;
  assign new_n2854 = ~new_n2850 & ~new_n2851;
  assign new_n2855 = ~new_n2852 & ~new_n2853;
  assign new_n2856 = new_n2854 & new_n2855;
  assign new_n2857 = ~shift6 & ~new_n2856;
  assign new_n2858 = new_n264 & ~new_n2244;
  assign new_n2859 = new_n309 & ~new_n2200;
  assign new_n2860 = new_n346 & ~new_n2260;
  assign new_n2861 = new_n383 & ~new_n2216;
  assign new_n2862 = ~new_n2858 & ~new_n2859;
  assign new_n2863 = ~new_n2860 & ~new_n2861;
  assign new_n2864 = new_n2862 & new_n2863;
  assign new_n2865 = shift6 & ~new_n2864;
  assign result46 = ~new_n2857 & ~new_n2865;
  assign new_n2867 = new_n264 & ~new_n2281;
  assign new_n2868 = new_n309 & ~new_n2309;
  assign new_n2869 = new_n346 & ~new_n2297;
  assign new_n2870 = new_n383 & ~new_n2325;
  assign new_n2871 = ~new_n2867 & ~new_n2868;
  assign new_n2872 = ~new_n2869 & ~new_n2870;
  assign new_n2873 = new_n2871 & new_n2872;
  assign new_n2874 = ~shift6 & ~new_n2873;
  assign new_n2875 = new_n264 & ~new_n2317;
  assign new_n2876 = new_n309 & ~new_n2273;
  assign new_n2877 = new_n346 & ~new_n2333;
  assign new_n2878 = new_n383 & ~new_n2289;
  assign new_n2879 = ~new_n2875 & ~new_n2876;
  assign new_n2880 = ~new_n2877 & ~new_n2878;
  assign new_n2881 = new_n2879 & new_n2880;
  assign new_n2882 = shift6 & ~new_n2881;
  assign result47 = ~new_n2874 & ~new_n2882;
  assign new_n2884 = new_n264 & ~new_n530;
  assign new_n2885 = new_n309 & ~new_n566;
  assign new_n2886 = ~new_n344 & new_n346;
  assign new_n2887 = new_n383 & ~new_n458;
  assign new_n2888 = ~new_n2884 & ~new_n2885;
  assign new_n2889 = ~new_n2886 & ~new_n2887;
  assign new_n2890 = new_n2888 & new_n2889;
  assign new_n2891 = ~shift6 & ~new_n2890;
  assign new_n2892 = new_n264 & ~new_n381;
  assign new_n2893 = new_n309 & ~new_n418;
  assign new_n2894 = new_n346 & ~new_n494;
  assign new_n2895 = ~new_n307 & new_n383;
  assign new_n2896 = ~new_n2892 & ~new_n2893;
  assign new_n2897 = ~new_n2894 & ~new_n2895;
  assign new_n2898 = new_n2896 & new_n2897;
  assign new_n2899 = shift6 & ~new_n2898;
  assign result48 = ~new_n2891 & ~new_n2899;
  assign new_n2901 = new_n264 & ~new_n827;
  assign new_n2902 = new_n309 & ~new_n863;
  assign new_n2903 = new_n346 & ~new_n643;
  assign new_n2904 = new_n383 & ~new_n755;
  assign new_n2905 = ~new_n2901 & ~new_n2902;
  assign new_n2906 = ~new_n2903 & ~new_n2904;
  assign new_n2907 = new_n2905 & new_n2906;
  assign new_n2908 = ~shift6 & ~new_n2907;
  assign new_n2909 = new_n264 & ~new_n679;
  assign new_n2910 = new_n309 & ~new_n715;
  assign new_n2911 = new_n346 & ~new_n791;
  assign new_n2912 = new_n383 & ~new_n607;
  assign new_n2913 = ~new_n2909 & ~new_n2910;
  assign new_n2914 = ~new_n2911 & ~new_n2912;
  assign new_n2915 = new_n2913 & new_n2914;
  assign new_n2916 = shift6 & ~new_n2915;
  assign result49 = ~new_n2908 & ~new_n2916;
  assign new_n2918 = new_n264 & ~new_n1124;
  assign new_n2919 = new_n309 & ~new_n1160;
  assign new_n2920 = new_n346 & ~new_n940;
  assign new_n2921 = new_n383 & ~new_n1052;
  assign new_n2922 = ~new_n2918 & ~new_n2919;
  assign new_n2923 = ~new_n2920 & ~new_n2921;
  assign new_n2924 = new_n2922 & new_n2923;
  assign new_n2925 = ~shift6 & ~new_n2924;
  assign new_n2926 = new_n264 & ~new_n976;
  assign new_n2927 = new_n309 & ~new_n1012;
  assign new_n2928 = new_n346 & ~new_n1088;
  assign new_n2929 = new_n383 & ~new_n904;
  assign new_n2930 = ~new_n2926 & ~new_n2927;
  assign new_n2931 = ~new_n2928 & ~new_n2929;
  assign new_n2932 = new_n2930 & new_n2931;
  assign new_n2933 = shift6 & ~new_n2932;
  assign result50 = ~new_n2925 & ~new_n2933;
  assign new_n2935 = new_n264 & ~new_n1421;
  assign new_n2936 = new_n309 & ~new_n1457;
  assign new_n2937 = new_n346 & ~new_n1237;
  assign new_n2938 = new_n383 & ~new_n1349;
  assign new_n2939 = ~new_n2935 & ~new_n2936;
  assign new_n2940 = ~new_n2937 & ~new_n2938;
  assign new_n2941 = new_n2939 & new_n2940;
  assign new_n2942 = ~shift6 & ~new_n2941;
  assign new_n2943 = new_n264 & ~new_n1273;
  assign new_n2944 = new_n309 & ~new_n1309;
  assign new_n2945 = new_n346 & ~new_n1385;
  assign new_n2946 = new_n383 & ~new_n1201;
  assign new_n2947 = ~new_n2943 & ~new_n2944;
  assign new_n2948 = ~new_n2945 & ~new_n2946;
  assign new_n2949 = new_n2947 & new_n2948;
  assign new_n2950 = shift6 & ~new_n2949;
  assign result51 = ~new_n2942 & ~new_n2950;
  assign new_n2952 = new_n264 & ~new_n1522;
  assign new_n2953 = new_n309 & ~new_n1530;
  assign new_n2954 = new_n346 & ~new_n1478;
  assign new_n2955 = new_n383 & ~new_n1506;
  assign new_n2956 = ~new_n2952 & ~new_n2953;
  assign new_n2957 = ~new_n2954 & ~new_n2955;
  assign new_n2958 = new_n2956 & new_n2957;
  assign new_n2959 = ~shift6 & ~new_n2958;
  assign new_n2960 = new_n264 & ~new_n1486;
  assign new_n2961 = new_n309 & ~new_n1494;
  assign new_n2962 = new_n346 & ~new_n1514;
  assign new_n2963 = new_n383 & ~new_n1470;
  assign new_n2964 = ~new_n2960 & ~new_n2961;
  assign new_n2965 = ~new_n2962 & ~new_n2963;
  assign new_n2966 = new_n2964 & new_n2965;
  assign new_n2967 = shift6 & ~new_n2966;
  assign result52 = ~new_n2959 & ~new_n2967;
  assign new_n2969 = new_n264 & ~new_n1595;
  assign new_n2970 = new_n309 & ~new_n1603;
  assign new_n2971 = new_n346 & ~new_n1551;
  assign new_n2972 = new_n383 & ~new_n1579;
  assign new_n2973 = ~new_n2969 & ~new_n2970;
  assign new_n2974 = ~new_n2971 & ~new_n2972;
  assign new_n2975 = new_n2973 & new_n2974;
  assign new_n2976 = ~shift6 & ~new_n2975;
  assign new_n2977 = new_n264 & ~new_n1559;
  assign new_n2978 = new_n309 & ~new_n1567;
  assign new_n2979 = new_n346 & ~new_n1587;
  assign new_n2980 = new_n383 & ~new_n1543;
  assign new_n2981 = ~new_n2977 & ~new_n2978;
  assign new_n2982 = ~new_n2979 & ~new_n2980;
  assign new_n2983 = new_n2981 & new_n2982;
  assign new_n2984 = shift6 & ~new_n2983;
  assign result53 = ~new_n2976 & ~new_n2984;
  assign new_n2986 = new_n264 & ~new_n1668;
  assign new_n2987 = new_n309 & ~new_n1676;
  assign new_n2988 = new_n346 & ~new_n1624;
  assign new_n2989 = new_n383 & ~new_n1652;
  assign new_n2990 = ~new_n2986 & ~new_n2987;
  assign new_n2991 = ~new_n2988 & ~new_n2989;
  assign new_n2992 = new_n2990 & new_n2991;
  assign new_n2993 = ~shift6 & ~new_n2992;
  assign new_n2994 = new_n264 & ~new_n1632;
  assign new_n2995 = new_n309 & ~new_n1640;
  assign new_n2996 = new_n346 & ~new_n1660;
  assign new_n2997 = new_n383 & ~new_n1616;
  assign new_n2998 = ~new_n2994 & ~new_n2995;
  assign new_n2999 = ~new_n2996 & ~new_n2997;
  assign new_n3000 = new_n2998 & new_n2999;
  assign new_n3001 = shift6 & ~new_n3000;
  assign result54 = ~new_n2993 & ~new_n3001;
  assign new_n3003 = new_n264 & ~new_n1741;
  assign new_n3004 = new_n309 & ~new_n1749;
  assign new_n3005 = new_n346 & ~new_n1697;
  assign new_n3006 = new_n383 & ~new_n1725;
  assign new_n3007 = ~new_n3003 & ~new_n3004;
  assign new_n3008 = ~new_n3005 & ~new_n3006;
  assign new_n3009 = new_n3007 & new_n3008;
  assign new_n3010 = ~shift6 & ~new_n3009;
  assign new_n3011 = new_n264 & ~new_n1705;
  assign new_n3012 = new_n309 & ~new_n1713;
  assign new_n3013 = new_n346 & ~new_n1733;
  assign new_n3014 = new_n383 & ~new_n1689;
  assign new_n3015 = ~new_n3011 & ~new_n3012;
  assign new_n3016 = ~new_n3013 & ~new_n3014;
  assign new_n3017 = new_n3015 & new_n3016;
  assign new_n3018 = shift6 & ~new_n3017;
  assign result55 = ~new_n3010 & ~new_n3018;
  assign new_n3020 = new_n264 & ~new_n1814;
  assign new_n3021 = new_n309 & ~new_n1822;
  assign new_n3022 = new_n346 & ~new_n1770;
  assign new_n3023 = new_n383 & ~new_n1798;
  assign new_n3024 = ~new_n3020 & ~new_n3021;
  assign new_n3025 = ~new_n3022 & ~new_n3023;
  assign new_n3026 = new_n3024 & new_n3025;
  assign new_n3027 = ~shift6 & ~new_n3026;
  assign new_n3028 = new_n264 & ~new_n1778;
  assign new_n3029 = new_n309 & ~new_n1786;
  assign new_n3030 = new_n346 & ~new_n1806;
  assign new_n3031 = new_n383 & ~new_n1762;
  assign new_n3032 = ~new_n3028 & ~new_n3029;
  assign new_n3033 = ~new_n3030 & ~new_n3031;
  assign new_n3034 = new_n3032 & new_n3033;
  assign new_n3035 = shift6 & ~new_n3034;
  assign result56 = ~new_n3027 & ~new_n3035;
  assign new_n3037 = new_n264 & ~new_n1887;
  assign new_n3038 = new_n309 & ~new_n1895;
  assign new_n3039 = new_n346 & ~new_n1843;
  assign new_n3040 = new_n383 & ~new_n1871;
  assign new_n3041 = ~new_n3037 & ~new_n3038;
  assign new_n3042 = ~new_n3039 & ~new_n3040;
  assign new_n3043 = new_n3041 & new_n3042;
  assign new_n3044 = ~shift6 & ~new_n3043;
  assign new_n3045 = new_n264 & ~new_n1851;
  assign new_n3046 = new_n309 & ~new_n1859;
  assign new_n3047 = new_n346 & ~new_n1879;
  assign new_n3048 = new_n383 & ~new_n1835;
  assign new_n3049 = ~new_n3045 & ~new_n3046;
  assign new_n3050 = ~new_n3047 & ~new_n3048;
  assign new_n3051 = new_n3049 & new_n3050;
  assign new_n3052 = shift6 & ~new_n3051;
  assign result57 = ~new_n3044 & ~new_n3052;
  assign new_n3054 = new_n264 & ~new_n1960;
  assign new_n3055 = new_n309 & ~new_n1968;
  assign new_n3056 = new_n346 & ~new_n1916;
  assign new_n3057 = new_n383 & ~new_n1944;
  assign new_n3058 = ~new_n3054 & ~new_n3055;
  assign new_n3059 = ~new_n3056 & ~new_n3057;
  assign new_n3060 = new_n3058 & new_n3059;
  assign new_n3061 = ~shift6 & ~new_n3060;
  assign new_n3062 = new_n264 & ~new_n1924;
  assign new_n3063 = new_n309 & ~new_n1932;
  assign new_n3064 = new_n346 & ~new_n1952;
  assign new_n3065 = new_n383 & ~new_n1908;
  assign new_n3066 = ~new_n3062 & ~new_n3063;
  assign new_n3067 = ~new_n3064 & ~new_n3065;
  assign new_n3068 = new_n3066 & new_n3067;
  assign new_n3069 = shift6 & ~new_n3068;
  assign result58 = ~new_n3061 & ~new_n3069;
  assign new_n3071 = new_n264 & ~new_n2033;
  assign new_n3072 = new_n309 & ~new_n2041;
  assign new_n3073 = new_n346 & ~new_n1989;
  assign new_n3074 = new_n383 & ~new_n2017;
  assign new_n3075 = ~new_n3071 & ~new_n3072;
  assign new_n3076 = ~new_n3073 & ~new_n3074;
  assign new_n3077 = new_n3075 & new_n3076;
  assign new_n3078 = ~shift6 & ~new_n3077;
  assign new_n3079 = new_n264 & ~new_n1997;
  assign new_n3080 = new_n309 & ~new_n2005;
  assign new_n3081 = new_n346 & ~new_n2025;
  assign new_n3082 = new_n383 & ~new_n1981;
  assign new_n3083 = ~new_n3079 & ~new_n3080;
  assign new_n3084 = ~new_n3081 & ~new_n3082;
  assign new_n3085 = new_n3083 & new_n3084;
  assign new_n3086 = shift6 & ~new_n3085;
  assign result59 = ~new_n3078 & ~new_n3086;
  assign new_n3088 = new_n264 & ~new_n2106;
  assign new_n3089 = new_n309 & ~new_n2114;
  assign new_n3090 = new_n346 & ~new_n2062;
  assign new_n3091 = new_n383 & ~new_n2090;
  assign new_n3092 = ~new_n3088 & ~new_n3089;
  assign new_n3093 = ~new_n3090 & ~new_n3091;
  assign new_n3094 = new_n3092 & new_n3093;
  assign new_n3095 = ~shift6 & ~new_n3094;
  assign new_n3096 = new_n264 & ~new_n2070;
  assign new_n3097 = new_n309 & ~new_n2078;
  assign new_n3098 = new_n346 & ~new_n2098;
  assign new_n3099 = new_n383 & ~new_n2054;
  assign new_n3100 = ~new_n3096 & ~new_n3097;
  assign new_n3101 = ~new_n3098 & ~new_n3099;
  assign new_n3102 = new_n3100 & new_n3101;
  assign new_n3103 = shift6 & ~new_n3102;
  assign result60 = ~new_n3095 & ~new_n3103;
  assign new_n3105 = new_n264 & ~new_n2179;
  assign new_n3106 = new_n309 & ~new_n2187;
  assign new_n3107 = new_n346 & ~new_n2135;
  assign new_n3108 = new_n383 & ~new_n2163;
  assign new_n3109 = ~new_n3105 & ~new_n3106;
  assign new_n3110 = ~new_n3107 & ~new_n3108;
  assign new_n3111 = new_n3109 & new_n3110;
  assign new_n3112 = ~shift6 & ~new_n3111;
  assign new_n3113 = new_n264 & ~new_n2143;
  assign new_n3114 = new_n309 & ~new_n2151;
  assign new_n3115 = new_n346 & ~new_n2171;
  assign new_n3116 = new_n383 & ~new_n2127;
  assign new_n3117 = ~new_n3113 & ~new_n3114;
  assign new_n3118 = ~new_n3115 & ~new_n3116;
  assign new_n3119 = new_n3117 & new_n3118;
  assign new_n3120 = shift6 & ~new_n3119;
  assign result61 = ~new_n3112 & ~new_n3120;
  assign new_n3122 = new_n264 & ~new_n2252;
  assign new_n3123 = new_n309 & ~new_n2260;
  assign new_n3124 = new_n346 & ~new_n2208;
  assign new_n3125 = new_n383 & ~new_n2236;
  assign new_n3126 = ~new_n3122 & ~new_n3123;
  assign new_n3127 = ~new_n3124 & ~new_n3125;
  assign new_n3128 = new_n3126 & new_n3127;
  assign new_n3129 = ~shift6 & ~new_n3128;
  assign new_n3130 = new_n264 & ~new_n2216;
  assign new_n3131 = new_n309 & ~new_n2224;
  assign new_n3132 = new_n346 & ~new_n2244;
  assign new_n3133 = new_n383 & ~new_n2200;
  assign new_n3134 = ~new_n3130 & ~new_n3131;
  assign new_n3135 = ~new_n3132 & ~new_n3133;
  assign new_n3136 = new_n3134 & new_n3135;
  assign new_n3137 = shift6 & ~new_n3136;
  assign result62 = ~new_n3129 & ~new_n3137;
  assign new_n3139 = new_n264 & ~new_n2325;
  assign new_n3140 = new_n309 & ~new_n2333;
  assign new_n3141 = new_n346 & ~new_n2281;
  assign new_n3142 = new_n383 & ~new_n2309;
  assign new_n3143 = ~new_n3139 & ~new_n3140;
  assign new_n3144 = ~new_n3141 & ~new_n3142;
  assign new_n3145 = new_n3143 & new_n3144;
  assign new_n3146 = ~shift6 & ~new_n3145;
  assign new_n3147 = new_n264 & ~new_n2289;
  assign new_n3148 = new_n309 & ~new_n2297;
  assign new_n3149 = new_n346 & ~new_n2317;
  assign new_n3150 = new_n383 & ~new_n2273;
  assign new_n3151 = ~new_n3147 & ~new_n3148;
  assign new_n3152 = ~new_n3149 & ~new_n3150;
  assign new_n3153 = new_n3151 & new_n3152;
  assign new_n3154 = shift6 & ~new_n3153;
  assign result63 = ~new_n3146 & ~new_n3154;
  assign new_n3156 = shift6 & ~new_n422;
  assign new_n3157 = ~shift6 & ~new_n570;
  assign result64 = ~new_n3156 & ~new_n3157;
  assign new_n3159 = shift6 & ~new_n719;
  assign new_n3160 = ~shift6 & ~new_n867;
  assign result65 = ~new_n3159 & ~new_n3160;
  assign new_n3162 = shift6 & ~new_n1016;
  assign new_n3163 = ~shift6 & ~new_n1164;
  assign result66 = ~new_n3162 & ~new_n3163;
  assign new_n3165 = shift6 & ~new_n1313;
  assign new_n3166 = ~shift6 & ~new_n1461;
  assign result67 = ~new_n3165 & ~new_n3166;
  assign new_n3168 = shift6 & ~new_n1498;
  assign new_n3169 = ~shift6 & ~new_n1534;
  assign result68 = ~new_n3168 & ~new_n3169;
  assign new_n3171 = shift6 & ~new_n1571;
  assign new_n3172 = ~shift6 & ~new_n1607;
  assign result69 = ~new_n3171 & ~new_n3172;
  assign new_n3174 = shift6 & ~new_n1644;
  assign new_n3175 = ~shift6 & ~new_n1680;
  assign result70 = ~new_n3174 & ~new_n3175;
  assign new_n3177 = shift6 & ~new_n1717;
  assign new_n3178 = ~shift6 & ~new_n1753;
  assign result71 = ~new_n3177 & ~new_n3178;
  assign new_n3180 = shift6 & ~new_n1790;
  assign new_n3181 = ~shift6 & ~new_n1826;
  assign result72 = ~new_n3180 & ~new_n3181;
  assign new_n3183 = shift6 & ~new_n1863;
  assign new_n3184 = ~shift6 & ~new_n1899;
  assign result73 = ~new_n3183 & ~new_n3184;
  assign new_n3186 = shift6 & ~new_n1936;
  assign new_n3187 = ~shift6 & ~new_n1972;
  assign result74 = ~new_n3186 & ~new_n3187;
  assign new_n3189 = shift6 & ~new_n2009;
  assign new_n3190 = ~shift6 & ~new_n2045;
  assign result75 = ~new_n3189 & ~new_n3190;
  assign new_n3192 = shift6 & ~new_n2082;
  assign new_n3193 = ~shift6 & ~new_n2118;
  assign result76 = ~new_n3192 & ~new_n3193;
  assign new_n3195 = shift6 & ~new_n2155;
  assign new_n3196 = ~shift6 & ~new_n2191;
  assign result77 = ~new_n3195 & ~new_n3196;
  assign new_n3198 = shift6 & ~new_n2228;
  assign new_n3199 = ~shift6 & ~new_n2264;
  assign result78 = ~new_n3198 & ~new_n3199;
  assign new_n3201 = shift6 & ~new_n2301;
  assign new_n3202 = ~shift6 & ~new_n2337;
  assign result79 = ~new_n3201 & ~new_n3202;
  assign new_n3204 = shift6 & ~new_n2346;
  assign new_n3205 = ~shift6 & ~new_n2354;
  assign result80 = ~new_n3204 & ~new_n3205;
  assign new_n3207 = shift6 & ~new_n2363;
  assign new_n3208 = ~shift6 & ~new_n2371;
  assign result81 = ~new_n3207 & ~new_n3208;
  assign new_n3210 = shift6 & ~new_n2380;
  assign new_n3211 = ~shift6 & ~new_n2388;
  assign result82 = ~new_n3210 & ~new_n3211;
  assign new_n3213 = shift6 & ~new_n2397;
  assign new_n3214 = ~shift6 & ~new_n2405;
  assign result83 = ~new_n3213 & ~new_n3214;
  assign new_n3216 = shift6 & ~new_n2414;
  assign new_n3217 = ~shift6 & ~new_n2422;
  assign result84 = ~new_n3216 & ~new_n3217;
  assign new_n3219 = shift6 & ~new_n2431;
  assign new_n3220 = ~shift6 & ~new_n2439;
  assign result85 = ~new_n3219 & ~new_n3220;
  assign new_n3222 = shift6 & ~new_n2448;
  assign new_n3223 = ~shift6 & ~new_n2456;
  assign result86 = ~new_n3222 & ~new_n3223;
  assign new_n3225 = shift6 & ~new_n2465;
  assign new_n3226 = ~shift6 & ~new_n2473;
  assign result87 = ~new_n3225 & ~new_n3226;
  assign new_n3228 = shift6 & ~new_n2482;
  assign new_n3229 = ~shift6 & ~new_n2490;
  assign result88 = ~new_n3228 & ~new_n3229;
  assign new_n3231 = shift6 & ~new_n2499;
  assign new_n3232 = ~shift6 & ~new_n2507;
  assign result89 = ~new_n3231 & ~new_n3232;
  assign new_n3234 = shift6 & ~new_n2516;
  assign new_n3235 = ~shift6 & ~new_n2524;
  assign result90 = ~new_n3234 & ~new_n3235;
  assign new_n3237 = shift6 & ~new_n2533;
  assign new_n3238 = ~shift6 & ~new_n2541;
  assign result91 = ~new_n3237 & ~new_n3238;
  assign new_n3240 = shift6 & ~new_n2550;
  assign new_n3241 = ~shift6 & ~new_n2558;
  assign result92 = ~new_n3240 & ~new_n3241;
  assign new_n3243 = shift6 & ~new_n2567;
  assign new_n3244 = ~shift6 & ~new_n2575;
  assign result93 = ~new_n3243 & ~new_n3244;
  assign new_n3246 = shift6 & ~new_n2584;
  assign new_n3247 = ~shift6 & ~new_n2592;
  assign result94 = ~new_n3246 & ~new_n3247;
  assign new_n3249 = shift6 & ~new_n2601;
  assign new_n3250 = ~shift6 & ~new_n2609;
  assign result95 = ~new_n3249 & ~new_n3250;
  assign new_n3252 = shift6 & ~new_n2618;
  assign new_n3253 = ~shift6 & ~new_n2626;
  assign result96 = ~new_n3252 & ~new_n3253;
  assign new_n3255 = shift6 & ~new_n2635;
  assign new_n3256 = ~shift6 & ~new_n2643;
  assign result97 = ~new_n3255 & ~new_n3256;
  assign new_n3258 = shift6 & ~new_n2652;
  assign new_n3259 = ~shift6 & ~new_n2660;
  assign result98 = ~new_n3258 & ~new_n3259;
  assign new_n3261 = shift6 & ~new_n2669;
  assign new_n3262 = ~shift6 & ~new_n2677;
  assign result99 = ~new_n3261 & ~new_n3262;
  assign new_n3264 = shift6 & ~new_n2686;
  assign new_n3265 = ~shift6 & ~new_n2694;
  assign result100 = ~new_n3264 & ~new_n3265;
  assign new_n3267 = shift6 & ~new_n2703;
  assign new_n3268 = ~shift6 & ~new_n2711;
  assign result101 = ~new_n3267 & ~new_n3268;
  assign new_n3270 = shift6 & ~new_n2720;
  assign new_n3271 = ~shift6 & ~new_n2728;
  assign result102 = ~new_n3270 & ~new_n3271;
  assign new_n3273 = shift6 & ~new_n2737;
  assign new_n3274 = ~shift6 & ~new_n2745;
  assign result103 = ~new_n3273 & ~new_n3274;
  assign new_n3276 = shift6 & ~new_n2754;
  assign new_n3277 = ~shift6 & ~new_n2762;
  assign result104 = ~new_n3276 & ~new_n3277;
  assign new_n3279 = shift6 & ~new_n2771;
  assign new_n3280 = ~shift6 & ~new_n2779;
  assign result105 = ~new_n3279 & ~new_n3280;
  assign new_n3282 = shift6 & ~new_n2788;
  assign new_n3283 = ~shift6 & ~new_n2796;
  assign result106 = ~new_n3282 & ~new_n3283;
  assign new_n3285 = shift6 & ~new_n2805;
  assign new_n3286 = ~shift6 & ~new_n2813;
  assign result107 = ~new_n3285 & ~new_n3286;
  assign new_n3288 = shift6 & ~new_n2822;
  assign new_n3289 = ~shift6 & ~new_n2830;
  assign result108 = ~new_n3288 & ~new_n3289;
  assign new_n3291 = shift6 & ~new_n2839;
  assign new_n3292 = ~shift6 & ~new_n2847;
  assign result109 = ~new_n3291 & ~new_n3292;
  assign new_n3294 = shift6 & ~new_n2856;
  assign new_n3295 = ~shift6 & ~new_n2864;
  assign result110 = ~new_n3294 & ~new_n3295;
  assign new_n3297 = shift6 & ~new_n2873;
  assign new_n3298 = ~shift6 & ~new_n2881;
  assign result111 = ~new_n3297 & ~new_n3298;
  assign new_n3300 = shift6 & ~new_n2890;
  assign new_n3301 = ~shift6 & ~new_n2898;
  assign result112 = ~new_n3300 & ~new_n3301;
  assign new_n3303 = shift6 & ~new_n2907;
  assign new_n3304 = ~shift6 & ~new_n2915;
  assign result113 = ~new_n3303 & ~new_n3304;
  assign new_n3306 = shift6 & ~new_n2924;
  assign new_n3307 = ~shift6 & ~new_n2932;
  assign result114 = ~new_n3306 & ~new_n3307;
  assign new_n3309 = shift6 & ~new_n2941;
  assign new_n3310 = ~shift6 & ~new_n2949;
  assign result115 = ~new_n3309 & ~new_n3310;
  assign new_n3312 = shift6 & ~new_n2958;
  assign new_n3313 = ~shift6 & ~new_n2966;
  assign result116 = ~new_n3312 & ~new_n3313;
  assign new_n3315 = shift6 & ~new_n2975;
  assign new_n3316 = ~shift6 & ~new_n2983;
  assign result117 = ~new_n3315 & ~new_n3316;
  assign new_n3318 = shift6 & ~new_n2992;
  assign new_n3319 = ~shift6 & ~new_n3000;
  assign result118 = ~new_n3318 & ~new_n3319;
  assign new_n3321 = shift6 & ~new_n3009;
  assign new_n3322 = ~shift6 & ~new_n3017;
  assign result119 = ~new_n3321 & ~new_n3322;
  assign new_n3324 = shift6 & ~new_n3026;
  assign new_n3325 = ~shift6 & ~new_n3034;
  assign result120 = ~new_n3324 & ~new_n3325;
  assign new_n3327 = shift6 & ~new_n3043;
  assign new_n3328 = ~shift6 & ~new_n3051;
  assign result121 = ~new_n3327 & ~new_n3328;
  assign new_n3330 = shift6 & ~new_n3060;
  assign new_n3331 = ~shift6 & ~new_n3068;
  assign result122 = ~new_n3330 & ~new_n3331;
  assign new_n3333 = shift6 & ~new_n3077;
  assign new_n3334 = ~shift6 & ~new_n3085;
  assign result123 = ~new_n3333 & ~new_n3334;
  assign new_n3336 = shift6 & ~new_n3094;
  assign new_n3337 = ~shift6 & ~new_n3102;
  assign result124 = ~new_n3336 & ~new_n3337;
  assign new_n3339 = shift6 & ~new_n3111;
  assign new_n3340 = ~shift6 & ~new_n3119;
  assign result125 = ~new_n3339 & ~new_n3340;
  assign new_n3342 = shift6 & ~new_n3128;
  assign new_n3343 = ~shift6 & ~new_n3136;
  assign result126 = ~new_n3342 & ~new_n3343;
  assign new_n3345 = shift6 & ~new_n3145;
  assign new_n3346 = ~shift6 & ~new_n3153;
  assign result127 = ~new_n3345 & ~new_n3346;
endmodule


