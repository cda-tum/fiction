// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pina0, pinb1, pinc2, pind3, pina1, pinb0, pinc3, pind2, pmusel1, pinc4,
    pind5, pmusel2, pinc5, pind4, pmusel3, pina4, pinb5, pina5, pinb4,
    pina2, pinb3, pinc0, pind1, pina3, pinb2, pinc1, pind0, pind15, pinc15,
    pind14, pinb15, pinc14, pind13, popsel3, popsel1, popsel2, pina11,
    pinb10, pina10, popsel0, pina15, pinb14, pinc13, pind12, pina14,
    pinb13, pinc12, pind11, pina13, pinb12, pinc11, pind10, pina12, pinb11,
    pinc10, pina8, pinb9, pina9, pinb8, pina6, pinb7, pina7, pinb6, psh0,
    pinc6, pind7, pmusel4, psh1, pinc7, pind6, psh2, pinc8, pind9, pinc9,
    pind8,
    po12, po11, po14, po13, po15, po9, po8, po7, po6, po5, po4, po3, po2,
    po1, po0, po10  );
  input  pina0, pinb1, pinc2, pind3, pina1, pinb0, pinc3, pind2, pmusel1,
    pinc4, pind5, pmusel2, pinc5, pind4, pmusel3, pina4, pinb5, pina5,
    pinb4, pina2, pinb3, pinc0, pind1, pina3, pinb2, pinc1, pind0, pind15,
    pinc15, pind14, pinb15, pinc14, pind13, popsel3, popsel1, popsel2,
    pina11, pinb10, pina10, popsel0, pina15, pinb14, pinc13, pind12,
    pina14, pinb13, pinc12, pind11, pina13, pinb12, pinc11, pind10, pina12,
    pinb11, pinc10, pina8, pinb9, pina9, pinb8, pina6, pinb7, pina7, pinb6,
    psh0, pinc6, pind7, pmusel4, psh1, pinc7, pind6, psh2, pinc8, pind9,
    pinc9, pind8;
  output po12, po11, po14, po13, po15, po9, po8, po7, po6, po5, po4, po3, po2,
    po1, po0, po10;
  wire new_n92, new_n93, new_n94, new_n95, new_n96, new_n97, new_n98,
    new_n99, new_n100, new_n101, new_n102, new_n103, new_n104, new_n105,
    new_n106, new_n107, new_n108, new_n109, new_n110, new_n111, new_n112,
    new_n113, new_n114, new_n115, new_n116, new_n117, new_n118, new_n119,
    new_n120, new_n121, new_n122, new_n123, new_n124, new_n125, new_n126,
    new_n127, new_n128, new_n129, new_n130, new_n131, new_n132, new_n133,
    new_n134, new_n135, new_n136, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n162, new_n163, new_n164, new_n165, new_n166, new_n167, new_n168,
    new_n169, new_n170, new_n171, new_n172, new_n173, new_n174, new_n175,
    new_n176, new_n177, new_n178, new_n179, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n290, new_n291, new_n292, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n474, new_n475, new_n476,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1607, new_n1608, new_n1609, new_n1610, new_n1611, new_n1612,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1640, new_n1641, new_n1642,
    new_n1643, new_n1644, new_n1645, new_n1646, new_n1647, new_n1648,
    new_n1649, new_n1650, new_n1651, new_n1652, new_n1653, new_n1654,
    new_n1655, new_n1656, new_n1657, new_n1658, new_n1659, new_n1660,
    new_n1661, new_n1662, new_n1663, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825;
  assign new_n92 = pmusel2 & pinc0;
  assign new_n93 = ~pmusel1 & new_n92;
  assign new_n94 = pina0 & ~pmusel2;
  assign new_n95 = pmusel1 & new_n94;
  assign new_n96 = ~new_n93 & ~new_n95;
  assign new_n97 = ~pmusel3 & pmusel4;
  assign new_n98 = ~new_n96 & new_n97;
  assign new_n99 = pmusel2 & pinc15;
  assign new_n100 = ~pmusel1 & new_n99;
  assign new_n101 = ~pmusel2 & pina15;
  assign new_n102 = pmusel1 & new_n101;
  assign new_n103 = ~new_n100 & ~new_n102;
  assign new_n104 = new_n97 & ~new_n103;
  assign new_n105 = new_n98 & ~new_n104;
  assign new_n106 = ~new_n98 & new_n104;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = pinc2 & pmusel2;
  assign new_n109 = ~pmusel1 & new_n108;
  assign new_n110 = ~pmusel2 & pina2;
  assign new_n111 = pmusel1 & new_n110;
  assign new_n112 = ~new_n109 & ~new_n111;
  assign new_n113 = new_n97 & ~new_n112;
  assign new_n114 = ~new_n104 & new_n113;
  assign new_n115 = new_n104 & ~new_n113;
  assign new_n116 = ~new_n114 & ~new_n115;
  assign new_n117 = pmusel2 & pinc1;
  assign new_n118 = ~pmusel1 & new_n117;
  assign new_n119 = pina1 & ~pmusel2;
  assign new_n120 = pmusel1 & new_n119;
  assign new_n121 = ~new_n118 & ~new_n120;
  assign new_n122 = new_n97 & ~new_n121;
  assign new_n123 = ~new_n104 & new_n122;
  assign new_n124 = new_n104 & ~new_n122;
  assign new_n125 = ~new_n123 & ~new_n124;
  assign new_n126 = pinc3 & pmusel2;
  assign new_n127 = ~pmusel1 & new_n126;
  assign new_n128 = ~pmusel2 & pina3;
  assign new_n129 = pmusel1 & new_n128;
  assign new_n130 = ~new_n127 & ~new_n129;
  assign new_n131 = new_n97 & ~new_n130;
  assign new_n132 = ~new_n104 & new_n131;
  assign new_n133 = new_n104 & ~new_n131;
  assign new_n134 = ~new_n132 & ~new_n133;
  assign new_n135 = ~new_n107 & ~new_n116;
  assign new_n136 = ~new_n125 & ~new_n134;
  assign new_n137 = new_n135 & new_n136;
  assign new_n138 = pmusel2 & pinc8;
  assign new_n139 = ~pmusel1 & new_n138;
  assign new_n140 = ~pmusel2 & pina8;
  assign new_n141 = pmusel1 & new_n140;
  assign new_n142 = ~new_n139 & ~new_n141;
  assign new_n143 = new_n97 & ~new_n142;
  assign new_n144 = ~new_n104 & new_n143;
  assign new_n145 = new_n104 & ~new_n143;
  assign new_n146 = ~new_n144 & ~new_n145;
  assign new_n147 = pmusel2 & pinc10;
  assign new_n148 = ~pmusel1 & new_n147;
  assign new_n149 = ~pmusel2 & pina10;
  assign new_n150 = pmusel1 & new_n149;
  assign new_n151 = ~new_n148 & ~new_n150;
  assign new_n152 = new_n97 & ~new_n151;
  assign new_n153 = ~new_n104 & new_n152;
  assign new_n154 = new_n104 & ~new_n152;
  assign new_n155 = ~new_n153 & ~new_n154;
  assign new_n156 = pmusel2 & pinc9;
  assign new_n157 = ~pmusel1 & new_n156;
  assign new_n158 = ~pmusel2 & pina9;
  assign new_n159 = pmusel1 & new_n158;
  assign new_n160 = ~new_n157 & ~new_n159;
  assign new_n161 = new_n97 & ~new_n160;
  assign new_n162 = ~new_n104 & new_n161;
  assign new_n163 = new_n104 & ~new_n161;
  assign new_n164 = ~new_n162 & ~new_n163;
  assign new_n165 = pmusel2 & pinc11;
  assign new_n166 = ~pmusel1 & new_n165;
  assign new_n167 = ~pmusel2 & pina11;
  assign new_n168 = pmusel1 & new_n167;
  assign new_n169 = ~new_n166 & ~new_n168;
  assign new_n170 = new_n97 & ~new_n169;
  assign new_n171 = ~new_n104 & new_n170;
  assign new_n172 = new_n104 & ~new_n170;
  assign new_n173 = ~new_n171 & ~new_n172;
  assign new_n174 = ~new_n146 & ~new_n155;
  assign new_n175 = ~new_n164 & ~new_n173;
  assign new_n176 = new_n174 & new_n175;
  assign new_n177 = pinc4 & pmusel2;
  assign new_n178 = ~pmusel1 & new_n177;
  assign new_n179 = ~pmusel2 & pina4;
  assign new_n180 = pmusel1 & new_n179;
  assign new_n181 = ~new_n178 & ~new_n180;
  assign new_n182 = new_n97 & ~new_n181;
  assign new_n183 = ~new_n104 & new_n182;
  assign new_n184 = new_n104 & ~new_n182;
  assign new_n185 = ~new_n183 & ~new_n184;
  assign new_n186 = pmusel2 & pinc6;
  assign new_n187 = ~pmusel1 & new_n186;
  assign new_n188 = ~pmusel2 & pina6;
  assign new_n189 = pmusel1 & new_n188;
  assign new_n190 = ~new_n187 & ~new_n189;
  assign new_n191 = new_n97 & ~new_n190;
  assign new_n192 = ~new_n104 & new_n191;
  assign new_n193 = new_n104 & ~new_n191;
  assign new_n194 = ~new_n192 & ~new_n193;
  assign new_n195 = pmusel2 & pinc5;
  assign new_n196 = ~pmusel1 & new_n195;
  assign new_n197 = ~pmusel2 & pina5;
  assign new_n198 = pmusel1 & new_n197;
  assign new_n199 = ~new_n196 & ~new_n198;
  assign new_n200 = new_n97 & ~new_n199;
  assign new_n201 = ~new_n104 & new_n200;
  assign new_n202 = new_n104 & ~new_n200;
  assign new_n203 = ~new_n201 & ~new_n202;
  assign new_n204 = pmusel2 & pinc7;
  assign new_n205 = ~pmusel1 & new_n204;
  assign new_n206 = ~pmusel2 & pina7;
  assign new_n207 = pmusel1 & new_n206;
  assign new_n208 = ~new_n205 & ~new_n207;
  assign new_n209 = new_n97 & ~new_n208;
  assign new_n210 = ~new_n104 & new_n209;
  assign new_n211 = new_n104 & ~new_n209;
  assign new_n212 = ~new_n210 & ~new_n211;
  assign new_n213 = ~new_n185 & ~new_n194;
  assign new_n214 = ~new_n203 & ~new_n212;
  assign new_n215 = new_n213 & new_n214;
  assign new_n216 = new_n137 & new_n176;
  assign new_n217 = new_n104 & new_n216;
  assign new_n218 = new_n215 & new_n217;
  assign new_n219 = pmusel2 & pinc12;
  assign new_n220 = ~pmusel1 & new_n219;
  assign new_n221 = ~pmusel2 & pina12;
  assign new_n222 = pmusel1 & new_n221;
  assign new_n223 = ~new_n220 & ~new_n222;
  assign new_n224 = new_n97 & ~new_n223;
  assign new_n225 = ~new_n104 & new_n224;
  assign new_n226 = new_n104 & ~new_n224;
  assign new_n227 = ~new_n225 & ~new_n226;
  assign new_n228 = new_n218 & new_n227;
  assign new_n229 = ~new_n218 & ~new_n227;
  assign new_n230 = ~new_n228 & ~new_n229;
  assign new_n231 = popsel2 & ~new_n230;
  assign new_n232 = ~popsel1 & ~popsel0;
  assign new_n233 = new_n231 & new_n232;
  assign new_n234 = ~popsel2 & new_n230;
  assign new_n235 = psh0 & psh1;
  assign new_n236 = pmusel3 & ~pmusel4;
  assign new_n237 = pmusel2 & pind15;
  assign new_n238 = ~pinb15 & ~new_n237;
  assign new_n239 = pmusel1 & ~pmusel2;
  assign new_n240 = ~pmusel1 & pmusel2;
  assign new_n241 = ~new_n239 & ~new_n240;
  assign new_n242 = ~new_n237 & new_n241;
  assign new_n243 = ~pmusel1 & ~pinb15;
  assign new_n244 = ~pmusel1 & new_n241;
  assign new_n245 = ~new_n238 & ~new_n242;
  assign new_n246 = ~new_n243 & ~new_n244;
  assign new_n247 = new_n245 & new_n246;
  assign new_n248 = new_n236 & new_n247;
  assign new_n249 = ~pmusel1 & ~pmusel2;
  assign new_n250 = pind15 & new_n249;
  assign new_n251 = new_n97 & new_n250;
  assign new_n252 = ~new_n248 & ~new_n251;
  assign new_n253 = new_n235 & ~new_n252;
  assign new_n254 = psh0 & ~psh1;
  assign new_n255 = pmusel2 & pind13;
  assign new_n256 = ~pinb13 & ~new_n255;
  assign new_n257 = new_n241 & ~new_n255;
  assign new_n258 = ~pmusel1 & ~pinb13;
  assign new_n259 = ~new_n256 & ~new_n257;
  assign new_n260 = ~new_n244 & ~new_n258;
  assign new_n261 = new_n259 & new_n260;
  assign new_n262 = new_n236 & new_n261;
  assign new_n263 = ~pmusel3 & pind13;
  assign new_n264 = pmusel4 & new_n249;
  assign new_n265 = new_n263 & new_n264;
  assign new_n266 = ~new_n262 & ~new_n265;
  assign new_n267 = new_n254 & ~new_n266;
  assign new_n268 = ~new_n253 & ~new_n267;
  assign new_n269 = pmusel2 & pind14;
  assign new_n270 = ~pinb14 & ~new_n269;
  assign new_n271 = new_n241 & ~new_n269;
  assign new_n272 = ~pmusel1 & ~pinb14;
  assign new_n273 = ~new_n270 & ~new_n271;
  assign new_n274 = ~new_n244 & ~new_n272;
  assign new_n275 = new_n273 & new_n274;
  assign new_n276 = new_n236 & new_n275;
  assign new_n277 = ~pmusel3 & pind14;
  assign new_n278 = new_n264 & new_n277;
  assign new_n279 = ~new_n276 & ~new_n278;
  assign new_n280 = psh1 & ~new_n279;
  assign new_n281 = pmusel2 & pind12;
  assign new_n282 = ~pinb12 & ~new_n281;
  assign new_n283 = new_n241 & ~new_n281;
  assign new_n284 = ~pmusel1 & ~pinb12;
  assign new_n285 = ~new_n282 & ~new_n283;
  assign new_n286 = ~new_n244 & ~new_n284;
  assign new_n287 = new_n285 & new_n286;
  assign new_n288 = new_n236 & new_n287;
  assign new_n289 = ~pmusel3 & pind12;
  assign new_n290 = new_n264 & new_n289;
  assign new_n291 = ~new_n288 & ~new_n290;
  assign new_n292 = ~psh1 & ~new_n291;
  assign new_n293 = ~new_n280 & ~new_n292;
  assign new_n294 = new_n268 & new_n293;
  assign new_n295 = psh0 & new_n268;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = ~psh2 & new_n296;
  assign new_n298 = ~new_n235 & new_n252;
  assign new_n299 = new_n235 & new_n291;
  assign new_n300 = new_n252 & new_n291;
  assign new_n301 = ~new_n299 & ~new_n300;
  assign new_n302 = ~new_n298 & new_n301;
  assign new_n303 = psh2 & new_n302;
  assign new_n304 = ~new_n297 & ~new_n303;
  assign new_n305 = new_n230 & new_n304;
  assign new_n306 = popsel2 & new_n304;
  assign new_n307 = ~new_n305 & ~new_n306;
  assign new_n308 = ~new_n234 & new_n307;
  assign new_n309 = ~new_n233 & ~new_n308;
  assign new_n310 = new_n232 & ~new_n233;
  assign new_n311 = ~new_n309 & ~new_n310;
  assign new_n312 = ~popsel3 & new_n311;
  assign new_n313 = popsel3 & ~popsel2;
  assign new_n314 = ~popsel1 & popsel0;
  assign new_n315 = popsel1 & ~popsel0;
  assign new_n316 = ~new_n314 & ~new_n315;
  assign new_n317 = ~new_n232 & new_n316;
  assign new_n318 = ~pmusel3 & pinb11;
  assign new_n319 = pmusel2 & new_n318;
  assign new_n320 = ~pmusel1 & new_n319;
  assign new_n321 = pmusel3 & pind11;
  assign new_n322 = ~pmusel2 & new_n321;
  assign new_n323 = ~pmusel1 & new_n322;
  assign new_n324 = ~new_n320 & ~new_n323;
  assign new_n325 = ~pina11 & ~pinc11;
  assign new_n326 = pmusel2 & ~pinc11;
  assign new_n327 = ~pmusel2 & ~pina11;
  assign new_n328 = ~new_n325 & ~new_n326;
  assign new_n329 = ~new_n327 & new_n328;
  assign new_n330 = pmusel1 & ~pmusel3;
  assign new_n331 = new_n329 & new_n330;
  assign new_n332 = new_n324 & ~new_n331;
  assign new_n333 = ~pmusel4 & ~new_n332;
  assign new_n334 = ~pmusel3 & pinb10;
  assign new_n335 = pmusel2 & new_n334;
  assign new_n336 = ~pmusel1 & new_n335;
  assign new_n337 = pmusel3 & pind10;
  assign new_n338 = ~pmusel2 & new_n337;
  assign new_n339 = ~pmusel1 & new_n338;
  assign new_n340 = ~new_n336 & ~new_n339;
  assign new_n341 = ~pina10 & ~pinc10;
  assign new_n342 = pmusel2 & ~pinc10;
  assign new_n343 = ~pmusel2 & ~pina10;
  assign new_n344 = ~new_n341 & ~new_n342;
  assign new_n345 = ~new_n343 & new_n344;
  assign new_n346 = new_n330 & new_n345;
  assign new_n347 = new_n340 & ~new_n346;
  assign new_n348 = ~pmusel4 & ~new_n347;
  assign new_n349 = popsel3 & popsel2;
  assign new_n350 = popsel1 & ~popsel2;
  assign new_n351 = ~popsel3 & ~popsel1;
  assign new_n352 = ~new_n350 & ~new_n351;
  assign new_n353 = ~popsel0 & ~new_n349;
  assign new_n354 = new_n352 & new_n353;
  assign new_n355 = ~pina10 & ~new_n147;
  assign new_n356 = ~new_n147 & new_n241;
  assign new_n357 = ~pmusel1 & ~pina10;
  assign new_n358 = ~new_n355 & ~new_n356;
  assign new_n359 = ~new_n244 & ~new_n357;
  assign new_n360 = new_n358 & new_n359;
  assign new_n361 = new_n236 & new_n360;
  assign new_n362 = pinc10 & pmusel4;
  assign new_n363 = ~pmusel1 & new_n362;
  assign new_n364 = ~pmusel2 & new_n363;
  assign new_n365 = ~pmusel3 & new_n364;
  assign new_n366 = ~new_n361 & ~new_n365;
  assign new_n367 = ~new_n354 & ~new_n366;
  assign new_n368 = new_n354 & new_n366;
  assign new_n369 = ~new_n367 & ~new_n368;
  assign new_n370 = new_n348 & ~new_n369;
  assign new_n371 = ~pmusel3 & pinb9;
  assign new_n372 = pmusel2 & new_n371;
  assign new_n373 = ~pmusel1 & new_n372;
  assign new_n374 = pmusel3 & pind9;
  assign new_n375 = ~pmusel2 & new_n374;
  assign new_n376 = ~pmusel1 & new_n375;
  assign new_n377 = ~new_n373 & ~new_n376;
  assign new_n378 = ~pina9 & ~pinc9;
  assign new_n379 = pmusel2 & ~pinc9;
  assign new_n380 = ~pmusel2 & ~pina9;
  assign new_n381 = ~new_n378 & ~new_n379;
  assign new_n382 = ~new_n380 & new_n381;
  assign new_n383 = new_n330 & new_n382;
  assign new_n384 = new_n377 & ~new_n383;
  assign new_n385 = ~pmusel4 & ~new_n384;
  assign new_n386 = ~pina9 & ~new_n156;
  assign new_n387 = ~new_n156 & new_n241;
  assign new_n388 = ~pmusel1 & ~pina9;
  assign new_n389 = ~new_n386 & ~new_n387;
  assign new_n390 = ~new_n244 & ~new_n388;
  assign new_n391 = new_n389 & new_n390;
  assign new_n392 = new_n236 & new_n391;
  assign new_n393 = pmusel4 & pinc9;
  assign new_n394 = ~pmusel1 & new_n393;
  assign new_n395 = ~pmusel2 & new_n394;
  assign new_n396 = ~pmusel3 & new_n395;
  assign new_n397 = ~new_n392 & ~new_n396;
  assign new_n398 = ~new_n354 & ~new_n397;
  assign new_n399 = new_n354 & new_n397;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = new_n385 & ~new_n400;
  assign new_n402 = ~pmusel3 & pinb8;
  assign new_n403 = pmusel2 & new_n402;
  assign new_n404 = ~pmusel1 & new_n403;
  assign new_n405 = pmusel3 & pind8;
  assign new_n406 = ~pmusel2 & new_n405;
  assign new_n407 = ~pmusel1 & new_n406;
  assign new_n408 = ~new_n404 & ~new_n407;
  assign new_n409 = ~pina8 & ~pinc8;
  assign new_n410 = pmusel2 & ~pinc8;
  assign new_n411 = ~pmusel2 & ~pina8;
  assign new_n412 = ~new_n409 & ~new_n410;
  assign new_n413 = ~new_n411 & new_n412;
  assign new_n414 = new_n330 & new_n413;
  assign new_n415 = new_n408 & ~new_n414;
  assign new_n416 = ~pmusel4 & ~new_n415;
  assign new_n417 = ~pina8 & ~new_n138;
  assign new_n418 = ~new_n138 & new_n241;
  assign new_n419 = ~pmusel1 & ~pina8;
  assign new_n420 = ~new_n417 & ~new_n418;
  assign new_n421 = ~new_n244 & ~new_n419;
  assign new_n422 = new_n420 & new_n421;
  assign new_n423 = new_n236 & new_n422;
  assign new_n424 = pmusel4 & pinc8;
  assign new_n425 = ~pmusel1 & new_n424;
  assign new_n426 = ~pmusel2 & new_n425;
  assign new_n427 = ~pmusel3 & new_n426;
  assign new_n428 = ~new_n423 & ~new_n427;
  assign new_n429 = ~new_n354 & ~new_n428;
  assign new_n430 = new_n354 & new_n428;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = new_n416 & ~new_n431;
  assign new_n433 = ~new_n400 & new_n432;
  assign new_n434 = new_n385 & new_n432;
  assign new_n435 = ~new_n433 & ~new_n434;
  assign new_n436 = ~new_n401 & new_n435;
  assign new_n437 = ~new_n348 & new_n369;
  assign new_n438 = ~new_n436 & ~new_n437;
  assign new_n439 = ~new_n370 & ~new_n438;
  assign new_n440 = ~new_n333 & new_n439;
  assign new_n441 = ~pina11 & ~new_n165;
  assign new_n442 = ~new_n165 & new_n241;
  assign new_n443 = ~pmusel1 & ~pina11;
  assign new_n444 = ~new_n441 & ~new_n442;
  assign new_n445 = ~new_n244 & ~new_n443;
  assign new_n446 = new_n444 & new_n445;
  assign new_n447 = new_n236 & new_n446;
  assign new_n448 = pinc11 & pmusel4;
  assign new_n449 = ~pmusel1 & new_n448;
  assign new_n450 = ~pmusel2 & new_n449;
  assign new_n451 = ~pmusel3 & new_n450;
  assign new_n452 = ~new_n447 & ~new_n451;
  assign new_n453 = ~new_n354 & ~new_n452;
  assign new_n454 = new_n354 & new_n452;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = new_n439 & new_n455;
  assign new_n457 = ~new_n333 & new_n455;
  assign new_n458 = ~new_n333 & new_n457;
  assign new_n459 = new_n455 & new_n457;
  assign new_n460 = ~new_n440 & ~new_n456;
  assign new_n461 = ~new_n458 & ~new_n459;
  assign new_n462 = new_n460 & new_n461;
  assign new_n463 = ~new_n369 & ~new_n455;
  assign new_n464 = new_n348 & ~new_n455;
  assign new_n465 = new_n333 & ~new_n369;
  assign new_n466 = new_n333 & new_n348;
  assign new_n467 = ~new_n463 & ~new_n464;
  assign new_n468 = ~new_n465 & ~new_n466;
  assign new_n469 = new_n467 & new_n468;
  assign new_n470 = ~new_n400 & ~new_n431;
  assign new_n471 = ~new_n400 & new_n416;
  assign new_n472 = new_n385 & ~new_n431;
  assign new_n473 = new_n385 & new_n416;
  assign new_n474 = ~new_n470 & ~new_n471;
  assign new_n475 = ~new_n472 & ~new_n473;
  assign new_n476 = new_n474 & new_n475;
  assign new_n477 = ~pina4 & ~new_n177;
  assign new_n478 = ~new_n177 & new_n241;
  assign new_n479 = ~pmusel1 & ~pina4;
  assign new_n480 = ~new_n477 & ~new_n478;
  assign new_n481 = ~new_n244 & ~new_n479;
  assign new_n482 = new_n480 & new_n481;
  assign new_n483 = new_n236 & new_n482;
  assign new_n484 = pinc4 & pmusel4;
  assign new_n485 = ~pmusel1 & new_n484;
  assign new_n486 = ~pmusel2 & new_n485;
  assign new_n487 = ~pmusel3 & new_n486;
  assign new_n488 = ~new_n483 & ~new_n487;
  assign new_n489 = ~new_n354 & ~new_n488;
  assign new_n490 = new_n354 & new_n488;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = ~pina5 & ~new_n195;
  assign new_n493 = ~new_n195 & new_n241;
  assign new_n494 = ~pmusel1 & ~pina5;
  assign new_n495 = ~new_n492 & ~new_n493;
  assign new_n496 = ~new_n244 & ~new_n494;
  assign new_n497 = new_n495 & new_n496;
  assign new_n498 = new_n236 & new_n497;
  assign new_n499 = pinc5 & pmusel4;
  assign new_n500 = ~pmusel1 & new_n499;
  assign new_n501 = ~pmusel2 & new_n500;
  assign new_n502 = ~pmusel3 & new_n501;
  assign new_n503 = ~new_n498 & ~new_n502;
  assign new_n504 = ~new_n354 & ~new_n503;
  assign new_n505 = new_n354 & new_n503;
  assign new_n506 = ~new_n504 & ~new_n505;
  assign new_n507 = ~new_n491 & ~new_n506;
  assign new_n508 = ~pmusel3 & pinb4;
  assign new_n509 = pmusel2 & new_n508;
  assign new_n510 = ~pmusel1 & new_n509;
  assign new_n511 = pind4 & pmusel3;
  assign new_n512 = ~pmusel2 & new_n511;
  assign new_n513 = ~pmusel1 & new_n512;
  assign new_n514 = ~new_n510 & ~new_n513;
  assign new_n515 = ~pinc4 & ~pina4;
  assign new_n516 = ~pinc4 & pmusel2;
  assign new_n517 = ~pmusel2 & ~pina4;
  assign new_n518 = ~new_n515 & ~new_n516;
  assign new_n519 = ~new_n517 & new_n518;
  assign new_n520 = new_n330 & new_n519;
  assign new_n521 = new_n514 & ~new_n520;
  assign new_n522 = ~pmusel4 & ~new_n521;
  assign new_n523 = ~new_n506 & new_n522;
  assign new_n524 = ~pmusel3 & pinb5;
  assign new_n525 = pmusel2 & new_n524;
  assign new_n526 = ~pmusel1 & new_n525;
  assign new_n527 = pind5 & pmusel3;
  assign new_n528 = ~pmusel2 & new_n527;
  assign new_n529 = ~pmusel1 & new_n528;
  assign new_n530 = ~new_n526 & ~new_n529;
  assign new_n531 = ~pinc5 & ~pina5;
  assign new_n532 = pmusel2 & ~pinc5;
  assign new_n533 = ~pmusel2 & ~pina5;
  assign new_n534 = ~new_n531 & ~new_n532;
  assign new_n535 = ~new_n533 & new_n534;
  assign new_n536 = new_n330 & new_n535;
  assign new_n537 = new_n530 & ~new_n536;
  assign new_n538 = ~pmusel4 & ~new_n537;
  assign new_n539 = ~new_n491 & new_n538;
  assign new_n540 = new_n522 & new_n538;
  assign new_n541 = ~new_n507 & ~new_n523;
  assign new_n542 = ~new_n539 & ~new_n540;
  assign new_n543 = new_n541 & new_n542;
  assign new_n544 = ~pina6 & ~new_n186;
  assign new_n545 = ~new_n186 & new_n241;
  assign new_n546 = ~pmusel1 & ~pina6;
  assign new_n547 = ~new_n544 & ~new_n545;
  assign new_n548 = ~new_n244 & ~new_n546;
  assign new_n549 = new_n547 & new_n548;
  assign new_n550 = new_n236 & new_n549;
  assign new_n551 = pinc6 & pmusel4;
  assign new_n552 = ~pmusel1 & new_n551;
  assign new_n553 = ~pmusel2 & new_n552;
  assign new_n554 = ~pmusel3 & new_n553;
  assign new_n555 = ~new_n550 & ~new_n554;
  assign new_n556 = ~new_n354 & ~new_n555;
  assign new_n557 = new_n354 & new_n555;
  assign new_n558 = ~new_n556 & ~new_n557;
  assign new_n559 = ~pina7 & ~new_n204;
  assign new_n560 = ~new_n204 & new_n241;
  assign new_n561 = ~pmusel1 & ~pina7;
  assign new_n562 = ~new_n559 & ~new_n560;
  assign new_n563 = ~new_n244 & ~new_n561;
  assign new_n564 = new_n562 & new_n563;
  assign new_n565 = new_n236 & new_n564;
  assign new_n566 = pmusel4 & pinc7;
  assign new_n567 = ~pmusel1 & new_n566;
  assign new_n568 = ~pmusel2 & new_n567;
  assign new_n569 = ~pmusel3 & new_n568;
  assign new_n570 = ~new_n565 & ~new_n569;
  assign new_n571 = ~new_n354 & ~new_n570;
  assign new_n572 = new_n354 & new_n570;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = ~new_n558 & ~new_n573;
  assign new_n575 = ~pmusel3 & pinb6;
  assign new_n576 = pmusel2 & new_n575;
  assign new_n577 = ~pmusel1 & new_n576;
  assign new_n578 = pmusel3 & pind6;
  assign new_n579 = ~pmusel2 & new_n578;
  assign new_n580 = ~pmusel1 & new_n579;
  assign new_n581 = ~new_n577 & ~new_n580;
  assign new_n582 = ~pina6 & ~pinc6;
  assign new_n583 = pmusel2 & ~pinc6;
  assign new_n584 = ~pmusel2 & ~pina6;
  assign new_n585 = ~new_n582 & ~new_n583;
  assign new_n586 = ~new_n584 & new_n585;
  assign new_n587 = new_n330 & new_n586;
  assign new_n588 = new_n581 & ~new_n587;
  assign new_n589 = ~pmusel4 & ~new_n588;
  assign new_n590 = ~new_n573 & new_n589;
  assign new_n591 = ~pmusel3 & pinb7;
  assign new_n592 = pmusel2 & new_n591;
  assign new_n593 = ~pmusel1 & new_n592;
  assign new_n594 = pmusel3 & pind7;
  assign new_n595 = ~pmusel2 & new_n594;
  assign new_n596 = ~pmusel1 & new_n595;
  assign new_n597 = ~new_n593 & ~new_n596;
  assign new_n598 = ~pina7 & ~pinc7;
  assign new_n599 = pmusel2 & ~pinc7;
  assign new_n600 = ~pmusel2 & ~pina7;
  assign new_n601 = ~new_n598 & ~new_n599;
  assign new_n602 = ~new_n600 & new_n601;
  assign new_n603 = new_n330 & new_n602;
  assign new_n604 = new_n597 & ~new_n603;
  assign new_n605 = ~pmusel4 & ~new_n604;
  assign new_n606 = ~new_n558 & new_n605;
  assign new_n607 = new_n589 & new_n605;
  assign new_n608 = ~new_n574 & ~new_n590;
  assign new_n609 = ~new_n606 & ~new_n607;
  assign new_n610 = new_n608 & new_n609;
  assign new_n611 = ~new_n543 & ~new_n610;
  assign new_n612 = ~pmusel3 & pinb3;
  assign new_n613 = pmusel2 & new_n612;
  assign new_n614 = ~pmusel1 & new_n613;
  assign new_n615 = pind3 & pmusel3;
  assign new_n616 = ~pmusel2 & new_n615;
  assign new_n617 = ~pmusel1 & new_n616;
  assign new_n618 = ~new_n614 & ~new_n617;
  assign new_n619 = ~pinc3 & ~pina3;
  assign new_n620 = ~pinc3 & pmusel2;
  assign new_n621 = ~pmusel2 & ~pina3;
  assign new_n622 = ~new_n619 & ~new_n620;
  assign new_n623 = ~new_n621 & new_n622;
  assign new_n624 = new_n330 & new_n623;
  assign new_n625 = new_n618 & ~new_n624;
  assign new_n626 = ~pmusel4 & ~new_n625;
  assign new_n627 = ~pina3 & ~new_n126;
  assign new_n628 = ~new_n126 & new_n241;
  assign new_n629 = ~pmusel1 & ~pina3;
  assign new_n630 = ~new_n627 & ~new_n628;
  assign new_n631 = ~new_n244 & ~new_n629;
  assign new_n632 = new_n630 & new_n631;
  assign new_n633 = new_n236 & new_n632;
  assign new_n634 = pinc3 & pmusel4;
  assign new_n635 = ~pmusel1 & new_n634;
  assign new_n636 = ~pmusel2 & new_n635;
  assign new_n637 = ~pmusel3 & new_n636;
  assign new_n638 = ~new_n633 & ~new_n637;
  assign new_n639 = ~new_n354 & ~new_n638;
  assign new_n640 = new_n354 & new_n638;
  assign new_n641 = ~new_n639 & ~new_n640;
  assign new_n642 = new_n626 & ~new_n641;
  assign new_n643 = ~pmusel3 & pinb2;
  assign new_n644 = pmusel2 & new_n643;
  assign new_n645 = ~pmusel1 & new_n644;
  assign new_n646 = pind2 & pmusel3;
  assign new_n647 = ~pmusel2 & new_n646;
  assign new_n648 = ~pmusel1 & new_n647;
  assign new_n649 = ~new_n645 & ~new_n648;
  assign new_n650 = ~pinc2 & ~pina2;
  assign new_n651 = ~pinc2 & pmusel2;
  assign new_n652 = ~pmusel2 & ~pina2;
  assign new_n653 = ~new_n650 & ~new_n651;
  assign new_n654 = ~new_n652 & new_n653;
  assign new_n655 = new_n330 & new_n654;
  assign new_n656 = new_n649 & ~new_n655;
  assign new_n657 = ~pmusel4 & ~new_n656;
  assign new_n658 = ~pina2 & ~new_n108;
  assign new_n659 = ~new_n108 & new_n241;
  assign new_n660 = ~pmusel1 & ~pina2;
  assign new_n661 = ~new_n658 & ~new_n659;
  assign new_n662 = ~new_n244 & ~new_n660;
  assign new_n663 = new_n661 & new_n662;
  assign new_n664 = new_n236 & new_n663;
  assign new_n665 = pinc2 & pmusel4;
  assign new_n666 = ~pmusel1 & new_n665;
  assign new_n667 = ~pmusel2 & new_n666;
  assign new_n668 = ~pmusel3 & new_n667;
  assign new_n669 = ~new_n664 & ~new_n668;
  assign new_n670 = ~new_n354 & ~new_n669;
  assign new_n671 = new_n354 & new_n669;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = new_n657 & ~new_n672;
  assign new_n674 = pinb1 & ~pmusel3;
  assign new_n675 = pmusel2 & new_n674;
  assign new_n676 = ~pmusel1 & new_n675;
  assign new_n677 = pmusel3 & pind1;
  assign new_n678 = ~pmusel2 & new_n677;
  assign new_n679 = ~pmusel1 & new_n678;
  assign new_n680 = ~new_n676 & ~new_n679;
  assign new_n681 = ~pina1 & ~pinc1;
  assign new_n682 = pmusel2 & ~pinc1;
  assign new_n683 = ~pina1 & ~pmusel2;
  assign new_n684 = ~new_n681 & ~new_n682;
  assign new_n685 = ~new_n683 & new_n684;
  assign new_n686 = new_n330 & new_n685;
  assign new_n687 = new_n680 & ~new_n686;
  assign new_n688 = ~pmusel4 & ~new_n687;
  assign new_n689 = ~pina1 & ~new_n117;
  assign new_n690 = ~new_n117 & new_n241;
  assign new_n691 = ~pina1 & ~pmusel1;
  assign new_n692 = ~new_n689 & ~new_n690;
  assign new_n693 = ~new_n244 & ~new_n691;
  assign new_n694 = new_n692 & new_n693;
  assign new_n695 = new_n236 & new_n694;
  assign new_n696 = pinc1 & pmusel4;
  assign new_n697 = ~pmusel1 & new_n696;
  assign new_n698 = ~pmusel2 & new_n697;
  assign new_n699 = ~pmusel3 & new_n698;
  assign new_n700 = ~new_n695 & ~new_n699;
  assign new_n701 = ~new_n354 & ~new_n700;
  assign new_n702 = new_n354 & new_n700;
  assign new_n703 = ~new_n701 & ~new_n702;
  assign new_n704 = new_n688 & ~new_n703;
  assign new_n705 = pinb0 & ~pmusel3;
  assign new_n706 = pmusel2 & new_n705;
  assign new_n707 = ~pmusel1 & new_n706;
  assign new_n708 = pmusel3 & pind0;
  assign new_n709 = ~pmusel2 & new_n708;
  assign new_n710 = ~pmusel1 & new_n709;
  assign new_n711 = ~new_n707 & ~new_n710;
  assign new_n712 = ~pina0 & ~pinc0;
  assign new_n713 = pmusel2 & ~pinc0;
  assign new_n714 = ~pina0 & ~pmusel2;
  assign new_n715 = ~new_n712 & ~new_n713;
  assign new_n716 = ~new_n714 & new_n715;
  assign new_n717 = new_n330 & new_n716;
  assign new_n718 = new_n711 & ~new_n717;
  assign new_n719 = ~pmusel4 & ~new_n718;
  assign new_n720 = ~pina0 & ~new_n92;
  assign new_n721 = ~new_n92 & new_n241;
  assign new_n722 = ~pina0 & ~pmusel1;
  assign new_n723 = ~new_n720 & ~new_n721;
  assign new_n724 = ~new_n244 & ~new_n722;
  assign new_n725 = new_n723 & new_n724;
  assign new_n726 = new_n236 & new_n725;
  assign new_n727 = pinc0 & pmusel4;
  assign new_n728 = ~pmusel1 & new_n727;
  assign new_n729 = ~pmusel2 & new_n728;
  assign new_n730 = ~pmusel3 & new_n729;
  assign new_n731 = ~new_n726 & ~new_n730;
  assign new_n732 = ~new_n354 & ~new_n731;
  assign new_n733 = new_n354 & new_n731;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = new_n719 & ~new_n734;
  assign new_n736 = ~new_n704 & ~new_n735;
  assign new_n737 = ~new_n688 & new_n703;
  assign new_n738 = ~new_n704 & new_n737;
  assign new_n739 = ~new_n736 & ~new_n738;
  assign new_n740 = ~new_n672 & new_n739;
  assign new_n741 = new_n657 & new_n739;
  assign new_n742 = ~new_n740 & ~new_n741;
  assign new_n743 = ~new_n673 & new_n742;
  assign new_n744 = ~new_n626 & new_n641;
  assign new_n745 = ~new_n743 & ~new_n744;
  assign new_n746 = ~new_n642 & ~new_n745;
  assign new_n747 = ~new_n703 & ~new_n734;
  assign new_n748 = ~new_n703 & new_n719;
  assign new_n749 = new_n688 & ~new_n734;
  assign new_n750 = new_n688 & new_n719;
  assign new_n751 = ~new_n747 & ~new_n748;
  assign new_n752 = ~new_n749 & ~new_n750;
  assign new_n753 = new_n751 & new_n752;
  assign new_n754 = ~new_n641 & ~new_n672;
  assign new_n755 = ~new_n641 & new_n657;
  assign new_n756 = new_n626 & ~new_n672;
  assign new_n757 = new_n626 & new_n657;
  assign new_n758 = ~new_n754 & ~new_n755;
  assign new_n759 = ~new_n756 & ~new_n757;
  assign new_n760 = new_n758 & new_n759;
  assign new_n761 = ~new_n753 & ~new_n760;
  assign new_n762 = ~popsel3 & popsel2;
  assign new_n763 = popsel1 & new_n762;
  assign new_n764 = ~popsel1 & new_n313;
  assign new_n765 = ~new_n763 & ~new_n764;
  assign new_n766 = ~popsel0 & ~new_n765;
  assign new_n767 = new_n761 & new_n766;
  assign new_n768 = new_n746 & ~new_n767;
  assign new_n769 = new_n611 & ~new_n768;
  assign new_n770 = ~new_n573 & new_n605;
  assign new_n771 = ~new_n558 & new_n589;
  assign new_n772 = ~new_n506 & new_n538;
  assign new_n773 = ~new_n491 & new_n522;
  assign new_n774 = ~new_n772 & ~new_n773;
  assign new_n775 = new_n506 & ~new_n538;
  assign new_n776 = ~new_n772 & new_n775;
  assign new_n777 = ~new_n774 & ~new_n776;
  assign new_n778 = ~new_n558 & new_n777;
  assign new_n779 = new_n589 & new_n777;
  assign new_n780 = ~new_n778 & ~new_n779;
  assign new_n781 = ~new_n771 & new_n780;
  assign new_n782 = new_n573 & ~new_n605;
  assign new_n783 = ~new_n781 & ~new_n782;
  assign new_n784 = ~new_n770 & ~new_n783;
  assign new_n785 = ~new_n769 & new_n784;
  assign new_n786 = ~new_n469 & ~new_n476;
  assign new_n787 = ~new_n785 & new_n786;
  assign new_n788 = ~new_n462 & ~new_n787;
  assign new_n789 = ~pina12 & ~new_n219;
  assign new_n790 = ~new_n219 & new_n241;
  assign new_n791 = ~pmusel1 & ~pina12;
  assign new_n792 = ~new_n789 & ~new_n790;
  assign new_n793 = ~new_n244 & ~new_n791;
  assign new_n794 = new_n792 & new_n793;
  assign new_n795 = new_n236 & new_n794;
  assign new_n796 = pinc12 & pmusel4;
  assign new_n797 = ~pmusel1 & new_n796;
  assign new_n798 = ~pmusel2 & new_n797;
  assign new_n799 = ~pmusel3 & new_n798;
  assign new_n800 = ~new_n795 & ~new_n799;
  assign new_n801 = ~new_n354 & ~new_n800;
  assign new_n802 = new_n354 & new_n800;
  assign new_n803 = ~new_n801 & ~new_n802;
  assign new_n804 = ~pmusel3 & pinb12;
  assign new_n805 = pmusel2 & new_n804;
  assign new_n806 = ~pmusel1 & new_n805;
  assign new_n807 = pmusel3 & pind12;
  assign new_n808 = ~pmusel2 & new_n807;
  assign new_n809 = ~pmusel1 & new_n808;
  assign new_n810 = ~new_n806 & ~new_n809;
  assign new_n811 = ~pinc12 & ~pina12;
  assign new_n812 = pmusel2 & ~pinc12;
  assign new_n813 = ~pmusel2 & ~pina12;
  assign new_n814 = ~new_n811 & ~new_n812;
  assign new_n815 = ~new_n813 & new_n814;
  assign new_n816 = new_n330 & new_n815;
  assign new_n817 = new_n810 & ~new_n816;
  assign new_n818 = ~pmusel4 & ~new_n817;
  assign new_n819 = new_n803 & new_n818;
  assign new_n820 = ~new_n803 & ~new_n818;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = new_n788 & ~new_n821;
  assign new_n823 = ~new_n788 & new_n821;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = ~new_n232 & new_n824;
  assign new_n826 = new_n304 & new_n316;
  assign new_n827 = new_n304 & new_n824;
  assign new_n828 = ~new_n317 & ~new_n825;
  assign new_n829 = ~new_n826 & ~new_n827;
  assign new_n830 = new_n828 & new_n829;
  assign new_n831 = new_n313 & new_n830;
  assign po12 = new_n312 | new_n831;
  assign new_n833 = ~new_n164 & new_n217;
  assign new_n834 = new_n174 & new_n833;
  assign new_n835 = new_n173 & new_n834;
  assign new_n836 = ~new_n173 & ~new_n834;
  assign new_n837 = ~new_n835 & ~new_n836;
  assign new_n838 = popsel2 & ~new_n837;
  assign new_n839 = new_n232 & new_n838;
  assign new_n840 = ~popsel2 & new_n837;
  assign new_n841 = ~psh2 & ~new_n279;
  assign new_n842 = ~psh2 & ~new_n841;
  assign new_n843 = pmusel2 & pind11;
  assign new_n844 = ~pinb11 & ~new_n843;
  assign new_n845 = new_n241 & ~new_n843;
  assign new_n846 = ~pmusel1 & ~pinb11;
  assign new_n847 = ~new_n844 & ~new_n845;
  assign new_n848 = ~new_n244 & ~new_n846;
  assign new_n849 = new_n847 & new_n848;
  assign new_n850 = new_n236 & new_n849;
  assign new_n851 = ~pmusel3 & pind11;
  assign new_n852 = new_n264 & new_n851;
  assign new_n853 = ~new_n850 & ~new_n852;
  assign new_n854 = ~new_n841 & new_n853;
  assign new_n855 = ~new_n842 & ~new_n854;
  assign new_n856 = new_n235 & new_n855;
  assign new_n857 = psh1 & ~new_n266;
  assign new_n858 = new_n853 & ~new_n857;
  assign new_n859 = psh1 & ~new_n857;
  assign new_n860 = ~new_n858 & ~new_n859;
  assign new_n861 = ~psh0 & new_n860;
  assign new_n862 = new_n254 & ~new_n291;
  assign new_n863 = ~new_n861 & ~new_n862;
  assign new_n864 = psh2 & ~new_n252;
  assign new_n865 = new_n863 & ~new_n864;
  assign new_n866 = psh2 & ~new_n864;
  assign new_n867 = new_n235 & new_n863;
  assign new_n868 = psh2 & new_n235;
  assign new_n869 = ~new_n865 & ~new_n866;
  assign new_n870 = ~new_n867 & ~new_n868;
  assign new_n871 = new_n869 & new_n870;
  assign new_n872 = ~new_n856 & ~new_n871;
  assign new_n873 = new_n837 & new_n872;
  assign new_n874 = popsel2 & new_n872;
  assign new_n875 = ~new_n873 & ~new_n874;
  assign new_n876 = ~new_n840 & new_n875;
  assign new_n877 = ~new_n839 & ~new_n876;
  assign new_n878 = new_n232 & ~new_n839;
  assign new_n879 = ~new_n877 & ~new_n878;
  assign new_n880 = ~popsel3 & new_n879;
  assign new_n881 = popsel1 & popsel0;
  assign new_n882 = ~new_n232 & ~new_n881;
  assign new_n883 = ~new_n333 & ~new_n455;
  assign new_n884 = new_n333 & new_n455;
  assign new_n885 = ~new_n883 & ~new_n884;
  assign new_n886 = ~new_n416 & new_n431;
  assign new_n887 = ~new_n432 & new_n886;
  assign new_n888 = ~new_n432 & new_n785;
  assign new_n889 = ~new_n887 & ~new_n888;
  assign new_n890 = ~new_n385 & new_n400;
  assign new_n891 = new_n889 & ~new_n890;
  assign new_n892 = ~new_n401 & ~new_n891;
  assign new_n893 = ~new_n437 & ~new_n892;
  assign new_n894 = new_n885 & new_n893;
  assign new_n895 = new_n370 & new_n885;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = ~new_n886 & ~new_n888;
  assign new_n898 = ~new_n890 & new_n897;
  assign new_n899 = new_n401 & ~new_n890;
  assign new_n900 = ~new_n898 & ~new_n899;
  assign new_n901 = ~new_n370 & new_n900;
  assign new_n902 = ~new_n437 & ~new_n901;
  assign new_n903 = new_n896 & new_n902;
  assign new_n904 = new_n885 & new_n896;
  assign new_n905 = ~new_n903 & ~new_n904;
  assign new_n906 = new_n882 & new_n905;
  assign new_n907 = new_n232 & ~new_n872;
  assign new_n908 = ~new_n906 & ~new_n907;
  assign new_n909 = new_n313 & ~new_n908;
  assign po11 = new_n880 | new_n909;
  assign new_n911 = pmusel2 & pinc13;
  assign new_n912 = ~pmusel1 & new_n911;
  assign new_n913 = ~pmusel2 & pina13;
  assign new_n914 = pmusel1 & new_n913;
  assign new_n915 = ~new_n912 & ~new_n914;
  assign new_n916 = new_n97 & ~new_n915;
  assign new_n917 = ~new_n104 & new_n916;
  assign new_n918 = new_n104 & ~new_n916;
  assign new_n919 = ~new_n917 & ~new_n918;
  assign new_n920 = ~new_n227 & ~new_n919;
  assign new_n921 = new_n218 & new_n920;
  assign new_n922 = pmusel2 & pinc14;
  assign new_n923 = ~pmusel1 & new_n922;
  assign new_n924 = ~pmusel2 & pina14;
  assign new_n925 = pmusel1 & new_n924;
  assign new_n926 = ~new_n923 & ~new_n925;
  assign new_n927 = new_n97 & ~new_n926;
  assign new_n928 = ~new_n104 & new_n927;
  assign new_n929 = new_n104 & ~new_n927;
  assign new_n930 = ~new_n928 & ~new_n929;
  assign new_n931 = new_n921 & new_n930;
  assign new_n932 = ~new_n921 & ~new_n930;
  assign new_n933 = ~new_n931 & ~new_n932;
  assign new_n934 = popsel2 & ~new_n933;
  assign new_n935 = new_n232 & new_n934;
  assign new_n936 = ~popsel2 & new_n933;
  assign new_n937 = psh1 & ~psh2;
  assign new_n938 = ~psh0 & ~psh2;
  assign new_n939 = ~new_n937 & ~new_n938;
  assign new_n940 = ~new_n235 & new_n939;
  assign new_n941 = ~new_n937 & ~new_n940;
  assign new_n942 = ~new_n279 & new_n941;
  assign new_n943 = ~new_n252 & ~new_n941;
  assign new_n944 = ~new_n942 & ~new_n943;
  assign new_n945 = new_n933 & new_n944;
  assign new_n946 = popsel2 & new_n944;
  assign new_n947 = ~new_n945 & ~new_n946;
  assign new_n948 = ~new_n936 & new_n947;
  assign new_n949 = ~new_n935 & ~new_n948;
  assign new_n950 = new_n232 & ~new_n935;
  assign new_n951 = ~new_n949 & ~new_n950;
  assign new_n952 = ~popsel3 & new_n951;
  assign new_n953 = ~pina14 & ~new_n922;
  assign new_n954 = new_n241 & ~new_n922;
  assign new_n955 = ~pmusel1 & ~pina14;
  assign new_n956 = ~new_n953 & ~new_n954;
  assign new_n957 = ~new_n244 & ~new_n955;
  assign new_n958 = new_n956 & new_n957;
  assign new_n959 = new_n236 & new_n958;
  assign new_n960 = pinc14 & pmusel4;
  assign new_n961 = ~pmusel1 & new_n960;
  assign new_n962 = ~pmusel2 & new_n961;
  assign new_n963 = ~pmusel3 & new_n962;
  assign new_n964 = ~new_n959 & ~new_n963;
  assign new_n965 = ~new_n354 & ~new_n964;
  assign new_n966 = new_n354 & new_n964;
  assign new_n967 = ~new_n965 & ~new_n966;
  assign new_n968 = ~pmusel3 & pinb14;
  assign new_n969 = pmusel2 & new_n968;
  assign new_n970 = ~pmusel1 & new_n969;
  assign new_n971 = pmusel3 & pind14;
  assign new_n972 = ~pmusel2 & new_n971;
  assign new_n973 = ~pmusel1 & new_n972;
  assign new_n974 = ~new_n970 & ~new_n973;
  assign new_n975 = ~pinc14 & ~pina14;
  assign new_n976 = pmusel2 & ~pinc14;
  assign new_n977 = ~pmusel2 & ~pina14;
  assign new_n978 = ~new_n975 & ~new_n976;
  assign new_n979 = ~new_n977 & new_n978;
  assign new_n980 = new_n330 & new_n979;
  assign new_n981 = new_n974 & ~new_n980;
  assign new_n982 = ~pmusel4 & ~new_n981;
  assign new_n983 = ~new_n967 & ~new_n982;
  assign new_n984 = new_n967 & new_n982;
  assign new_n985 = ~new_n983 & ~new_n984;
  assign new_n986 = new_n803 & ~new_n818;
  assign new_n987 = ~new_n788 & ~new_n986;
  assign new_n988 = ~new_n803 & new_n818;
  assign new_n989 = ~new_n987 & ~new_n988;
  assign new_n990 = ~pina13 & ~new_n911;
  assign new_n991 = new_n241 & ~new_n911;
  assign new_n992 = ~pmusel1 & ~pina13;
  assign new_n993 = ~new_n990 & ~new_n991;
  assign new_n994 = ~new_n244 & ~new_n992;
  assign new_n995 = new_n993 & new_n994;
  assign new_n996 = new_n236 & new_n995;
  assign new_n997 = pinc13 & pmusel4;
  assign new_n998 = ~pmusel1 & new_n997;
  assign new_n999 = ~pmusel2 & new_n998;
  assign new_n1000 = ~pmusel3 & new_n999;
  assign new_n1001 = ~new_n996 & ~new_n1000;
  assign new_n1002 = ~new_n354 & ~new_n1001;
  assign new_n1003 = new_n354 & new_n1001;
  assign new_n1004 = ~new_n1002 & ~new_n1003;
  assign new_n1005 = ~pmusel3 & pinb13;
  assign new_n1006 = pmusel2 & new_n1005;
  assign new_n1007 = ~pmusel1 & new_n1006;
  assign new_n1008 = pmusel3 & pind13;
  assign new_n1009 = ~pmusel2 & new_n1008;
  assign new_n1010 = ~pmusel1 & new_n1009;
  assign new_n1011 = ~new_n1007 & ~new_n1010;
  assign new_n1012 = ~pinc13 & ~pina13;
  assign new_n1013 = pmusel2 & ~pinc13;
  assign new_n1014 = ~pmusel2 & ~pina13;
  assign new_n1015 = ~new_n1012 & ~new_n1013;
  assign new_n1016 = ~new_n1014 & new_n1015;
  assign new_n1017 = new_n330 & new_n1016;
  assign new_n1018 = new_n1011 & ~new_n1017;
  assign new_n1019 = ~pmusel4 & ~new_n1018;
  assign new_n1020 = new_n1004 & ~new_n1019;
  assign new_n1021 = ~new_n989 & ~new_n1020;
  assign new_n1022 = new_n985 & new_n1021;
  assign new_n1023 = ~new_n1004 & new_n1019;
  assign new_n1024 = new_n985 & new_n1023;
  assign new_n1025 = ~new_n1022 & ~new_n1024;
  assign new_n1026 = new_n985 & new_n1025;
  assign new_n1027 = new_n788 & ~new_n988;
  assign new_n1028 = ~new_n986 & ~new_n1027;
  assign new_n1029 = ~new_n1023 & ~new_n1028;
  assign new_n1030 = ~new_n1020 & ~new_n1029;
  assign new_n1031 = new_n1025 & new_n1030;
  assign new_n1032 = ~new_n1026 & ~new_n1031;
  assign new_n1033 = new_n882 & new_n1032;
  assign new_n1034 = new_n232 & ~new_n944;
  assign new_n1035 = ~new_n1033 & ~new_n1034;
  assign new_n1036 = new_n313 & ~new_n1035;
  assign po14 = new_n952 | new_n1036;
  assign new_n1038 = new_n218 & ~new_n227;
  assign new_n1039 = new_n919 & new_n1038;
  assign new_n1040 = ~new_n919 & ~new_n1038;
  assign new_n1041 = ~new_n1039 & ~new_n1040;
  assign new_n1042 = popsel2 & ~new_n1041;
  assign new_n1043 = new_n232 & new_n1042;
  assign new_n1044 = ~popsel2 & new_n1041;
  assign new_n1045 = psh0 & psh2;
  assign new_n1046 = new_n857 & new_n1045;
  assign new_n1047 = ~psh1 & ~psh2;
  assign new_n1048 = ~psh1 & psh2;
  assign new_n1049 = psh1 & ~new_n1045;
  assign new_n1050 = ~new_n1048 & ~new_n1049;
  assign new_n1051 = ~new_n1047 & new_n1050;
  assign new_n1052 = psh0 & ~new_n279;
  assign new_n1053 = ~psh0 & ~new_n266;
  assign new_n1054 = ~new_n1052 & ~new_n1053;
  assign new_n1055 = new_n1050 & new_n1054;
  assign new_n1056 = new_n252 & ~new_n1047;
  assign new_n1057 = new_n252 & new_n1054;
  assign new_n1058 = ~new_n1051 & ~new_n1055;
  assign new_n1059 = ~new_n1056 & ~new_n1057;
  assign new_n1060 = new_n1058 & new_n1059;
  assign new_n1061 = ~new_n1046 & ~new_n1060;
  assign new_n1062 = new_n1041 & new_n1061;
  assign new_n1063 = popsel2 & new_n1061;
  assign new_n1064 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = ~new_n1044 & new_n1064;
  assign new_n1066 = ~new_n1043 & ~new_n1065;
  assign new_n1067 = new_n232 & ~new_n1043;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = ~popsel3 & new_n1068;
  assign new_n1070 = ~new_n1004 & ~new_n1019;
  assign new_n1071 = new_n1004 & new_n1019;
  assign new_n1072 = ~new_n1070 & ~new_n1071;
  assign new_n1073 = new_n987 & new_n1072;
  assign new_n1074 = new_n988 & new_n1072;
  assign new_n1075 = ~new_n1073 & ~new_n1074;
  assign new_n1076 = new_n1072 & new_n1075;
  assign new_n1077 = new_n1028 & new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = new_n882 & new_n1078;
  assign new_n1080 = new_n232 & ~new_n1061;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign new_n1082 = new_n313 & ~new_n1081;
  assign po13 = new_n1069 | new_n1082;
  assign new_n1084 = new_n218 & ~new_n919;
  assign new_n1085 = ~new_n227 & ~new_n930;
  assign new_n1086 = new_n1084 & new_n1085;
  assign new_n1087 = popsel2 & new_n1086;
  assign new_n1088 = new_n232 & new_n1087;
  assign new_n1089 = ~popsel2 & new_n1086;
  assign new_n1090 = popsel2 & ~new_n252;
  assign new_n1091 = ~new_n1089 & ~new_n1090;
  assign new_n1092 = ~new_n1088 & new_n1091;
  assign new_n1093 = new_n232 & ~new_n1088;
  assign new_n1094 = ~new_n1092 & ~new_n1093;
  assign new_n1095 = ~popsel3 & new_n1094;
  assign new_n1096 = ~pina15 & ~new_n99;
  assign new_n1097 = ~new_n99 & new_n241;
  assign new_n1098 = ~pmusel1 & ~pina15;
  assign new_n1099 = ~new_n1096 & ~new_n1097;
  assign new_n1100 = ~new_n244 & ~new_n1098;
  assign new_n1101 = new_n1099 & new_n1100;
  assign new_n1102 = new_n236 & new_n1101;
  assign new_n1103 = pinc15 & pmusel4;
  assign new_n1104 = ~pmusel1 & new_n1103;
  assign new_n1105 = ~pmusel2 & new_n1104;
  assign new_n1106 = ~pmusel3 & new_n1105;
  assign new_n1107 = ~new_n1102 & ~new_n1106;
  assign new_n1108 = ~new_n354 & ~new_n1107;
  assign new_n1109 = new_n354 & new_n1107;
  assign new_n1110 = ~new_n1108 & ~new_n1109;
  assign new_n1111 = ~pmusel3 & pinb15;
  assign new_n1112 = pmusel2 & new_n1111;
  assign new_n1113 = ~pmusel1 & new_n1112;
  assign new_n1114 = pmusel3 & pind15;
  assign new_n1115 = ~pmusel2 & new_n1114;
  assign new_n1116 = ~pmusel1 & new_n1115;
  assign new_n1117 = ~new_n1113 & ~new_n1116;
  assign new_n1118 = ~pinc15 & ~pina15;
  assign new_n1119 = pmusel2 & ~pinc15;
  assign new_n1120 = ~pmusel2 & ~pina15;
  assign new_n1121 = ~new_n1118 & ~new_n1119;
  assign new_n1122 = ~new_n1120 & new_n1121;
  assign new_n1123 = new_n330 & new_n1122;
  assign new_n1124 = new_n1117 & ~new_n1123;
  assign new_n1125 = ~pmusel4 & ~new_n1124;
  assign new_n1126 = new_n1110 & new_n1125;
  assign new_n1127 = ~new_n1110 & ~new_n1125;
  assign new_n1128 = ~new_n1126 & ~new_n1127;
  assign new_n1129 = new_n986 & ~new_n988;
  assign new_n1130 = ~new_n1027 & ~new_n1129;
  assign new_n1131 = ~new_n1020 & new_n1130;
  assign new_n1132 = ~new_n1023 & ~new_n1131;
  assign new_n1133 = new_n967 & ~new_n982;
  assign new_n1134 = ~new_n1132 & ~new_n1133;
  assign new_n1135 = new_n1128 & new_n1134;
  assign new_n1136 = ~new_n967 & new_n982;
  assign new_n1137 = new_n1128 & new_n1136;
  assign new_n1138 = ~new_n1135 & ~new_n1137;
  assign new_n1139 = ~new_n1020 & new_n1028;
  assign new_n1140 = ~new_n1020 & new_n1023;
  assign new_n1141 = ~new_n1139 & ~new_n1140;
  assign new_n1142 = ~new_n1136 & new_n1141;
  assign new_n1143 = ~new_n1133 & ~new_n1142;
  assign new_n1144 = new_n1138 & new_n1143;
  assign new_n1145 = new_n1128 & new_n1138;
  assign new_n1146 = ~new_n1144 & ~new_n1145;
  assign new_n1147 = new_n882 & new_n1146;
  assign new_n1148 = new_n232 & ~new_n252;
  assign new_n1149 = ~new_n1147 & ~new_n1148;
  assign new_n1150 = new_n313 & ~new_n1149;
  assign po15 = new_n1095 | new_n1150;
  assign new_n1152 = ~new_n146 & new_n217;
  assign new_n1153 = new_n164 & new_n1152;
  assign new_n1154 = ~new_n164 & ~new_n1152;
  assign new_n1155 = ~new_n1153 & ~new_n1154;
  assign new_n1156 = popsel2 & ~new_n1155;
  assign new_n1157 = new_n232 & new_n1156;
  assign new_n1158 = ~popsel2 & new_n1155;
  assign new_n1159 = psh2 & ~new_n266;
  assign new_n1160 = pmusel2 & pind9;
  assign new_n1161 = ~pinb9 & ~new_n1160;
  assign new_n1162 = new_n241 & ~new_n1160;
  assign new_n1163 = ~pmusel1 & ~pinb9;
  assign new_n1164 = ~new_n1161 & ~new_n1162;
  assign new_n1165 = ~new_n244 & ~new_n1163;
  assign new_n1166 = new_n1164 & new_n1165;
  assign new_n1167 = new_n236 & new_n1166;
  assign new_n1168 = ~pmusel3 & pind9;
  assign new_n1169 = new_n264 & new_n1168;
  assign new_n1170 = ~new_n1167 & ~new_n1169;
  assign new_n1171 = ~psh2 & ~new_n1170;
  assign new_n1172 = ~new_n1159 & ~new_n1171;
  assign new_n1173 = ~psh1 & new_n1172;
  assign new_n1174 = ~psh2 & ~new_n853;
  assign new_n1175 = ~new_n864 & ~new_n1174;
  assign new_n1176 = new_n1172 & new_n1175;
  assign new_n1177 = psh1 & new_n1175;
  assign new_n1178 = ~new_n1176 & ~new_n1177;
  assign new_n1179 = ~new_n1173 & new_n1178;
  assign new_n1180 = ~psh0 & new_n1179;
  assign new_n1181 = psh2 & ~new_n279;
  assign new_n1182 = pmusel2 & pind10;
  assign new_n1183 = ~pinb10 & ~new_n1182;
  assign new_n1184 = new_n241 & ~new_n1182;
  assign new_n1185 = ~pmusel1 & ~pinb10;
  assign new_n1186 = ~new_n1183 & ~new_n1184;
  assign new_n1187 = ~new_n244 & ~new_n1185;
  assign new_n1188 = new_n1186 & new_n1187;
  assign new_n1189 = new_n236 & new_n1188;
  assign new_n1190 = ~pmusel3 & pind10;
  assign new_n1191 = new_n264 & new_n1190;
  assign new_n1192 = ~new_n1189 & ~new_n1191;
  assign new_n1193 = ~psh2 & ~new_n1192;
  assign new_n1194 = ~new_n1181 & ~new_n1193;
  assign new_n1195 = ~psh1 & new_n1194;
  assign new_n1196 = ~psh2 & ~new_n291;
  assign new_n1197 = psh2 & ~new_n1170;
  assign new_n1198 = ~new_n1196 & ~new_n1197;
  assign new_n1199 = new_n1194 & new_n1198;
  assign new_n1200 = psh1 & new_n1198;
  assign new_n1201 = ~new_n1199 & ~new_n1200;
  assign new_n1202 = ~new_n1195 & new_n1201;
  assign new_n1203 = psh0 & new_n1202;
  assign new_n1204 = ~new_n1180 & ~new_n1203;
  assign new_n1205 = new_n1155 & new_n1204;
  assign new_n1206 = popsel2 & new_n1204;
  assign new_n1207 = ~new_n1205 & ~new_n1206;
  assign new_n1208 = ~new_n1158 & new_n1207;
  assign new_n1209 = ~new_n1157 & ~new_n1208;
  assign new_n1210 = new_n232 & ~new_n1157;
  assign new_n1211 = ~new_n1209 & ~new_n1210;
  assign new_n1212 = ~popsel3 & new_n1211;
  assign new_n1213 = ~new_n385 & ~new_n400;
  assign new_n1214 = new_n385 & new_n400;
  assign new_n1215 = ~new_n1213 & ~new_n1214;
  assign new_n1216 = ~new_n785 & ~new_n886;
  assign new_n1217 = new_n1215 & new_n1216;
  assign new_n1218 = new_n432 & new_n1215;
  assign new_n1219 = ~new_n1217 & ~new_n1218;
  assign new_n1220 = new_n1215 & new_n1219;
  assign new_n1221 = new_n897 & new_n1219;
  assign new_n1222 = ~new_n1220 & ~new_n1221;
  assign new_n1223 = new_n882 & new_n1222;
  assign new_n1224 = new_n232 & ~new_n1204;
  assign new_n1225 = ~new_n1223 & ~new_n1224;
  assign new_n1226 = new_n313 & ~new_n1225;
  assign po9 = new_n1212 | new_n1226;
  assign new_n1228 = new_n146 & new_n217;
  assign new_n1229 = ~new_n146 & ~new_n217;
  assign new_n1230 = ~new_n1228 & ~new_n1229;
  assign new_n1231 = popsel2 & ~new_n1230;
  assign new_n1232 = new_n232 & new_n1231;
  assign new_n1233 = ~popsel2 & new_n1230;
  assign new_n1234 = psh2 & ~new_n291;
  assign new_n1235 = pmusel2 & pind8;
  assign new_n1236 = ~pinb8 & ~new_n1235;
  assign new_n1237 = new_n241 & ~new_n1235;
  assign new_n1238 = ~pmusel1 & ~pinb8;
  assign new_n1239 = ~new_n1236 & ~new_n1237;
  assign new_n1240 = ~new_n244 & ~new_n1238;
  assign new_n1241 = new_n1239 & new_n1240;
  assign new_n1242 = new_n236 & new_n1241;
  assign new_n1243 = ~pmusel3 & pind8;
  assign new_n1244 = new_n264 & new_n1243;
  assign new_n1245 = ~new_n1242 & ~new_n1244;
  assign new_n1246 = ~psh2 & ~new_n1245;
  assign new_n1247 = ~new_n1234 & ~new_n1246;
  assign new_n1248 = ~psh1 & new_n1247;
  assign new_n1249 = ~new_n864 & ~new_n1193;
  assign new_n1250 = new_n1247 & new_n1249;
  assign new_n1251 = psh1 & new_n1249;
  assign new_n1252 = ~new_n1250 & ~new_n1251;
  assign new_n1253 = ~new_n1248 & new_n1252;
  assign new_n1254 = ~psh0 & new_n1253;
  assign new_n1255 = psh2 & ~new_n1245;
  assign new_n1256 = ~new_n1174 & ~new_n1255;
  assign new_n1257 = new_n1172 & new_n1256;
  assign new_n1258 = psh1 & new_n1256;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = ~new_n1173 & new_n1259;
  assign new_n1261 = psh0 & new_n1260;
  assign new_n1262 = ~new_n1254 & ~new_n1261;
  assign new_n1263 = new_n1230 & new_n1262;
  assign new_n1264 = popsel2 & new_n1262;
  assign new_n1265 = ~new_n1263 & ~new_n1264;
  assign new_n1266 = ~new_n1233 & new_n1265;
  assign new_n1267 = ~new_n1232 & ~new_n1266;
  assign new_n1268 = new_n232 & ~new_n1232;
  assign new_n1269 = ~new_n1267 & ~new_n1268;
  assign new_n1270 = ~popsel3 & new_n1269;
  assign new_n1271 = ~new_n416 & ~new_n431;
  assign new_n1272 = new_n416 & new_n431;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = new_n785 & ~new_n1273;
  assign new_n1275 = ~new_n785 & new_n1273;
  assign new_n1276 = ~new_n1274 & ~new_n1275;
  assign new_n1277 = ~new_n232 & new_n1276;
  assign new_n1278 = new_n316 & new_n1262;
  assign new_n1279 = new_n1262 & new_n1276;
  assign new_n1280 = ~new_n317 & ~new_n1277;
  assign new_n1281 = ~new_n1278 & ~new_n1279;
  assign new_n1282 = new_n1280 & new_n1281;
  assign new_n1283 = new_n313 & new_n1282;
  assign po8 = new_n1270 | new_n1283;
  assign new_n1285 = new_n104 & new_n137;
  assign new_n1286 = ~new_n203 & new_n1285;
  assign new_n1287 = new_n213 & new_n1286;
  assign new_n1288 = new_n212 & new_n1287;
  assign new_n1289 = ~new_n212 & ~new_n1287;
  assign new_n1290 = ~new_n1288 & ~new_n1289;
  assign new_n1291 = popsel2 & ~new_n1290;
  assign new_n1292 = new_n232 & new_n1291;
  assign new_n1293 = ~popsel2 & new_n1290;
  assign new_n1294 = psh2 & ~new_n853;
  assign new_n1295 = pmusel2 & pind7;
  assign new_n1296 = ~pinb7 & ~new_n1295;
  assign new_n1297 = new_n241 & ~new_n1295;
  assign new_n1298 = ~pmusel1 & ~pinb7;
  assign new_n1299 = ~new_n1296 & ~new_n1297;
  assign new_n1300 = ~new_n244 & ~new_n1298;
  assign new_n1301 = new_n1299 & new_n1300;
  assign new_n1302 = new_n236 & new_n1301;
  assign new_n1303 = ~pmusel3 & pind7;
  assign new_n1304 = new_n264 & new_n1303;
  assign new_n1305 = ~new_n1302 & ~new_n1304;
  assign new_n1306 = ~psh2 & ~new_n1305;
  assign new_n1307 = ~new_n1294 & ~new_n1306;
  assign new_n1308 = ~psh1 & new_n1307;
  assign new_n1309 = ~new_n864 & ~new_n1171;
  assign new_n1310 = new_n1307 & new_n1309;
  assign new_n1311 = psh1 & new_n1309;
  assign new_n1312 = ~new_n1310 & ~new_n1311;
  assign new_n1313 = ~new_n1308 & new_n1312;
  assign new_n1314 = ~psh0 & new_n1313;
  assign new_n1315 = psh2 & ~new_n1305;
  assign new_n1316 = ~new_n1193 & ~new_n1315;
  assign new_n1317 = new_n1247 & new_n1316;
  assign new_n1318 = psh1 & new_n1316;
  assign new_n1319 = ~new_n1317 & ~new_n1318;
  assign new_n1320 = ~new_n1248 & new_n1319;
  assign new_n1321 = psh0 & new_n1320;
  assign new_n1322 = ~new_n1314 & ~new_n1321;
  assign new_n1323 = new_n1290 & new_n1322;
  assign new_n1324 = popsel2 & new_n1322;
  assign new_n1325 = ~new_n1323 & ~new_n1324;
  assign new_n1326 = ~new_n1293 & new_n1325;
  assign new_n1327 = ~new_n1292 & ~new_n1326;
  assign new_n1328 = new_n232 & ~new_n1292;
  assign new_n1329 = ~new_n1327 & ~new_n1328;
  assign new_n1330 = ~popsel3 & new_n1329;
  assign new_n1331 = ~new_n573 & ~new_n605;
  assign new_n1332 = new_n573 & new_n605;
  assign new_n1333 = ~new_n1331 & ~new_n1332;
  assign new_n1334 = new_n491 & ~new_n522;
  assign new_n1335 = ~new_n773 & new_n1334;
  assign new_n1336 = new_n768 & ~new_n773;
  assign new_n1337 = ~new_n1335 & ~new_n1336;
  assign new_n1338 = ~new_n775 & new_n1337;
  assign new_n1339 = ~new_n772 & ~new_n1338;
  assign new_n1340 = new_n558 & ~new_n589;
  assign new_n1341 = ~new_n1339 & ~new_n1340;
  assign new_n1342 = new_n1333 & new_n1341;
  assign new_n1343 = new_n771 & new_n1333;
  assign new_n1344 = ~new_n1342 & ~new_n1343;
  assign new_n1345 = ~new_n1334 & ~new_n1336;
  assign new_n1346 = ~new_n775 & new_n1345;
  assign new_n1347 = new_n772 & ~new_n775;
  assign new_n1348 = ~new_n1346 & ~new_n1347;
  assign new_n1349 = ~new_n771 & new_n1348;
  assign new_n1350 = ~new_n1340 & ~new_n1349;
  assign new_n1351 = new_n1344 & new_n1350;
  assign new_n1352 = new_n1333 & new_n1344;
  assign new_n1353 = ~new_n1351 & ~new_n1352;
  assign new_n1354 = new_n882 & new_n1353;
  assign new_n1355 = new_n232 & ~new_n1322;
  assign new_n1356 = ~new_n1354 & ~new_n1355;
  assign new_n1357 = new_n313 & ~new_n1356;
  assign po7 = new_n1330 | new_n1357;
  assign new_n1359 = ~new_n185 & ~new_n203;
  assign new_n1360 = new_n1285 & new_n1359;
  assign new_n1361 = new_n194 & new_n1360;
  assign new_n1362 = ~new_n194 & ~new_n1360;
  assign new_n1363 = ~new_n1361 & ~new_n1362;
  assign new_n1364 = popsel2 & ~new_n1363;
  assign new_n1365 = new_n232 & new_n1364;
  assign new_n1366 = ~popsel2 & new_n1363;
  assign new_n1367 = psh2 & ~new_n1192;
  assign new_n1368 = pmusel2 & pind6;
  assign new_n1369 = ~pinb6 & ~new_n1368;
  assign new_n1370 = new_n241 & ~new_n1368;
  assign new_n1371 = ~pmusel1 & ~pinb6;
  assign new_n1372 = ~new_n1369 & ~new_n1370;
  assign new_n1373 = ~new_n244 & ~new_n1371;
  assign new_n1374 = new_n1372 & new_n1373;
  assign new_n1375 = new_n236 & new_n1374;
  assign new_n1376 = ~pmusel3 & pind6;
  assign new_n1377 = new_n264 & new_n1376;
  assign new_n1378 = ~new_n1375 & ~new_n1377;
  assign new_n1379 = ~psh2 & ~new_n1378;
  assign new_n1380 = ~new_n1367 & ~new_n1379;
  assign new_n1381 = ~psh1 & new_n1380;
  assign new_n1382 = ~new_n1181 & ~new_n1246;
  assign new_n1383 = new_n1380 & new_n1382;
  assign new_n1384 = psh1 & new_n1382;
  assign new_n1385 = ~new_n1383 & ~new_n1384;
  assign new_n1386 = ~new_n1381 & new_n1385;
  assign new_n1387 = ~psh0 & new_n1386;
  assign new_n1388 = psh2 & ~new_n1378;
  assign new_n1389 = ~new_n1171 & ~new_n1388;
  assign new_n1390 = new_n1307 & new_n1389;
  assign new_n1391 = psh1 & new_n1389;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = ~new_n1308 & new_n1392;
  assign new_n1394 = psh0 & new_n1393;
  assign new_n1395 = ~new_n1387 & ~new_n1394;
  assign new_n1396 = new_n1363 & new_n1395;
  assign new_n1397 = popsel2 & new_n1395;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = ~new_n1366 & new_n1398;
  assign new_n1400 = ~new_n1365 & ~new_n1399;
  assign new_n1401 = new_n232 & ~new_n1365;
  assign new_n1402 = ~new_n1400 & ~new_n1401;
  assign new_n1403 = ~popsel3 & new_n1402;
  assign new_n1404 = ~new_n558 & ~new_n589;
  assign new_n1405 = new_n558 & new_n589;
  assign new_n1406 = ~new_n1404 & ~new_n1405;
  assign new_n1407 = ~new_n768 & ~new_n1334;
  assign new_n1408 = ~new_n773 & ~new_n1407;
  assign new_n1409 = ~new_n775 & ~new_n1408;
  assign new_n1410 = new_n1406 & new_n1409;
  assign new_n1411 = new_n772 & new_n1406;
  assign new_n1412 = ~new_n1410 & ~new_n1411;
  assign new_n1413 = new_n1406 & new_n1412;
  assign new_n1414 = ~new_n772 & ~new_n1345;
  assign new_n1415 = ~new_n775 & ~new_n1414;
  assign new_n1416 = new_n1412 & new_n1415;
  assign new_n1417 = ~new_n1413 & ~new_n1416;
  assign new_n1418 = new_n882 & new_n1417;
  assign new_n1419 = new_n232 & ~new_n1395;
  assign new_n1420 = ~new_n1418 & ~new_n1419;
  assign new_n1421 = new_n313 & ~new_n1420;
  assign po6 = new_n1403 | new_n1421;
  assign new_n1423 = ~new_n185 & new_n1285;
  assign new_n1424 = new_n203 & new_n1423;
  assign new_n1425 = ~new_n203 & ~new_n1423;
  assign new_n1426 = ~new_n1424 & ~new_n1425;
  assign new_n1427 = popsel2 & ~new_n1426;
  assign new_n1428 = new_n232 & new_n1427;
  assign new_n1429 = ~popsel2 & new_n1426;
  assign new_n1430 = pind5 & pmusel2;
  assign new_n1431 = ~pinb5 & ~new_n1430;
  assign new_n1432 = new_n241 & ~new_n1430;
  assign new_n1433 = ~pmusel1 & ~pinb5;
  assign new_n1434 = ~new_n1431 & ~new_n1432;
  assign new_n1435 = ~new_n244 & ~new_n1433;
  assign new_n1436 = new_n1434 & new_n1435;
  assign new_n1437 = new_n236 & new_n1436;
  assign new_n1438 = pind5 & ~pmusel3;
  assign new_n1439 = new_n264 & new_n1438;
  assign new_n1440 = ~new_n1437 & ~new_n1439;
  assign new_n1441 = ~psh2 & ~new_n1440;
  assign new_n1442 = ~new_n1197 & ~new_n1441;
  assign new_n1443 = ~psh1 & new_n1442;
  assign new_n1444 = ~new_n1159 & ~new_n1306;
  assign new_n1445 = new_n1442 & new_n1444;
  assign new_n1446 = psh1 & new_n1444;
  assign new_n1447 = ~new_n1445 & ~new_n1446;
  assign new_n1448 = ~new_n1443 & new_n1447;
  assign new_n1449 = ~psh0 & new_n1448;
  assign new_n1450 = psh2 & ~new_n1440;
  assign new_n1451 = ~new_n1246 & ~new_n1450;
  assign new_n1452 = new_n1380 & new_n1451;
  assign new_n1453 = psh1 & new_n1451;
  assign new_n1454 = ~new_n1452 & ~new_n1453;
  assign new_n1455 = ~new_n1381 & new_n1454;
  assign new_n1456 = psh0 & new_n1455;
  assign new_n1457 = ~new_n1449 & ~new_n1456;
  assign new_n1458 = new_n1426 & new_n1457;
  assign new_n1459 = popsel2 & new_n1457;
  assign new_n1460 = ~new_n1458 & ~new_n1459;
  assign new_n1461 = ~new_n1429 & new_n1460;
  assign new_n1462 = ~new_n1428 & ~new_n1461;
  assign new_n1463 = new_n232 & ~new_n1428;
  assign new_n1464 = ~new_n1462 & ~new_n1463;
  assign new_n1465 = ~popsel3 & new_n1464;
  assign new_n1466 = ~new_n506 & ~new_n538;
  assign new_n1467 = new_n506 & new_n538;
  assign new_n1468 = ~new_n1466 & ~new_n1467;
  assign new_n1469 = new_n1407 & new_n1468;
  assign new_n1470 = new_n773 & new_n1468;
  assign new_n1471 = ~new_n1469 & ~new_n1470;
  assign new_n1472 = new_n1468 & new_n1471;
  assign new_n1473 = new_n1345 & new_n1471;
  assign new_n1474 = ~new_n1472 & ~new_n1473;
  assign new_n1475 = new_n882 & new_n1474;
  assign new_n1476 = new_n232 & ~new_n1457;
  assign new_n1477 = ~new_n1475 & ~new_n1476;
  assign new_n1478 = new_n313 & ~new_n1477;
  assign po5 = new_n1465 | new_n1478;
  assign new_n1480 = new_n185 & new_n1285;
  assign new_n1481 = ~new_n185 & ~new_n1285;
  assign new_n1482 = ~new_n1480 & ~new_n1481;
  assign new_n1483 = popsel2 & ~new_n1482;
  assign new_n1484 = new_n232 & new_n1483;
  assign new_n1485 = ~popsel2 & new_n1482;
  assign new_n1486 = pmusel2 & pind4;
  assign new_n1487 = ~pinb4 & ~new_n1486;
  assign new_n1488 = new_n241 & ~new_n1486;
  assign new_n1489 = ~pmusel1 & ~pinb4;
  assign new_n1490 = ~new_n1487 & ~new_n1488;
  assign new_n1491 = ~new_n244 & ~new_n1489;
  assign new_n1492 = new_n1490 & new_n1491;
  assign new_n1493 = new_n236 & new_n1492;
  assign new_n1494 = pind4 & ~pmusel3;
  assign new_n1495 = new_n264 & new_n1494;
  assign new_n1496 = ~new_n1493 & ~new_n1495;
  assign new_n1497 = ~psh2 & ~new_n1496;
  assign new_n1498 = ~new_n1255 & ~new_n1497;
  assign new_n1499 = ~psh1 & new_n1498;
  assign new_n1500 = ~new_n1234 & ~new_n1379;
  assign new_n1501 = new_n1498 & new_n1500;
  assign new_n1502 = psh1 & new_n1500;
  assign new_n1503 = ~new_n1501 & ~new_n1502;
  assign new_n1504 = ~new_n1499 & new_n1503;
  assign new_n1505 = ~psh0 & new_n1504;
  assign new_n1506 = psh2 & ~new_n1496;
  assign new_n1507 = ~new_n1306 & ~new_n1506;
  assign new_n1508 = new_n1442 & new_n1507;
  assign new_n1509 = psh1 & new_n1507;
  assign new_n1510 = ~new_n1508 & ~new_n1509;
  assign new_n1511 = ~new_n1443 & new_n1510;
  assign new_n1512 = psh0 & new_n1511;
  assign new_n1513 = ~new_n1505 & ~new_n1512;
  assign new_n1514 = new_n1482 & new_n1513;
  assign new_n1515 = popsel2 & new_n1513;
  assign new_n1516 = ~new_n1514 & ~new_n1515;
  assign new_n1517 = ~new_n1485 & new_n1516;
  assign new_n1518 = ~new_n1484 & ~new_n1517;
  assign new_n1519 = new_n232 & ~new_n1484;
  assign new_n1520 = ~new_n1518 & ~new_n1519;
  assign new_n1521 = ~popsel3 & new_n1520;
  assign new_n1522 = new_n491 & new_n522;
  assign new_n1523 = ~new_n491 & ~new_n522;
  assign new_n1524 = ~new_n1522 & ~new_n1523;
  assign new_n1525 = new_n768 & ~new_n1524;
  assign new_n1526 = ~new_n768 & new_n1524;
  assign new_n1527 = ~new_n1525 & ~new_n1526;
  assign new_n1528 = ~new_n232 & new_n1527;
  assign new_n1529 = new_n316 & new_n1513;
  assign new_n1530 = new_n1513 & new_n1527;
  assign new_n1531 = ~new_n317 & ~new_n1528;
  assign new_n1532 = ~new_n1529 & ~new_n1530;
  assign new_n1533 = new_n1531 & new_n1532;
  assign new_n1534 = new_n313 & new_n1533;
  assign po4 = new_n1521 | new_n1534;
  assign new_n1536 = new_n104 & ~new_n125;
  assign new_n1537 = new_n135 & new_n1536;
  assign new_n1538 = new_n134 & new_n1537;
  assign new_n1539 = ~new_n134 & ~new_n1537;
  assign new_n1540 = ~new_n1538 & ~new_n1539;
  assign new_n1541 = popsel2 & ~new_n1540;
  assign new_n1542 = new_n232 & new_n1541;
  assign new_n1543 = ~popsel2 & new_n1540;
  assign new_n1544 = pind3 & pmusel2;
  assign new_n1545 = ~pinb3 & ~new_n1544;
  assign new_n1546 = new_n241 & ~new_n1544;
  assign new_n1547 = ~pmusel1 & ~pinb3;
  assign new_n1548 = ~new_n1545 & ~new_n1546;
  assign new_n1549 = ~new_n244 & ~new_n1547;
  assign new_n1550 = new_n1548 & new_n1549;
  assign new_n1551 = new_n236 & new_n1550;
  assign new_n1552 = pind3 & ~pmusel3;
  assign new_n1553 = new_n264 & new_n1552;
  assign new_n1554 = ~new_n1551 & ~new_n1553;
  assign new_n1555 = ~psh2 & ~new_n1554;
  assign new_n1556 = ~new_n1315 & ~new_n1555;
  assign new_n1557 = ~psh1 & new_n1556;
  assign new_n1558 = ~new_n1294 & ~new_n1441;
  assign new_n1559 = new_n1556 & new_n1558;
  assign new_n1560 = psh1 & new_n1558;
  assign new_n1561 = ~new_n1559 & ~new_n1560;
  assign new_n1562 = ~new_n1557 & new_n1561;
  assign new_n1563 = ~psh0 & new_n1562;
  assign new_n1564 = psh2 & ~new_n1554;
  assign new_n1565 = ~new_n1379 & ~new_n1564;
  assign new_n1566 = new_n1498 & new_n1565;
  assign new_n1567 = psh1 & new_n1565;
  assign new_n1568 = ~new_n1566 & ~new_n1567;
  assign new_n1569 = ~new_n1499 & new_n1568;
  assign new_n1570 = psh0 & new_n1569;
  assign new_n1571 = ~new_n1563 & ~new_n1570;
  assign new_n1572 = new_n1540 & new_n1571;
  assign new_n1573 = popsel2 & new_n1571;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = ~new_n1543 & new_n1574;
  assign new_n1576 = ~new_n1542 & ~new_n1575;
  assign new_n1577 = new_n232 & ~new_n1542;
  assign new_n1578 = ~new_n1576 & ~new_n1577;
  assign new_n1579 = ~popsel3 & new_n1578;
  assign new_n1580 = ~new_n626 & ~new_n641;
  assign new_n1581 = new_n626 & new_n641;
  assign new_n1582 = ~new_n1580 & ~new_n1581;
  assign new_n1583 = ~new_n719 & new_n734;
  assign new_n1584 = new_n766 & ~new_n1583;
  assign new_n1585 = ~new_n735 & ~new_n1584;
  assign new_n1586 = ~new_n737 & ~new_n1585;
  assign new_n1587 = ~new_n704 & ~new_n1586;
  assign new_n1588 = ~new_n657 & new_n672;
  assign new_n1589 = ~new_n1587 & ~new_n1588;
  assign new_n1590 = new_n1582 & new_n1589;
  assign new_n1591 = new_n673 & new_n1582;
  assign new_n1592 = ~new_n1590 & ~new_n1591;
  assign new_n1593 = new_n735 & ~new_n1583;
  assign new_n1594 = ~new_n1584 & ~new_n1593;
  assign new_n1595 = ~new_n704 & new_n1594;
  assign new_n1596 = ~new_n737 & ~new_n1595;
  assign new_n1597 = ~new_n673 & ~new_n1596;
  assign new_n1598 = ~new_n1588 & ~new_n1597;
  assign new_n1599 = new_n1592 & new_n1598;
  assign new_n1600 = new_n1582 & new_n1592;
  assign new_n1601 = ~new_n1599 & ~new_n1600;
  assign new_n1602 = new_n882 & new_n1601;
  assign new_n1603 = new_n232 & ~new_n1571;
  assign new_n1604 = ~new_n1602 & ~new_n1603;
  assign new_n1605 = new_n313 & ~new_n1604;
  assign po3 = new_n1579 | new_n1605;
  assign new_n1607 = ~new_n107 & ~new_n125;
  assign new_n1608 = new_n104 & new_n1607;
  assign new_n1609 = new_n116 & new_n1608;
  assign new_n1610 = ~new_n116 & ~new_n1608;
  assign new_n1611 = ~new_n1609 & ~new_n1610;
  assign new_n1612 = popsel2 & ~new_n1611;
  assign new_n1613 = new_n232 & new_n1612;
  assign new_n1614 = ~popsel2 & new_n1611;
  assign new_n1615 = pind2 & pmusel2;
  assign new_n1616 = ~pinb2 & ~new_n1615;
  assign new_n1617 = new_n241 & ~new_n1615;
  assign new_n1618 = ~pmusel1 & ~pinb2;
  assign new_n1619 = ~new_n1616 & ~new_n1617;
  assign new_n1620 = ~new_n244 & ~new_n1618;
  assign new_n1621 = new_n1619 & new_n1620;
  assign new_n1622 = new_n236 & new_n1621;
  assign new_n1623 = pind2 & ~pmusel3;
  assign new_n1624 = new_n264 & new_n1623;
  assign new_n1625 = ~new_n1622 & ~new_n1624;
  assign new_n1626 = ~psh2 & ~new_n1625;
  assign new_n1627 = ~new_n1388 & ~new_n1626;
  assign new_n1628 = ~psh1 & new_n1627;
  assign new_n1629 = ~new_n1367 & ~new_n1497;
  assign new_n1630 = new_n1627 & new_n1629;
  assign new_n1631 = psh1 & new_n1629;
  assign new_n1632 = ~new_n1630 & ~new_n1631;
  assign new_n1633 = ~new_n1628 & new_n1632;
  assign new_n1634 = ~psh0 & new_n1633;
  assign new_n1635 = psh2 & ~new_n1625;
  assign new_n1636 = ~new_n1441 & ~new_n1635;
  assign new_n1637 = new_n1556 & new_n1636;
  assign new_n1638 = psh1 & new_n1636;
  assign new_n1639 = ~new_n1637 & ~new_n1638;
  assign new_n1640 = ~new_n1557 & new_n1639;
  assign new_n1641 = psh0 & new_n1640;
  assign new_n1642 = ~new_n1634 & ~new_n1641;
  assign new_n1643 = new_n1611 & new_n1642;
  assign new_n1644 = popsel2 & new_n1642;
  assign new_n1645 = ~new_n1643 & ~new_n1644;
  assign new_n1646 = ~new_n1614 & new_n1645;
  assign new_n1647 = ~new_n1613 & ~new_n1646;
  assign new_n1648 = new_n232 & ~new_n1613;
  assign new_n1649 = ~new_n1647 & ~new_n1648;
  assign new_n1650 = ~popsel3 & new_n1649;
  assign new_n1651 = ~new_n657 & ~new_n672;
  assign new_n1652 = new_n657 & new_n672;
  assign new_n1653 = ~new_n1651 & ~new_n1652;
  assign new_n1654 = new_n1586 & new_n1653;
  assign new_n1655 = new_n704 & new_n1653;
  assign new_n1656 = ~new_n1654 & ~new_n1655;
  assign new_n1657 = new_n1653 & new_n1656;
  assign new_n1658 = new_n1596 & new_n1656;
  assign new_n1659 = ~new_n1657 & ~new_n1658;
  assign new_n1660 = new_n882 & new_n1659;
  assign new_n1661 = new_n232 & ~new_n1642;
  assign new_n1662 = ~new_n1660 & ~new_n1661;
  assign new_n1663 = new_n313 & ~new_n1662;
  assign po2 = new_n1650 | new_n1663;
  assign new_n1665 = new_n104 & ~new_n107;
  assign new_n1666 = new_n125 & new_n1665;
  assign new_n1667 = ~new_n125 & ~new_n1665;
  assign new_n1668 = ~new_n1666 & ~new_n1667;
  assign new_n1669 = popsel2 & ~new_n1668;
  assign new_n1670 = new_n232 & new_n1669;
  assign new_n1671 = ~popsel2 & new_n1668;
  assign new_n1672 = pmusel2 & pind1;
  assign new_n1673 = ~pinb1 & ~new_n1672;
  assign new_n1674 = new_n241 & ~new_n1672;
  assign new_n1675 = ~pinb1 & ~pmusel1;
  assign new_n1676 = ~new_n1673 & ~new_n1674;
  assign new_n1677 = ~new_n244 & ~new_n1675;
  assign new_n1678 = new_n1676 & new_n1677;
  assign new_n1679 = new_n236 & new_n1678;
  assign new_n1680 = ~pmusel3 & pind1;
  assign new_n1681 = new_n264 & new_n1680;
  assign new_n1682 = ~new_n1679 & ~new_n1681;
  assign new_n1683 = ~psh2 & ~new_n1682;
  assign new_n1684 = ~new_n1450 & ~new_n1683;
  assign new_n1685 = ~psh1 & new_n1684;
  assign new_n1686 = ~new_n1197 & ~new_n1555;
  assign new_n1687 = new_n1684 & new_n1686;
  assign new_n1688 = psh1 & new_n1686;
  assign new_n1689 = ~new_n1687 & ~new_n1688;
  assign new_n1690 = ~new_n1685 & new_n1689;
  assign new_n1691 = ~psh0 & new_n1690;
  assign new_n1692 = psh2 & ~new_n1682;
  assign new_n1693 = ~new_n1497 & ~new_n1692;
  assign new_n1694 = new_n1627 & new_n1693;
  assign new_n1695 = psh1 & new_n1693;
  assign new_n1696 = ~new_n1694 & ~new_n1695;
  assign new_n1697 = ~new_n1628 & new_n1696;
  assign new_n1698 = psh0 & new_n1697;
  assign new_n1699 = ~new_n1691 & ~new_n1698;
  assign new_n1700 = new_n1668 & new_n1699;
  assign new_n1701 = popsel2 & new_n1699;
  assign new_n1702 = ~new_n1700 & ~new_n1701;
  assign new_n1703 = ~new_n1671 & new_n1702;
  assign new_n1704 = ~new_n1670 & ~new_n1703;
  assign new_n1705 = new_n232 & ~new_n1670;
  assign new_n1706 = ~new_n1704 & ~new_n1705;
  assign new_n1707 = ~popsel3 & new_n1706;
  assign new_n1708 = ~new_n688 & ~new_n703;
  assign new_n1709 = new_n688 & new_n703;
  assign new_n1710 = ~new_n1708 & ~new_n1709;
  assign new_n1711 = new_n1584 & new_n1710;
  assign new_n1712 = new_n735 & new_n1710;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = new_n1710 & new_n1713;
  assign new_n1715 = ~new_n735 & ~new_n766;
  assign new_n1716 = ~new_n1583 & ~new_n1715;
  assign new_n1717 = new_n1713 & new_n1716;
  assign new_n1718 = ~new_n1714 & ~new_n1717;
  assign new_n1719 = new_n882 & new_n1718;
  assign new_n1720 = new_n232 & ~new_n1699;
  assign new_n1721 = ~new_n1719 & ~new_n1720;
  assign new_n1722 = new_n313 & ~new_n1721;
  assign po1 = new_n1707 | new_n1722;
  assign new_n1724 = new_n104 & new_n107;
  assign new_n1725 = ~new_n104 & ~new_n107;
  assign new_n1726 = ~new_n1724 & ~new_n1725;
  assign new_n1727 = popsel2 & ~new_n1726;
  assign new_n1728 = new_n232 & new_n1727;
  assign new_n1729 = ~popsel2 & new_n1726;
  assign new_n1730 = pmusel2 & pind0;
  assign new_n1731 = ~pinb0 & ~new_n1730;
  assign new_n1732 = new_n241 & ~new_n1730;
  assign new_n1733 = ~pinb0 & ~pmusel1;
  assign new_n1734 = ~new_n1731 & ~new_n1732;
  assign new_n1735 = ~new_n244 & ~new_n1733;
  assign new_n1736 = new_n1734 & new_n1735;
  assign new_n1737 = new_n236 & new_n1736;
  assign new_n1738 = ~pmusel3 & pind0;
  assign new_n1739 = new_n264 & new_n1738;
  assign new_n1740 = ~new_n1737 & ~new_n1739;
  assign new_n1741 = ~psh2 & ~new_n1740;
  assign new_n1742 = ~new_n1506 & ~new_n1741;
  assign new_n1743 = ~psh1 & new_n1742;
  assign new_n1744 = ~new_n1255 & ~new_n1626;
  assign new_n1745 = new_n1742 & new_n1744;
  assign new_n1746 = psh1 & new_n1744;
  assign new_n1747 = ~new_n1745 & ~new_n1746;
  assign new_n1748 = ~new_n1743 & new_n1747;
  assign new_n1749 = ~psh0 & new_n1748;
  assign new_n1750 = psh2 & ~new_n1740;
  assign new_n1751 = ~new_n1555 & ~new_n1750;
  assign new_n1752 = new_n1684 & new_n1751;
  assign new_n1753 = psh1 & new_n1751;
  assign new_n1754 = ~new_n1752 & ~new_n1753;
  assign new_n1755 = ~new_n1685 & new_n1754;
  assign new_n1756 = psh0 & new_n1755;
  assign new_n1757 = ~new_n1749 & ~new_n1756;
  assign new_n1758 = new_n1726 & new_n1757;
  assign new_n1759 = popsel2 & new_n1757;
  assign new_n1760 = ~new_n1758 & ~new_n1759;
  assign new_n1761 = ~new_n1729 & new_n1760;
  assign new_n1762 = ~new_n1728 & ~new_n1761;
  assign new_n1763 = new_n232 & ~new_n1728;
  assign new_n1764 = ~new_n1762 & ~new_n1763;
  assign new_n1765 = ~popsel3 & new_n1764;
  assign new_n1766 = new_n719 & new_n734;
  assign new_n1767 = ~new_n719 & ~new_n734;
  assign new_n1768 = ~new_n1766 & ~new_n1767;
  assign new_n1769 = new_n766 & new_n1768;
  assign new_n1770 = new_n1768 & ~new_n1769;
  assign new_n1771 = new_n766 & ~new_n1769;
  assign new_n1772 = ~new_n1770 & ~new_n1771;
  assign new_n1773 = new_n882 & new_n1772;
  assign new_n1774 = new_n232 & ~new_n1757;
  assign new_n1775 = ~new_n1773 & ~new_n1774;
  assign new_n1776 = new_n313 & ~new_n1775;
  assign po0 = new_n1765 | new_n1776;
  assign new_n1778 = ~new_n146 & ~new_n164;
  assign new_n1779 = new_n217 & new_n1778;
  assign new_n1780 = new_n155 & new_n1779;
  assign new_n1781 = ~new_n155 & ~new_n1779;
  assign new_n1782 = ~new_n1780 & ~new_n1781;
  assign new_n1783 = popsel2 & ~new_n1782;
  assign new_n1784 = new_n232 & new_n1783;
  assign new_n1785 = ~popsel2 & new_n1782;
  assign new_n1786 = ~new_n864 & ~new_n1196;
  assign new_n1787 = new_n1194 & new_n1786;
  assign new_n1788 = psh1 & new_n1786;
  assign new_n1789 = ~new_n1787 & ~new_n1788;
  assign new_n1790 = ~new_n1195 & new_n1789;
  assign new_n1791 = ~psh0 & new_n1790;
  assign new_n1792 = ~psh1 & new_n1175;
  assign new_n1793 = ~psh2 & ~new_n266;
  assign new_n1794 = ~new_n1367 & ~new_n1793;
  assign new_n1795 = new_n1175 & new_n1794;
  assign new_n1796 = psh1 & new_n1794;
  assign new_n1797 = ~new_n1795 & ~new_n1796;
  assign new_n1798 = ~new_n1792 & new_n1797;
  assign new_n1799 = psh0 & new_n1798;
  assign new_n1800 = ~new_n1791 & ~new_n1799;
  assign new_n1801 = new_n1782 & new_n1800;
  assign new_n1802 = popsel2 & new_n1800;
  assign new_n1803 = ~new_n1801 & ~new_n1802;
  assign new_n1804 = ~new_n1785 & new_n1803;
  assign new_n1805 = ~new_n1784 & ~new_n1804;
  assign new_n1806 = new_n232 & ~new_n1784;
  assign new_n1807 = ~new_n1805 & ~new_n1806;
  assign new_n1808 = ~popsel3 & new_n1807;
  assign new_n1809 = ~new_n348 & ~new_n369;
  assign new_n1810 = new_n348 & new_n369;
  assign new_n1811 = ~new_n1809 & ~new_n1810;
  assign new_n1812 = ~new_n432 & ~new_n1216;
  assign new_n1813 = ~new_n890 & ~new_n1812;
  assign new_n1814 = new_n1811 & new_n1813;
  assign new_n1815 = new_n401 & new_n1811;
  assign new_n1816 = ~new_n1814 & ~new_n1815;
  assign new_n1817 = new_n1811 & new_n1816;
  assign new_n1818 = ~new_n401 & ~new_n897;
  assign new_n1819 = ~new_n890 & ~new_n1818;
  assign new_n1820 = new_n1816 & new_n1819;
  assign new_n1821 = ~new_n1817 & ~new_n1820;
  assign new_n1822 = new_n882 & new_n1821;
  assign new_n1823 = new_n232 & ~new_n1800;
  assign new_n1824 = ~new_n1822 & ~new_n1823;
  assign new_n1825 = new_n313 & ~new_n1824;
  assign po10 = new_n1808 | new_n1825;
endmodule


