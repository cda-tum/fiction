// Benchmark "b20" written by ABC on Wed Sep  5 10:17:23 2018

module b20 ( clock, 
    SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_,
    SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_,
    SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_,
    SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123  );
  input  clock;
  input  SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_,
    SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_,
    SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_,
    SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123;
  reg P1_IR_REG_0_, P1_IR_REG_1_, P1_IR_REG_2_, P1_IR_REG_3_, P1_IR_REG_4_,
    P1_IR_REG_5_, P1_IR_REG_6_, P1_IR_REG_7_, P1_IR_REG_8_, P1_IR_REG_9_,
    P1_IR_REG_10_, P1_IR_REG_11_, P1_IR_REG_12_, P1_IR_REG_13_,
    P1_IR_REG_14_, P1_IR_REG_15_, P1_IR_REG_16_, P1_IR_REG_17_,
    P1_IR_REG_18_, P1_IR_REG_19_, P1_IR_REG_20_, P1_IR_REG_21_,
    P1_IR_REG_22_, P1_IR_REG_23_, P1_IR_REG_24_, P1_IR_REG_25_,
    P1_IR_REG_26_, P1_IR_REG_27_, P1_IR_REG_28_, P1_IR_REG_29_,
    P1_IR_REG_30_, P1_IR_REG_31_, P1_D_REG_0_, P1_D_REG_1_, P1_D_REG_2_,
    P1_D_REG_3_, P1_D_REG_4_, P1_D_REG_5_, P1_D_REG_6_, P1_D_REG_7_,
    P1_D_REG_8_, P1_D_REG_9_, P1_D_REG_10_, P1_D_REG_11_, P1_D_REG_12_,
    P1_D_REG_13_, P1_D_REG_14_, P1_D_REG_15_, P1_D_REG_16_, P1_D_REG_17_,
    P1_D_REG_18_, P1_D_REG_19_, P1_D_REG_20_, P1_D_REG_21_, P1_D_REG_22_,
    P1_D_REG_23_, P1_D_REG_24_, P1_D_REG_25_, P1_D_REG_26_, P1_D_REG_27_,
    P1_D_REG_28_, P1_D_REG_29_, P1_D_REG_30_, P1_D_REG_31_, P1_REG0_REG_0_,
    P1_REG0_REG_1_, P1_REG0_REG_2_, P1_REG0_REG_3_, P1_REG0_REG_4_,
    P1_REG0_REG_5_, P1_REG0_REG_6_, P1_REG0_REG_7_, P1_REG0_REG_8_,
    P1_REG0_REG_9_, P1_REG0_REG_10_, P1_REG0_REG_11_, P1_REG0_REG_12_,
    P1_REG0_REG_13_, P1_REG0_REG_14_, P1_REG0_REG_15_, P1_REG0_REG_16_,
    P1_REG0_REG_17_, P1_REG0_REG_18_, P1_REG0_REG_19_, P1_REG0_REG_20_,
    P1_REG0_REG_21_, P1_REG0_REG_22_, P1_REG0_REG_23_, P1_REG0_REG_24_,
    P1_REG0_REG_25_, P1_REG0_REG_26_, P1_REG0_REG_27_, P1_REG0_REG_28_,
    P1_REG0_REG_29_, P1_REG0_REG_30_, P1_REG0_REG_31_, P1_REG1_REG_0_,
    P1_REG1_REG_1_, P1_REG1_REG_2_, P1_REG1_REG_3_, P1_REG1_REG_4_,
    P1_REG1_REG_5_, P1_REG1_REG_6_, P1_REG1_REG_7_, P1_REG1_REG_8_,
    P1_REG1_REG_9_, P1_REG1_REG_10_, P1_REG1_REG_11_, P1_REG1_REG_12_,
    P1_REG1_REG_13_, P1_REG1_REG_14_, P1_REG1_REG_15_, P1_REG1_REG_16_,
    P1_REG1_REG_17_, P1_REG1_REG_18_, P1_REG1_REG_19_, P1_REG1_REG_20_,
    P1_REG1_REG_21_, P1_REG1_REG_22_, P1_REG1_REG_23_, P1_REG1_REG_24_,
    P1_REG1_REG_25_, P1_REG1_REG_26_, P1_REG1_REG_27_, P1_REG1_REG_28_,
    P1_REG1_REG_29_, P1_REG1_REG_30_, P1_REG1_REG_31_, P1_REG2_REG_0_,
    P1_REG2_REG_1_, P1_REG2_REG_2_, P1_REG2_REG_3_, P1_REG2_REG_4_,
    P1_REG2_REG_5_, P1_REG2_REG_6_, P1_REG2_REG_7_, P1_REG2_REG_8_,
    P1_REG2_REG_9_, P1_REG2_REG_10_, P1_REG2_REG_11_, P1_REG2_REG_12_,
    P1_REG2_REG_13_, P1_REG2_REG_14_, P1_REG2_REG_15_, P1_REG2_REG_16_,
    P1_REG2_REG_17_, P1_REG2_REG_18_, P1_REG2_REG_19_, P1_REG2_REG_20_,
    P1_REG2_REG_21_, P1_REG2_REG_22_, P1_REG2_REG_23_, P1_REG2_REG_24_,
    P1_REG2_REG_25_, P1_REG2_REG_26_, P1_REG2_REG_27_, P1_REG2_REG_28_,
    P1_REG2_REG_29_, P1_REG2_REG_30_, P1_REG2_REG_31_, P1_ADDR_REG_19_,
    P1_ADDR_REG_18_, P1_ADDR_REG_17_, P1_ADDR_REG_16_, P1_ADDR_REG_15_,
    P1_ADDR_REG_14_, P1_ADDR_REG_13_, P1_ADDR_REG_12_, P1_ADDR_REG_11_,
    P1_ADDR_REG_10_, P1_ADDR_REG_9_, P1_ADDR_REG_8_, P1_ADDR_REG_7_,
    P1_ADDR_REG_6_, P1_ADDR_REG_5_, P1_ADDR_REG_4_, P1_ADDR_REG_3_,
    P1_ADDR_REG_2_, P1_ADDR_REG_1_, P1_ADDR_REG_0_, P1_DATAO_REG_0_,
    P1_DATAO_REG_1_, P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_,
    P1_DATAO_REG_5_, P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_,
    P1_DATAO_REG_9_, P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_,
    P1_DATAO_REG_13_, P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_,
    P1_DATAO_REG_17_, P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_,
    P1_DATAO_REG_21_, P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_,
    P1_DATAO_REG_25_, P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_,
    P1_DATAO_REG_29_, P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_B_REG,
    P1_REG3_REG_15_, P1_REG3_REG_26_, P1_REG3_REG_6_, P1_REG3_REG_18_,
    P1_REG3_REG_2_, P1_REG3_REG_11_, P1_REG3_REG_22_, P1_REG3_REG_13_,
    P1_REG3_REG_20_, P1_REG3_REG_0_, P1_REG3_REG_9_, P1_REG3_REG_4_,
    P1_REG3_REG_24_, P1_REG3_REG_17_, P1_REG3_REG_5_, P1_REG3_REG_16_,
    P1_REG3_REG_25_, P1_REG3_REG_12_, P1_REG3_REG_21_, P1_REG3_REG_1_,
    P1_REG3_REG_8_, P1_REG3_REG_28_, P1_REG3_REG_19_, P1_REG3_REG_3_,
    P1_REG3_REG_10_, P1_REG3_REG_23_, P1_REG3_REG_14_, P1_REG3_REG_27_,
    P1_REG3_REG_7_, P1_STATE_REG, P1_RD_REG, P1_WR_REG, P2_IR_REG_0_,
    P2_IR_REG_1_, P2_IR_REG_2_, P2_IR_REG_3_, P2_IR_REG_4_, P2_IR_REG_5_,
    P2_IR_REG_6_, P2_IR_REG_7_, P2_IR_REG_8_, P2_IR_REG_9_, P2_IR_REG_10_,
    P2_IR_REG_11_, P2_IR_REG_12_, P2_IR_REG_13_, P2_IR_REG_14_,
    P2_IR_REG_15_, P2_IR_REG_16_, P2_IR_REG_17_, P2_IR_REG_18_,
    P2_IR_REG_19_, P2_IR_REG_20_, P2_IR_REG_21_, P2_IR_REG_22_,
    P2_IR_REG_23_, P2_IR_REG_24_, P2_IR_REG_25_, P2_IR_REG_26_,
    P2_IR_REG_27_, P2_IR_REG_28_, P2_IR_REG_29_, P2_IR_REG_30_,
    P2_IR_REG_31_, P2_D_REG_0_, P2_D_REG_1_, P2_D_REG_2_, P2_D_REG_3_,
    P2_D_REG_4_, P2_D_REG_5_, P2_D_REG_6_, P2_D_REG_7_, P2_D_REG_8_,
    P2_D_REG_9_, P2_D_REG_10_, P2_D_REG_11_, P2_D_REG_12_, P2_D_REG_13_,
    P2_D_REG_14_, P2_D_REG_15_, P2_D_REG_16_, P2_D_REG_17_, P2_D_REG_18_,
    P2_D_REG_19_, P2_D_REG_20_, P2_D_REG_21_, P2_D_REG_22_, P2_D_REG_23_,
    P2_D_REG_24_, P2_D_REG_25_, P2_D_REG_26_, P2_D_REG_27_, P2_D_REG_28_,
    P2_D_REG_29_, P2_D_REG_30_, P2_D_REG_31_, P2_REG0_REG_0_,
    P2_REG0_REG_1_, P2_REG0_REG_2_, P2_REG0_REG_3_, P2_REG0_REG_4_,
    P2_REG0_REG_5_, P2_REG0_REG_6_, P2_REG0_REG_7_, P2_REG0_REG_8_,
    P2_REG0_REG_9_, P2_REG0_REG_10_, P2_REG0_REG_11_, P2_REG0_REG_12_,
    P2_REG0_REG_13_, P2_REG0_REG_14_, P2_REG0_REG_15_, P2_REG0_REG_16_,
    P2_REG0_REG_17_, P2_REG0_REG_18_, P2_REG0_REG_19_, P2_REG0_REG_20_,
    P2_REG0_REG_21_, P2_REG0_REG_22_, P2_REG0_REG_23_, P2_REG0_REG_24_,
    P2_REG0_REG_25_, P2_REG0_REG_26_, P2_REG0_REG_27_, P2_REG0_REG_28_,
    P2_REG0_REG_29_, P2_REG0_REG_30_, P2_REG0_REG_31_, P2_REG1_REG_0_,
    P2_REG1_REG_1_, P2_REG1_REG_2_, P2_REG1_REG_3_, P2_REG1_REG_4_,
    P2_REG1_REG_5_, P2_REG1_REG_6_, P2_REG1_REG_7_, P2_REG1_REG_8_,
    P2_REG1_REG_9_, P2_REG1_REG_10_, P2_REG1_REG_11_, P2_REG1_REG_12_,
    P2_REG1_REG_13_, P2_REG1_REG_14_, P2_REG1_REG_15_, P2_REG1_REG_16_,
    P2_REG1_REG_17_, P2_REG1_REG_18_, P2_REG1_REG_19_, P2_REG1_REG_20_,
    P2_REG1_REG_21_, P2_REG1_REG_22_, P2_REG1_REG_23_, P2_REG1_REG_24_,
    P2_REG1_REG_25_, P2_REG1_REG_26_, P2_REG1_REG_27_, P2_REG1_REG_28_,
    P2_REG1_REG_29_, P2_REG1_REG_30_, P2_REG1_REG_31_, P2_REG2_REG_0_,
    P2_REG2_REG_1_, P2_REG2_REG_2_, P2_REG2_REG_3_, P2_REG2_REG_4_,
    P2_REG2_REG_5_, P2_REG2_REG_6_, P2_REG2_REG_7_, P2_REG2_REG_8_,
    P2_REG2_REG_9_, P2_REG2_REG_10_, P2_REG2_REG_11_, P2_REG2_REG_12_,
    P2_REG2_REG_13_, P2_REG2_REG_14_, P2_REG2_REG_15_, P2_REG2_REG_16_,
    P2_REG2_REG_17_, P2_REG2_REG_18_, P2_REG2_REG_19_, P2_REG2_REG_20_,
    P2_REG2_REG_21_, P2_REG2_REG_22_, P2_REG2_REG_23_, P2_REG2_REG_24_,
    P2_REG2_REG_25_, P2_REG2_REG_26_, P2_REG2_REG_27_, P2_REG2_REG_28_,
    P2_REG2_REG_29_, P2_REG2_REG_30_, P2_REG2_REG_31_, P2_ADDR_REG_19_,
    P2_ADDR_REG_18_, P2_ADDR_REG_17_, P2_ADDR_REG_16_, P2_ADDR_REG_15_,
    P2_ADDR_REG_14_, P2_ADDR_REG_13_, P2_ADDR_REG_12_, P2_ADDR_REG_11_,
    P2_ADDR_REG_10_, P2_ADDR_REG_9_, P2_ADDR_REG_8_, P2_ADDR_REG_7_,
    P2_ADDR_REG_6_, P2_ADDR_REG_5_, P2_ADDR_REG_4_, P2_ADDR_REG_3_,
    P2_ADDR_REG_2_, P2_ADDR_REG_1_, P2_ADDR_REG_0_, P2_DATAO_REG_0_,
    P2_DATAO_REG_1_, P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_,
    P2_DATAO_REG_5_, P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_,
    P2_DATAO_REG_9_, P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_,
    P2_DATAO_REG_13_, P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_,
    P2_DATAO_REG_17_, P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_,
    P2_DATAO_REG_21_, P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_,
    P2_DATAO_REG_25_, P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_,
    P2_DATAO_REG_29_, P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_B_REG,
    P2_REG3_REG_15_, P2_REG3_REG_26_, P2_REG3_REG_6_, P2_REG3_REG_18_,
    P2_REG3_REG_2_, P2_REG3_REG_11_, P2_REG3_REG_22_, P2_REG3_REG_13_,
    P2_REG3_REG_20_, P2_REG3_REG_0_, P2_REG3_REG_9_, P2_REG3_REG_4_,
    P2_REG3_REG_24_, P2_REG3_REG_17_, P2_REG3_REG_5_, P2_REG3_REG_16_,
    P2_REG3_REG_25_, P2_REG3_REG_12_, P2_REG3_REG_21_, P2_REG3_REG_1_,
    P2_REG3_REG_8_, P2_REG3_REG_28_, P2_REG3_REG_19_, P2_REG3_REG_3_,
    P2_REG3_REG_10_, P2_REG3_REG_23_, P2_REG3_REG_14_, P2_REG3_REG_27_,
    P2_REG3_REG_7_, P2_STATE_REG, P2_RD_REG, P2_WR_REG;
  wire n1525_1, n1526, n1527, n1528, n1529, n1530_1, n1531, n1532, n1533,
    n1534, n1535_1, n1536, n1537, n1538, n1539, n1540_1, n1541, n1542,
    n1543, n1544, n1545_1, n1546, n1547, n1548, n1549, n1550_1, n1551,
    n1552, n1553, n1554, n1555_1, n1556, n1557, n1558, n1559, n1560_1,
    n1561, n1562, n1563, n1564, n1565_1, n1566, n1567, n1568, n1569,
    n1570_1, n1571, n1572, n1573, n1574, n1575_1, n1576, n1577, n1578,
    n1579, n1580_1, n1581, n1582, n1583, n1584, n1585_1, n1586, n1587,
    n1588, n1589, n1590_1, n1591, n1592, n1593, n1594, n1595_1, n1596,
    n1597, n1598, n1599, n1600_1, n1601, n1602, n1603, n1604, n1606, n1607,
    n1608, n1609, n1610_1, n1612, n1613, n1614, n1615_1, n1616, n1618,
    n1619, n1620_1, n1621, n1622, n1624, n1625_1, n1626, n1627, n1628,
    n1630_1, n1631, n1632, n1633, n1634, n1636, n1637, n1638, n1639,
    n1640_1, n1642, n1643, n1644, n1645_1, n1646, n1648, n1649, n1650_1,
    n1651, n1652, n1654, n1655_1, n1656, n1657, n1658, n1660_1, n1661,
    n1662, n1663, n1664, n1666, n1667, n1668, n1669, n1670_1, n1672, n1673,
    n1674, n1675_1, n1676, n1678, n1679, n1680_1, n1681, n1682, n1684,
    n1685_1, n1686, n1687, n1688, n1690_1, n1691, n1692, n1693, n1694,
    n1696, n1697, n1698, n1699, n1700_1, n1702, n1703, n1704, n1705_1,
    n1706, n1708, n1709, n1710_1, n1711, n1712, n1713, n1714, n1715_1,
    n1717, n1718, n1720_1, n1721, n1723, n1724, n1726, n1727, n1728, n1729,
    n1730_1, n1731, n1732, n1733, n1734, n1735_1, n1736, n1737, n1738,
    n1739, n1740_1, n1741, n1742, n1743, n1744, n1745_1, n1747, n1748,
    n1749, n1750_1, n1751, n1752, n1753, n1754, n1755_1, n1756, n1757,
    n1758, n1759, n1760_1, n1761, n1762, n1763, n1764, n1765_1, n1766,
    n1767, n1768, n1769, n1770_1, n1771, n1773, n1774, n1775_1, n1776,
    n1777, n1778, n1779, n1780_1, n1781, n1782, n1783, n1784, n1785_1,
    n1786, n1787, n1788, n1789, n1790_1, n1791, n1792, n1793, n1794,
    n1795_1, n1796, n1798, n1799, n1800_1, n1801, n1802, n1803, n1804,
    n1805_1, n1806, n1807, n1808, n1809, n1810_1, n1811, n1812, n1813,
    n1814, n1815_1, n1816, n1817, n1818, n1819, n1820_1, n1822, n1823,
    n1824, n1825_1, n1826, n1827, n1828, n1829, n1830_1, n1831, n1832,
    n1833, n1834, n1835_1, n1836, n1837, n1838, n1839, n1840_1, n1841,
    n1842, n1843, n1844, n1845_1, n1846, n1847, n1848, n1850_1, n1851,
    n1852, n1853, n1854, n1855_1, n1856, n1857, n1858, n1859, n1860_1,
    n1861, n1862, n1863, n1864, n1865_1, n1866, n1867, n1868, n1869,
    n1870_1, n1871, n1872, n1874, n1875_1, n1876, n1877, n1878, n1879,
    n1880_1, n1881, n1882, n1883, n1884, n1885_1, n1886, n1887, n1888,
    n1889, n1890_1, n1891, n1892, n1893, n1894, n1895_1, n1896, n1897,
    n1898, n1899, n1900_1, n1902, n1903, n1904, n1905_1, n1906, n1907,
    n1908, n1909, n1910_1, n1911, n1912, n1913, n1914, n1915_1, n1916,
    n1917, n1918, n1919, n1920_1, n1921, n1922, n1923, n1924, n1925_1,
    n1926, n1927, n1929, n1930_1, n1931, n1932, n1933, n1934, n1935_1,
    n1936, n1937, n1938, n1939, n1940_1, n1941, n1942, n1943, n1944,
    n1945_1, n1946, n1947, n1948, n1949, n1950_1, n1951, n1952, n1953,
    n1954, n1955_1, n1957, n1958, n1959, n1960_1, n1961, n1962, n1963,
    n1964, n1965_1, n1966, n1967, n1968, n1969, n1970_1, n1971, n1972,
    n1973, n1974, n1975_1, n1976, n1977, n1978, n1979, n1980_1, n1981,
    n1982, n1984, n1985_1, n1986, n1987, n1988, n1989, n1990_1, n1991,
    n1992, n1993, n1994, n1995_1, n1996, n1997, n1998, n1999, n2000_1,
    n2001, n2002, n2003, n2004, n2005_1, n2006, n2007, n2008, n2009,
    n2010_1, n2012, n2013, n2014, n2015_1, n2016, n2017, n2018, n2019,
    n2020_1, n2021, n2022, n2023, n2024, n2025_1, n2026, n2027, n2028,
    n2029, n2030_1, n2031, n2032, n2033, n2034, n2035_1, n2036, n2037,
    n2039, n2040_1, n2041, n2042, n2043, n2044, n2045_1, n2046, n2047,
    n2048, n2049, n2050_1, n2051, n2052, n2053, n2054, n2055_1, n2056,
    n2057, n2058, n2059, n2060_1, n2061, n2062, n2063, n2064, n2066, n2067,
    n2068, n2069, n2070_1, n2071, n2072, n2073, n2074, n2075_1, n2076,
    n2077, n2078, n2079, n2080_1, n2081, n2082, n2083, n2084, n2085_1,
    n2086, n2087, n2088, n2089, n2090_1, n2091, n2093, n2094, n2095_1,
    n2096, n2097, n2098, n2099, n2100_1, n2101, n2102, n2103, n2104,
    n2105_1, n2106, n2107, n2108, n2109, n2110_1, n2111, n2112, n2113,
    n2114, n2115_1, n2116, n2117, n2118, n2119, n2121, n2122, n2123, n2124,
    n2125_1, n2126, n2127, n2128, n2129, n2130_1, n2131, n2132, n2133,
    n2134, n2135_1, n2136, n2137, n2138, n2139, n2140_1, n2141, n2142,
    n2143, n2144, n2145_1, n2146, n2148, n2149, n2150_1, n2151, n2152,
    n2153, n2154, n2155_1, n2156, n2157, n2158, n2159, n2160_1, n2161,
    n2162, n2163, n2164, n2165_1, n2166, n2167, n2168, n2169, n2170_1,
    n2171, n2172, n2173, n2174, n2175_1, n2176, n2177, n2178, n2179,
    n2180_1, n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189,
    n2190_1, n2191, n2192, n2193, n2194, n2195_1, n2196, n2197, n2198,
    n2199, n2200_1, n2201, n2202, n2203, n2204, n2205_1, n2206, n2207,
    n2208, n2210_1, n2211, n2212, n2213, n2214, n2215_1, n2216, n2217,
    n2218, n2219, n2220_1, n2221, n2222, n2223, n2224, n2225_1, n2226,
    n2227, n2228, n2229, n2230_1, n2231, n2232, n2233, n2234, n2235_1,
    n2236, n2237, n2238, n2239, n2240_1, n2241, n2242, n2244, n2245_1,
    n2246, n2247, n2248, n2249, n2250_1, n2251, n2252, n2253, n2254,
    n2255_1, n2256, n2257, n2258, n2259, n2260_1, n2261, n2262, n2263,
    n2264, n2265_1, n2266, n2267, n2268, n2269, n2270_1, n2271, n2272,
    n2273, n2274, n2275_1, n2276, n2277, n2278, n2279, n2281, n2282, n2283,
    n2284, n2285_1, n2286, n2287, n2288, n2289, n2290_1, n2291, n2292,
    n2293, n2294, n2295_1, n2296, n2297, n2298, n2299, n2300_1, n2301,
    n2302, n2303, n2304, n2305_1, n2306, n2307, n2308, n2309, n2310_1,
    n2311, n2312, n2313, n2314, n2315_1, n2316, n2318, n2319, n2320_1,
    n2321, n2322, n2323, n2324, n2325_1, n2326, n2327, n2328, n2329,
    n2330_1, n2331, n2332, n2333, n2334, n2335_1, n2336, n2337, n2338,
    n2339, n2340_1, n2342, n2343, n2344, n2345_1, n2346, n2347, n2348,
    n2349, n2350_1, n2351, n2352, n2353, n2354, n2355_1, n2356, n2357,
    n2358, n2359, n2360_1, n2361, n2362, n2363, n2364, n2365_1, n2366,
    n2367, n2368, n2369, n2370_1, n2371, n2372, n2373, n2374, n2375_1,
    n2376, n2377, n2379, n2380_1, n2381, n2382, n2383, n2384, n2385_1,
    n2386, n2387, n2388, n2389, n2390_1, n2391, n2392, n2393, n2394,
    n2395_1, n2396, n2397, n2398, n2399, n2400_1, n2401, n2402, n2403,
    n2404, n2405_1, n2406, n2407, n2408, n2409, n2410_1, n2411, n2412,
    n2413, n2414, n2415_1, n2416, n2417, n2418, n2419, n2421, n2422, n2423,
    n2424, n2425_1, n2426, n2427, n2428, n2429, n2430_1, n2431, n2432,
    n2433, n2434, n2435_1, n2436, n2437, n2438, n2439, n2440_1, n2441,
    n2442, n2443, n2444, n2445_1, n2446, n2447, n2448, n2449, n2450_1,
    n2451, n2452, n2453, n2454, n2455_1, n2456, n2457, n2458, n2459, n2461,
    n2462, n2463, n2464, n2465_1, n2466, n2467, n2468, n2469, n2470_1,
    n2471, n2472, n2473, n2474, n2475_1, n2476, n2477, n2478, n2479,
    n2480_1, n2481, n2482, n2483, n2485_1, n2486, n2487, n2488, n2489,
    n2490_1, n2491, n2492, n2493, n2494, n2495_1, n2496, n2497, n2498,
    n2499, n2500_1, n2501, n2502, n2503, n2504, n2505_1, n2506, n2507,
    n2508, n2509, n2510_1, n2511, n2512, n2513, n2514, n2515_1, n2516,
    n2517, n2518, n2519, n2520_1, n2521, n2522, n2523, n2524, n2525_1,
    n2526, n2528, n2529, n2530_1, n2531, n2532, n2533, n2534, n2535_1,
    n2536, n2537, n2538, n2539, n2540_1, n2541, n2542, n2543, n2544,
    n2545_1, n2546, n2547, n2548, n2549, n2550_1, n2552, n2553, n2554,
    n2555_1, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2708, n2709,
    n2710, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
    n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
    n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
    n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
    n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
    n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
    n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
    n3703, n3704, n3705, n3706, n3707, n3708, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
    n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
    n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
    n4577, n4578, n4579, n4580, n4581, n4582, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
    n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
    n4638, n4639, n4640, n4641, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4791, n4792,
    n4793, n4794, n4796, n4797, n4799, n4800, n4802, n4803, n4805, n4806,
    n4808, n4809, n4811, n4812, n4814, n4815, n4817, n4818, n4820, n4821,
    n4823, n4824, n4826, n4827, n4829, n4830, n4832, n4833, n4835, n4836,
    n4838, n4839, n4841, n4842, n4844, n4845, n4847, n4848, n4850, n4851,
    n4853, n4854, n4856, n4857, n4859, n4860, n4862, n4863, n4865, n4866,
    n4868, n4869, n4871, n4872, n4874, n4875, n4877, n4878, n4880, n4881,
    n4883, n4884, n4886, n4887, n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
    n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5296, n5297, n5298, n5299, n5300, n5301, n5303, n5304, n5305,
    n5306, n5307, n5309, n5310, n5311, n5312, n5313, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
    n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
    n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
    n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
    n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
    n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
    n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
    n6167, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6191, n6192, n6194, n6195, n6197, n6198, n6200, n6201,
    n6203, n6204, n6206, n6207, n6209, n6210, n6212, n6213, n6215, n6216,
    n6218, n6219, n6221, n6222, n6224, n6225, n6227, n6228, n6230, n6231,
    n6233, n6234, n6236, n6237, n6239, n6240, n6242, n6243, n6245, n6246,
    n6248, n6249, n6251, n6252, n6254, n6255, n6257, n6258, n6260, n6261,
    n6263, n6264, n6266, n6267, n6269, n6270, n6272, n6273, n6275, n6276,
    n6278, n6279, n6281, n6282, n6284, n6285, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
    n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
    n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
    n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
    n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
    n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
    n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
    n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
    n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
    n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
    n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7415, n7416, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
    n7656, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
    n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8323, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
    n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8459, n8460, n8461, n8462, n8463,
    n8464, n8465, n8466, n8467, n8468, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
    n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
    n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8556, n8557, n8558, n8559, n8560, n8561,
    n8562, n8563, n8564, n8565, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8594, n8595, n8596, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8864, n8865, n8866,
    n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
    n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
    n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
    n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
    n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
    n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
    n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
    n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
    n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
    n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
    n9232, n9233, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9364,
    n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
    n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725, n9727, n9728, n9729, n9730,
    n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
    n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
    n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9913,
    n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
    n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
    n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
    n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
    n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10185, n10186, n10187,
    n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
    n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
    n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
    n10398, n10399, n10400, n10401, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
    n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10531, n10532, n10533, n10534, n10535, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552, n10554, n10555, n10557,
    n10558, n10560, n10561, n10563, n10564, n10566, n10567, n10569, n10570,
    n10572, n10573, n10575, n10576, n10578, n10579, n10581, n10582, n10584,
    n10585, n10587, n10588, n10590, n10591, n10593, n10594, n10596, n10597,
    n10599, n10600, n10602, n10603, n10605, n10606, n10608, n10609, n10611,
    n10612, n10614, n10615, n10617, n10618, n10620, n10621, n10623, n10624,
    n10626, n10627, n10629, n10630, n10632, n10633, n10635, n10636, n10638,
    n10639, n10641, n10642, n10644, n10645, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
    n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
    n10738, n10739, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
    n10837, n10838, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
    n10936, n10937, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10958, n10959, n10961, n10962, n10963, n10964, n10965,
    n10966, n10967, n10968, n10969, n10970, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981, n10983, n10984, n10985,
    n10986, n10987, n10988, n10989, n10990, n10992, n10993, n10994, n10995,
    n10996, n10998, n10999, n11000, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
    n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
    n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
    n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
    n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11809, n11810, n11811, n11812, n11813, n11814,
    n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
    n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
    n11833, n11834, n11835, n11836, n11837, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11874, n11875, n11876, n11877, n11878, n11879,
    n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11904, n11905, n11906, n11907,
    n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
    n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
    n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
    n11935, n11936, n11937, n11938, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
    n11964, n11965, n11967, n11968, n11970, n11971, n11973, n11974, n11976,
    n11977, n11979, n11980, n11982, n11983, n11985, n11986, n11988, n11989,
    n11991, n11992, n11994, n11995, n11997, n11998, n12000, n12001, n12003,
    n12004, n12006, n12007, n12009, n12010, n12012, n12013, n12015, n12016,
    n12018, n12019, n12021, n12022, n12024, n12025, n12027, n12028, n12030,
    n12031, n12033, n12034, n12036, n12037, n12039, n12040, n12042, n12043,
    n12045, n12046, n12048, n12049, n12051, n12052, n12054, n12055, n12057,
    n12058, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
    n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
    n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
    n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
    n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
    n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
    n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
    n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
    n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
    n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
    n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
    n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
    n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
    n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
    n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
    n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
    n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
    n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
    n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
    n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
    n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
    n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
    n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
    n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
    n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
    n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
    n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
    n13226, n13227, n13228, n13229, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13251, n13252, n13253, n13254,
    n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
    n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
    n13273, n13274, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
    n13330, n13331, n13332, n13333, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13372, n13373, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13438, n13439, n13440, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458, n13460, n13461, n13462,
    n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13592, n13593,
    n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
    n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13741, n13742, n110, n115,
    n120, n125, n130, n135, n140, n145, n150, n155, n160, n165, n170, n175,
    n180, n185, n190, n195, n200, n205, n210, n215, n220, n225, n230, n235,
    n240, n245, n250, n255, n260, n265, n270, n275, n280, n285, n290, n295,
    n300, n305, n310, n315, n320, n325, n330, n335, n340, n345, n350, n355,
    n360, n365, n370, n375, n380, n385, n390, n395, n400, n405, n410, n415,
    n420, n425, n430, n435, n440, n445, n450, n455, n460, n465, n470, n475,
    n480, n485, n490, n495, n500, n505, n510, n515, n520, n525, n530, n535,
    n540, n545, n550, n555, n560, n565, n570, n575, n580, n585, n590, n595,
    n600, n605, n610, n615, n620, n625, n630, n635, n640, n645, n650, n655,
    n660, n665, n670, n675, n680, n685, n690, n695, n700, n705, n710, n715,
    n720, n725, n730, n735, n740, n745, n750, n755, n760, n765, n770, n775,
    n780, n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835,
    n840, n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895,
    n900, n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955,
    n960, n965, n970, n975, n980, n985, n990, n995, n1000, n1005, n1010,
    n1015, n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060,
    n1065, n1070, n1075, n1080, n1085, n1090, n1095, n1100, n1105, n1110,
    n1115, n1120, n1125, n1130, n1135, n1140, n1145, n1150, n1155, n1160,
    n1165, n1170, n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210,
    n1215, n1220, n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260,
    n1265, n1270, n1275, n1280, n1285, n1290, n1295, n1300, n1305, n1310,
    n1315, n1320, n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360,
    n1365, n1370, n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410,
    n1415, n1420, n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460,
    n1465, n1470, n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510,
    n1515, n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560,
    n1565, n1570, n1575, n1580, n1585, n1590, n1595, n1600, n1605, n1610,
    n1615, n1620, n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660,
    n1665, n1670, n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710,
    n1715, n1720, n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760,
    n1765, n1770, n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810,
    n1815, n1820, n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860,
    n1865, n1870, n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910,
    n1915, n1920, n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960,
    n1965, n1970, n1975, n1980, n1985, n1990, n1995, n2000, n2005, n2010,
    n2015, n2020, n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060,
    n2065, n2070, n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110,
    n2115, n2120, n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160,
    n2165, n2170, n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210,
    n2215, n2220, n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260,
    n2265, n2270, n2275, n2280, n2285, n2290, n2295, n2300, n2305, n2310,
    n2315, n2320, n2325, n2330, n2335, n2340, n2345, n2350, n2355, n2360,
    n2365, n2370, n2375, n2380, n2385, n2390, n2395, n2400, n2405, n2410,
    n2415, n2420, n2425, n2430, n2435, n2440, n2445, n2450, n2455, n2460,
    n2465, n2470, n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510,
    n2515, n2520, n2525, n2530, n2535, n2540, n2545, n2550, n2555;
  assign n1525_1 = ~P1_ADDR_REG_18_ & ~P2_ADDR_REG_18_;
  assign n1526 = P1_ADDR_REG_19_ & ~P2_ADDR_REG_19_;
  assign n1527 = ~P1_ADDR_REG_19_ & P2_ADDR_REG_19_;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = P1_ADDR_REG_17_ & P2_ADDR_REG_17_;
  assign n1530_1 = ~P1_ADDR_REG_17_ & ~P2_ADDR_REG_17_;
  assign n1531 = P1_ADDR_REG_16_ & P2_ADDR_REG_16_;
  assign n1532 = ~P1_ADDR_REG_16_ & ~P2_ADDR_REG_16_;
  assign n1533 = P1_ADDR_REG_15_ & P2_ADDR_REG_15_;
  assign n1534 = ~P1_ADDR_REG_15_ & ~P2_ADDR_REG_15_;
  assign n1535_1 = P1_ADDR_REG_14_ & P2_ADDR_REG_14_;
  assign n1536 = ~P1_ADDR_REG_14_ & ~P2_ADDR_REG_14_;
  assign n1537 = P1_ADDR_REG_13_ & P2_ADDR_REG_13_;
  assign n1538 = ~P1_ADDR_REG_13_ & ~P2_ADDR_REG_13_;
  assign n1539 = P1_ADDR_REG_12_ & P2_ADDR_REG_12_;
  assign n1540_1 = ~P1_ADDR_REG_12_ & ~P2_ADDR_REG_12_;
  assign n1541 = P1_ADDR_REG_11_ & P2_ADDR_REG_11_;
  assign n1542 = ~P1_ADDR_REG_11_ & ~P2_ADDR_REG_11_;
  assign n1543 = P1_ADDR_REG_10_ & P2_ADDR_REG_10_;
  assign n1544 = ~P1_ADDR_REG_10_ & ~P2_ADDR_REG_10_;
  assign n1545_1 = P1_ADDR_REG_9_ & P2_ADDR_REG_9_;
  assign n1546 = ~P1_ADDR_REG_9_ & ~P2_ADDR_REG_9_;
  assign n1547 = P1_ADDR_REG_8_ & P2_ADDR_REG_8_;
  assign n1548 = ~P1_ADDR_REG_8_ & ~P2_ADDR_REG_8_;
  assign n1549 = P1_ADDR_REG_7_ & P2_ADDR_REG_7_;
  assign n1550_1 = ~P1_ADDR_REG_7_ & ~P2_ADDR_REG_7_;
  assign n1551 = P1_ADDR_REG_6_ & P2_ADDR_REG_6_;
  assign n1552 = ~P1_ADDR_REG_6_ & ~P2_ADDR_REG_6_;
  assign n1553 = P1_ADDR_REG_5_ & P2_ADDR_REG_5_;
  assign n1554 = ~P1_ADDR_REG_5_ & ~P2_ADDR_REG_5_;
  assign n1555_1 = P1_ADDR_REG_4_ & P2_ADDR_REG_4_;
  assign n1556 = ~P1_ADDR_REG_4_ & ~P2_ADDR_REG_4_;
  assign n1557 = P1_ADDR_REG_3_ & P2_ADDR_REG_3_;
  assign n1558 = ~P1_ADDR_REG_3_ & ~P2_ADDR_REG_3_;
  assign n1559 = P1_ADDR_REG_2_ & P2_ADDR_REG_2_;
  assign n1560_1 = ~P1_ADDR_REG_2_ & ~P2_ADDR_REG_2_;
  assign n1561 = P1_ADDR_REG_0_ & P2_ADDR_REG_0_;
  assign n1562 = P1_ADDR_REG_1_ & n1561;
  assign n1563 = ~P1_ADDR_REG_1_ & ~n1561;
  assign n1564 = P2_ADDR_REG_1_ & ~n1563;
  assign n1565_1 = ~n1562 & ~n1564;
  assign n1566 = ~n1560_1 & ~n1565_1;
  assign n1567 = ~n1559 & ~n1566;
  assign n1568 = ~n1558 & ~n1567;
  assign n1569 = ~n1557 & ~n1568;
  assign n1570_1 = ~n1556 & ~n1569;
  assign n1571 = ~n1555_1 & ~n1570_1;
  assign n1572 = ~n1554 & ~n1571;
  assign n1573 = ~n1553 & ~n1572;
  assign n1574 = ~n1552 & ~n1573;
  assign n1575_1 = ~n1551 & ~n1574;
  assign n1576 = ~n1550_1 & ~n1575_1;
  assign n1577 = ~n1549 & ~n1576;
  assign n1578 = ~n1548 & ~n1577;
  assign n1579 = ~n1547 & ~n1578;
  assign n1580_1 = ~n1546 & ~n1579;
  assign n1581 = ~n1545_1 & ~n1580_1;
  assign n1582 = ~n1544 & ~n1581;
  assign n1583 = ~n1543 & ~n1582;
  assign n1584 = ~n1542 & ~n1583;
  assign n1585_1 = ~n1541 & ~n1584;
  assign n1586 = ~n1540_1 & ~n1585_1;
  assign n1587 = ~n1539 & ~n1586;
  assign n1588 = ~n1538 & ~n1587;
  assign n1589 = ~n1537 & ~n1588;
  assign n1590_1 = ~n1536 & ~n1589;
  assign n1591 = ~n1535_1 & ~n1590_1;
  assign n1592 = ~n1534 & ~n1591;
  assign n1593 = ~n1533 & ~n1592;
  assign n1594 = ~n1532 & ~n1593;
  assign n1595_1 = ~n1531 & ~n1594;
  assign n1596 = ~n1530_1 & ~n1595_1;
  assign n1597 = ~n1529 & ~n1596;
  assign n1598 = P1_ADDR_REG_18_ & P2_ADDR_REG_18_;
  assign n1599 = n1597 & ~n1598;
  assign n1600_1 = ~n1525_1 & ~n1528;
  assign n1601 = ~n1599 & n1600_1;
  assign n1602 = ~n1525_1 & ~n1597;
  assign n1603 = n1528 & ~n1598;
  assign n1604 = ~n1602 & n1603;
  assign ADD_1068_U4 = ~n1601 & ~n1604;
  assign n1606 = P1_ADDR_REG_18_ & ~P2_ADDR_REG_18_;
  assign n1607 = ~P1_ADDR_REG_18_ & P2_ADDR_REG_18_;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = n1597 & ~n1608;
  assign n1610_1 = ~n1597 & n1608;
  assign ADD_1068_U55 = n1609 | n1610_1;
  assign n1612 = P1_ADDR_REG_17_ & ~P2_ADDR_REG_17_;
  assign n1613 = ~P1_ADDR_REG_17_ & P2_ADDR_REG_17_;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615_1 = n1595_1 & ~n1614;
  assign n1616 = ~n1595_1 & n1614;
  assign ADD_1068_U56 = n1615_1 | n1616;
  assign n1618 = P1_ADDR_REG_16_ & ~P2_ADDR_REG_16_;
  assign n1619 = ~P1_ADDR_REG_16_ & P2_ADDR_REG_16_;
  assign n1620_1 = ~n1618 & ~n1619;
  assign n1621 = n1593 & ~n1620_1;
  assign n1622 = ~n1593 & n1620_1;
  assign ADD_1068_U57 = n1621 | n1622;
  assign n1624 = P1_ADDR_REG_15_ & ~P2_ADDR_REG_15_;
  assign n1625_1 = ~P1_ADDR_REG_15_ & P2_ADDR_REG_15_;
  assign n1626 = ~n1624 & ~n1625_1;
  assign n1627 = n1591 & ~n1626;
  assign n1628 = ~n1591 & n1626;
  assign ADD_1068_U58 = n1627 | n1628;
  assign n1630_1 = P1_ADDR_REG_14_ & ~P2_ADDR_REG_14_;
  assign n1631 = ~P1_ADDR_REG_14_ & P2_ADDR_REG_14_;
  assign n1632 = ~n1630_1 & ~n1631;
  assign n1633 = n1589 & ~n1632;
  assign n1634 = ~n1589 & n1632;
  assign ADD_1068_U59 = n1633 | n1634;
  assign n1636 = P1_ADDR_REG_13_ & ~P2_ADDR_REG_13_;
  assign n1637 = ~P1_ADDR_REG_13_ & P2_ADDR_REG_13_;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = n1587 & ~n1638;
  assign n1640_1 = ~n1587 & n1638;
  assign ADD_1068_U60 = n1639 | n1640_1;
  assign n1642 = P1_ADDR_REG_12_ & ~P2_ADDR_REG_12_;
  assign n1643 = ~P1_ADDR_REG_12_ & P2_ADDR_REG_12_;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645_1 = n1585_1 & ~n1644;
  assign n1646 = ~n1585_1 & n1644;
  assign ADD_1068_U61 = n1645_1 | n1646;
  assign n1648 = P1_ADDR_REG_11_ & ~P2_ADDR_REG_11_;
  assign n1649 = ~P1_ADDR_REG_11_ & P2_ADDR_REG_11_;
  assign n1650_1 = ~n1648 & ~n1649;
  assign n1651 = n1583 & ~n1650_1;
  assign n1652 = ~n1583 & n1650_1;
  assign ADD_1068_U62 = n1651 | n1652;
  assign n1654 = P1_ADDR_REG_10_ & ~P2_ADDR_REG_10_;
  assign n1655_1 = ~P1_ADDR_REG_10_ & P2_ADDR_REG_10_;
  assign n1656 = ~n1654 & ~n1655_1;
  assign n1657 = n1581 & ~n1656;
  assign n1658 = ~n1581 & n1656;
  assign ADD_1068_U63 = n1657 | n1658;
  assign n1660_1 = P1_ADDR_REG_9_ & ~P2_ADDR_REG_9_;
  assign n1661 = ~P1_ADDR_REG_9_ & P2_ADDR_REG_9_;
  assign n1662 = ~n1660_1 & ~n1661;
  assign n1663 = n1579 & ~n1662;
  assign n1664 = ~n1579 & n1662;
  assign ADD_1068_U47 = n1663 | n1664;
  assign n1666 = P1_ADDR_REG_8_ & ~P2_ADDR_REG_8_;
  assign n1667 = ~P1_ADDR_REG_8_ & P2_ADDR_REG_8_;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = n1577 & ~n1668;
  assign n1670_1 = ~n1577 & n1668;
  assign ADD_1068_U48 = n1669 | n1670_1;
  assign n1672 = P1_ADDR_REG_7_ & ~P2_ADDR_REG_7_;
  assign n1673 = ~P1_ADDR_REG_7_ & P2_ADDR_REG_7_;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675_1 = n1575_1 & ~n1674;
  assign n1676 = ~n1575_1 & n1674;
  assign ADD_1068_U49 = n1675_1 | n1676;
  assign n1678 = P1_ADDR_REG_6_ & ~P2_ADDR_REG_6_;
  assign n1679 = ~P1_ADDR_REG_6_ & P2_ADDR_REG_6_;
  assign n1680_1 = ~n1678 & ~n1679;
  assign n1681 = n1573 & ~n1680_1;
  assign n1682 = ~n1573 & n1680_1;
  assign ADD_1068_U50 = n1681 | n1682;
  assign n1684 = P1_ADDR_REG_5_ & ~P2_ADDR_REG_5_;
  assign n1685_1 = ~P1_ADDR_REG_5_ & P2_ADDR_REG_5_;
  assign n1686 = ~n1684 & ~n1685_1;
  assign n1687 = n1571 & ~n1686;
  assign n1688 = ~n1571 & n1686;
  assign ADD_1068_U51 = n1687 | n1688;
  assign n1690_1 = P1_ADDR_REG_4_ & ~P2_ADDR_REG_4_;
  assign n1691 = ~P1_ADDR_REG_4_ & P2_ADDR_REG_4_;
  assign n1692 = ~n1690_1 & ~n1691;
  assign n1693 = n1569 & ~n1692;
  assign n1694 = ~n1569 & n1692;
  assign ADD_1068_U52 = n1693 | n1694;
  assign n1696 = P1_ADDR_REG_3_ & ~P2_ADDR_REG_3_;
  assign n1697 = ~P1_ADDR_REG_3_ & P2_ADDR_REG_3_;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = n1567 & ~n1698;
  assign n1700_1 = ~n1567 & n1698;
  assign ADD_1068_U53 = n1699 | n1700_1;
  assign n1702 = P1_ADDR_REG_2_ & ~P2_ADDR_REG_2_;
  assign n1703 = ~P1_ADDR_REG_2_ & P2_ADDR_REG_2_;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705_1 = n1565_1 & ~n1704;
  assign n1706 = ~n1565_1 & n1704;
  assign ADD_1068_U54 = n1705_1 | n1706;
  assign n1708 = P2_ADDR_REG_1_ & n1562;
  assign n1709 = P1_ADDR_REG_1_ & ~n1561;
  assign n1710_1 = ~P2_ADDR_REG_1_ & n1709;
  assign n1711 = ~P2_ADDR_REG_1_ & n1561;
  assign n1712 = P2_ADDR_REG_1_ & ~n1561;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = ~P1_ADDR_REG_1_ & ~n1713;
  assign n1715_1 = ~n1708 & ~n1710_1;
  assign ADD_1068_U5 = n1714 | ~n1715_1;
  assign n1717 = P1_ADDR_REG_0_ & ~P2_ADDR_REG_0_;
  assign n1718 = ~P1_ADDR_REG_0_ & P2_ADDR_REG_0_;
  assign ADD_1068_U46 = n1717 | n1718;
  assign n1720_1 = P1_RD_REG & ~P2_RD_REG;
  assign n1721 = ~P1_RD_REG & P2_RD_REG;
  assign U126 = ~n1720_1 & ~n1721;
  assign n1723 = P1_WR_REG & ~P2_WR_REG;
  assign n1724 = ~P1_WR_REG & P2_WR_REG;
  assign U123 = ~n1723 & ~n1724;
  assign n1726 = ~P1_IR_REG_31_ & P1_STATE_REG;
  assign n1727 = P1_STATE_REG & ~n1726;
  assign n1728 = P1_IR_REG_0_ & n1727;
  assign n1729 = P1_IR_REG_0_ & n1726;
  assign n1730_1 = P1_ADDR_REG_19_ & ~P2_RD_REG;
  assign n1731 = P2_ADDR_REG_19_ & n1730_1;
  assign n1732 = ~P1_ADDR_REG_19_ & ~P1_RD_REG;
  assign n1733 = ~P2_ADDR_REG_19_ & n1732;
  assign n1734 = ~n1731 & ~n1733;
  assign n1735_1 = P2_DATAO_REG_0_ & n1734;
  assign n1736 = P1_DATAO_REG_0_ & n1734;
  assign n1737 = P2_DATAO_REG_0_ & ~n1734;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = SI_0_ & n1738;
  assign n1740_1 = ~SI_0_ & ~n1738;
  assign n1741 = ~n1739 & ~n1740_1;
  assign n1742 = ~n1734 & ~n1741;
  assign n1743 = ~n1735_1 & ~n1742;
  assign n1744 = ~P1_STATE_REG & ~n1743;
  assign n1745_1 = ~n1728 & ~n1729;
  assign n110 = n1744 | ~n1745_1;
  assign n1747 = P1_IR_REG_0_ & ~P1_IR_REG_1_;
  assign n1748 = ~P1_IR_REG_0_ & P1_IR_REG_1_;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750_1 = n1727 & ~n1749;
  assign n1751 = P1_IR_REG_1_ & n1726;
  assign n1752 = P2_DATAO_REG_1_ & n1734;
  assign n1753 = SI_0_ & ~n1738;
  assign n1754 = P1_DATAO_REG_1_ & n1734;
  assign n1755_1 = P2_DATAO_REG_1_ & ~n1734;
  assign n1756 = ~n1754 & ~n1755_1;
  assign n1757 = n1753 & n1756;
  assign n1758 = ~n1753 & ~n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760_1 = ~SI_1_ & ~n1759;
  assign n1761 = ~n1753 & n1756;
  assign n1762 = SI_1_ & n1761;
  assign n1763 = SI_1_ & SI_0_;
  assign n1764 = ~n1738 & n1763;
  assign n1765_1 = ~n1756 & n1764;
  assign n1766 = ~n1760_1 & ~n1762;
  assign n1767 = ~n1765_1 & n1766;
  assign n1768 = ~n1734 & ~n1767;
  assign n1769 = ~n1752 & ~n1768;
  assign n1770_1 = ~P1_STATE_REG & ~n1769;
  assign n1771 = ~n1750_1 & ~n1751;
  assign n115 = n1770_1 | ~n1771;
  assign n1773 = ~P1_IR_REG_0_ & ~P1_IR_REG_1_;
  assign n1774 = P1_IR_REG_2_ & ~n1773;
  assign n1775_1 = ~P1_IR_REG_2_ & n1773;
  assign n1776 = ~n1774 & ~n1775_1;
  assign n1777 = n1727 & n1776;
  assign n1778 = P1_IR_REG_2_ & n1726;
  assign n1779 = P2_DATAO_REG_2_ & n1734;
  assign n1780_1 = SI_1_ & ~n1756;
  assign n1781 = n1753 & ~n1756;
  assign n1782 = ~n1764 & ~n1780_1;
  assign n1783 = ~n1781 & n1782;
  assign n1784 = P1_DATAO_REG_2_ & n1734;
  assign n1785_1 = P2_DATAO_REG_2_ & ~n1734;
  assign n1786 = ~n1784 & ~n1785_1;
  assign n1787 = SI_2_ & n1786;
  assign n1788 = ~SI_2_ & ~n1786;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790_1 = n1783 & ~n1789;
  assign n1791 = ~n1783 & n1789;
  assign n1792 = ~n1790_1 & ~n1791;
  assign n1793 = ~n1734 & ~n1792;
  assign n1794 = ~n1779 & ~n1793;
  assign n1795_1 = ~P1_STATE_REG & ~n1794;
  assign n1796 = ~n1777 & ~n1778;
  assign n120 = n1795_1 | ~n1796;
  assign n1798 = P1_IR_REG_3_ & ~n1775_1;
  assign n1799 = ~P1_IR_REG_3_ & n1775_1;
  assign n1800_1 = ~n1798 & ~n1799;
  assign n1801 = n1727 & n1800_1;
  assign n1802 = P1_IR_REG_3_ & n1726;
  assign n1803 = P2_DATAO_REG_3_ & n1734;
  assign n1804 = SI_2_ & ~n1786;
  assign n1805_1 = ~SI_2_ & n1786;
  assign n1806 = ~n1783 & ~n1805_1;
  assign n1807 = ~n1804 & ~n1806;
  assign n1808 = P1_DATAO_REG_3_ & n1734;
  assign n1809 = P2_DATAO_REG_3_ & ~n1734;
  assign n1810_1 = ~n1808 & ~n1809;
  assign n1811 = SI_3_ & n1810_1;
  assign n1812 = ~SI_3_ & ~n1810_1;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = n1807 & ~n1813;
  assign n1815_1 = ~n1807 & n1813;
  assign n1816 = ~n1814 & ~n1815_1;
  assign n1817 = ~n1734 & ~n1816;
  assign n1818 = ~n1803 & ~n1817;
  assign n1819 = ~P1_STATE_REG & ~n1818;
  assign n1820_1 = ~n1801 & ~n1802;
  assign n125 = n1819 | ~n1820_1;
  assign n1822 = P1_IR_REG_4_ & ~n1799;
  assign n1823 = ~P1_IR_REG_3_ & ~P1_IR_REG_4_;
  assign n1824 = n1775_1 & n1823;
  assign n1825_1 = ~n1822 & ~n1824;
  assign n1826 = n1727 & n1825_1;
  assign n1827 = P1_IR_REG_4_ & n1726;
  assign n1828 = P2_DATAO_REG_4_ & n1734;
  assign n1829 = ~SI_3_ & n1810_1;
  assign n1830_1 = n1804 & ~n1829;
  assign n1831 = SI_3_ & ~n1810_1;
  assign n1832 = ~n1830_1 & ~n1831;
  assign n1833 = ~n1805_1 & ~n1829;
  assign n1834 = ~n1783 & n1833;
  assign n1835_1 = n1832 & ~n1834;
  assign n1836 = P1_DATAO_REG_4_ & n1734;
  assign n1837 = P2_DATAO_REG_4_ & ~n1734;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = SI_4_ & n1838;
  assign n1840_1 = ~SI_4_ & ~n1838;
  assign n1841 = ~n1839 & ~n1840_1;
  assign n1842 = n1835_1 & ~n1841;
  assign n1843 = ~n1835_1 & n1841;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845_1 = ~n1734 & ~n1844;
  assign n1846 = ~n1828 & ~n1845_1;
  assign n1847 = ~P1_STATE_REG & ~n1846;
  assign n1848 = ~n1826 & ~n1827;
  assign n130 = n1847 | ~n1848;
  assign n1850_1 = ~P1_IR_REG_5_ & n1824;
  assign n1851 = P1_IR_REG_5_ & ~n1824;
  assign n1852 = ~n1850_1 & ~n1851;
  assign n1853 = n1727 & n1852;
  assign n1854 = P1_IR_REG_5_ & n1726;
  assign n1855_1 = P2_DATAO_REG_5_ & n1734;
  assign n1856 = ~SI_4_ & n1838;
  assign n1857 = ~n1835_1 & ~n1856;
  assign n1858 = SI_4_ & ~n1838;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860_1 = P1_DATAO_REG_5_ & n1734;
  assign n1861 = P2_DATAO_REG_5_ & ~n1734;
  assign n1862 = ~n1860_1 & ~n1861;
  assign n1863 = SI_5_ & n1862;
  assign n1864 = ~SI_5_ & ~n1862;
  assign n1865_1 = ~n1863 & ~n1864;
  assign n1866 = n1859 & ~n1865_1;
  assign n1867 = ~n1859 & n1865_1;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = ~n1734 & ~n1868;
  assign n1870_1 = ~n1855_1 & ~n1869;
  assign n1871 = ~P1_STATE_REG & ~n1870_1;
  assign n1872 = ~n1853 & ~n1854;
  assign n135 = n1871 | ~n1872;
  assign n1874 = P1_IR_REG_6_ & ~n1850_1;
  assign n1875_1 = ~P1_IR_REG_5_ & ~P1_IR_REG_6_;
  assign n1876 = n1824 & n1875_1;
  assign n1877 = ~n1874 & ~n1876;
  assign n1878 = n1727 & n1877;
  assign n1879 = P1_IR_REG_6_ & n1726;
  assign n1880_1 = P2_DATAO_REG_6_ & n1734;
  assign n1881 = ~SI_5_ & n1862;
  assign n1882 = n1858 & ~n1881;
  assign n1883 = SI_5_ & ~n1862;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885_1 = ~n1856 & ~n1881;
  assign n1886 = ~n1835_1 & n1885_1;
  assign n1887 = n1884 & ~n1886;
  assign n1888 = P1_DATAO_REG_6_ & n1734;
  assign n1889 = P2_DATAO_REG_6_ & ~n1734;
  assign n1890_1 = ~n1888 & ~n1889;
  assign n1891 = SI_6_ & n1890_1;
  assign n1892 = ~SI_6_ & ~n1890_1;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = n1887 & ~n1893;
  assign n1895_1 = ~n1887 & n1893;
  assign n1896 = ~n1894 & ~n1895_1;
  assign n1897 = ~n1734 & ~n1896;
  assign n1898 = ~n1880_1 & ~n1897;
  assign n1899 = ~P1_STATE_REG & ~n1898;
  assign n1900_1 = ~n1878 & ~n1879;
  assign n140 = n1899 | ~n1900_1;
  assign n1902 = P1_IR_REG_7_ & ~n1876;
  assign n1903 = ~P1_IR_REG_7_ & n1876;
  assign n1904 = ~n1902 & ~n1903;
  assign n1905_1 = n1727 & n1904;
  assign n1906 = P1_IR_REG_7_ & n1726;
  assign n1907 = P2_DATAO_REG_7_ & n1734;
  assign n1908 = ~SI_6_ & n1890_1;
  assign n1909 = ~n1884 & ~n1908;
  assign n1910_1 = SI_6_ & ~n1890_1;
  assign n1911 = ~n1909 & ~n1910_1;
  assign n1912 = n1885_1 & ~n1908;
  assign n1913 = ~n1835_1 & n1912;
  assign n1914 = n1911 & ~n1913;
  assign n1915_1 = P1_DATAO_REG_7_ & n1734;
  assign n1916 = P2_DATAO_REG_7_ & ~n1734;
  assign n1917 = ~n1915_1 & ~n1916;
  assign n1918 = SI_7_ & n1917;
  assign n1919 = ~SI_7_ & ~n1917;
  assign n1920_1 = ~n1918 & ~n1919;
  assign n1921 = n1914 & ~n1920_1;
  assign n1922 = ~n1914 & n1920_1;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~n1734 & ~n1923;
  assign n1925_1 = ~n1907 & ~n1924;
  assign n1926 = ~P1_STATE_REG & ~n1925_1;
  assign n1927 = ~n1905_1 & ~n1906;
  assign n145 = n1926 | ~n1927;
  assign n1929 = P1_IR_REG_8_ & ~n1903;
  assign n1930_1 = ~P1_IR_REG_7_ & ~P1_IR_REG_8_;
  assign n1931 = ~P1_IR_REG_5_ & n1823;
  assign n1932 = ~P1_IR_REG_6_ & n1931;
  assign n1933 = n1775_1 & n1930_1;
  assign n1934 = n1932 & n1933;
  assign n1935_1 = ~n1929 & ~n1934;
  assign n1936 = n1727 & n1935_1;
  assign n1937 = P1_IR_REG_8_ & n1726;
  assign n1938 = P2_DATAO_REG_8_ & n1734;
  assign n1939 = ~SI_7_ & n1917;
  assign n1940_1 = ~n1914 & ~n1939;
  assign n1941 = SI_7_ & ~n1917;
  assign n1942 = ~n1940_1 & ~n1941;
  assign n1943 = P1_DATAO_REG_8_ & n1734;
  assign n1944 = P2_DATAO_REG_8_ & ~n1734;
  assign n1945_1 = ~n1943 & ~n1944;
  assign n1946 = SI_8_ & n1945_1;
  assign n1947 = ~SI_8_ & ~n1945_1;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = n1942 & ~n1948;
  assign n1950_1 = ~n1942 & n1948;
  assign n1951 = ~n1949 & ~n1950_1;
  assign n1952 = ~n1734 & ~n1951;
  assign n1953 = ~n1938 & ~n1952;
  assign n1954 = ~P1_STATE_REG & ~n1953;
  assign n1955_1 = ~n1936 & ~n1937;
  assign n150 = n1954 | ~n1955_1;
  assign n1957 = ~P1_IR_REG_9_ & n1934;
  assign n1958 = P1_IR_REG_9_ & ~n1934;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960_1 = n1727 & n1959;
  assign n1961 = P1_IR_REG_9_ & n1726;
  assign n1962 = P2_DATAO_REG_9_ & n1734;
  assign n1963 = ~SI_8_ & n1945_1;
  assign n1964 = n1941 & ~n1963;
  assign n1965_1 = SI_8_ & ~n1945_1;
  assign n1966 = ~n1964 & ~n1965_1;
  assign n1967 = ~n1939 & ~n1963;
  assign n1968 = ~n1914 & n1967;
  assign n1969 = n1966 & ~n1968;
  assign n1970_1 = P1_DATAO_REG_9_ & n1734;
  assign n1971 = P2_DATAO_REG_9_ & ~n1734;
  assign n1972 = ~n1970_1 & ~n1971;
  assign n1973 = SI_9_ & n1972;
  assign n1974 = ~SI_9_ & ~n1972;
  assign n1975_1 = ~n1973 & ~n1974;
  assign n1976 = n1969 & ~n1975_1;
  assign n1977 = ~n1969 & n1975_1;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1734 & ~n1978;
  assign n1980_1 = ~n1962 & ~n1979;
  assign n1981 = ~P1_STATE_REG & ~n1980_1;
  assign n1982 = ~n1960_1 & ~n1961;
  assign n155 = n1981 | ~n1982;
  assign n1984 = P1_IR_REG_10_ & ~n1957;
  assign n1985_1 = ~P1_IR_REG_9_ & ~P1_IR_REG_10_;
  assign n1986 = n1934 & n1985_1;
  assign n1987 = ~n1984 & ~n1986;
  assign n1988 = n1727 & n1987;
  assign n1989 = P1_IR_REG_10_ & n1726;
  assign n1990_1 = P2_DATAO_REG_10_ & n1734;
  assign n1991 = ~SI_9_ & n1972;
  assign n1992 = ~n1966 & ~n1991;
  assign n1993 = SI_9_ & ~n1972;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995_1 = n1967 & ~n1991;
  assign n1996 = ~n1914 & n1995_1;
  assign n1997 = n1994 & ~n1996;
  assign n1998 = P1_DATAO_REG_10_ & n1734;
  assign n1999 = P2_DATAO_REG_10_ & ~n1734;
  assign n2000_1 = ~n1998 & ~n1999;
  assign n2001 = SI_10_ & n2000_1;
  assign n2002 = ~SI_10_ & ~n2000_1;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = n1997 & ~n2003;
  assign n2005_1 = ~n1997 & n2003;
  assign n2006 = ~n2004 & ~n2005_1;
  assign n2007 = ~n1734 & ~n2006;
  assign n2008 = ~n1990_1 & ~n2007;
  assign n2009 = ~P1_STATE_REG & ~n2008;
  assign n2010_1 = ~n1988 & ~n1989;
  assign n160 = n2009 | ~n2010_1;
  assign n2012 = P1_IR_REG_11_ & ~n1986;
  assign n2013 = ~P1_IR_REG_11_ & n1986;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015_1 = n1727 & n2014;
  assign n2016 = P1_IR_REG_11_ & n1726;
  assign n2017 = P2_DATAO_REG_11_ & n1734;
  assign n2018 = ~SI_10_ & n2000_1;
  assign n2019 = ~n1994 & ~n2018;
  assign n2020_1 = SI_10_ & ~n2000_1;
  assign n2021 = ~n2019 & ~n2020_1;
  assign n2022 = n1995_1 & ~n2018;
  assign n2023 = ~n1914 & n2022;
  assign n2024 = n2021 & ~n2023;
  assign n2025_1 = P1_DATAO_REG_11_ & n1734;
  assign n2026 = P2_DATAO_REG_11_ & ~n1734;
  assign n2027 = ~n2025_1 & ~n2026;
  assign n2028 = SI_11_ & n2027;
  assign n2029 = ~SI_11_ & ~n2027;
  assign n2030_1 = ~n2028 & ~n2029;
  assign n2031 = n2024 & ~n2030_1;
  assign n2032 = ~n2024 & n2030_1;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n1734 & ~n2033;
  assign n2035_1 = ~n2017 & ~n2034;
  assign n2036 = ~P1_STATE_REG & ~n2035_1;
  assign n2037 = ~n2015_1 & ~n2016;
  assign n165 = n2036 | ~n2037;
  assign n2039 = P1_IR_REG_12_ & ~n2013;
  assign n2040_1 = ~P1_IR_REG_10_ & ~P1_IR_REG_11_;
  assign n2041 = ~P1_IR_REG_12_ & n2040_1;
  assign n2042 = ~P1_IR_REG_9_ & n2041;
  assign n2043 = n1934 & n2042;
  assign n2044 = ~n2039 & ~n2043;
  assign n2045_1 = n1727 & n2044;
  assign n2046 = P1_IR_REG_12_ & n1726;
  assign n2047 = P2_DATAO_REG_12_ & n1734;
  assign n2048 = SI_11_ & ~n2027;
  assign n2049 = ~SI_11_ & n2027;
  assign n2050_1 = ~n2024 & ~n2049;
  assign n2051 = ~n2048 & ~n2050_1;
  assign n2052 = P1_DATAO_REG_12_ & n1734;
  assign n2053 = P2_DATAO_REG_12_ & ~n1734;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055_1 = SI_12_ & n2054;
  assign n2056 = ~SI_12_ & ~n2054;
  assign n2057 = ~n2055_1 & ~n2056;
  assign n2058 = n2051 & ~n2057;
  assign n2059 = ~n2051 & n2057;
  assign n2060_1 = ~n2058 & ~n2059;
  assign n2061 = ~n1734 & ~n2060_1;
  assign n2062 = ~n2047 & ~n2061;
  assign n2063 = ~P1_STATE_REG & ~n2062;
  assign n2064 = ~n2045_1 & ~n2046;
  assign n170 = n2063 | ~n2064;
  assign n2066 = ~P1_IR_REG_13_ & n2043;
  assign n2067 = P1_IR_REG_13_ & ~n2043;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = n1727 & n2068;
  assign n2070_1 = P1_IR_REG_13_ & n1726;
  assign n2071 = P2_DATAO_REG_13_ & n1734;
  assign n2072 = ~SI_12_ & n2054;
  assign n2073 = n2048 & ~n2072;
  assign n2074 = SI_12_ & ~n2054;
  assign n2075_1 = ~n2073 & ~n2074;
  assign n2076 = ~n2049 & ~n2072;
  assign n2077 = ~n2024 & n2076;
  assign n2078 = n2075_1 & ~n2077;
  assign n2079 = P1_DATAO_REG_13_ & n1734;
  assign n2080_1 = P2_DATAO_REG_13_ & ~n1734;
  assign n2081 = ~n2079 & ~n2080_1;
  assign n2082 = SI_13_ & n2081;
  assign n2083 = ~SI_13_ & ~n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085_1 = n2078 & ~n2084;
  assign n2086 = ~n2078 & n2084;
  assign n2087 = ~n2085_1 & ~n2086;
  assign n2088 = ~n1734 & ~n2087;
  assign n2089 = ~n2071 & ~n2088;
  assign n2090_1 = ~P1_STATE_REG & ~n2089;
  assign n2091 = ~n2069 & ~n2070_1;
  assign n175 = n2090_1 | ~n2091;
  assign n2093 = P1_IR_REG_14_ & ~n2066;
  assign n2094 = ~P1_IR_REG_13_ & ~P1_IR_REG_14_;
  assign n2095_1 = n2043 & n2094;
  assign n2096 = ~n2093 & ~n2095_1;
  assign n2097 = n1727 & n2096;
  assign n2098 = P1_IR_REG_14_ & n1726;
  assign n2099 = P2_DATAO_REG_14_ & n1734;
  assign n2100_1 = ~SI_13_ & n2081;
  assign n2101 = ~n2075_1 & ~n2100_1;
  assign n2102 = SI_13_ & ~n2081;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = n2076 & ~n2100_1;
  assign n2105_1 = ~n2024 & n2104;
  assign n2106 = n2103 & ~n2105_1;
  assign n2107 = P1_DATAO_REG_14_ & n1734;
  assign n2108 = P2_DATAO_REG_14_ & ~n1734;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110_1 = SI_14_ & n2109;
  assign n2111 = ~SI_14_ & ~n2109;
  assign n2112 = ~n2110_1 & ~n2111;
  assign n2113 = n2106 & ~n2112;
  assign n2114 = ~n2106 & n2112;
  assign n2115_1 = ~n2113 & ~n2114;
  assign n2116 = ~n1734 & ~n2115_1;
  assign n2117 = ~n2099 & ~n2116;
  assign n2118 = ~P1_STATE_REG & ~n2117;
  assign n2119 = ~n2097 & ~n2098;
  assign n180 = n2118 | ~n2119;
  assign n2121 = P1_IR_REG_15_ & ~n2095_1;
  assign n2122 = ~P1_IR_REG_15_ & n2095_1;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = n1727 & n2123;
  assign n2125_1 = P1_IR_REG_15_ & n1726;
  assign n2126 = P2_DATAO_REG_15_ & n1734;
  assign n2127 = ~SI_14_ & n2109;
  assign n2128 = ~n2103 & ~n2127;
  assign n2129 = SI_14_ & ~n2109;
  assign n2130_1 = ~n2128 & ~n2129;
  assign n2131 = n2104 & ~n2127;
  assign n2132 = ~n2024 & n2131;
  assign n2133 = n2130_1 & ~n2132;
  assign n2134 = P1_DATAO_REG_15_ & n1734;
  assign n2135_1 = P2_DATAO_REG_15_ & ~n1734;
  assign n2136 = ~n2134 & ~n2135_1;
  assign n2137 = SI_15_ & n2136;
  assign n2138 = ~SI_15_ & ~n2136;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140_1 = n2133 & ~n2139;
  assign n2141 = ~n2133 & n2139;
  assign n2142 = ~n2140_1 & ~n2141;
  assign n2143 = ~n1734 & ~n2142;
  assign n2144 = ~n2126 & ~n2143;
  assign n2145_1 = ~P1_STATE_REG & ~n2144;
  assign n2146 = ~n2124 & ~n2125_1;
  assign n185 = n2145_1 | ~n2146;
  assign n2148 = P1_IR_REG_16_ & ~n2122;
  assign n2149 = ~P1_IR_REG_6_ & ~P1_IR_REG_7_;
  assign n2150_1 = ~P1_IR_REG_8_ & n2149;
  assign n2151 = ~P1_IR_REG_9_ & n2150_1;
  assign n2152 = ~P1_IR_REG_2_ & ~P1_IR_REG_3_;
  assign n2153 = ~P1_IR_REG_4_ & n2152;
  assign n2154 = ~P1_IR_REG_5_ & n2153;
  assign n2155_1 = ~P1_IR_REG_15_ & ~P1_IR_REG_16_;
  assign n2156 = ~P1_IR_REG_1_ & n2155_1;
  assign n2157 = ~P1_IR_REG_0_ & n2156;
  assign n2158 = ~P1_IR_REG_12_ & n2094;
  assign n2159 = ~P1_IR_REG_10_ & n2158;
  assign n2160_1 = ~P1_IR_REG_11_ & n2159;
  assign n2161 = n2151 & n2154;
  assign n2162 = n2157 & n2161;
  assign n2163 = n2160_1 & n2162;
  assign n2164 = ~n2148 & ~n2163;
  assign n2165_1 = n1727 & n2164;
  assign n2166 = P1_IR_REG_16_ & n1726;
  assign n2167 = P2_DATAO_REG_16_ & n1734;
  assign n2168 = SI_15_ & ~n2136;
  assign n2169 = ~SI_15_ & n2136;
  assign n2170_1 = ~n2133 & ~n2169;
  assign n2171 = ~n2168 & ~n2170_1;
  assign n2172 = P1_DATAO_REG_16_ & n1734;
  assign n2173 = P2_DATAO_REG_16_ & ~n1734;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175_1 = SI_16_ & n2174;
  assign n2176 = ~SI_16_ & ~n2174;
  assign n2177 = ~n2175_1 & ~n2176;
  assign n2178 = n2171 & ~n2177;
  assign n2179 = ~n2171 & n2177;
  assign n2180_1 = ~n2178 & ~n2179;
  assign n2181 = ~n1734 & ~n2180_1;
  assign n2182 = ~n2167 & ~n2181;
  assign n2183 = ~P1_STATE_REG & ~n2182;
  assign n2184 = ~n2165_1 & ~n2166;
  assign n190 = n2183 | ~n2184;
  assign n2186 = ~P1_IR_REG_17_ & n2163;
  assign n2187 = P1_IR_REG_17_ & ~n2163;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n1727 & n2188;
  assign n2190_1 = P1_IR_REG_17_ & n1726;
  assign n2191 = P2_DATAO_REG_17_ & n1734;
  assign n2192 = SI_16_ & ~n2174;
  assign n2193 = ~SI_16_ & n2174;
  assign n2194 = ~n2171 & ~n2193;
  assign n2195_1 = ~n2192 & ~n2194;
  assign n2196 = P1_DATAO_REG_17_ & n1734;
  assign n2197 = P2_DATAO_REG_17_ & ~n1734;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = SI_17_ & n2198;
  assign n2200_1 = ~SI_17_ & ~n2198;
  assign n2201 = ~n2199 & ~n2200_1;
  assign n2202 = n2195_1 & ~n2201;
  assign n2203 = ~n2195_1 & n2201;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205_1 = ~n1734 & ~n2204;
  assign n2206 = ~n2191 & ~n2205_1;
  assign n2207 = ~P1_STATE_REG & ~n2206;
  assign n2208 = ~n2189 & ~n2190_1;
  assign n195 = n2207 | ~n2208;
  assign n2210_1 = P1_IR_REG_18_ & ~n2186;
  assign n2211 = ~P1_IR_REG_4_ & ~P1_IR_REG_5_;
  assign n2212 = ~P1_IR_REG_3_ & n2211;
  assign n2213 = ~P1_IR_REG_0_ & n2212;
  assign n2214 = ~P1_IR_REG_2_ & n2213;
  assign n2215_1 = ~P1_IR_REG_1_ & ~P1_IR_REG_18_;
  assign n2216 = ~P1_IR_REG_17_ & n2215_1;
  assign n2217 = ~P1_IR_REG_15_ & n2216;
  assign n2218 = ~P1_IR_REG_16_ & n2217;
  assign n2219 = n2151 & n2214;
  assign n2220_1 = n2218 & n2219;
  assign n2221 = n2160_1 & n2220_1;
  assign n2222 = ~n2210_1 & ~n2221;
  assign n2223 = n1727 & n2222;
  assign n2224 = P1_IR_REG_18_ & n1726;
  assign n2225_1 = P2_DATAO_REG_18_ & n1734;
  assign n2226 = SI_17_ & ~n2198;
  assign n2227 = ~SI_17_ & n2198;
  assign n2228 = ~n2195_1 & ~n2227;
  assign n2229 = ~n2226 & ~n2228;
  assign n2230_1 = P1_DATAO_REG_18_ & n1734;
  assign n2231 = P2_DATAO_REG_18_ & ~n1734;
  assign n2232 = ~n2230_1 & ~n2231;
  assign n2233 = SI_18_ & n2232;
  assign n2234 = ~SI_18_ & ~n2232;
  assign n2235_1 = ~n2233 & ~n2234;
  assign n2236 = n2229 & ~n2235_1;
  assign n2237 = ~n2229 & n2235_1;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n1734 & ~n2238;
  assign n2240_1 = ~n2225_1 & ~n2239;
  assign n2241 = ~P1_STATE_REG & ~n2240_1;
  assign n2242 = ~n2223 & ~n2224;
  assign n200 = n2241 | ~n2242;
  assign n2244 = P1_IR_REG_19_ & ~n2221;
  assign n2245_1 = ~P1_IR_REG_8_ & ~P1_IR_REG_9_;
  assign n2246 = ~P1_IR_REG_7_ & n2245_1;
  assign n2247 = ~P1_IR_REG_5_ & n2246;
  assign n2248 = ~P1_IR_REG_6_ & n2247;
  assign n2249 = ~P1_IR_REG_2_ & n1823;
  assign n2250_1 = ~P1_IR_REG_1_ & n2249;
  assign n2251 = ~P1_IR_REG_0_ & n2250_1;
  assign n2252 = ~P1_IR_REG_18_ & ~P1_IR_REG_19_;
  assign n2253 = ~P1_IR_REG_17_ & n2252;
  assign n2254 = ~P1_IR_REG_15_ & n2253;
  assign n2255_1 = ~P1_IR_REG_16_ & n2254;
  assign n2256 = n2248 & n2251;
  assign n2257 = n2255_1 & n2256;
  assign n2258 = n2160_1 & n2257;
  assign n2259 = ~n2244 & ~n2258;
  assign n2260_1 = n1727 & n2259;
  assign n2261 = P1_IR_REG_19_ & n1726;
  assign n2262 = P2_DATAO_REG_19_ & n1734;
  assign n2263 = SI_18_ & ~n2232;
  assign n2264 = ~SI_18_ & n2232;
  assign n2265_1 = ~n2229 & ~n2264;
  assign n2266 = ~n2263 & ~n2265_1;
  assign n2267 = P1_DATAO_REG_19_ & n1734;
  assign n2268 = P2_DATAO_REG_19_ & ~n1734;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270_1 = SI_19_ & n2269;
  assign n2271 = ~SI_19_ & ~n2269;
  assign n2272 = ~n2270_1 & ~n2271;
  assign n2273 = n2266 & ~n2272;
  assign n2274 = ~n2266 & n2272;
  assign n2275_1 = ~n2273 & ~n2274;
  assign n2276 = ~n1734 & ~n2275_1;
  assign n2277 = ~n2262 & ~n2276;
  assign n2278 = ~P1_STATE_REG & ~n2277;
  assign n2279 = ~n2260_1 & ~n2261;
  assign n205 = n2278 | ~n2279;
  assign n2281 = P1_IR_REG_20_ & ~n2258;
  assign n2282 = ~P1_IR_REG_13_ & ~P1_IR_REG_15_;
  assign n2283 = ~P1_IR_REG_14_ & n2282;
  assign n2284 = ~P1_IR_REG_10_ & ~P1_IR_REG_12_;
  assign n2285_1 = ~P1_IR_REG_11_ & n2284;
  assign n2286 = ~P1_IR_REG_1_ & ~P1_IR_REG_19_;
  assign n2287 = ~P1_IR_REG_18_ & n2286;
  assign n2288 = ~P1_IR_REG_16_ & n2287;
  assign n2289 = ~P1_IR_REG_17_ & n2288;
  assign n2290_1 = ~P1_IR_REG_0_ & n2249;
  assign n2291 = ~P1_IR_REG_20_ & n2290_1;
  assign n2292 = n2283 & n2285_1;
  assign n2293 = n2289 & n2292;
  assign n2294 = n2248 & n2293;
  assign n2295_1 = n2291 & n2294;
  assign n2296 = ~n2281 & ~n2295_1;
  assign n2297 = n1727 & n2296;
  assign n2298 = P1_IR_REG_20_ & n1726;
  assign n2299 = P2_DATAO_REG_20_ & n1734;
  assign n2300_1 = SI_19_ & ~n2269;
  assign n2301 = ~SI_19_ & n2269;
  assign n2302 = ~n2266 & ~n2301;
  assign n2303 = ~n2300_1 & ~n2302;
  assign n2304 = P1_DATAO_REG_20_ & n1734;
  assign n2305_1 = P2_DATAO_REG_20_ & ~n1734;
  assign n2306 = ~n2304 & ~n2305_1;
  assign n2307 = SI_20_ & n2306;
  assign n2308 = ~SI_20_ & ~n2306;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310_1 = n2303 & ~n2309;
  assign n2311 = ~n2303 & n2309;
  assign n2312 = ~n2310_1 & ~n2311;
  assign n2313 = ~n1734 & ~n2312;
  assign n2314 = ~n2299 & ~n2313;
  assign n2315_1 = ~P1_STATE_REG & ~n2314;
  assign n2316 = ~n2297 & ~n2298;
  assign n210 = n2315_1 | ~n2316;
  assign n2318 = ~P1_IR_REG_21_ & n2295_1;
  assign n2319 = P1_IR_REG_21_ & ~n2295_1;
  assign n2320_1 = ~n2318 & ~n2319;
  assign n2321 = n1727 & n2320_1;
  assign n2322 = P1_IR_REG_21_ & n1726;
  assign n2323 = P2_DATAO_REG_21_ & n1734;
  assign n2324 = SI_20_ & ~n2306;
  assign n2325_1 = ~SI_20_ & n2306;
  assign n2326 = ~n2303 & ~n2325_1;
  assign n2327 = ~n2324 & ~n2326;
  assign n2328 = P1_DATAO_REG_21_ & n1734;
  assign n2329 = P2_DATAO_REG_21_ & ~n1734;
  assign n2330_1 = ~n2328 & ~n2329;
  assign n2331 = SI_21_ & n2330_1;
  assign n2332 = ~SI_21_ & ~n2330_1;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = n2327 & ~n2333;
  assign n2335_1 = ~n2327 & n2333;
  assign n2336 = ~n2334 & ~n2335_1;
  assign n2337 = ~n1734 & ~n2336;
  assign n2338 = ~n2323 & ~n2337;
  assign n2339 = ~P1_STATE_REG & ~n2338;
  assign n2340_1 = ~n2321 & ~n2322;
  assign n215 = n2339 | ~n2340_1;
  assign n2342 = ~P1_IR_REG_2_ & ~P1_IR_REG_4_;
  assign n2343 = ~P1_IR_REG_3_ & n2342;
  assign n2344 = ~P1_IR_REG_0_ & ~P1_IR_REG_21_;
  assign n2345_1 = ~P1_IR_REG_20_ & n2344;
  assign n2346 = n2343 & n2345_1;
  assign n2347 = n2248 & n2346;
  assign n2348 = n2289 & n2347;
  assign n2349 = n2292 & n2348;
  assign n2350_1 = P1_IR_REG_22_ & ~n2349;
  assign n2351 = ~P1_IR_REG_19_ & ~P1_IR_REG_20_;
  assign n2352 = ~P1_IR_REG_17_ & ~P1_IR_REG_18_;
  assign n2353 = ~P1_IR_REG_21_ & ~P1_IR_REG_22_;
  assign n2354 = n2351 & n2352;
  assign n2355_1 = n2353 & n2354;
  assign n2356 = n2163 & n2355_1;
  assign n2357 = ~n2350_1 & ~n2356;
  assign n2358 = n1727 & n2357;
  assign n2359 = P1_IR_REG_22_ & n1726;
  assign n2360_1 = P2_DATAO_REG_22_ & n1734;
  assign n2361 = SI_21_ & ~n2330_1;
  assign n2362 = ~SI_21_ & n2330_1;
  assign n2363 = ~n2327 & ~n2362;
  assign n2364 = ~n2361 & ~n2363;
  assign n2365_1 = P1_DATAO_REG_22_ & n1734;
  assign n2366 = P2_DATAO_REG_22_ & ~n1734;
  assign n2367 = ~n2365_1 & ~n2366;
  assign n2368 = SI_22_ & n2367;
  assign n2369 = ~SI_22_ & ~n2367;
  assign n2370_1 = ~n2368 & ~n2369;
  assign n2371 = n2364 & ~n2370_1;
  assign n2372 = ~n2364 & n2370_1;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~n1734 & ~n2373;
  assign n2375_1 = ~n2360_1 & ~n2374;
  assign n2376 = ~P1_STATE_REG & ~n2375_1;
  assign n2377 = ~n2358 & ~n2359;
  assign n220 = n2376 | ~n2377;
  assign n2379 = P1_IR_REG_23_ & ~n2356;
  assign n2380_1 = ~P1_IR_REG_7_ & ~P1_IR_REG_9_;
  assign n2381 = ~P1_IR_REG_8_ & n2380_1;
  assign n2382 = ~P1_IR_REG_4_ & ~P1_IR_REG_6_;
  assign n2383 = ~P1_IR_REG_5_ & n2382;
  assign n2384 = ~P1_IR_REG_3_ & ~P1_IR_REG_23_;
  assign n2385_1 = ~P1_IR_REG_2_ & n2384;
  assign n2386 = ~P1_IR_REG_20_ & ~P1_IR_REG_22_;
  assign n2387 = ~P1_IR_REG_21_ & n2386;
  assign n2388 = n2381 & n2383;
  assign n2389 = n2385_1 & n2388;
  assign n2390_1 = n2387 & n2389;
  assign n2391 = ~P1_IR_REG_0_ & ~P1_IR_REG_19_;
  assign n2392 = ~P1_IR_REG_1_ & n2391;
  assign n2393 = ~P1_IR_REG_16_ & ~P1_IR_REG_18_;
  assign n2394 = ~P1_IR_REG_17_ & n2393;
  assign n2395_1 = n2392 & n2394;
  assign n2396 = n2283 & n2395_1;
  assign n2397 = n2285_1 & n2396;
  assign n2398 = n2390_1 & n2397;
  assign n2399 = ~n2379 & ~n2398;
  assign n2400_1 = n1727 & n2399;
  assign n2401 = P1_IR_REG_23_ & n1726;
  assign n2402 = P2_DATAO_REG_23_ & n1734;
  assign n2403 = SI_22_ & ~n2367;
  assign n2404 = ~SI_22_ & n2367;
  assign n2405_1 = ~n2364 & ~n2404;
  assign n2406 = ~n2403 & ~n2405_1;
  assign n2407 = P1_DATAO_REG_23_ & n1734;
  assign n2408 = P2_DATAO_REG_23_ & ~n1734;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410_1 = SI_23_ & n2409;
  assign n2411 = ~SI_23_ & ~n2409;
  assign n2412 = ~n2410_1 & ~n2411;
  assign n2413 = n2406 & ~n2412;
  assign n2414 = ~n2406 & n2412;
  assign n2415_1 = ~n2413 & ~n2414;
  assign n2416 = ~n1734 & ~n2415_1;
  assign n2417 = ~n2402 & ~n2416;
  assign n2418 = ~P1_STATE_REG & ~n2417;
  assign n2419 = ~n2400_1 & ~n2401;
  assign n225 = n2418 | ~n2419;
  assign n2421 = P1_IR_REG_24_ & ~n2398;
  assign n2422 = ~P1_IR_REG_3_ & ~P1_IR_REG_24_;
  assign n2423 = ~P1_IR_REG_2_ & n2422;
  assign n2424 = ~P1_IR_REG_21_ & ~P1_IR_REG_23_;
  assign n2425_1 = ~P1_IR_REG_22_ & n2424;
  assign n2426 = n2388 & n2423;
  assign n2427 = n2425_1 & n2426;
  assign n2428 = ~P1_IR_REG_1_ & ~P1_IR_REG_20_;
  assign n2429 = ~P1_IR_REG_0_ & n2428;
  assign n2430_1 = ~P1_IR_REG_17_ & ~P1_IR_REG_19_;
  assign n2431 = ~P1_IR_REG_18_ & n2430_1;
  assign n2432 = ~P1_IR_REG_14_ & ~P1_IR_REG_16_;
  assign n2433 = ~P1_IR_REG_15_ & n2432;
  assign n2434 = ~P1_IR_REG_13_ & n2041;
  assign n2435_1 = n2429 & n2431;
  assign n2436 = n2433 & n2435_1;
  assign n2437 = n2434 & n2436;
  assign n2438 = n2427 & n2437;
  assign n2439 = ~n2421 & ~n2438;
  assign n2440_1 = n1727 & n2439;
  assign n2441 = P1_IR_REG_24_ & n1726;
  assign n2442 = P2_DATAO_REG_24_ & n1734;
  assign n2443 = SI_23_ & ~n2409;
  assign n2444 = ~SI_23_ & n2409;
  assign n2445_1 = ~n2406 & ~n2444;
  assign n2446 = ~n2443 & ~n2445_1;
  assign n2447 = P1_DATAO_REG_24_ & n1734;
  assign n2448 = P2_DATAO_REG_24_ & ~n1734;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450_1 = SI_24_ & n2449;
  assign n2451 = ~SI_24_ & ~n2449;
  assign n2452 = ~n2450_1 & ~n2451;
  assign n2453 = n2446 & ~n2452;
  assign n2454 = ~n2446 & n2452;
  assign n2455_1 = ~n2453 & ~n2454;
  assign n2456 = ~n1734 & ~n2455_1;
  assign n2457 = ~n2442 & ~n2456;
  assign n2458 = ~P1_STATE_REG & ~n2457;
  assign n2459 = ~n2440_1 & ~n2441;
  assign n230 = n2458 | ~n2459;
  assign n2461 = ~P1_IR_REG_25_ & n2438;
  assign n2462 = P1_IR_REG_25_ & ~n2438;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = n1727 & n2463;
  assign n2465_1 = P1_IR_REG_25_ & n1726;
  assign n2466 = P2_DATAO_REG_25_ & n1734;
  assign n2467 = SI_24_ & ~n2449;
  assign n2468 = ~SI_24_ & n2449;
  assign n2469 = ~n2446 & ~n2468;
  assign n2470_1 = ~n2467 & ~n2469;
  assign n2471 = P1_DATAO_REG_25_ & n1734;
  assign n2472 = P2_DATAO_REG_25_ & ~n1734;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = SI_25_ & n2473;
  assign n2475_1 = ~SI_25_ & ~n2473;
  assign n2476 = ~n2474 & ~n2475_1;
  assign n2477 = n2470_1 & ~n2476;
  assign n2478 = ~n2470_1 & n2476;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480_1 = ~n1734 & ~n2479;
  assign n2481 = ~n2466 & ~n2480_1;
  assign n2482 = ~P1_STATE_REG & ~n2481;
  assign n2483 = ~n2464 & ~n2465_1;
  assign n235 = n2482 | ~n2483;
  assign n2485_1 = ~P1_IR_REG_3_ & ~P1_IR_REG_25_;
  assign n2486 = ~P1_IR_REG_2_ & n2485_1;
  assign n2487 = ~P1_IR_REG_23_ & n2353;
  assign n2488 = ~P1_IR_REG_24_ & n2487;
  assign n2489 = n2388 & n2486;
  assign n2490_1 = n2488 & n2489;
  assign n2491 = n2437 & n2490_1;
  assign n2492 = P1_IR_REG_26_ & ~n2491;
  assign n2493 = ~P1_IR_REG_3_ & ~P1_IR_REG_26_;
  assign n2494 = ~P1_IR_REG_2_ & n2493;
  assign n2495_1 = ~P1_IR_REG_22_ & ~P1_IR_REG_23_;
  assign n2496 = ~P1_IR_REG_24_ & n2495_1;
  assign n2497 = ~P1_IR_REG_25_ & n2496;
  assign n2498 = n2388 & n2494;
  assign n2499 = n2497 & n2498;
  assign n2500_1 = ~P1_IR_REG_19_ & n2352;
  assign n2501 = ~P1_IR_REG_1_ & n2500_1;
  assign n2502 = n2345_1 & n2501;
  assign n2503 = n2433 & n2502;
  assign n2504 = n2434 & n2503;
  assign n2505_1 = n2499 & n2504;
  assign n2506 = ~n2492 & ~n2505_1;
  assign n2507 = n1727 & n2506;
  assign n2508 = P1_IR_REG_26_ & n1726;
  assign n2509 = P2_DATAO_REG_26_ & n1734;
  assign n2510_1 = SI_25_ & ~n2473;
  assign n2511 = ~SI_25_ & n2473;
  assign n2512 = ~n2470_1 & ~n2511;
  assign n2513 = ~n2510_1 & ~n2512;
  assign n2514 = P1_DATAO_REG_26_ & n1734;
  assign n2515_1 = P2_DATAO_REG_26_ & ~n1734;
  assign n2516 = ~n2514 & ~n2515_1;
  assign n2517 = SI_26_ & n2516;
  assign n2518 = ~SI_26_ & ~n2516;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520_1 = n2513 & ~n2519;
  assign n2521 = ~n2513 & n2519;
  assign n2522 = ~n2520_1 & ~n2521;
  assign n2523 = ~n1734 & ~n2522;
  assign n2524 = ~n2509 & ~n2523;
  assign n2525_1 = ~P1_STATE_REG & ~n2524;
  assign n2526 = ~n2507 & ~n2508;
  assign n240 = n2525_1 | ~n2526;
  assign n2528 = ~P1_IR_REG_27_ & ~n2505_1;
  assign n2529 = P1_IR_REG_27_ & n2505_1;
  assign n2530_1 = ~n2528 & ~n2529;
  assign n2531 = n1727 & ~n2530_1;
  assign n2532 = P1_IR_REG_27_ & n1726;
  assign n2533 = P2_DATAO_REG_27_ & n1734;
  assign n2534 = SI_26_ & ~n2516;
  assign n2535_1 = ~SI_26_ & n2516;
  assign n2536 = ~n2513 & ~n2535_1;
  assign n2537 = ~n2534 & ~n2536;
  assign n2538 = P1_DATAO_REG_27_ & n1734;
  assign n2539 = P2_DATAO_REG_27_ & ~n1734;
  assign n2540_1 = ~n2538 & ~n2539;
  assign n2541 = SI_27_ & n2540_1;
  assign n2542 = ~SI_27_ & ~n2540_1;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = n2537 & ~n2543;
  assign n2545_1 = ~n2537 & n2543;
  assign n2546 = ~n2544 & ~n2545_1;
  assign n2547 = ~n1734 & ~n2546;
  assign n2548 = ~n2533 & ~n2547;
  assign n2549 = ~P1_STATE_REG & ~n2548;
  assign n2550_1 = ~n2531 & ~n2532;
  assign n245 = n2549 | ~n2550_1;
  assign n2552 = ~P1_IR_REG_2_ & ~P1_IR_REG_26_;
  assign n2553 = ~P1_IR_REG_27_ & n2552;
  assign n2554 = n1932 & n2381;
  assign n2555_1 = n2553 & n2554;
  assign n2556 = n2497 & n2555_1;
  assign n2557 = n2504 & n2556;
  assign n2558 = P1_IR_REG_28_ & ~n2557;
  assign n2559 = ~P1_IR_REG_2_ & ~P1_IR_REG_27_;
  assign n2560 = ~P1_IR_REG_28_ & n2559;
  assign n2561 = ~P1_IR_REG_23_ & ~P1_IR_REG_24_;
  assign n2562 = ~P1_IR_REG_25_ & n2561;
  assign n2563 = ~P1_IR_REG_26_ & n2562;
  assign n2564 = n2554 & n2560;
  assign n2565 = n2563 & n2564;
  assign n2566 = ~P1_IR_REG_1_ & n2252;
  assign n2567 = ~P1_IR_REG_0_ & n2566;
  assign n2568 = ~P1_IR_REG_14_ & ~P1_IR_REG_15_;
  assign n2569 = ~P1_IR_REG_16_ & n2568;
  assign n2570 = ~P1_IR_REG_17_ & n2569;
  assign n2571 = n2387 & n2567;
  assign n2572 = n2570 & n2571;
  assign n2573 = n2434 & n2572;
  assign n2574 = n2565 & n2573;
  assign n2575 = ~n2558 & ~n2574;
  assign n2576 = n1727 & n2575;
  assign n2577 = P1_IR_REG_28_ & n1726;
  assign n2578 = P2_DATAO_REG_28_ & n1734;
  assign n2579 = SI_27_ & ~n2540_1;
  assign n2580 = ~SI_27_ & n2540_1;
  assign n2581 = ~n2537 & ~n2580;
  assign n2582 = ~n2579 & ~n2581;
  assign n2583 = P1_DATAO_REG_28_ & n1734;
  assign n2584 = P2_DATAO_REG_28_ & ~n1734;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = SI_28_ & n2585;
  assign n2587 = ~SI_28_ & ~n2585;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = n2582 & ~n2588;
  assign n2590 = ~n2582 & n2588;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = ~n1734 & ~n2591;
  assign n2593 = ~n2578 & ~n2592;
  assign n2594 = ~P1_STATE_REG & ~n2593;
  assign n2595 = ~n2576 & ~n2577;
  assign n250 = n2594 | ~n2595;
  assign n2597 = P1_IR_REG_29_ & ~n2574;
  assign n2598 = ~P1_IR_REG_27_ & ~P1_IR_REG_28_;
  assign n2599 = ~P1_IR_REG_29_ & n2598;
  assign n2600 = ~P1_IR_REG_2_ & n2599;
  assign n2601 = n2554 & n2600;
  assign n2602 = n2563 & n2601;
  assign n2603 = n2573 & n2602;
  assign n2604 = ~n2597 & ~n2603;
  assign n2605 = n1727 & n2604;
  assign n2606 = P1_IR_REG_29_ & n1726;
  assign n2607 = P2_DATAO_REG_29_ & n1734;
  assign n2608 = SI_28_ & ~n2585;
  assign n2609 = ~SI_28_ & n2585;
  assign n2610 = ~n2582 & ~n2609;
  assign n2611 = ~n2608 & ~n2610;
  assign n2612 = P1_DATAO_REG_29_ & n1734;
  assign n2613 = P2_DATAO_REG_29_ & ~n1734;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = SI_29_ & n2614;
  assign n2616 = ~SI_29_ & ~n2614;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = n2611 & ~n2617;
  assign n2619 = ~n2611 & n2617;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = ~n1734 & ~n2620;
  assign n2622 = ~n2607 & ~n2621;
  assign n2623 = ~P1_STATE_REG & ~n2622;
  assign n2624 = ~n2605 & ~n2606;
  assign n255 = n2623 | ~n2624;
  assign n2626 = ~P1_IR_REG_30_ & n2603;
  assign n2627 = P1_IR_REG_30_ & ~n2603;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n1727 & n2628;
  assign n2630 = P1_IR_REG_30_ & n1726;
  assign n2631 = P2_DATAO_REG_30_ & n1734;
  assign n2632 = SI_29_ & ~n2614;
  assign n2633 = ~SI_29_ & n2614;
  assign n2634 = ~n2611 & ~n2633;
  assign n2635 = ~n2632 & ~n2634;
  assign n2636 = P1_DATAO_REG_30_ & n1734;
  assign n2637 = P2_DATAO_REG_30_ & ~n1734;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = SI_30_ & n2638;
  assign n2640 = ~SI_30_ & ~n2638;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = n2635 & ~n2641;
  assign n2643 = ~n2635 & n2641;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = ~n1734 & ~n2644;
  assign n2646 = ~n2631 & ~n2645;
  assign n2647 = ~P1_STATE_REG & ~n2646;
  assign n2648 = ~n2629 & ~n2630;
  assign n260 = n2647 | ~n2648;
  assign n2650 = P1_IR_REG_31_ & n2626;
  assign n2651 = ~P1_IR_REG_31_ & ~n2626;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = n1727 & ~n2652;
  assign n2654 = P1_IR_REG_31_ & n1726;
  assign n2655 = P2_DATAO_REG_31_ & n1734;
  assign n2656 = P1_DATAO_REG_31_ & n1734;
  assign n2657 = P2_DATAO_REG_31_ & ~n1734;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = SI_31_ & n2658;
  assign n2660 = ~SI_31_ & ~n2658;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = SI_30_ & ~n2661;
  assign n2663 = ~n2638 & n2662;
  assign n2664 = ~SI_30_ & n2661;
  assign n2665 = n2638 & n2664;
  assign n2666 = ~n2663 & ~n2665;
  assign n2667 = SI_30_ & ~n2638;
  assign n2668 = n2661 & ~n2667;
  assign n2669 = ~n2632 & n2668;
  assign n2670 = ~n2634 & n2669;
  assign n2671 = n2666 & ~n2670;
  assign n2672 = ~SI_30_ & n2638;
  assign n2673 = ~n2661 & ~n2672;
  assign n2674 = ~n2635 & n2673;
  assign n2675 = n2671 & ~n2674;
  assign n2676 = ~n1734 & n2675;
  assign n2677 = ~n2655 & ~n2676;
  assign n2678 = ~P1_STATE_REG & ~n2677;
  assign n2679 = ~n2653 & ~n2654;
  assign n265 = n2678 | ~n2679;
  assign n2681 = P1_IR_REG_31_ & n2399;
  assign n2682 = P1_IR_REG_23_ & ~P1_IR_REG_31_;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = P1_IR_REG_31_ & n2439;
  assign n2685 = P1_IR_REG_24_ & ~P1_IR_REG_31_;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = P1_IR_REG_31_ & n2506;
  assign n2688 = P1_IR_REG_26_ & ~P1_IR_REG_31_;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2686 & ~n2689;
  assign n2691 = P1_IR_REG_31_ & n2463;
  assign n2692 = P1_IR_REG_25_ & ~P1_IR_REG_31_;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = n2690 & ~n2693;
  assign n2695 = n2683 & ~n2694;
  assign n2696 = P1_STATE_REG & n2695;
  assign n2697 = ~n2689 & n2693;
  assign n2698 = n2686 & n2697;
  assign n2699 = P1_B_REG & n2698;
  assign n2700 = ~P1_B_REG & n2690;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = ~n2689 & n2701;
  assign n2703 = n2696 & ~n2702;
  assign n2704 = n2686 & ~n2697;
  assign n2705 = n2703 & ~n2704;
  assign n2706 = P1_D_REG_0_ & ~n2703;
  assign n270 = n2705 | n2706;
  assign n2708 = n2693 & ~n2697;
  assign n2709 = n2703 & ~n2708;
  assign n2710 = P1_D_REG_1_ & ~n2703;
  assign n275 = n2709 | n2710;
  assign n280 = P1_D_REG_2_ & ~n2703;
  assign n285 = P1_D_REG_3_ & ~n2703;
  assign n290 = P1_D_REG_4_ & ~n2703;
  assign n295 = P1_D_REG_5_ & ~n2703;
  assign n300 = P1_D_REG_6_ & ~n2703;
  assign n305 = P1_D_REG_7_ & ~n2703;
  assign n310 = P1_D_REG_8_ & ~n2703;
  assign n315 = P1_D_REG_9_ & ~n2703;
  assign n320 = P1_D_REG_10_ & ~n2703;
  assign n325 = P1_D_REG_11_ & ~n2703;
  assign n330 = P1_D_REG_12_ & ~n2703;
  assign n335 = P1_D_REG_13_ & ~n2703;
  assign n340 = P1_D_REG_14_ & ~n2703;
  assign n345 = P1_D_REG_15_ & ~n2703;
  assign n350 = P1_D_REG_16_ & ~n2703;
  assign n355 = P1_D_REG_17_ & ~n2703;
  assign n360 = P1_D_REG_18_ & ~n2703;
  assign n365 = P1_D_REG_19_ & ~n2703;
  assign n370 = P1_D_REG_20_ & ~n2703;
  assign n375 = P1_D_REG_21_ & ~n2703;
  assign n380 = P1_D_REG_22_ & ~n2703;
  assign n385 = P1_D_REG_23_ & ~n2703;
  assign n390 = P1_D_REG_24_ & ~n2703;
  assign n395 = P1_D_REG_25_ & ~n2703;
  assign n400 = P1_D_REG_26_ & ~n2703;
  assign n405 = P1_D_REG_27_ & ~n2703;
  assign n410 = P1_D_REG_28_ & ~n2703;
  assign n415 = P1_D_REG_29_ & ~n2703;
  assign n420 = P1_D_REG_30_ & ~n2703;
  assign n425 = P1_D_REG_31_ & ~n2703;
  assign n2742 = P1_D_REG_0_ & n2702;
  assign n2743 = n2686 & n2689;
  assign n2744 = ~n2702 & ~n2743;
  assign n2745 = ~n2742 & ~n2744;
  assign n2746 = n2696 & n2745;
  assign n2747 = ~n2702 & ~n2708;
  assign n2748 = P1_D_REG_1_ & n2702;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = P1_IR_REG_31_ & n2357;
  assign n2751 = P1_IR_REG_22_ & ~P1_IR_REG_31_;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = P1_IR_REG_31_ & n2296;
  assign n2754 = P1_IR_REG_20_ & ~P1_IR_REG_31_;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = P1_IR_REG_31_ & n2320_1;
  assign n2757 = P1_IR_REG_21_ & ~P1_IR_REG_31_;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = n2755 & n2758;
  assign n2760 = n2752 & ~n2759;
  assign n2761 = ~n2752 & n2758;
  assign n2762 = P1_IR_REG_31_ & n2259;
  assign n2763 = P1_IR_REG_19_ & ~P1_IR_REG_31_;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n2755 & n2764;
  assign n2766 = ~n2760 & ~n2761;
  assign n2767 = ~n2765 & n2766;
  assign n2768 = n2749 & ~n2767;
  assign n2769 = P1_D_REG_8_ & n2702;
  assign n2770 = P1_D_REG_7_ & n2702;
  assign n2771 = P1_D_REG_9_ & n2702;
  assign n2772 = ~n2769 & ~n2770;
  assign n2773 = ~n2771 & n2772;
  assign n2774 = P1_D_REG_6_ & n2702;
  assign n2775 = P1_D_REG_5_ & n2702;
  assign n2776 = P1_D_REG_4_ & n2702;
  assign n2777 = P1_D_REG_3_ & n2702;
  assign n2778 = ~n2774 & ~n2775;
  assign n2779 = ~n2776 & n2778;
  assign n2780 = ~n2777 & n2779;
  assign n2781 = P1_D_REG_31_ & n2702;
  assign n2782 = P1_D_REG_30_ & n2702;
  assign n2783 = P1_D_REG_2_ & n2702;
  assign n2784 = P1_D_REG_29_ & n2702;
  assign n2785 = ~n2781 & ~n2782;
  assign n2786 = ~n2783 & n2785;
  assign n2787 = ~n2784 & n2786;
  assign n2788 = P1_D_REG_28_ & n2702;
  assign n2789 = P1_D_REG_27_ & n2702;
  assign n2790 = P1_D_REG_26_ & n2702;
  assign n2791 = P1_D_REG_25_ & n2702;
  assign n2792 = ~n2788 & ~n2789;
  assign n2793 = ~n2790 & n2792;
  assign n2794 = ~n2791 & n2793;
  assign n2795 = n2773 & n2780;
  assign n2796 = n2787 & n2795;
  assign n2797 = n2794 & n2796;
  assign n2798 = P1_D_REG_23_ & n2702;
  assign n2799 = P1_D_REG_22_ & n2702;
  assign n2800 = P1_D_REG_24_ & n2702;
  assign n2801 = ~n2798 & ~n2799;
  assign n2802 = ~n2800 & n2801;
  assign n2803 = P1_D_REG_21_ & n2702;
  assign n2804 = P1_D_REG_20_ & n2702;
  assign n2805 = P1_D_REG_19_ & n2702;
  assign n2806 = P1_D_REG_18_ & n2702;
  assign n2807 = ~n2803 & ~n2804;
  assign n2808 = ~n2805 & n2807;
  assign n2809 = ~n2806 & n2808;
  assign n2810 = P1_D_REG_17_ & n2702;
  assign n2811 = P1_D_REG_16_ & n2702;
  assign n2812 = P1_D_REG_15_ & n2702;
  assign n2813 = P1_D_REG_14_ & n2702;
  assign n2814 = ~n2810 & ~n2811;
  assign n2815 = ~n2812 & n2814;
  assign n2816 = ~n2813 & n2815;
  assign n2817 = P1_D_REG_13_ & n2702;
  assign n2818 = P1_D_REG_12_ & n2702;
  assign n2819 = P1_D_REG_11_ & n2702;
  assign n2820 = P1_D_REG_10_ & n2702;
  assign n2821 = ~n2817 & ~n2818;
  assign n2822 = ~n2819 & n2821;
  assign n2823 = ~n2820 & n2822;
  assign n2824 = n2802 & n2809;
  assign n2825 = n2816 & n2824;
  assign n2826 = n2823 & n2825;
  assign n2827 = n2797 & n2826;
  assign n2828 = n2768 & n2827;
  assign n2829 = n2746 & n2828;
  assign n2830 = ~n2752 & ~n2758;
  assign n2831 = P1_IR_REG_31_ & n2575;
  assign n2832 = P1_IR_REG_28_ & ~P1_IR_REG_31_;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = n2830 & n2833;
  assign n2835 = P1_IR_REG_31_ & n2628;
  assign n2836 = P1_IR_REG_30_ & ~P1_IR_REG_31_;
  assign n2837 = ~n2835 & ~n2836;
  assign n2838 = P1_IR_REG_31_ & n2604;
  assign n2839 = P1_IR_REG_29_ & ~P1_IR_REG_31_;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = ~n2837 & ~n2840;
  assign n2842 = P1_REG3_REG_1_ & n2841;
  assign n2843 = n2837 & n2840;
  assign n2844 = P1_REG0_REG_1_ & n2843;
  assign n2845 = n2837 & ~n2840;
  assign n2846 = P1_REG1_REG_1_ & n2845;
  assign n2847 = ~n2837 & n2840;
  assign n2848 = P1_REG2_REG_1_ & n2847;
  assign n2849 = ~n2842 & ~n2844;
  assign n2850 = ~n2846 & n2849;
  assign n2851 = ~n2848 & n2850;
  assign n2852 = n2834 & ~n2851;
  assign n2853 = P1_IR_REG_31_ & ~n2530_1;
  assign n2854 = P1_IR_REG_27_ & ~P1_IR_REG_31_;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = n2833 & n2855;
  assign n2857 = P1_IR_REG_0_ & P1_IR_REG_31_;
  assign n2858 = P1_IR_REG_0_ & ~P1_IR_REG_31_;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = n2856 & ~n2859;
  assign n2861 = ~n1743 & ~n2856;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n2752 & n2758;
  assign n2864 = n2755 & n2863;
  assign n2865 = ~n2862 & n2864;
  assign n2866 = ~n2755 & n2764;
  assign n2867 = n2863 & n2866;
  assign n2868 = n2752 & ~n2764;
  assign n2869 = n2758 & n2868;
  assign n2870 = ~n2867 & ~n2869;
  assign n2871 = ~n2862 & ~n2870;
  assign n2872 = P1_REG3_REG_0_ & n2841;
  assign n2873 = P1_REG2_REG_0_ & n2847;
  assign n2874 = P1_REG1_REG_0_ & n2845;
  assign n2875 = P1_REG0_REG_0_ & n2843;
  assign n2876 = ~n2872 & ~n2873;
  assign n2877 = ~n2874 & n2876;
  assign n2878 = ~n2875 & n2877;
  assign n2879 = ~n2862 & n2878;
  assign n2880 = n2862 & ~n2878;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = n2755 & n2868;
  assign n2883 = ~n2881 & n2882;
  assign n2884 = ~n2852 & ~n2865;
  assign n2885 = ~n2871 & n2884;
  assign n2886 = ~n2883 & n2885;
  assign n2887 = ~n2752 & n2765;
  assign n2888 = n2758 & n2887;
  assign n2889 = ~n2881 & n2888;
  assign n2890 = ~n2758 & n2866;
  assign n2891 = ~n2881 & n2890;
  assign n2892 = ~n2758 & n2765;
  assign n2893 = n2752 & n2892;
  assign n2894 = ~n2881 & n2893;
  assign n2895 = ~n2755 & ~n2764;
  assign n2896 = ~n2758 & n2895;
  assign n2897 = ~n2881 & n2896;
  assign n2898 = ~n2752 & n2866;
  assign n2899 = ~n2881 & n2898;
  assign n2900 = ~n2897 & ~n2899;
  assign n2901 = ~n2752 & n2895;
  assign n2902 = ~n2881 & n2901;
  assign n2903 = n2755 & ~n2764;
  assign n2904 = ~n2752 & n2903;
  assign n2905 = ~n2881 & n2904;
  assign n2906 = ~n2902 & ~n2905;
  assign n2907 = ~n2889 & ~n2891;
  assign n2908 = ~n2894 & n2907;
  assign n2909 = n2900 & n2908;
  assign n2910 = n2906 & n2909;
  assign n2911 = n2886 & n2910;
  assign n2912 = n2829 & ~n2911;
  assign n2913 = P1_REG0_REG_0_ & ~n2829;
  assign n430 = n2912 | n2913;
  assign n2915 = P1_REG3_REG_2_ & n2841;
  assign n2916 = P1_REG0_REG_2_ & n2843;
  assign n2917 = P1_REG1_REG_2_ & n2845;
  assign n2918 = P1_REG2_REG_2_ & n2847;
  assign n2919 = ~n2915 & ~n2916;
  assign n2920 = ~n2917 & n2919;
  assign n2921 = ~n2918 & n2920;
  assign n2922 = n2834 & ~n2921;
  assign n2923 = P1_IR_REG_31_ & ~n1749;
  assign n2924 = P1_IR_REG_1_ & ~P1_IR_REG_31_;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = n2856 & ~n2925;
  assign n2927 = ~n1769 & ~n2856;
  assign n2928 = ~n2926 & ~n2927;
  assign n2929 = ~n2862 & n2928;
  assign n2930 = n2862 & ~n2928;
  assign n2931 = ~n2929 & ~n2930;
  assign n2932 = n2864 & ~n2931;
  assign n2933 = ~n2870 & ~n2928;
  assign n2934 = ~n2851 & ~n2928;
  assign n2935 = n2851 & n2928;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = ~n2862 & ~n2878;
  assign n2938 = n2936 & ~n2937;
  assign n2939 = ~n2936 & n2937;
  assign n2940 = ~n2938 & ~n2939;
  assign n2941 = n2882 & ~n2940;
  assign n2942 = ~n2922 & ~n2932;
  assign n2943 = ~n2933 & n2942;
  assign n2944 = ~n2941 & n2943;
  assign n2945 = ~n2851 & ~n2879;
  assign n2946 = n2851 & n2879;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = n2928 & ~n2947;
  assign n2949 = ~n2928 & n2947;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n2904 & ~n2950;
  assign n2952 = n2830 & ~n2833;
  assign n2953 = ~n2878 & n2952;
  assign n2954 = n2898 & ~n2940;
  assign n2955 = n2901 & ~n2950;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = n2893 & ~n2940;
  assign n2958 = n2888 & ~n2940;
  assign n2959 = n2890 & ~n2950;
  assign n2960 = n2896 & ~n2950;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = ~n2957 & ~n2958;
  assign n2963 = n2961 & n2962;
  assign n2964 = ~n2951 & ~n2953;
  assign n2965 = n2956 & n2964;
  assign n2966 = n2963 & n2965;
  assign n2967 = n2944 & n2966;
  assign n2968 = n2829 & ~n2967;
  assign n2969 = P1_REG0_REG_1_ & ~n2829;
  assign n435 = n2968 | n2969;
  assign n2971 = ~P1_REG3_REG_3_ & n2841;
  assign n2972 = P1_REG0_REG_3_ & n2843;
  assign n2973 = P1_REG1_REG_3_ & n2845;
  assign n2974 = P1_REG2_REG_3_ & n2847;
  assign n2975 = ~n2971 & ~n2972;
  assign n2976 = ~n2973 & n2975;
  assign n2977 = ~n2974 & n2976;
  assign n2978 = n2834 & ~n2977;
  assign n2979 = P1_IR_REG_31_ & n1776;
  assign n2980 = P1_IR_REG_2_ & ~P1_IR_REG_31_;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = n2856 & ~n2981;
  assign n2983 = ~n1794 & ~n2856;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = n2862 & n2928;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = n2862 & n2984;
  assign n2988 = n2928 & n2987;
  assign n2989 = ~n2986 & ~n2988;
  assign n2990 = n2864 & n2989;
  assign n2991 = ~n2870 & ~n2984;
  assign n2992 = ~n2921 & ~n2984;
  assign n2993 = n2921 & n2984;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2935 & n2937;
  assign n2996 = ~n2934 & ~n2995;
  assign n2997 = n2994 & ~n2996;
  assign n2998 = n2921 & ~n2984;
  assign n2999 = ~n2921 & n2984;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = ~n2934 & n3000;
  assign n3002 = ~n2995 & n3001;
  assign n3003 = ~n2997 & ~n3002;
  assign n3004 = n2882 & n3003;
  assign n3005 = ~n2978 & ~n2990;
  assign n3006 = ~n2991 & n3005;
  assign n3007 = ~n3004 & n3006;
  assign n3008 = n2928 & ~n2946;
  assign n3009 = ~n2945 & ~n3008;
  assign n3010 = n3000 & n3009;
  assign n3011 = ~n3000 & ~n3009;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = n2904 & ~n3012;
  assign n3014 = ~n2851 & n2952;
  assign n3015 = n2898 & n3003;
  assign n3016 = n2901 & ~n3012;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = n2893 & n3003;
  assign n3019 = n2888 & n3003;
  assign n3020 = n2890 & ~n3012;
  assign n3021 = n2896 & ~n3012;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = ~n3018 & ~n3019;
  assign n3024 = n3022 & n3023;
  assign n3025 = ~n3013 & ~n3014;
  assign n3026 = n3017 & n3025;
  assign n3027 = n3024 & n3026;
  assign n3028 = n3007 & n3027;
  assign n3029 = n2829 & ~n3028;
  assign n3030 = P1_REG0_REG_2_ & ~n2829;
  assign n440 = n3029 | n3030;
  assign n3032 = ~P1_REG3_REG_4_ & P1_REG3_REG_3_;
  assign n3033 = P1_REG3_REG_4_ & ~P1_REG3_REG_3_;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = n2841 & ~n3034;
  assign n3036 = P1_REG0_REG_4_ & n2843;
  assign n3037 = P1_REG1_REG_4_ & n2845;
  assign n3038 = P1_REG2_REG_4_ & n2847;
  assign n3039 = ~n3035 & ~n3036;
  assign n3040 = ~n3037 & n3039;
  assign n3041 = ~n3038 & n3040;
  assign n3042 = n2834 & ~n3041;
  assign n3043 = P1_IR_REG_31_ & n1800_1;
  assign n3044 = P1_IR_REG_3_ & ~P1_IR_REG_31_;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n2856 & ~n3045;
  assign n3047 = ~n1818 & ~n2856;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = ~n2988 & ~n3048;
  assign n3050 = n2988 & n3048;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n2864 & n3051;
  assign n3053 = ~n2870 & ~n3048;
  assign n3054 = n2934 & ~n2993;
  assign n3055 = ~n2992 & ~n3054;
  assign n3056 = ~n2993 & n2995;
  assign n3057 = n3055 & ~n3056;
  assign n3058 = n2977 & ~n3048;
  assign n3059 = ~n2977 & n3048;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = n3057 & ~n3060;
  assign n3062 = ~n2977 & ~n3048;
  assign n3063 = n2977 & n3048;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = ~n3057 & ~n3064;
  assign n3066 = ~n3061 & ~n3065;
  assign n3067 = n2882 & ~n3066;
  assign n3068 = ~n3042 & ~n3052;
  assign n3069 = ~n3053 & n3068;
  assign n3070 = ~n3067 & n3069;
  assign n3071 = ~n2998 & ~n3060;
  assign n3072 = ~n2999 & n3009;
  assign n3073 = n3071 & ~n3072;
  assign n3074 = ~n2999 & n3060;
  assign n3075 = ~n2998 & ~n3009;
  assign n3076 = n3074 & ~n3075;
  assign n3077 = ~n3073 & ~n3076;
  assign n3078 = n2904 & ~n3077;
  assign n3079 = ~n2921 & n2952;
  assign n3080 = n2901 & ~n3077;
  assign n3081 = n2898 & ~n3066;
  assign n3082 = n2893 & ~n3066;
  assign n3083 = n2888 & ~n3066;
  assign n3084 = n2890 & ~n3077;
  assign n3085 = n2896 & ~n3077;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~n3082 & ~n3083;
  assign n3088 = n3086 & n3087;
  assign n3089 = ~n3078 & ~n3079;
  assign n3090 = ~n3080 & n3089;
  assign n3091 = ~n3081 & n3090;
  assign n3092 = n3088 & n3091;
  assign n3093 = n3070 & n3092;
  assign n3094 = n2829 & ~n3093;
  assign n3095 = P1_REG0_REG_3_ & ~n2829;
  assign n445 = n3094 | n3095;
  assign n3097 = P1_REG3_REG_4_ & P1_REG3_REG_3_;
  assign n3098 = ~P1_REG3_REG_5_ & n3097;
  assign n3099 = P1_REG3_REG_5_ & ~n3097;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = n2841 & ~n3100;
  assign n3102 = P1_REG0_REG_5_ & n2843;
  assign n3103 = P1_REG1_REG_5_ & n2845;
  assign n3104 = P1_REG2_REG_5_ & n2847;
  assign n3105 = ~n3101 & ~n3102;
  assign n3106 = ~n3103 & n3105;
  assign n3107 = ~n3104 & n3106;
  assign n3108 = n2834 & ~n3107;
  assign n3109 = P1_IR_REG_31_ & n1825_1;
  assign n3110 = P1_IR_REG_4_ & ~P1_IR_REG_31_;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = n2856 & ~n3111;
  assign n3113 = ~n1846 & ~n2856;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~n3050 & ~n3114;
  assign n3116 = n3050 & n3114;
  assign n3117 = ~n3115 & ~n3116;
  assign n3118 = n2864 & n3117;
  assign n3119 = ~n2870 & ~n3114;
  assign n3120 = n3041 & ~n3114;
  assign n3121 = ~n3041 & n3114;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = ~n2993 & ~n3063;
  assign n3124 = n2995 & n3123;
  assign n3125 = ~n3062 & ~n3124;
  assign n3126 = ~n3055 & ~n3063;
  assign n3127 = n3125 & ~n3126;
  assign n3128 = ~n3122 & n3127;
  assign n3129 = n3041 & n3114;
  assign n3130 = ~n3041 & ~n3114;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = ~n3127 & ~n3131;
  assign n3133 = ~n3128 & ~n3132;
  assign n3134 = n2882 & ~n3133;
  assign n3135 = ~n3108 & ~n3118;
  assign n3136 = ~n3119 & n3135;
  assign n3137 = ~n3134 & n3136;
  assign n3138 = n2977 & ~n2999;
  assign n3139 = n3048 & ~n3138;
  assign n3140 = ~n2977 & n2999;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n3058 & n3075;
  assign n3143 = n3141 & ~n3142;
  assign n3144 = n3122 & n3143;
  assign n3145 = ~n3122 & ~n3143;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = n2904 & ~n3146;
  assign n3148 = n2952 & ~n2977;
  assign n3149 = n2901 & ~n3146;
  assign n3150 = n2898 & ~n3133;
  assign n3151 = n2893 & ~n3133;
  assign n3152 = n2888 & ~n3133;
  assign n3153 = n2890 & ~n3146;
  assign n3154 = n2896 & ~n3146;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3151 & ~n3152;
  assign n3157 = n3155 & n3156;
  assign n3158 = ~n3147 & ~n3148;
  assign n3159 = ~n3149 & n3158;
  assign n3160 = ~n3150 & n3159;
  assign n3161 = n3157 & n3160;
  assign n3162 = n3137 & n3161;
  assign n3163 = n2829 & ~n3162;
  assign n3164 = P1_REG0_REG_4_ & ~n2829;
  assign n450 = n3163 | n3164;
  assign n3166 = P1_REG3_REG_5_ & n3097;
  assign n3167 = ~P1_REG3_REG_6_ & n3166;
  assign n3168 = P1_REG3_REG_6_ & ~n3166;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = n2841 & ~n3169;
  assign n3171 = P1_REG0_REG_6_ & n2843;
  assign n3172 = P1_REG1_REG_6_ & n2845;
  assign n3173 = P1_REG2_REG_6_ & n2847;
  assign n3174 = ~n3170 & ~n3171;
  assign n3175 = ~n3172 & n3174;
  assign n3176 = ~n3173 & n3175;
  assign n3177 = n2834 & ~n3176;
  assign n3178 = P1_IR_REG_31_ & n1852;
  assign n3179 = P1_IR_REG_5_ & ~P1_IR_REG_31_;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = n2856 & ~n3180;
  assign n3182 = ~n1870_1 & ~n2856;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = n3116 & n3183;
  assign n3185 = ~n3116 & ~n3183;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = n2864 & n3186;
  assign n3188 = ~n2870 & ~n3183;
  assign n3189 = ~n3107 & ~n3183;
  assign n3190 = n3107 & n3183;
  assign n3191 = ~n3129 & ~n3190;
  assign n3192 = ~n3189 & n3191;
  assign n3193 = n3127 & ~n3130;
  assign n3194 = n3192 & ~n3193;
  assign n3195 = n3107 & ~n3183;
  assign n3196 = ~n3107 & n3183;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3130 & n3197;
  assign n3199 = ~n3127 & ~n3129;
  assign n3200 = n3198 & ~n3199;
  assign n3201 = ~n3194 & ~n3200;
  assign n3202 = n2882 & n3201;
  assign n3203 = ~n3177 & ~n3187;
  assign n3204 = ~n3188 & n3203;
  assign n3205 = ~n3202 & n3204;
  assign n3206 = ~n3120 & ~n3143;
  assign n3207 = ~n3121 & ~n3206;
  assign n3208 = n3197 & n3207;
  assign n3209 = ~n3197 & ~n3207;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n2904 & ~n3210;
  assign n3212 = n2952 & ~n3041;
  assign n3213 = n2898 & n3201;
  assign n3214 = n2901 & ~n3210;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = n2893 & n3201;
  assign n3217 = n2888 & n3201;
  assign n3218 = n2890 & ~n3210;
  assign n3219 = n2896 & ~n3210;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = ~n3216 & ~n3217;
  assign n3222 = n3220 & n3221;
  assign n3223 = ~n3211 & ~n3212;
  assign n3224 = n3215 & n3223;
  assign n3225 = n3222 & n3224;
  assign n3226 = n3205 & n3225;
  assign n3227 = n2829 & ~n3226;
  assign n3228 = P1_REG0_REG_5_ & ~n2829;
  assign n455 = n3227 | n3228;
  assign n3230 = P1_REG3_REG_6_ & n3166;
  assign n3231 = ~P1_REG3_REG_7_ & n3230;
  assign n3232 = P1_REG3_REG_7_ & ~n3230;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = n2841 & ~n3233;
  assign n3235 = P1_REG0_REG_7_ & n2843;
  assign n3236 = P1_REG1_REG_7_ & n2845;
  assign n3237 = P1_REG2_REG_7_ & n2847;
  assign n3238 = ~n3234 & ~n3235;
  assign n3239 = ~n3236 & n3238;
  assign n3240 = ~n3237 & n3239;
  assign n3241 = n2834 & ~n3240;
  assign n3242 = P1_IR_REG_31_ & n1877;
  assign n3243 = P1_IR_REG_6_ & ~P1_IR_REG_31_;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = n2856 & ~n3244;
  assign n3246 = ~n1898 & ~n2856;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = ~n3184 & ~n3247;
  assign n3249 = n3183 & n3247;
  assign n3250 = n3116 & n3249;
  assign n3251 = ~n3248 & ~n3250;
  assign n3252 = n2864 & n3251;
  assign n3253 = ~n2870 & ~n3247;
  assign n3254 = n3176 & ~n3247;
  assign n3255 = ~n3176 & n3247;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = n3130 & ~n3183;
  assign n3258 = ~n3130 & n3183;
  assign n3259 = ~n3107 & ~n3258;
  assign n3260 = ~n3257 & ~n3259;
  assign n3261 = n2992 & ~n3063;
  assign n3262 = ~n3062 & ~n3261;
  assign n3263 = ~n2996 & n3123;
  assign n3264 = n3262 & ~n3263;
  assign n3265 = n3191 & ~n3264;
  assign n3266 = n3260 & ~n3265;
  assign n3267 = ~n3256 & n3266;
  assign n3268 = n3176 & n3247;
  assign n3269 = ~n3176 & ~n3247;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~n3266 & ~n3270;
  assign n3272 = ~n3267 & ~n3271;
  assign n3273 = n2882 & ~n3272;
  assign n3274 = ~n3241 & ~n3252;
  assign n3275 = ~n3253 & n3274;
  assign n3276 = ~n3273 & n3275;
  assign n3277 = ~n3195 & ~n3256;
  assign n3278 = ~n3196 & n3207;
  assign n3279 = n3277 & ~n3278;
  assign n3280 = ~n3196 & ~n3255;
  assign n3281 = ~n3254 & n3280;
  assign n3282 = ~n3195 & ~n3207;
  assign n3283 = n3281 & ~n3282;
  assign n3284 = ~n3279 & ~n3283;
  assign n3285 = n2904 & ~n3284;
  assign n3286 = n2952 & ~n3107;
  assign n3287 = n2898 & ~n3272;
  assign n3288 = n2901 & ~n3284;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = n2893 & ~n3272;
  assign n3291 = n2888 & ~n3272;
  assign n3292 = n2890 & ~n3284;
  assign n3293 = n2896 & ~n3284;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = ~n3290 & ~n3291;
  assign n3296 = n3294 & n3295;
  assign n3297 = ~n3285 & ~n3286;
  assign n3298 = n3289 & n3297;
  assign n3299 = n3296 & n3298;
  assign n3300 = n3276 & n3299;
  assign n3301 = n2829 & ~n3300;
  assign n3302 = P1_REG0_REG_6_ & ~n2829;
  assign n460 = n3301 | n3302;
  assign n3304 = P1_REG3_REG_7_ & n3230;
  assign n3305 = ~P1_REG3_REG_8_ & n3304;
  assign n3306 = P1_REG3_REG_8_ & ~n3304;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = n2841 & ~n3307;
  assign n3309 = P1_REG0_REG_8_ & n2843;
  assign n3310 = P1_REG1_REG_8_ & n2845;
  assign n3311 = P1_REG2_REG_8_ & n2847;
  assign n3312 = ~n3308 & ~n3309;
  assign n3313 = ~n3310 & n3312;
  assign n3314 = ~n3311 & n3313;
  assign n3315 = n2834 & ~n3314;
  assign n3316 = P1_IR_REG_31_ & n1904;
  assign n3317 = P1_IR_REG_7_ & ~P1_IR_REG_31_;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = n2856 & ~n3318;
  assign n3320 = ~n1925_1 & ~n2856;
  assign n3321 = ~n3319 & ~n3320;
  assign n3322 = ~n3250 & ~n3321;
  assign n3323 = n3250 & n3321;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = n2864 & n3324;
  assign n3326 = ~n2870 & ~n3321;
  assign n3327 = ~n3240 & ~n3321;
  assign n3328 = n3240 & n3321;
  assign n3329 = ~n3268 & ~n3328;
  assign n3330 = ~n3327 & n3329;
  assign n3331 = n3266 & ~n3269;
  assign n3332 = n3330 & ~n3331;
  assign n3333 = n3240 & ~n3321;
  assign n3334 = ~n3240 & n3321;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3269 & n3335;
  assign n3337 = ~n3266 & ~n3268;
  assign n3338 = n3336 & ~n3337;
  assign n3339 = ~n3332 & ~n3338;
  assign n3340 = n2882 & n3339;
  assign n3341 = ~n3315 & ~n3325;
  assign n3342 = ~n3326 & n3341;
  assign n3343 = ~n3340 & n3342;
  assign n3344 = n3121 & ~n3195;
  assign n3345 = n3280 & ~n3344;
  assign n3346 = ~n3254 & ~n3345;
  assign n3347 = ~n3120 & ~n3254;
  assign n3348 = ~n3143 & ~n3195;
  assign n3349 = n3347 & n3348;
  assign n3350 = ~n3346 & ~n3349;
  assign n3351 = n3335 & n3350;
  assign n3352 = ~n3335 & ~n3350;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = n2904 & ~n3353;
  assign n3355 = n2952 & ~n3176;
  assign n3356 = n2898 & n3339;
  assign n3357 = n2901 & ~n3353;
  assign n3358 = ~n3356 & ~n3357;
  assign n3359 = n2893 & n3339;
  assign n3360 = n2888 & n3339;
  assign n3361 = n2890 & ~n3353;
  assign n3362 = n2896 & ~n3353;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = ~n3359 & ~n3360;
  assign n3365 = n3363 & n3364;
  assign n3366 = ~n3354 & ~n3355;
  assign n3367 = n3358 & n3366;
  assign n3368 = n3365 & n3367;
  assign n3369 = n3343 & n3368;
  assign n3370 = n2829 & ~n3369;
  assign n3371 = P1_REG0_REG_7_ & ~n2829;
  assign n465 = n3370 | n3371;
  assign n3373 = P1_REG1_REG_9_ & n2845;
  assign n3374 = P1_REG0_REG_9_ & n2843;
  assign n3375 = P1_REG2_REG_9_ & n2847;
  assign n3376 = P1_REG3_REG_8_ & n3304;
  assign n3377 = ~P1_REG3_REG_9_ & n3376;
  assign n3378 = P1_REG3_REG_9_ & ~n3376;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = n2841 & ~n3379;
  assign n3381 = ~n3373 & ~n3374;
  assign n3382 = ~n3375 & n3381;
  assign n3383 = ~n3380 & n3382;
  assign n3384 = n2834 & ~n3383;
  assign n3385 = P1_IR_REG_31_ & n1935_1;
  assign n3386 = P1_IR_REG_8_ & ~P1_IR_REG_31_;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = n2856 & ~n3387;
  assign n3389 = ~n1953 & ~n2856;
  assign n3390 = ~n3388 & ~n3389;
  assign n3391 = ~n3323 & ~n3390;
  assign n3392 = n3323 & n3390;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = n2864 & n3393;
  assign n3395 = ~n2870 & ~n3390;
  assign n3396 = n3269 & ~n3321;
  assign n3397 = ~n3269 & n3321;
  assign n3398 = ~n3240 & ~n3397;
  assign n3399 = ~n3396 & ~n3398;
  assign n3400 = ~n3266 & n3329;
  assign n3401 = n3399 & ~n3400;
  assign n3402 = n3314 & ~n3390;
  assign n3403 = ~n3314 & n3390;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3401 & ~n3404;
  assign n3406 = n3314 & n3390;
  assign n3407 = ~n3314 & ~n3390;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = ~n3401 & ~n3408;
  assign n3410 = ~n3405 & ~n3409;
  assign n3411 = n2882 & ~n3410;
  assign n3412 = ~n3384 & ~n3394;
  assign n3413 = ~n3395 & n3412;
  assign n3414 = ~n3411 & n3413;
  assign n3415 = ~n3333 & ~n3404;
  assign n3416 = ~n3334 & n3350;
  assign n3417 = n3415 & ~n3416;
  assign n3418 = ~n3334 & n3404;
  assign n3419 = ~n3333 & ~n3350;
  assign n3420 = n3418 & ~n3419;
  assign n3421 = ~n3417 & ~n3420;
  assign n3422 = n2904 & ~n3421;
  assign n3423 = n2952 & ~n3240;
  assign n3424 = n2898 & ~n3410;
  assign n3425 = n2901 & ~n3421;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = n2893 & ~n3410;
  assign n3428 = n2888 & ~n3410;
  assign n3429 = n2890 & ~n3421;
  assign n3430 = n2896 & ~n3421;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = ~n3427 & ~n3428;
  assign n3433 = n3431 & n3432;
  assign n3434 = ~n3422 & ~n3423;
  assign n3435 = n3426 & n3434;
  assign n3436 = n3433 & n3435;
  assign n3437 = n3414 & n3436;
  assign n3438 = n2829 & ~n3437;
  assign n3439 = P1_REG0_REG_8_ & ~n2829;
  assign n470 = n3438 | n3439;
  assign n3441 = P1_REG1_REG_10_ & n2845;
  assign n3442 = P1_REG0_REG_10_ & n2843;
  assign n3443 = P1_REG2_REG_10_ & n2847;
  assign n3444 = P1_REG3_REG_9_ & n3376;
  assign n3445 = ~P1_REG3_REG_10_ & n3444;
  assign n3446 = P1_REG3_REG_10_ & ~n3444;
  assign n3447 = ~n3445 & ~n3446;
  assign n3448 = n2841 & ~n3447;
  assign n3449 = ~n3441 & ~n3442;
  assign n3450 = ~n3443 & n3449;
  assign n3451 = ~n3448 & n3450;
  assign n3452 = n2834 & ~n3451;
  assign n3453 = P1_IR_REG_31_ & n1959;
  assign n3454 = P1_IR_REG_9_ & ~P1_IR_REG_31_;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = n2856 & ~n3455;
  assign n3457 = ~n1980_1 & ~n2856;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = n3392 & n3458;
  assign n3460 = ~n3392 & ~n3458;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = n2864 & n3461;
  assign n3463 = ~n2870 & ~n3458;
  assign n3464 = n3383 & ~n3458;
  assign n3465 = ~n3383 & n3458;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = ~n3401 & ~n3406;
  assign n3468 = ~n3407 & ~n3467;
  assign n3469 = ~n3466 & n3468;
  assign n3470 = n3383 & n3458;
  assign n3471 = ~n3383 & ~n3458;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = ~n3468 & ~n3472;
  assign n3474 = ~n3469 & ~n3473;
  assign n3475 = n2882 & ~n3474;
  assign n3476 = ~n3452 & ~n3462;
  assign n3477 = ~n3463 & n3476;
  assign n3478 = ~n3475 & n3477;
  assign n3479 = n3314 & ~n3334;
  assign n3480 = n3390 & ~n3479;
  assign n3481 = ~n3314 & n3334;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = ~n3333 & ~n3402;
  assign n3484 = ~n3350 & n3483;
  assign n3485 = n3482 & ~n3484;
  assign n3486 = n3466 & n3485;
  assign n3487 = ~n3466 & ~n3485;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = n2904 & ~n3488;
  assign n3490 = n2952 & ~n3314;
  assign n3491 = n2898 & ~n3474;
  assign n3492 = n2901 & ~n3488;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = n2893 & ~n3474;
  assign n3495 = n2888 & ~n3474;
  assign n3496 = n2890 & ~n3488;
  assign n3497 = n2896 & ~n3488;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = ~n3494 & ~n3495;
  assign n3500 = n3498 & n3499;
  assign n3501 = ~n3489 & ~n3490;
  assign n3502 = n3493 & n3501;
  assign n3503 = n3500 & n3502;
  assign n3504 = n3478 & n3503;
  assign n3505 = n2829 & ~n3504;
  assign n3506 = P1_REG0_REG_9_ & ~n2829;
  assign n475 = n3505 | n3506;
  assign n3508 = P1_REG1_REG_11_ & n2845;
  assign n3509 = P1_REG0_REG_11_ & n2843;
  assign n3510 = P1_REG2_REG_11_ & n2847;
  assign n3511 = P1_REG3_REG_10_ & n3444;
  assign n3512 = ~P1_REG3_REG_11_ & n3511;
  assign n3513 = P1_REG3_REG_11_ & ~n3511;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n2841 & ~n3514;
  assign n3516 = ~n3508 & ~n3509;
  assign n3517 = ~n3510 & n3516;
  assign n3518 = ~n3515 & n3517;
  assign n3519 = n2834 & ~n3518;
  assign n3520 = P1_IR_REG_31_ & n1987;
  assign n3521 = P1_IR_REG_10_ & ~P1_IR_REG_31_;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n2856 & ~n3522;
  assign n3524 = ~n2008 & ~n2856;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = ~n3459 & ~n3525;
  assign n3527 = n3458 & n3525;
  assign n3528 = n3392 & n3527;
  assign n3529 = ~n3526 & ~n3528;
  assign n3530 = n2864 & n3529;
  assign n3531 = ~n2870 & ~n3525;
  assign n3532 = ~n3451 & ~n3525;
  assign n3533 = n3451 & n3525;
  assign n3534 = ~n3470 & ~n3533;
  assign n3535 = ~n3532 & n3534;
  assign n3536 = n3468 & ~n3471;
  assign n3537 = n3535 & ~n3536;
  assign n3538 = n3451 & ~n3525;
  assign n3539 = ~n3451 & n3525;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~n3471 & n3540;
  assign n3542 = ~n3468 & ~n3470;
  assign n3543 = n3541 & ~n3542;
  assign n3544 = ~n3537 & ~n3543;
  assign n3545 = n2882 & n3544;
  assign n3546 = ~n3519 & ~n3530;
  assign n3547 = ~n3531 & n3546;
  assign n3548 = ~n3545 & n3547;
  assign n3549 = ~n3464 & ~n3485;
  assign n3550 = ~n3465 & ~n3549;
  assign n3551 = n3540 & n3550;
  assign n3552 = ~n3540 & ~n3550;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = n2904 & ~n3553;
  assign n3555 = n2952 & ~n3383;
  assign n3556 = n2898 & n3544;
  assign n3557 = n2901 & ~n3553;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = n2893 & n3544;
  assign n3560 = n2888 & n3544;
  assign n3561 = n2890 & ~n3553;
  assign n3562 = n2896 & ~n3553;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n3559 & ~n3560;
  assign n3565 = n3563 & n3564;
  assign n3566 = ~n3554 & ~n3555;
  assign n3567 = n3558 & n3566;
  assign n3568 = n3565 & n3567;
  assign n3569 = n3548 & n3568;
  assign n3570 = n2829 & ~n3569;
  assign n3571 = P1_REG0_REG_10_ & ~n2829;
  assign n480 = n3570 | n3571;
  assign n3573 = P1_IR_REG_31_ & n2014;
  assign n3574 = P1_IR_REG_11_ & ~P1_IR_REG_31_;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = n2856 & ~n3575;
  assign n3577 = ~n2035_1 & ~n2856;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = ~n2870 & ~n3578;
  assign n3580 = ~n3471 & ~n3532;
  assign n3581 = n3407 & n3534;
  assign n3582 = n3580 & ~n3581;
  assign n3583 = ~n3533 & ~n3582;
  assign n3584 = ~n3406 & n3534;
  assign n3585 = ~n3401 & n3584;
  assign n3586 = ~n3583 & ~n3585;
  assign n3587 = n3518 & ~n3578;
  assign n3588 = ~n3518 & n3578;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = n3586 & ~n3589;
  assign n3591 = n3518 & n3578;
  assign n3592 = ~n3518 & ~n3578;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = ~n3586 & ~n3593;
  assign n3595 = ~n3590 & ~n3594;
  assign n3596 = n2882 & ~n3595;
  assign n3597 = P1_REG1_REG_12_ & n2845;
  assign n3598 = P1_REG0_REG_12_ & n2843;
  assign n3599 = P1_REG2_REG_12_ & n2847;
  assign n3600 = P1_REG3_REG_11_ & n3511;
  assign n3601 = ~P1_REG3_REG_12_ & n3600;
  assign n3602 = P1_REG3_REG_12_ & ~n3600;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = n2841 & ~n3603;
  assign n3605 = ~n3597 & ~n3598;
  assign n3606 = ~n3599 & n3605;
  assign n3607 = ~n3604 & n3606;
  assign n3608 = n2834 & ~n3607;
  assign n3609 = ~n3528 & ~n3578;
  assign n3610 = n3528 & n3578;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = n2864 & n3611;
  assign n3613 = ~n3579 & ~n3596;
  assign n3614 = ~n3608 & n3613;
  assign n3615 = ~n3612 & n3614;
  assign n3616 = ~n3538 & ~n3589;
  assign n3617 = ~n3539 & n3550;
  assign n3618 = n3616 & ~n3617;
  assign n3619 = ~n3539 & ~n3588;
  assign n3620 = ~n3587 & n3619;
  assign n3621 = ~n3538 & ~n3550;
  assign n3622 = n3620 & ~n3621;
  assign n3623 = ~n3618 & ~n3622;
  assign n3624 = n2904 & ~n3623;
  assign n3625 = n2952 & ~n3451;
  assign n3626 = n2898 & ~n3595;
  assign n3627 = n2901 & ~n3623;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = n2893 & ~n3595;
  assign n3630 = n2888 & ~n3595;
  assign n3631 = n2890 & ~n3623;
  assign n3632 = n2896 & ~n3623;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = ~n3629 & ~n3630;
  assign n3635 = n3633 & n3634;
  assign n3636 = ~n3624 & ~n3625;
  assign n3637 = n3628 & n3636;
  assign n3638 = n3635 & n3637;
  assign n3639 = n3615 & n3638;
  assign n3640 = n2829 & ~n3639;
  assign n3641 = P1_REG0_REG_11_ & ~n2829;
  assign n485 = n3640 | n3641;
  assign n3643 = P1_IR_REG_31_ & n2044;
  assign n3644 = P1_IR_REG_12_ & ~P1_IR_REG_31_;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = n2856 & ~n3645;
  assign n3647 = ~n2062 & ~n2856;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = ~n2870 & ~n3648;
  assign n3650 = n3607 & ~n3648;
  assign n3651 = ~n3607 & n3648;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = ~n3586 & ~n3591;
  assign n3654 = ~n3592 & ~n3653;
  assign n3655 = ~n3652 & n3654;
  assign n3656 = n3607 & n3648;
  assign n3657 = ~n3607 & ~n3648;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = ~n3654 & ~n3658;
  assign n3660 = ~n3655 & ~n3659;
  assign n3661 = n2882 & ~n3660;
  assign n3662 = P1_REG1_REG_13_ & n2845;
  assign n3663 = P1_REG0_REG_13_ & n2843;
  assign n3664 = P1_REG2_REG_13_ & n2847;
  assign n3665 = P1_REG3_REG_12_ & n3600;
  assign n3666 = ~P1_REG3_REG_13_ & n3665;
  assign n3667 = P1_REG3_REG_13_ & ~n3665;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = n2841 & ~n3668;
  assign n3670 = ~n3662 & ~n3663;
  assign n3671 = ~n3664 & n3670;
  assign n3672 = ~n3669 & n3671;
  assign n3673 = n2834 & ~n3672;
  assign n3674 = ~n3610 & ~n3648;
  assign n3675 = n3610 & n3648;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = n2864 & n3676;
  assign n3678 = ~n3649 & ~n3661;
  assign n3679 = ~n3673 & n3678;
  assign n3680 = ~n3677 & n3679;
  assign n3681 = n3465 & ~n3538;
  assign n3682 = n3619 & ~n3681;
  assign n3683 = ~n3587 & ~n3682;
  assign n3684 = ~n3464 & ~n3587;
  assign n3685 = ~n3538 & n3684;
  assign n3686 = ~n3485 & n3685;
  assign n3687 = ~n3683 & ~n3686;
  assign n3688 = ~n3652 & ~n3687;
  assign n3689 = n3652 & n3687;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = n2904 & ~n3690;
  assign n3692 = n2952 & ~n3518;
  assign n3693 = n2898 & ~n3660;
  assign n3694 = n2901 & ~n3690;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = n2893 & ~n3660;
  assign n3697 = n2888 & ~n3660;
  assign n3698 = n2890 & ~n3690;
  assign n3699 = n2896 & ~n3690;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3696 & ~n3697;
  assign n3702 = n3700 & n3701;
  assign n3703 = ~n3691 & ~n3692;
  assign n3704 = n3695 & n3703;
  assign n3705 = n3702 & n3704;
  assign n3706 = n3680 & n3705;
  assign n3707 = n2829 & ~n3706;
  assign n3708 = P1_REG0_REG_12_ & ~n2829;
  assign n490 = n3707 | n3708;
  assign n3710 = P1_IR_REG_31_ & n2068;
  assign n3711 = P1_IR_REG_13_ & ~P1_IR_REG_31_;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = n2856 & ~n3712;
  assign n3714 = ~n2089 & ~n2856;
  assign n3715 = ~n3713 & ~n3714;
  assign n3716 = ~n2870 & ~n3715;
  assign n3717 = n3675 & n3715;
  assign n3718 = ~n3675 & ~n3715;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = n2864 & n3719;
  assign n3721 = P1_REG1_REG_14_ & n2845;
  assign n3722 = P1_REG0_REG_14_ & n2843;
  assign n3723 = P1_REG2_REG_14_ & n2847;
  assign n3724 = P1_REG3_REG_13_ & n3665;
  assign n3725 = ~P1_REG3_REG_14_ & n3724;
  assign n3726 = P1_REG3_REG_14_ & ~n3724;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = n2841 & ~n3727;
  assign n3729 = ~n3721 & ~n3722;
  assign n3730 = ~n3723 & n3729;
  assign n3731 = ~n3728 & n3730;
  assign n3732 = n2834 & ~n3731;
  assign n3733 = ~n3672 & ~n3715;
  assign n3734 = n3672 & n3715;
  assign n3735 = ~n3656 & ~n3734;
  assign n3736 = ~n3733 & n3735;
  assign n3737 = n3654 & ~n3657;
  assign n3738 = n3736 & ~n3737;
  assign n3739 = n3672 & ~n3715;
  assign n3740 = ~n3672 & n3715;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = ~n3657 & n3741;
  assign n3743 = ~n3654 & ~n3656;
  assign n3744 = n3742 & ~n3743;
  assign n3745 = ~n3738 & ~n3744;
  assign n3746 = n2882 & n3745;
  assign n3747 = ~n3716 & ~n3720;
  assign n3748 = ~n3732 & n3747;
  assign n3749 = ~n3746 & n3748;
  assign n3750 = ~n3650 & ~n3687;
  assign n3751 = ~n3651 & ~n3750;
  assign n3752 = ~n3741 & ~n3751;
  assign n3753 = n3741 & n3751;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = n2904 & ~n3754;
  assign n3756 = n2952 & ~n3607;
  assign n3757 = n2898 & n3745;
  assign n3758 = n2901 & ~n3754;
  assign n3759 = ~n3757 & ~n3758;
  assign n3760 = n2893 & n3745;
  assign n3761 = n2888 & n3745;
  assign n3762 = n2890 & ~n3754;
  assign n3763 = n2896 & ~n3754;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = ~n3760 & ~n3761;
  assign n3766 = n3764 & n3765;
  assign n3767 = ~n3755 & ~n3756;
  assign n3768 = n3759 & n3767;
  assign n3769 = n3766 & n3768;
  assign n3770 = n3749 & n3769;
  assign n3771 = n2829 & ~n3770;
  assign n3772 = P1_REG0_REG_13_ & ~n2829;
  assign n495 = n3771 | n3772;
  assign n3774 = P1_REG1_REG_15_ & n2845;
  assign n3775 = P1_REG0_REG_15_ & n2843;
  assign n3776 = P1_REG2_REG_15_ & n2847;
  assign n3777 = P1_REG3_REG_14_ & n3724;
  assign n3778 = ~P1_REG3_REG_15_ & n3777;
  assign n3779 = P1_REG3_REG_15_ & ~n3777;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = n2841 & ~n3780;
  assign n3782 = ~n3774 & ~n3775;
  assign n3783 = ~n3776 & n3782;
  assign n3784 = ~n3781 & n3783;
  assign n3785 = n2834 & ~n3784;
  assign n3786 = ~n3657 & ~n3733;
  assign n3787 = n3592 & n3735;
  assign n3788 = n3786 & ~n3787;
  assign n3789 = ~n3734 & ~n3788;
  assign n3790 = ~n3591 & n3735;
  assign n3791 = ~n3586 & n3790;
  assign n3792 = ~n3789 & ~n3791;
  assign n3793 = P1_IR_REG_31_ & n2096;
  assign n3794 = P1_IR_REG_14_ & ~P1_IR_REG_31_;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n2856 & ~n3795;
  assign n3797 = ~n2117 & ~n2856;
  assign n3798 = ~n3796 & ~n3797;
  assign n3799 = n3731 & ~n3798;
  assign n3800 = ~n3731 & n3798;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = n3792 & ~n3801;
  assign n3803 = ~n3792 & n3801;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = n2882 & ~n3804;
  assign n3806 = ~n2870 & ~n3798;
  assign n3807 = ~n3717 & ~n3798;
  assign n3808 = n3715 & n3798;
  assign n3809 = n3675 & n3808;
  assign n3810 = ~n3807 & ~n3809;
  assign n3811 = n2864 & n3810;
  assign n3812 = ~n3785 & ~n3805;
  assign n3813 = ~n3806 & n3812;
  assign n3814 = ~n3811 & n3813;
  assign n3815 = ~n3739 & ~n3751;
  assign n3816 = ~n3740 & ~n3815;
  assign n3817 = n3801 & n3816;
  assign n3818 = ~n3801 & ~n3816;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = n2904 & ~n3819;
  assign n3821 = n2952 & ~n3672;
  assign n3822 = n2898 & ~n3804;
  assign n3823 = n2901 & ~n3819;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n2893 & ~n3804;
  assign n3826 = n2888 & ~n3804;
  assign n3827 = n2890 & ~n3819;
  assign n3828 = n2896 & ~n3819;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~n3825 & ~n3826;
  assign n3831 = n3829 & n3830;
  assign n3832 = ~n3820 & ~n3821;
  assign n3833 = n3824 & n3832;
  assign n3834 = n3831 & n3833;
  assign n3835 = n3814 & n3834;
  assign n3836 = n2829 & ~n3835;
  assign n3837 = P1_REG0_REG_14_ & ~n2829;
  assign n500 = n3836 | n3837;
  assign n3839 = P1_REG1_REG_16_ & n2845;
  assign n3840 = P1_REG0_REG_16_ & n2843;
  assign n3841 = P1_REG2_REG_16_ & n2847;
  assign n3842 = P1_REG3_REG_15_ & n3777;
  assign n3843 = ~P1_REG3_REG_16_ & n3842;
  assign n3844 = P1_REG3_REG_16_ & ~n3842;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = n2841 & ~n3845;
  assign n3847 = ~n3839 & ~n3840;
  assign n3848 = ~n3841 & n3847;
  assign n3849 = ~n3846 & n3848;
  assign n3850 = n2834 & ~n3849;
  assign n3851 = ~n3731 & ~n3798;
  assign n3852 = n3731 & n3798;
  assign n3853 = ~n3792 & ~n3852;
  assign n3854 = ~n3851 & ~n3853;
  assign n3855 = P1_IR_REG_31_ & n2123;
  assign n3856 = P1_IR_REG_15_ & ~P1_IR_REG_31_;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = n2856 & ~n3857;
  assign n3859 = ~n2144 & ~n2856;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = n3784 & ~n3860;
  assign n3862 = ~n3784 & n3860;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = n3854 & ~n3863;
  assign n3865 = ~n3854 & n3863;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n2882 & ~n3866;
  assign n3868 = ~n2870 & ~n3860;
  assign n3869 = ~n3809 & ~n3860;
  assign n3870 = n3809 & n3860;
  assign n3871 = ~n3869 & ~n3870;
  assign n3872 = n2864 & n3871;
  assign n3873 = ~n3850 & ~n3867;
  assign n3874 = ~n3868 & n3873;
  assign n3875 = ~n3872 & n3874;
  assign n3876 = ~n3799 & ~n3816;
  assign n3877 = ~n3800 & ~n3876;
  assign n3878 = n3863 & n3877;
  assign n3879 = ~n3863 & ~n3877;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = n2904 & ~n3880;
  assign n3882 = n2952 & ~n3731;
  assign n3883 = n2898 & ~n3866;
  assign n3884 = n2901 & ~n3880;
  assign n3885 = ~n3883 & ~n3884;
  assign n3886 = n2893 & ~n3866;
  assign n3887 = n2888 & ~n3866;
  assign n3888 = n2890 & ~n3880;
  assign n3889 = n2896 & ~n3880;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~n3886 & ~n3887;
  assign n3892 = n3890 & n3891;
  assign n3893 = ~n3881 & ~n3882;
  assign n3894 = n3885 & n3893;
  assign n3895 = n3892 & n3894;
  assign n3896 = n3875 & n3895;
  assign n3897 = n2829 & ~n3896;
  assign n3898 = P1_REG0_REG_15_ & ~n2829;
  assign n505 = n3897 | n3898;
  assign n3900 = P1_REG1_REG_17_ & n2845;
  assign n3901 = P1_REG0_REG_17_ & n2843;
  assign n3902 = P1_REG2_REG_17_ & n2847;
  assign n3903 = P1_REG3_REG_16_ & n3842;
  assign n3904 = ~P1_REG3_REG_17_ & n3903;
  assign n3905 = P1_REG3_REG_17_ & ~n3903;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = n2841 & ~n3906;
  assign n3908 = ~n3900 & ~n3901;
  assign n3909 = ~n3902 & n3908;
  assign n3910 = ~n3907 & n3909;
  assign n3911 = n2834 & ~n3910;
  assign n3912 = P1_IR_REG_31_ & n2164;
  assign n3913 = P1_IR_REG_16_ & ~P1_IR_REG_31_;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = n2856 & ~n3914;
  assign n3916 = ~n2182 & ~n2856;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = n3849 & ~n3917;
  assign n3919 = ~n3849 & n3917;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = ~n3784 & ~n3860;
  assign n3922 = n3784 & n3860;
  assign n3923 = ~n3854 & ~n3922;
  assign n3924 = ~n3921 & ~n3923;
  assign n3925 = ~n3920 & n3924;
  assign n3926 = n3849 & n3917;
  assign n3927 = ~n3849 & ~n3917;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = ~n3924 & ~n3928;
  assign n3930 = ~n3925 & ~n3929;
  assign n3931 = n2882 & ~n3930;
  assign n3932 = ~n2870 & ~n3917;
  assign n3933 = ~n3870 & ~n3917;
  assign n3934 = n3870 & n3917;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = n2864 & n3935;
  assign n3937 = ~n3911 & ~n3931;
  assign n3938 = ~n3932 & n3937;
  assign n3939 = ~n3936 & n3938;
  assign n3940 = ~n3861 & ~n3920;
  assign n3941 = ~n3862 & n3877;
  assign n3942 = n3940 & ~n3941;
  assign n3943 = ~n3862 & ~n3919;
  assign n3944 = ~n3918 & n3943;
  assign n3945 = ~n3861 & ~n3877;
  assign n3946 = n3944 & ~n3945;
  assign n3947 = ~n3942 & ~n3946;
  assign n3948 = n2904 & ~n3947;
  assign n3949 = n2952 & ~n3784;
  assign n3950 = n2898 & ~n3930;
  assign n3951 = n2901 & ~n3947;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = n2893 & ~n3930;
  assign n3954 = n2888 & ~n3930;
  assign n3955 = n2890 & ~n3947;
  assign n3956 = n2896 & ~n3947;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3953 & ~n3954;
  assign n3959 = n3957 & n3958;
  assign n3960 = ~n3948 & ~n3949;
  assign n3961 = n3952 & n3960;
  assign n3962 = n3959 & n3961;
  assign n3963 = n3939 & n3962;
  assign n3964 = n2829 & ~n3963;
  assign n3965 = P1_REG0_REG_16_ & ~n2829;
  assign n510 = n3964 | n3965;
  assign n3967 = P1_REG1_REG_18_ & n2845;
  assign n3968 = P1_REG0_REG_18_ & n2843;
  assign n3969 = P1_REG2_REG_18_ & n2847;
  assign n3970 = P1_REG3_REG_17_ & n3903;
  assign n3971 = ~P1_REG3_REG_18_ & n3970;
  assign n3972 = P1_REG3_REG_18_ & ~n3970;
  assign n3973 = ~n3971 & ~n3972;
  assign n3974 = n2841 & ~n3973;
  assign n3975 = ~n3967 & ~n3968;
  assign n3976 = ~n3969 & n3975;
  assign n3977 = ~n3974 & n3976;
  assign n3978 = n2834 & ~n3977;
  assign n3979 = P1_IR_REG_31_ & n2188;
  assign n3980 = P1_IR_REG_17_ & ~P1_IR_REG_31_;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n2856 & ~n3981;
  assign n3983 = ~n2206 & ~n2856;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = ~n3910 & ~n3984;
  assign n3986 = n3910 & n3984;
  assign n3987 = ~n3926 & ~n3986;
  assign n3988 = ~n3985 & n3987;
  assign n3989 = n3924 & ~n3927;
  assign n3990 = n3988 & ~n3989;
  assign n3991 = n3910 & ~n3984;
  assign n3992 = ~n3910 & n3984;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~n3927 & n3993;
  assign n3995 = ~n3924 & ~n3926;
  assign n3996 = n3994 & ~n3995;
  assign n3997 = ~n3990 & ~n3996;
  assign n3998 = n2882 & n3997;
  assign n3999 = ~n2870 & ~n3984;
  assign n4000 = n3934 & n3984;
  assign n4001 = ~n3934 & ~n3984;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = n2864 & n4002;
  assign n4004 = ~n3978 & ~n3998;
  assign n4005 = ~n3999 & n4004;
  assign n4006 = ~n4003 & n4005;
  assign n4007 = n3800 & ~n3861;
  assign n4008 = n3943 & ~n4007;
  assign n4009 = ~n3918 & ~n4008;
  assign n4010 = ~n3799 & ~n3861;
  assign n4011 = ~n3918 & n4010;
  assign n4012 = ~n3816 & n4011;
  assign n4013 = ~n4009 & ~n4012;
  assign n4014 = ~n3993 & ~n4013;
  assign n4015 = n3993 & n4013;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = n2904 & ~n4016;
  assign n4018 = n2952 & ~n3849;
  assign n4019 = n2898 & n3997;
  assign n4020 = n2901 & ~n4016;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = n2893 & n3997;
  assign n4023 = n2888 & n3997;
  assign n4024 = n2890 & ~n4016;
  assign n4025 = n2896 & ~n4016;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = ~n4022 & ~n4023;
  assign n4028 = n4026 & n4027;
  assign n4029 = ~n4017 & ~n4018;
  assign n4030 = n4021 & n4029;
  assign n4031 = n4028 & n4030;
  assign n4032 = n4006 & n4031;
  assign n4033 = n2829 & ~n4032;
  assign n4034 = P1_REG0_REG_17_ & ~n2829;
  assign n515 = n4033 | n4034;
  assign n4036 = P1_REG1_REG_19_ & n2845;
  assign n4037 = P1_REG0_REG_19_ & n2843;
  assign n4038 = P1_REG2_REG_19_ & n2847;
  assign n4039 = P1_REG3_REG_18_ & n3970;
  assign n4040 = ~P1_REG3_REG_19_ & n4039;
  assign n4041 = P1_REG3_REG_19_ & ~n4039;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = n2841 & ~n4042;
  assign n4044 = ~n4036 & ~n4037;
  assign n4045 = ~n4038 & n4044;
  assign n4046 = ~n4043 & n4045;
  assign n4047 = n2834 & ~n4046;
  assign n4048 = n3927 & ~n3984;
  assign n4049 = ~n3927 & n3984;
  assign n4050 = ~n3910 & ~n4049;
  assign n4051 = ~n4048 & ~n4050;
  assign n4052 = ~n3924 & n3987;
  assign n4053 = n4051 & ~n4052;
  assign n4054 = P1_IR_REG_31_ & n2222;
  assign n4055 = P1_IR_REG_18_ & ~P1_IR_REG_31_;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n2856 & ~n4056;
  assign n4058 = ~n2240_1 & ~n2856;
  assign n4059 = ~n4057 & ~n4058;
  assign n4060 = n3977 & ~n4059;
  assign n4061 = ~n3977 & n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n4053 & ~n4062;
  assign n4064 = n3977 & n4059;
  assign n4065 = ~n3977 & ~n4059;
  assign n4066 = ~n4064 & ~n4065;
  assign n4067 = ~n4053 & ~n4066;
  assign n4068 = ~n4063 & ~n4067;
  assign n4069 = n2882 & ~n4068;
  assign n4070 = ~n2870 & ~n4059;
  assign n4071 = ~n4000 & ~n4059;
  assign n4072 = n3984 & n4059;
  assign n4073 = n3934 & n4072;
  assign n4074 = ~n4071 & ~n4073;
  assign n4075 = n2864 & n4074;
  assign n4076 = ~n4047 & ~n4069;
  assign n4077 = ~n4070 & n4076;
  assign n4078 = ~n4075 & n4077;
  assign n4079 = ~n3991 & ~n4013;
  assign n4080 = ~n3992 & ~n4079;
  assign n4081 = ~n4062 & ~n4080;
  assign n4082 = n4062 & n4080;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = n2904 & ~n4083;
  assign n4085 = n2952 & ~n3910;
  assign n4086 = n2898 & ~n4068;
  assign n4087 = n2901 & ~n4083;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = n2893 & ~n4068;
  assign n4090 = n2888 & ~n4068;
  assign n4091 = n2890 & ~n4083;
  assign n4092 = n2896 & ~n4083;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = ~n4089 & ~n4090;
  assign n4095 = n4093 & n4094;
  assign n4096 = ~n4084 & ~n4085;
  assign n4097 = n4088 & n4096;
  assign n4098 = n4095 & n4097;
  assign n4099 = n4078 & n4098;
  assign n4100 = n2829 & ~n4099;
  assign n4101 = P1_REG0_REG_18_ & ~n2829;
  assign n520 = n4100 | n4101;
  assign n4103 = P1_REG1_REG_20_ & n2845;
  assign n4104 = P1_REG0_REG_20_ & n2843;
  assign n4105 = P1_REG2_REG_20_ & n2847;
  assign n4106 = P1_REG3_REG_19_ & n4039;
  assign n4107 = ~P1_REG3_REG_20_ & n4106;
  assign n4108 = P1_REG3_REG_20_ & ~n4106;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = n2841 & ~n4109;
  assign n4111 = ~n4103 & ~n4104;
  assign n4112 = ~n4105 & n4111;
  assign n4113 = ~n4110 & n4112;
  assign n4114 = n2834 & ~n4113;
  assign n4115 = ~n2764 & n2856;
  assign n4116 = ~n2277 & ~n2856;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = n4046 & ~n4117;
  assign n4119 = ~n4046 & n4117;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = ~n4053 & ~n4064;
  assign n4122 = ~n4065 & ~n4121;
  assign n4123 = ~n4120 & n4122;
  assign n4124 = n4046 & n4117;
  assign n4125 = ~n4046 & ~n4117;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~n4122 & ~n4126;
  assign n4128 = ~n4123 & ~n4127;
  assign n4129 = n2882 & ~n4128;
  assign n4130 = ~n2870 & ~n4117;
  assign n4131 = n4073 & n4117;
  assign n4132 = ~n4073 & ~n4117;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = n2864 & n4133;
  assign n4135 = ~n4114 & ~n4129;
  assign n4136 = ~n4130 & n4135;
  assign n4137 = ~n4134 & n4136;
  assign n4138 = ~n3977 & ~n4080;
  assign n4139 = n3977 & n4080;
  assign n4140 = n4059 & ~n4139;
  assign n4141 = ~n4138 & ~n4140;
  assign n4142 = ~n4120 & ~n4141;
  assign n4143 = n4120 & n4141;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = n2904 & ~n4144;
  assign n4146 = n2952 & ~n3977;
  assign n4147 = n2898 & ~n4128;
  assign n4148 = n2901 & ~n4144;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = n2893 & ~n4128;
  assign n4151 = n2888 & ~n4128;
  assign n4152 = n2890 & ~n4144;
  assign n4153 = n2896 & ~n4144;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = ~n4150 & ~n4151;
  assign n4156 = n4154 & n4155;
  assign n4157 = ~n4145 & ~n4146;
  assign n4158 = n4149 & n4157;
  assign n4159 = n4156 & n4158;
  assign n4160 = n4137 & n4159;
  assign n4161 = n2829 & ~n4160;
  assign n4162 = P1_REG0_REG_19_ & ~n2829;
  assign n525 = n4161 | n4162;
  assign n4164 = ~n2314 & ~n2856;
  assign n4165 = ~n2870 & n4164;
  assign n4166 = ~n4131 & n4164;
  assign n4167 = n4131 & ~n4164;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = n2864 & n4168;
  assign n4170 = P1_REG1_REG_21_ & n2845;
  assign n4171 = P1_REG0_REG_21_ & n2843;
  assign n4172 = P1_REG2_REG_21_ & n2847;
  assign n4173 = P1_REG3_REG_20_ & n4106;
  assign n4174 = ~P1_REG3_REG_21_ & n4173;
  assign n4175 = P1_REG3_REG_21_ & ~n4173;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n2841 & ~n4176;
  assign n4178 = ~n4170 & ~n4171;
  assign n4179 = ~n4172 & n4178;
  assign n4180 = ~n4177 & n4179;
  assign n4181 = n2834 & ~n4180;
  assign n4182 = ~n4113 & n4164;
  assign n4183 = n4122 & ~n4125;
  assign n4184 = n4113 & ~n4164;
  assign n4185 = ~n4124 & ~n4184;
  assign n4186 = ~n4182 & ~n4183;
  assign n4187 = n4185 & n4186;
  assign n4188 = n4113 & n4164;
  assign n4189 = ~n4113 & ~n4164;
  assign n4190 = ~n4188 & ~n4189;
  assign n4191 = ~n4125 & n4190;
  assign n4192 = ~n4122 & ~n4124;
  assign n4193 = n4191 & ~n4192;
  assign n4194 = ~n4187 & ~n4193;
  assign n4195 = n2882 & n4194;
  assign n4196 = ~n4165 & ~n4169;
  assign n4197 = ~n4181 & n4196;
  assign n4198 = ~n4195 & n4197;
  assign n4199 = ~n4118 & ~n4141;
  assign n4200 = ~n4119 & ~n4199;
  assign n4201 = ~n4190 & ~n4200;
  assign n4202 = n4190 & n4200;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = n2904 & ~n4203;
  assign n4205 = n2952 & ~n4046;
  assign n4206 = n2898 & n4194;
  assign n4207 = n2901 & ~n4203;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = n2893 & n4194;
  assign n4210 = n2888 & n4194;
  assign n4211 = n2890 & ~n4203;
  assign n4212 = n2896 & ~n4203;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = ~n4209 & ~n4210;
  assign n4215 = n4213 & n4214;
  assign n4216 = ~n4204 & ~n4205;
  assign n4217 = n4208 & n4216;
  assign n4218 = n4215 & n4217;
  assign n4219 = n4198 & n4218;
  assign n4220 = n2829 & ~n4219;
  assign n4221 = P1_REG0_REG_20_ & ~n2829;
  assign n530 = n4220 | n4221;
  assign n4223 = P1_REG1_REG_22_ & n2845;
  assign n4224 = P1_REG0_REG_22_ & n2843;
  assign n4225 = P1_REG2_REG_22_ & n2847;
  assign n4226 = P1_REG3_REG_21_ & n4173;
  assign n4227 = ~P1_REG3_REG_22_ & n4226;
  assign n4228 = P1_REG3_REG_22_ & ~n4226;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = n2841 & ~n4229;
  assign n4231 = ~n4223 & ~n4224;
  assign n4232 = ~n4225 & n4231;
  assign n4233 = ~n4230 & n4232;
  assign n4234 = n2834 & ~n4233;
  assign n4235 = ~n2338 & ~n2856;
  assign n4236 = n4180 & n4235;
  assign n4237 = ~n4180 & ~n4235;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~n4122 & n4185;
  assign n4240 = ~n4125 & ~n4164;
  assign n4241 = n4125 & n4164;
  assign n4242 = n4113 & ~n4241;
  assign n4243 = ~n4240 & ~n4242;
  assign n4244 = ~n4239 & ~n4243;
  assign n4245 = ~n4238 & ~n4244;
  assign n4246 = n4238 & ~n4243;
  assign n4247 = ~n4239 & n4246;
  assign n4248 = ~n4245 & ~n4247;
  assign n4249 = n2882 & n4248;
  assign n4250 = ~n2870 & n4235;
  assign n4251 = n4167 & ~n4235;
  assign n4252 = ~n4167 & n4235;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = n2864 & n4253;
  assign n4255 = ~n4234 & ~n4249;
  assign n4256 = ~n4250 & n4255;
  assign n4257 = ~n4254 & n4256;
  assign n4258 = ~n4188 & ~n4200;
  assign n4259 = ~n4189 & ~n4258;
  assign n4260 = n4238 & n4259;
  assign n4261 = ~n4238 & ~n4259;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = n2904 & ~n4262;
  assign n4264 = n2952 & ~n4113;
  assign n4265 = n2898 & n4248;
  assign n4266 = n2901 & ~n4262;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = n2893 & n4248;
  assign n4269 = n2888 & n4248;
  assign n4270 = n2890 & ~n4262;
  assign n4271 = n2896 & ~n4262;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = ~n4268 & ~n4269;
  assign n4274 = n4272 & n4273;
  assign n4275 = ~n4263 & ~n4264;
  assign n4276 = n4267 & n4275;
  assign n4277 = n4274 & n4276;
  assign n4278 = n4257 & n4277;
  assign n4279 = n2829 & ~n4278;
  assign n4280 = P1_REG0_REG_21_ & ~n2829;
  assign n535 = n4279 | n4280;
  assign n4282 = ~n2375_1 & ~n2856;
  assign n4283 = ~n2870 & n4282;
  assign n4284 = ~n4251 & n4282;
  assign n4285 = n4251 & ~n4282;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = n2864 & n4286;
  assign n4288 = P1_REG1_REG_23_ & n2845;
  assign n4289 = P1_REG0_REG_23_ & n2843;
  assign n4290 = P1_REG2_REG_23_ & n2847;
  assign n4291 = P1_REG3_REG_22_ & n4226;
  assign n4292 = ~P1_REG3_REG_23_ & n4291;
  assign n4293 = P1_REG3_REG_23_ & ~n4291;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = n2841 & ~n4294;
  assign n4296 = ~n4288 & ~n4289;
  assign n4297 = ~n4290 & n4296;
  assign n4298 = ~n4295 & n4297;
  assign n4299 = n2834 & ~n4298;
  assign n4300 = n4180 & ~n4235;
  assign n4301 = n4065 & n4185;
  assign n4302 = ~n4243 & ~n4301;
  assign n4303 = ~n4300 & ~n4302;
  assign n4304 = ~n4180 & n4235;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = ~n4064 & n4185;
  assign n4307 = ~n4053 & ~n4300;
  assign n4308 = n4306 & n4307;
  assign n4309 = n4305 & ~n4308;
  assign n4310 = n4233 & n4282;
  assign n4311 = ~n4233 & ~n4282;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = n4309 & ~n4312;
  assign n4314 = ~n4309 & n4312;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = n2882 & ~n4315;
  assign n4317 = ~n4283 & ~n4287;
  assign n4318 = ~n4299 & n4317;
  assign n4319 = ~n4316 & n4318;
  assign n4320 = ~n4236 & ~n4259;
  assign n4321 = ~n4237 & ~n4320;
  assign n4322 = n4312 & n4321;
  assign n4323 = ~n4312 & ~n4321;
  assign n4324 = ~n4322 & ~n4323;
  assign n4325 = n2904 & ~n4324;
  assign n4326 = n2952 & ~n4180;
  assign n4327 = n2898 & ~n4315;
  assign n4328 = n2901 & ~n4324;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = n2893 & ~n4315;
  assign n4331 = n2888 & ~n4315;
  assign n4332 = n2890 & ~n4324;
  assign n4333 = n2896 & ~n4324;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = ~n4330 & ~n4331;
  assign n4336 = n4334 & n4335;
  assign n4337 = ~n4325 & ~n4326;
  assign n4338 = n4329 & n4337;
  assign n4339 = n4336 & n4338;
  assign n4340 = n4319 & n4339;
  assign n4341 = n2829 & ~n4340;
  assign n4342 = P1_REG0_REG_22_ & ~n2829;
  assign n540 = n4341 | n4342;
  assign n4344 = ~n2417 & ~n2856;
  assign n4345 = ~n2870 & n4344;
  assign n4346 = ~n4233 & n4282;
  assign n4347 = n4233 & ~n4282;
  assign n4348 = ~n4309 & ~n4347;
  assign n4349 = ~n4346 & ~n4348;
  assign n4350 = n4298 & n4344;
  assign n4351 = ~n4298 & ~n4344;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = n4349 & ~n4352;
  assign n4354 = ~n4349 & n4352;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = n2882 & ~n4355;
  assign n4357 = P1_REG1_REG_24_ & n2845;
  assign n4358 = P1_REG0_REG_24_ & n2843;
  assign n4359 = P1_REG2_REG_24_ & n2847;
  assign n4360 = P1_REG3_REG_23_ & n4291;
  assign n4361 = ~P1_REG3_REG_24_ & n4360;
  assign n4362 = P1_REG3_REG_24_ & ~n4360;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = n2841 & ~n4363;
  assign n4365 = ~n4357 & ~n4358;
  assign n4366 = ~n4359 & n4365;
  assign n4367 = ~n4364 & n4366;
  assign n4368 = n2834 & ~n4367;
  assign n4369 = n4285 & ~n4344;
  assign n4370 = ~n4285 & n4344;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = n2864 & n4371;
  assign n4373 = ~n4345 & ~n4356;
  assign n4374 = ~n4368 & n4373;
  assign n4375 = ~n4372 & n4374;
  assign n4376 = ~n4310 & ~n4352;
  assign n4377 = ~n4311 & n4321;
  assign n4378 = n4376 & ~n4377;
  assign n4379 = ~n4310 & ~n4321;
  assign n4380 = ~n4311 & ~n4351;
  assign n4381 = ~n4350 & ~n4379;
  assign n4382 = n4380 & n4381;
  assign n4383 = ~n4378 & ~n4382;
  assign n4384 = n2904 & ~n4383;
  assign n4385 = n2952 & ~n4233;
  assign n4386 = n2898 & ~n4355;
  assign n4387 = n2901 & ~n4383;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = n2893 & ~n4355;
  assign n4390 = n2888 & ~n4355;
  assign n4391 = n2890 & ~n4383;
  assign n4392 = n2896 & ~n4383;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = ~n4389 & ~n4390;
  assign n4395 = n4393 & n4394;
  assign n4396 = ~n4384 & ~n4385;
  assign n4397 = n4388 & n4396;
  assign n4398 = n4395 & n4397;
  assign n4399 = n4375 & n4398;
  assign n4400 = n2829 & ~n4399;
  assign n4401 = P1_REG0_REG_23_ & ~n2829;
  assign n545 = n4400 | n4401;
  assign n4403 = P1_REG1_REG_25_ & n2845;
  assign n4404 = P1_REG0_REG_25_ & n2843;
  assign n4405 = P1_REG2_REG_25_ & n2847;
  assign n4406 = P1_REG3_REG_24_ & n4360;
  assign n4407 = ~P1_REG3_REG_25_ & n4406;
  assign n4408 = P1_REG3_REG_25_ & ~n4406;
  assign n4409 = ~n4407 & ~n4408;
  assign n4410 = n2841 & ~n4409;
  assign n4411 = ~n4403 & ~n4404;
  assign n4412 = ~n4405 & n4411;
  assign n4413 = ~n4410 & n4412;
  assign n4414 = n2834 & ~n4413;
  assign n4415 = ~n2457 & ~n2856;
  assign n4416 = ~n4369 & n4415;
  assign n4417 = n4369 & ~n4415;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = n2864 & n4418;
  assign n4420 = ~n2870 & n4415;
  assign n4421 = ~n4298 & n4344;
  assign n4422 = n4298 & ~n4344;
  assign n4423 = ~n4349 & ~n4422;
  assign n4424 = ~n4421 & ~n4423;
  assign n4425 = n4367 & n4415;
  assign n4426 = ~n4367 & ~n4415;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = n4424 & ~n4427;
  assign n4429 = n4367 & ~n4415;
  assign n4430 = ~n4367 & n4415;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = ~n4424 & ~n4431;
  assign n4433 = ~n4428 & ~n4432;
  assign n4434 = n2882 & ~n4433;
  assign n4435 = ~n4414 & ~n4419;
  assign n4436 = ~n4420 & n4435;
  assign n4437 = ~n4434 & n4436;
  assign n4438 = n4237 & ~n4310;
  assign n4439 = n4380 & ~n4438;
  assign n4440 = ~n4350 & ~n4439;
  assign n4441 = ~n4236 & ~n4310;
  assign n4442 = ~n4259 & n4441;
  assign n4443 = ~n4350 & n4442;
  assign n4444 = ~n4440 & ~n4443;
  assign n4445 = ~n4427 & ~n4444;
  assign n4446 = n4427 & n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n2904 & ~n4447;
  assign n4449 = n2952 & ~n4298;
  assign n4450 = n2898 & ~n4433;
  assign n4451 = n2901 & ~n4447;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = n2893 & ~n4433;
  assign n4454 = n2888 & ~n4433;
  assign n4455 = n2890 & ~n4447;
  assign n4456 = n2896 & ~n4447;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n4453 & ~n4454;
  assign n4459 = n4457 & n4458;
  assign n4460 = ~n4448 & ~n4449;
  assign n4461 = n4452 & n4460;
  assign n4462 = n4459 & n4461;
  assign n4463 = n4437 & n4462;
  assign n4464 = n2829 & ~n4463;
  assign n4465 = P1_REG0_REG_24_ & ~n2829;
  assign n550 = n4464 | n4465;
  assign n4467 = P1_REG1_REG_26_ & n2845;
  assign n4468 = P1_REG0_REG_26_ & n2843;
  assign n4469 = P1_REG2_REG_26_ & n2847;
  assign n4470 = P1_REG3_REG_25_ & n4406;
  assign n4471 = ~P1_REG3_REG_26_ & n4470;
  assign n4472 = P1_REG3_REG_26_ & ~n4470;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = n2841 & ~n4473;
  assign n4475 = ~n4467 & ~n4468;
  assign n4476 = ~n4469 & n4475;
  assign n4477 = ~n4474 & n4476;
  assign n4478 = n2834 & ~n4477;
  assign n4479 = ~n2481 & ~n2856;
  assign n4480 = n4417 & ~n4479;
  assign n4481 = ~n4417 & n4479;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n2864 & n4482;
  assign n4484 = ~n2870 & n4479;
  assign n4485 = n4413 & n4479;
  assign n4486 = ~n4413 & ~n4479;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~n4424 & ~n4429;
  assign n4489 = ~n4430 & ~n4488;
  assign n4490 = ~n4487 & n4489;
  assign n4491 = n4413 & ~n4479;
  assign n4492 = ~n4413 & n4479;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~n4489 & ~n4493;
  assign n4495 = ~n4490 & ~n4494;
  assign n4496 = n2882 & ~n4495;
  assign n4497 = ~n4478 & ~n4483;
  assign n4498 = ~n4484 & n4497;
  assign n4499 = ~n4496 & n4498;
  assign n4500 = ~n4425 & ~n4444;
  assign n4501 = ~n4426 & ~n4500;
  assign n4502 = ~n4487 & ~n4501;
  assign n4503 = n4487 & n4501;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = n2904 & ~n4504;
  assign n4506 = n2952 & ~n4367;
  assign n4507 = n2898 & ~n4495;
  assign n4508 = n2901 & ~n4504;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = n2893 & ~n4495;
  assign n4511 = n2888 & ~n4495;
  assign n4512 = n2890 & ~n4504;
  assign n4513 = n2896 & ~n4504;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4510 & ~n4511;
  assign n4516 = n4514 & n4515;
  assign n4517 = ~n4505 & ~n4506;
  assign n4518 = n4509 & n4517;
  assign n4519 = n4516 & n4518;
  assign n4520 = n4499 & n4519;
  assign n4521 = n2829 & ~n4520;
  assign n4522 = P1_REG0_REG_25_ & ~n2829;
  assign n555 = n4521 | n4522;
  assign n4524 = P1_REG1_REG_27_ & n2845;
  assign n4525 = P1_REG0_REG_27_ & n2843;
  assign n4526 = P1_REG2_REG_27_ & n2847;
  assign n4527 = P1_REG3_REG_26_ & n4470;
  assign n4528 = ~P1_REG3_REG_27_ & n4527;
  assign n4529 = P1_REG3_REG_27_ & ~n4527;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = n2841 & ~n4530;
  assign n4532 = ~n4524 & ~n4525;
  assign n4533 = ~n4526 & n4532;
  assign n4534 = ~n4531 & n4533;
  assign n4535 = n2834 & ~n4534;
  assign n4536 = ~n2524 & ~n2856;
  assign n4537 = ~n4480 & n4536;
  assign n4538 = n4480 & ~n4536;
  assign n4539 = ~n4537 & ~n4538;
  assign n4540 = n2864 & n4539;
  assign n4541 = ~n2870 & n4536;
  assign n4542 = n4489 & ~n4492;
  assign n4543 = ~n4477 & n4536;
  assign n4544 = ~n4491 & n4536;
  assign n4545 = ~n4477 & ~n4491;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~n4542 & ~n4543;
  assign n4548 = ~n4546 & n4547;
  assign n4549 = ~n4489 & ~n4491;
  assign n4550 = n4477 & n4536;
  assign n4551 = ~n4477 & ~n4536;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4492 & ~n4549;
  assign n4554 = n4552 & n4553;
  assign n4555 = ~n4548 & ~n4554;
  assign n4556 = n2882 & n4555;
  assign n4557 = ~n4535 & ~n4540;
  assign n4558 = ~n4541 & n4557;
  assign n4559 = ~n4556 & n4558;
  assign n4560 = ~n4485 & ~n4501;
  assign n4561 = ~n4486 & ~n4560;
  assign n4562 = n4552 & n4561;
  assign n4563 = ~n4552 & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = n2904 & ~n4564;
  assign n4566 = n2952 & ~n4413;
  assign n4567 = n2898 & n4555;
  assign n4568 = n2901 & ~n4564;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = n2893 & n4555;
  assign n4571 = n2888 & n4555;
  assign n4572 = n2890 & ~n4564;
  assign n4573 = n2896 & ~n4564;
  assign n4574 = ~n4572 & ~n4573;
  assign n4575 = ~n4570 & ~n4571;
  assign n4576 = n4574 & n4575;
  assign n4577 = ~n4565 & ~n4566;
  assign n4578 = n4569 & n4577;
  assign n4579 = n4576 & n4578;
  assign n4580 = n4559 & n4579;
  assign n4581 = n2829 & ~n4580;
  assign n4582 = P1_REG0_REG_26_ & ~n2829;
  assign n560 = n4581 | n4582;
  assign n4584 = P1_REG1_REG_28_ & n2845;
  assign n4585 = P1_REG0_REG_28_ & n2843;
  assign n4586 = P1_REG2_REG_28_ & n2847;
  assign n4587 = P1_REG3_REG_27_ & n4527;
  assign n4588 = ~P1_REG3_REG_28_ & n4587;
  assign n4589 = P1_REG3_REG_28_ & ~n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n2841 & ~n4590;
  assign n4592 = ~n4584 & ~n4585;
  assign n4593 = ~n4586 & n4592;
  assign n4594 = ~n4591 & n4593;
  assign n4595 = n2834 & ~n4594;
  assign n4596 = ~n2548 & ~n2856;
  assign n4597 = n4538 & ~n4596;
  assign n4598 = ~n4538 & n4596;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = n2864 & n4599;
  assign n4601 = ~n2870 & n4596;
  assign n4602 = ~n4430 & ~n4492;
  assign n4603 = ~n4546 & ~n4602;
  assign n4604 = n4488 & ~n4546;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = ~n4543 & n4605;
  assign n4607 = n4534 & n4596;
  assign n4608 = ~n4534 & ~n4596;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = n4606 & ~n4609;
  assign n4611 = ~n4606 & n4609;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = n2882 & ~n4612;
  assign n4614 = ~n4595 & ~n4600;
  assign n4615 = ~n4601 & n4614;
  assign n4616 = ~n4613 & n4615;
  assign n4617 = ~n4550 & ~n4609;
  assign n4618 = ~n4551 & n4561;
  assign n4619 = n4617 & ~n4618;
  assign n4620 = ~n4551 & n4609;
  assign n4621 = ~n4550 & ~n4561;
  assign n4622 = n4620 & ~n4621;
  assign n4623 = ~n4619 & ~n4622;
  assign n4624 = n2904 & ~n4623;
  assign n4625 = n2952 & ~n4477;
  assign n4626 = n2898 & ~n4612;
  assign n4627 = n2901 & ~n4623;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = n2893 & ~n4612;
  assign n4630 = n2888 & ~n4612;
  assign n4631 = n2890 & ~n4623;
  assign n4632 = n2896 & ~n4623;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n4629 & ~n4630;
  assign n4635 = n4633 & n4634;
  assign n4636 = ~n4624 & ~n4625;
  assign n4637 = n4628 & n4636;
  assign n4638 = n4635 & n4637;
  assign n4639 = n4616 & n4638;
  assign n4640 = n2829 & ~n4639;
  assign n4641 = P1_REG0_REG_27_ & ~n2829;
  assign n565 = n4640 | n4641;
  assign n4643 = P1_REG0_REG_29_ & n2843;
  assign n4644 = P1_REG1_REG_29_ & n2845;
  assign n4645 = P1_REG2_REG_29_ & n2847;
  assign n4646 = P1_REG3_REG_28_ & P1_REG3_REG_27_;
  assign n4647 = n4527 & n4646;
  assign n4648 = n2841 & n4647;
  assign n4649 = ~n4643 & ~n4644;
  assign n4650 = ~n4645 & n4649;
  assign n4651 = ~n4648 & n4650;
  assign n4652 = n2834 & ~n4651;
  assign n4653 = ~n2593 & ~n2856;
  assign n4654 = ~n4597 & n4653;
  assign n4655 = n4597 & ~n4653;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = n2864 & n4656;
  assign n4658 = ~n2870 & n4653;
  assign n4659 = n4534 & ~n4596;
  assign n4660 = n4543 & ~n4659;
  assign n4661 = ~n4429 & ~n4659;
  assign n4662 = ~n4424 & ~n4546;
  assign n4663 = n4661 & n4662;
  assign n4664 = n4603 & ~n4659;
  assign n4665 = ~n4534 & n4596;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = ~n4660 & ~n4663;
  assign n4668 = n4666 & n4667;
  assign n4669 = n4594 & n4653;
  assign n4670 = ~n4594 & ~n4653;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = n4668 & ~n4671;
  assign n4673 = ~n4668 & n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = n2882 & ~n4674;
  assign n4676 = ~n4652 & ~n4657;
  assign n4677 = ~n4658 & n4676;
  assign n4678 = ~n4675 & n4677;
  assign n4679 = n4534 & ~n4551;
  assign n4680 = ~n4596 & ~n4679;
  assign n4681 = ~n4534 & n4551;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = ~n4607 & n4621;
  assign n4684 = n4682 & ~n4683;
  assign n4685 = ~n4671 & ~n4684;
  assign n4686 = n4671 & n4684;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = n2904 & ~n4687;
  assign n4689 = n2952 & ~n4534;
  assign n4690 = n2898 & ~n4674;
  assign n4691 = n2901 & ~n4687;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = n2893 & ~n4674;
  assign n4694 = n2888 & ~n4674;
  assign n4695 = n2890 & ~n4687;
  assign n4696 = n2896 & ~n4687;
  assign n4697 = ~n4695 & ~n4696;
  assign n4698 = ~n4693 & ~n4694;
  assign n4699 = n4697 & n4698;
  assign n4700 = ~n4688 & ~n4689;
  assign n4701 = n4692 & n4700;
  assign n4702 = n4699 & n4701;
  assign n4703 = n4678 & n4702;
  assign n4704 = n2829 & ~n4703;
  assign n4705 = P1_REG0_REG_28_ & ~n2829;
  assign n570 = n4704 | n4705;
  assign n4707 = ~n2622 & ~n2856;
  assign n4708 = n4655 & ~n4707;
  assign n4709 = ~n4655 & n4707;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = n2864 & n4710;
  assign n4712 = ~n2870 & n4707;
  assign n4713 = n4653 & ~n4668;
  assign n4714 = ~n4594 & ~n4668;
  assign n4715 = ~n4594 & n4653;
  assign n4716 = ~n4713 & ~n4714;
  assign n4717 = ~n4715 & n4716;
  assign n4718 = n4651 & n4707;
  assign n4719 = ~n4651 & ~n4707;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = n4717 & ~n4720;
  assign n4722 = ~n4717 & n4720;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = n2882 & ~n4723;
  assign n4725 = ~n4711 & ~n4712;
  assign n4726 = ~n4724 & n4725;
  assign n4727 = n2888 & ~n4723;
  assign n4728 = n2898 & ~n4723;
  assign n4729 = n2952 & ~n4594;
  assign n4730 = ~P1_B_REG & n2833;
  assign n4731 = ~n2856 & ~n4730;
  assign n4732 = n2830 & ~n4731;
  assign n4733 = P1_REG1_REG_30_ & n2845;
  assign n4734 = P1_REG0_REG_30_ & n2843;
  assign n4735 = P1_REG2_REG_30_ & n2847;
  assign n4736 = ~n4733 & ~n4734;
  assign n4737 = ~n4735 & n4736;
  assign n4738 = n4732 & ~n4737;
  assign n4739 = ~n4727 & ~n4728;
  assign n4740 = ~n4729 & n4739;
  assign n4741 = ~n4738 & n4740;
  assign n4742 = n2893 & ~n4723;
  assign n4743 = ~n4670 & n4684;
  assign n4744 = ~n4669 & ~n4743;
  assign n4745 = ~n4720 & n4744;
  assign n4746 = ~n4669 & ~n4684;
  assign n4747 = ~n4670 & ~n4746;
  assign n4748 = n4720 & n4747;
  assign n4749 = ~n4745 & ~n4748;
  assign n4750 = n2890 & ~n4749;
  assign n4751 = ~n4742 & ~n4750;
  assign n4752 = n2901 & ~n4749;
  assign n4753 = n2904 & ~n4749;
  assign n4754 = n2896 & ~n4749;
  assign n4755 = ~n4752 & ~n4753;
  assign n4756 = ~n4754 & n4755;
  assign n4757 = n4726 & n4741;
  assign n4758 = n4751 & n4757;
  assign n4759 = n4756 & n4758;
  assign n4760 = n2829 & ~n4759;
  assign n4761 = P1_REG0_REG_29_ & ~n2829;
  assign n575 = n4760 | n4761;
  assign n4763 = ~n2646 & ~n2856;
  assign n4764 = ~n2870 & n4763;
  assign n4765 = P1_REG1_REG_31_ & n2845;
  assign n4766 = P1_REG0_REG_31_ & n2843;
  assign n4767 = P1_REG2_REG_31_ & n2847;
  assign n4768 = ~n4765 & ~n4766;
  assign n4769 = ~n4767 & n4768;
  assign n4770 = n4732 & ~n4769;
  assign n4771 = ~n4708 & n4763;
  assign n4772 = n4708 & ~n4763;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = n2864 & n4773;
  assign n4775 = ~n4764 & ~n4770;
  assign n4776 = ~n4774 & n4775;
  assign n4777 = n2829 & ~n4776;
  assign n4778 = P1_REG0_REG_30_ & ~n2829;
  assign n580 = n4777 | n4778;
  assign n4780 = ~n2677 & ~n2856;
  assign n4781 = ~n2870 & n4780;
  assign n4782 = n4772 & ~n4780;
  assign n4783 = ~n4772 & n4780;
  assign n4784 = ~n4782 & ~n4783;
  assign n4785 = n2864 & n4784;
  assign n4786 = ~n4770 & ~n4781;
  assign n4787 = ~n4785 & n4786;
  assign n4788 = n2829 & ~n4787;
  assign n4789 = P1_REG0_REG_31_ & ~n2829;
  assign n585 = n4788 | n4789;
  assign n4791 = n2696 & ~n2745;
  assign n4792 = n2828 & n4791;
  assign n4793 = ~n2911 & n4792;
  assign n4794 = P1_REG1_REG_0_ & ~n4792;
  assign n590 = n4793 | n4794;
  assign n4796 = ~n2967 & n4792;
  assign n4797 = P1_REG1_REG_1_ & ~n4792;
  assign n595 = n4796 | n4797;
  assign n4799 = ~n3028 & n4792;
  assign n4800 = P1_REG1_REG_2_ & ~n4792;
  assign n600 = n4799 | n4800;
  assign n4802 = ~n3093 & n4792;
  assign n4803 = P1_REG1_REG_3_ & ~n4792;
  assign n605 = n4802 | n4803;
  assign n4805 = ~n3162 & n4792;
  assign n4806 = P1_REG1_REG_4_ & ~n4792;
  assign n610 = n4805 | n4806;
  assign n4808 = ~n3226 & n4792;
  assign n4809 = P1_REG1_REG_5_ & ~n4792;
  assign n615 = n4808 | n4809;
  assign n4811 = ~n3300 & n4792;
  assign n4812 = P1_REG1_REG_6_ & ~n4792;
  assign n620 = n4811 | n4812;
  assign n4814 = ~n3369 & n4792;
  assign n4815 = P1_REG1_REG_7_ & ~n4792;
  assign n625 = n4814 | n4815;
  assign n4817 = ~n3437 & n4792;
  assign n4818 = P1_REG1_REG_8_ & ~n4792;
  assign n630 = n4817 | n4818;
  assign n4820 = ~n3504 & n4792;
  assign n4821 = P1_REG1_REG_9_ & ~n4792;
  assign n635 = n4820 | n4821;
  assign n4823 = ~n3569 & n4792;
  assign n4824 = P1_REG1_REG_10_ & ~n4792;
  assign n640 = n4823 | n4824;
  assign n4826 = ~n3639 & n4792;
  assign n4827 = P1_REG1_REG_11_ & ~n4792;
  assign n645 = n4826 | n4827;
  assign n4829 = ~n3706 & n4792;
  assign n4830 = P1_REG1_REG_12_ & ~n4792;
  assign n650 = n4829 | n4830;
  assign n4832 = ~n3770 & n4792;
  assign n4833 = P1_REG1_REG_13_ & ~n4792;
  assign n655 = n4832 | n4833;
  assign n4835 = ~n3835 & n4792;
  assign n4836 = P1_REG1_REG_14_ & ~n4792;
  assign n660 = n4835 | n4836;
  assign n4838 = ~n3896 & n4792;
  assign n4839 = P1_REG1_REG_15_ & ~n4792;
  assign n665 = n4838 | n4839;
  assign n4841 = ~n3963 & n4792;
  assign n4842 = P1_REG1_REG_16_ & ~n4792;
  assign n670 = n4841 | n4842;
  assign n4844 = ~n4032 & n4792;
  assign n4845 = P1_REG1_REG_17_ & ~n4792;
  assign n675 = n4844 | n4845;
  assign n4847 = ~n4099 & n4792;
  assign n4848 = P1_REG1_REG_18_ & ~n4792;
  assign n680 = n4847 | n4848;
  assign n4850 = ~n4160 & n4792;
  assign n4851 = P1_REG1_REG_19_ & ~n4792;
  assign n685 = n4850 | n4851;
  assign n4853 = ~n4219 & n4792;
  assign n4854 = P1_REG1_REG_20_ & ~n4792;
  assign n690 = n4853 | n4854;
  assign n4856 = ~n4278 & n4792;
  assign n4857 = P1_REG1_REG_21_ & ~n4792;
  assign n695 = n4856 | n4857;
  assign n4859 = ~n4340 & n4792;
  assign n4860 = P1_REG1_REG_22_ & ~n4792;
  assign n700 = n4859 | n4860;
  assign n4862 = ~n4399 & n4792;
  assign n4863 = P1_REG1_REG_23_ & ~n4792;
  assign n705 = n4862 | n4863;
  assign n4865 = ~n4463 & n4792;
  assign n4866 = P1_REG1_REG_24_ & ~n4792;
  assign n710 = n4865 | n4866;
  assign n4868 = ~n4520 & n4792;
  assign n4869 = P1_REG1_REG_25_ & ~n4792;
  assign n715 = n4868 | n4869;
  assign n4871 = ~n4580 & n4792;
  assign n4872 = P1_REG1_REG_26_ & ~n4792;
  assign n720 = n4871 | n4872;
  assign n4874 = ~n4639 & n4792;
  assign n4875 = P1_REG1_REG_27_ & ~n4792;
  assign n725 = n4874 | n4875;
  assign n4877 = ~n4703 & n4792;
  assign n4878 = P1_REG1_REG_28_ & ~n4792;
  assign n730 = n4877 | n4878;
  assign n4880 = ~n4759 & n4792;
  assign n4881 = P1_REG1_REG_29_ & ~n4792;
  assign n735 = n4880 | n4881;
  assign n4883 = ~n4776 & n4792;
  assign n4884 = P1_REG1_REG_30_ & ~n4792;
  assign n740 = n4883 | n4884;
  assign n4886 = ~n4787 & n4792;
  assign n4887 = P1_REG1_REG_31_ & ~n4792;
  assign n745 = n4886 | n4887;
  assign n4889 = n2764 & n2864;
  assign n4890 = n2755 & n2869;
  assign n4891 = ~n2765 & n2830;
  assign n4892 = n2745 & ~n4891;
  assign n4893 = ~n2749 & n4892;
  assign n4894 = n2827 & n4893;
  assign n4895 = ~n4890 & ~n4894;
  assign n4896 = n2696 & ~n4895;
  assign n4897 = n4889 & n4896;
  assign n4898 = ~n2862 & n4897;
  assign n4899 = ~n2755 & n2869;
  assign n4900 = ~n2867 & ~n4899;
  assign n4901 = n4896 & ~n4900;
  assign n4902 = ~n2862 & n4901;
  assign n4903 = ~n2910 & n4896;
  assign n4904 = P1_REG2_REG_0_ & ~n4896;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = ~n4898 & ~n4902;
  assign n4907 = n4905 & n4906;
  assign n4908 = n4890 & n4896;
  assign n4909 = P1_REG3_REG_0_ & n4908;
  assign n4910 = n2834 & n4896;
  assign n4911 = ~n2851 & n4910;
  assign n4912 = ~n2758 & n2903;
  assign n4913 = n4896 & n4912;
  assign n4914 = ~n2881 & n4913;
  assign n4915 = ~n4909 & ~n4911;
  assign n4916 = ~n4914 & n4915;
  assign n750 = ~n4907 | ~n4916;
  assign n4918 = ~n2931 & n4897;
  assign n4919 = ~n2928 & n4901;
  assign n4920 = ~n2966 & n4896;
  assign n4921 = P1_REG2_REG_1_ & ~n4896;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = ~n4918 & ~n4919;
  assign n4924 = n4922 & n4923;
  assign n4925 = P1_REG3_REG_1_ & n4908;
  assign n4926 = ~n2921 & n4910;
  assign n4927 = ~n2940 & n4913;
  assign n4928 = ~n4925 & ~n4926;
  assign n4929 = ~n4927 & n4928;
  assign n755 = ~n4924 | ~n4929;
  assign n4931 = n2989 & n4897;
  assign n4932 = ~n2984 & n4901;
  assign n4933 = ~n3027 & n4896;
  assign n4934 = P1_REG2_REG_2_ & ~n4896;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = ~n4931 & ~n4932;
  assign n4937 = n4935 & n4936;
  assign n4938 = P1_REG3_REG_2_ & n4908;
  assign n4939 = ~n2977 & n4910;
  assign n4940 = n3003 & n4913;
  assign n4941 = ~n4938 & ~n4939;
  assign n4942 = ~n4940 & n4941;
  assign n760 = ~n4937 | ~n4942;
  assign n4944 = n3051 & n4897;
  assign n4945 = ~n3048 & n4901;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = ~P1_REG3_REG_3_ & n4908;
  assign n4948 = ~n3041 & n4910;
  assign n4949 = ~n3066 & n4913;
  assign n4950 = ~n4947 & ~n4948;
  assign n4951 = ~n4949 & n4950;
  assign n4952 = ~n3092 & n4896;
  assign n4953 = P1_REG2_REG_3_ & ~n4896;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = n4946 & n4951;
  assign n765 = ~n4954 | ~n4955;
  assign n4957 = ~n3034 & n4908;
  assign n4958 = ~n3107 & n4910;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = n3117 & n4897;
  assign n4961 = ~n3114 & n4901;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~n3133 & n4913;
  assign n4964 = ~n3161 & n4896;
  assign n4965 = P1_REG2_REG_4_ & ~n4896;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = n4959 & n4962;
  assign n4968 = ~n4963 & n4967;
  assign n770 = ~n4966 | ~n4968;
  assign n4970 = ~n3100 & n4908;
  assign n4971 = ~n3176 & n4910;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = n3186 & n4897;
  assign n4974 = ~n3183 & n4901;
  assign n4975 = ~n4973 & ~n4974;
  assign n4976 = n3201 & n4913;
  assign n4977 = ~n3225 & n4896;
  assign n4978 = P1_REG2_REG_5_ & ~n4896;
  assign n4979 = ~n4977 & ~n4978;
  assign n4980 = n4972 & n4975;
  assign n4981 = ~n4976 & n4980;
  assign n775 = ~n4979 | ~n4981;
  assign n4983 = ~n3169 & n4908;
  assign n4984 = ~n3240 & n4910;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = n3251 & n4897;
  assign n4987 = ~n3247 & n4901;
  assign n4988 = ~n4986 & ~n4987;
  assign n4989 = ~n3272 & n4913;
  assign n4990 = ~n3299 & n4896;
  assign n4991 = P1_REG2_REG_6_ & ~n4896;
  assign n4992 = ~n4990 & ~n4991;
  assign n4993 = n4985 & n4988;
  assign n4994 = ~n4989 & n4993;
  assign n780 = ~n4992 | ~n4994;
  assign n4996 = ~n3233 & n4908;
  assign n4997 = ~n3314 & n4910;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n3324 & n4897;
  assign n5000 = ~n3321 & n4901;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = n3339 & n4913;
  assign n5003 = ~n3368 & n4896;
  assign n5004 = P1_REG2_REG_7_ & ~n4896;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = n4998 & n5001;
  assign n5007 = ~n5002 & n5006;
  assign n785 = ~n5005 | ~n5007;
  assign n5009 = ~n3307 & n4908;
  assign n5010 = ~n3383 & n4910;
  assign n5011 = ~n5009 & ~n5010;
  assign n5012 = n3393 & n4897;
  assign n5013 = ~n3390 & n4901;
  assign n5014 = ~n5012 & ~n5013;
  assign n5015 = ~n3410 & n4913;
  assign n5016 = ~n3436 & n4896;
  assign n5017 = P1_REG2_REG_8_ & ~n4896;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = n5011 & n5014;
  assign n5020 = ~n5015 & n5019;
  assign n790 = ~n5018 | ~n5020;
  assign n5022 = ~n3379 & n4908;
  assign n5023 = ~n3451 & n4910;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = n3461 & n4897;
  assign n5026 = ~n3458 & n4901;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~n3474 & n4913;
  assign n5029 = ~n3503 & n4896;
  assign n5030 = P1_REG2_REG_9_ & ~n4896;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = n5024 & n5027;
  assign n5033 = ~n5028 & n5032;
  assign n795 = ~n5031 | ~n5033;
  assign n5035 = ~n3447 & n4908;
  assign n5036 = ~n3518 & n4910;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = n3529 & n4897;
  assign n5039 = ~n3525 & n4901;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = n3544 & n4913;
  assign n5042 = ~n3568 & n4896;
  assign n5043 = P1_REG2_REG_10_ & ~n4896;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = n5037 & n5040;
  assign n5046 = ~n5041 & n5045;
  assign n800 = ~n5044 | ~n5046;
  assign n5048 = n3611 & n4897;
  assign n5049 = ~n3578 & n4901;
  assign n5050 = ~n5048 & ~n5049;
  assign n5051 = ~n3514 & n4908;
  assign n5052 = ~n3607 & n4910;
  assign n5053 = ~n3595 & n4913;
  assign n5054 = ~n5051 & ~n5052;
  assign n5055 = ~n5053 & n5054;
  assign n5056 = ~n3638 & n4896;
  assign n5057 = P1_REG2_REG_11_ & ~n4896;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = n5050 & n5055;
  assign n805 = ~n5058 | ~n5059;
  assign n5061 = n3676 & n4897;
  assign n5062 = ~n3648 & n4901;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = ~n3603 & n4908;
  assign n5065 = ~n3672 & n4910;
  assign n5066 = ~n3660 & n4913;
  assign n5067 = ~n5064 & ~n5065;
  assign n5068 = ~n5066 & n5067;
  assign n5069 = ~n3705 & n4896;
  assign n5070 = P1_REG2_REG_12_ & ~n4896;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = n5063 & n5068;
  assign n810 = ~n5071 | ~n5072;
  assign n5074 = n3719 & n4897;
  assign n5075 = ~n3715 & n4901;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~n3668 & n4908;
  assign n5078 = ~n3731 & n4910;
  assign n5079 = n3745 & n4913;
  assign n5080 = ~n5077 & ~n5078;
  assign n5081 = ~n5079 & n5080;
  assign n5082 = ~n3769 & n4896;
  assign n5083 = P1_REG2_REG_13_ & ~n4896;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = n5076 & n5081;
  assign n815 = ~n5084 | ~n5085;
  assign n5087 = ~n3727 & n4908;
  assign n5088 = ~n3784 & n4910;
  assign n5089 = ~n3804 & n4913;
  assign n5090 = ~n3798 & n4901;
  assign n5091 = n3810 & n4897;
  assign n5092 = ~n5087 & ~n5088;
  assign n5093 = ~n5089 & n5092;
  assign n5094 = ~n5090 & n5093;
  assign n5095 = ~n5091 & n5094;
  assign n5096 = ~n3834 & n4896;
  assign n5097 = P1_REG2_REG_14_ & ~n4896;
  assign n5098 = ~n5096 & ~n5097;
  assign n820 = ~n5095 | ~n5098;
  assign n5100 = ~n3780 & n4908;
  assign n5101 = ~n3849 & n4910;
  assign n5102 = ~n3866 & n4913;
  assign n5103 = ~n3860 & n4901;
  assign n5104 = n3871 & n4897;
  assign n5105 = ~n5100 & ~n5101;
  assign n5106 = ~n5102 & n5105;
  assign n5107 = ~n5103 & n5106;
  assign n5108 = ~n5104 & n5107;
  assign n5109 = ~n3895 & n4896;
  assign n5110 = P1_REG2_REG_15_ & ~n4896;
  assign n5111 = ~n5109 & ~n5110;
  assign n825 = ~n5108 | ~n5111;
  assign n5113 = ~n3845 & n4908;
  assign n5114 = ~n3910 & n4910;
  assign n5115 = ~n3930 & n4913;
  assign n5116 = ~n3917 & n4901;
  assign n5117 = n3935 & n4897;
  assign n5118 = ~n5113 & ~n5114;
  assign n5119 = ~n5115 & n5118;
  assign n5120 = ~n5116 & n5119;
  assign n5121 = ~n5117 & n5120;
  assign n5122 = ~n3962 & n4896;
  assign n5123 = P1_REG2_REG_16_ & ~n4896;
  assign n5124 = ~n5122 & ~n5123;
  assign n830 = ~n5121 | ~n5124;
  assign n5126 = ~n3906 & n4908;
  assign n5127 = ~n3977 & n4910;
  assign n5128 = n3997 & n4913;
  assign n5129 = ~n3984 & n4901;
  assign n5130 = n4002 & n4897;
  assign n5131 = ~n5126 & ~n5127;
  assign n5132 = ~n5128 & n5131;
  assign n5133 = ~n5129 & n5132;
  assign n5134 = ~n5130 & n5133;
  assign n5135 = ~n4031 & n4896;
  assign n5136 = P1_REG2_REG_17_ & ~n4896;
  assign n5137 = ~n5135 & ~n5136;
  assign n835 = ~n5134 | ~n5137;
  assign n5139 = ~n3973 & n4908;
  assign n5140 = ~n4046 & n4910;
  assign n5141 = ~n4068 & n4913;
  assign n5142 = ~n4059 & n4901;
  assign n5143 = n4074 & n4897;
  assign n5144 = ~n5139 & ~n5140;
  assign n5145 = ~n5141 & n5144;
  assign n5146 = ~n5142 & n5145;
  assign n5147 = ~n5143 & n5146;
  assign n5148 = ~n4098 & n4896;
  assign n5149 = P1_REG2_REG_18_ & ~n4896;
  assign n5150 = ~n5148 & ~n5149;
  assign n840 = ~n5147 | ~n5150;
  assign n5152 = ~n4042 & n4908;
  assign n5153 = ~n4113 & n4910;
  assign n5154 = ~n4128 & n4913;
  assign n5155 = ~n4117 & n4901;
  assign n5156 = n4133 & n4897;
  assign n5157 = ~n5152 & ~n5153;
  assign n5158 = ~n5154 & n5157;
  assign n5159 = ~n5155 & n5158;
  assign n5160 = ~n5156 & n5159;
  assign n5161 = ~n4159 & n4896;
  assign n5162 = P1_REG2_REG_19_ & ~n4896;
  assign n5163 = ~n5161 & ~n5162;
  assign n845 = ~n5160 | ~n5163;
  assign n5165 = n4168 & n4897;
  assign n5166 = n4164 & n4901;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n4109 & n4908;
  assign n5169 = ~n4180 & n4910;
  assign n5170 = n4194 & n4913;
  assign n5171 = ~n5168 & ~n5169;
  assign n5172 = ~n5170 & n5171;
  assign n5173 = ~n4218 & n4896;
  assign n5174 = P1_REG2_REG_20_ & ~n4896;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = n5167 & n5172;
  assign n850 = ~n5175 | ~n5176;
  assign n5178 = ~n4176 & n4908;
  assign n5179 = ~n4233 & n4910;
  assign n5180 = n4248 & n4913;
  assign n5181 = n4235 & n4901;
  assign n5182 = n4253 & n4897;
  assign n5183 = ~n5178 & ~n5179;
  assign n5184 = ~n5180 & n5183;
  assign n5185 = ~n5181 & n5184;
  assign n5186 = ~n5182 & n5185;
  assign n5187 = ~n4277 & n4896;
  assign n5188 = P1_REG2_REG_21_ & ~n4896;
  assign n5189 = ~n5187 & ~n5188;
  assign n855 = ~n5186 | ~n5189;
  assign n5191 = n4286 & n4897;
  assign n5192 = n4282 & n4901;
  assign n5193 = ~n5191 & ~n5192;
  assign n5194 = ~n4229 & n4908;
  assign n5195 = ~n4298 & n4910;
  assign n5196 = ~n4315 & n4913;
  assign n5197 = ~n5194 & ~n5195;
  assign n5198 = ~n5196 & n5197;
  assign n5199 = ~n4339 & n4896;
  assign n5200 = P1_REG2_REG_22_ & ~n4896;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = n5193 & n5198;
  assign n860 = ~n5201 | ~n5202;
  assign n5204 = n4371 & n4897;
  assign n5205 = n4344 & n4901;
  assign n5206 = ~n5204 & ~n5205;
  assign n5207 = ~n4294 & n4908;
  assign n5208 = ~n4367 & n4910;
  assign n5209 = ~n4355 & n4913;
  assign n5210 = ~n5207 & ~n5208;
  assign n5211 = ~n5209 & n5210;
  assign n5212 = ~n4398 & n4896;
  assign n5213 = P1_REG2_REG_23_ & ~n4896;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = n5206 & n5211;
  assign n865 = ~n5214 | ~n5215;
  assign n5217 = ~n4363 & n4908;
  assign n5218 = ~n4413 & n4910;
  assign n5219 = ~n5217 & ~n5218;
  assign n5220 = n4418 & n4897;
  assign n5221 = n4415 & n4901;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = ~n4433 & n4913;
  assign n5224 = ~n4462 & n4896;
  assign n5225 = P1_REG2_REG_24_ & ~n4896;
  assign n5226 = ~n5224 & ~n5225;
  assign n5227 = n5219 & n5222;
  assign n5228 = ~n5223 & n5227;
  assign n870 = ~n5226 | ~n5228;
  assign n5230 = ~n4409 & n4908;
  assign n5231 = ~n4477 & n4910;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = n4482 & n4897;
  assign n5234 = n4479 & n4901;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~n4495 & n4913;
  assign n5237 = ~n4519 & n4896;
  assign n5238 = P1_REG2_REG_25_ & ~n4896;
  assign n5239 = ~n5237 & ~n5238;
  assign n5240 = n5232 & n5235;
  assign n5241 = ~n5236 & n5240;
  assign n875 = ~n5239 | ~n5241;
  assign n5243 = ~n4473 & n4908;
  assign n5244 = ~n4534 & n4910;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = n4539 & n4897;
  assign n5247 = n4536 & n4901;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n4555 & n4913;
  assign n5250 = ~n4579 & n4896;
  assign n5251 = P1_REG2_REG_26_ & ~n4896;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = n5245 & n5248;
  assign n5254 = ~n5249 & n5253;
  assign n880 = ~n5252 | ~n5254;
  assign n5256 = ~n4530 & n4908;
  assign n5257 = ~n4594 & n4910;
  assign n5258 = ~n5256 & ~n5257;
  assign n5259 = n4599 & n4897;
  assign n5260 = n4596 & n4901;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n4612 & n4913;
  assign n5263 = ~n4638 & n4896;
  assign n5264 = P1_REG2_REG_27_ & ~n4896;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = n5258 & n5261;
  assign n5267 = ~n5262 & n5266;
  assign n885 = ~n5265 | ~n5267;
  assign n5269 = ~n4590 & n4908;
  assign n5270 = ~n4651 & n4910;
  assign n5271 = ~n5269 & ~n5270;
  assign n5272 = n4656 & n4897;
  assign n5273 = n4653 & n4901;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = ~n4674 & n4913;
  assign n5276 = ~n4702 & n4896;
  assign n5277 = P1_REG2_REG_28_ & ~n4896;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = n5271 & n5274;
  assign n5280 = ~n5275 & n5279;
  assign n890 = ~n5278 | ~n5280;
  assign n5282 = n4707 & n4901;
  assign n5283 = n4647 & n4908;
  assign n5284 = n4710 & n4897;
  assign n5285 = ~n4723 & n4913;
  assign n5286 = n4751 & ~n4754;
  assign n5287 = n4741 & n4755;
  assign n5288 = n5286 & n5287;
  assign n5289 = n4896 & ~n5288;
  assign n5290 = P1_REG2_REG_29_ & ~n4896;
  assign n5291 = ~n5289 & ~n5290;
  assign n5292 = ~n5282 & ~n5283;
  assign n5293 = ~n5284 & n5292;
  assign n5294 = ~n5285 & n5293;
  assign n895 = ~n5291 | ~n5294;
  assign n5296 = n4770 & n4896;
  assign n5297 = P1_REG2_REG_30_ & ~n4896;
  assign n5298 = ~n5296 & ~n5297;
  assign n5299 = n4763 & n4901;
  assign n5300 = n4773 & n4897;
  assign n5301 = n5298 & ~n5299;
  assign n900 = n5300 | ~n5301;
  assign n5303 = P1_REG2_REG_31_ & ~n4896;
  assign n5304 = ~n5296 & ~n5303;
  assign n5305 = n4780 & n4901;
  assign n5306 = n4784 & n4897;
  assign n5307 = n5304 & ~n5305;
  assign n905 = n5306 | ~n5307;
  assign n5309 = P1_STATE_REG & ~n2683;
  assign n5310 = n2683 & n2694;
  assign n5311 = n2695 & ~n2830;
  assign n5312 = n2683 & ~n5311;
  assign n5313 = ~n2856 & ~n5312;
  assign n1325 = ~P1_STATE_REG | n5313;
  assign n5315 = ~n5310 & ~n1325;
  assign n5316 = n5309 & ~n5315;
  assign n5317 = ~n2833 & ~n2855;
  assign n5318 = n5316 & n5317;
  assign n5319 = ~P1_REG2_REG_18_ & n4056;
  assign n5320 = P1_REG2_REG_19_ & n2764;
  assign n5321 = ~P1_REG2_REG_19_ & ~n2764;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = P1_REG2_REG_16_ & ~n3914;
  assign n5324 = P1_REG2_REG_17_ & n5323;
  assign n5325 = ~P1_REG2_REG_17_ & ~n5323;
  assign n5326 = ~n3981 & ~n5325;
  assign n5327 = ~P1_REG2_REG_16_ & n3914;
  assign n5328 = ~P1_REG2_REG_17_ & n3981;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = P1_REG2_REG_15_ & ~n3857;
  assign n5331 = ~P1_REG2_REG_15_ & n3857;
  assign n5332 = P1_REG2_REG_14_ & ~n3795;
  assign n5333 = ~P1_REG2_REG_14_ & n3795;
  assign n5334 = ~P1_REG2_REG_13_ & n3712;
  assign n5335 = P1_REG2_REG_13_ & ~n3712;
  assign n5336 = P1_REG2_REG_12_ & ~n3645;
  assign n5337 = P1_REG2_REG_11_ & ~n3575;
  assign n5338 = ~P1_REG2_REG_12_ & n3645;
  assign n5339 = ~n5334 & ~n5338;
  assign n5340 = n5337 & n5339;
  assign n5341 = ~n5335 & ~n5336;
  assign n5342 = ~n5340 & n5341;
  assign n5343 = ~n5334 & ~n5342;
  assign n5344 = ~P1_REG2_REG_11_ & n3575;
  assign n5345 = ~P1_REG2_REG_10_ & n3522;
  assign n5346 = P1_REG2_REG_10_ & ~n3522;
  assign n5347 = P1_REG2_REG_9_ & ~n3455;
  assign n5348 = P1_REG2_REG_8_ & ~n3387;
  assign n5349 = ~P1_REG2_REG_9_ & n3455;
  assign n5350 = ~n5345 & ~n5349;
  assign n5351 = n5348 & n5350;
  assign n5352 = ~n5346 & ~n5347;
  assign n5353 = ~n5351 & n5352;
  assign n5354 = ~n5345 & ~n5353;
  assign n5355 = ~P1_REG2_REG_8_ & n3387;
  assign n5356 = P1_REG2_REG_6_ & ~n3244;
  assign n5357 = P1_REG2_REG_7_ & n5356;
  assign n5358 = ~P1_REG2_REG_7_ & ~n5356;
  assign n5359 = ~n3318 & ~n5358;
  assign n5360 = ~P1_REG2_REG_6_ & n3244;
  assign n5361 = ~P1_REG2_REG_7_ & n3318;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = P1_REG2_REG_4_ & ~n3111;
  assign n5364 = P1_REG2_REG_5_ & n5363;
  assign n5365 = ~P1_REG2_REG_5_ & ~n5363;
  assign n5366 = ~n3180 & ~n5365;
  assign n5367 = ~P1_REG2_REG_4_ & n3111;
  assign n5368 = ~P1_REG2_REG_5_ & n3180;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = P1_REG2_REG_3_ & ~n3045;
  assign n5371 = ~P1_REG2_REG_3_ & n3045;
  assign n5372 = P1_REG2_REG_2_ & ~n2981;
  assign n5373 = ~n5371 & n5372;
  assign n5374 = ~P1_REG2_REG_2_ & n2981;
  assign n5375 = ~n5371 & ~n5374;
  assign n5376 = P1_REG2_REG_0_ & ~n2859;
  assign n5377 = ~P1_REG2_REG_1_ & n2925;
  assign n5378 = n5376 & ~n5377;
  assign n5379 = P1_REG2_REG_1_ & ~n2925;
  assign n5380 = ~n5378 & ~n5379;
  assign n5381 = n5375 & ~n5380;
  assign n5382 = ~n5370 & ~n5373;
  assign n5383 = ~n5381 & n5382;
  assign n5384 = n5369 & ~n5383;
  assign n5385 = ~n5364 & ~n5366;
  assign n5386 = ~n5384 & n5385;
  assign n5387 = n5362 & ~n5386;
  assign n5388 = ~n5357 & ~n5359;
  assign n5389 = ~n5387 & n5388;
  assign n5390 = n5350 & ~n5355;
  assign n5391 = ~n5389 & n5390;
  assign n5392 = ~n5354 & ~n5391;
  assign n5393 = n5339 & ~n5344;
  assign n5394 = ~n5392 & n5393;
  assign n5395 = ~n5343 & ~n5394;
  assign n5396 = ~n5333 & ~n5395;
  assign n5397 = ~n5332 & ~n5396;
  assign n5398 = ~n5331 & ~n5397;
  assign n5399 = ~n5330 & ~n5398;
  assign n5400 = n5329 & ~n5399;
  assign n5401 = ~n5324 & ~n5326;
  assign n5402 = ~n5400 & n5401;
  assign n5403 = P1_REG2_REG_18_ & ~n4056;
  assign n5404 = n5402 & ~n5403;
  assign n5405 = ~n5319 & ~n5322;
  assign n5406 = ~n5404 & n5405;
  assign n5407 = ~n5319 & ~n5402;
  assign n5408 = n5322 & ~n5403;
  assign n5409 = ~n5407 & n5408;
  assign n5410 = ~n5406 & ~n5409;
  assign n5411 = n5318 & n5410;
  assign n5412 = P1_REG3_REG_19_ & ~P1_STATE_REG;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = P1_ADDR_REG_19_ & n5315;
  assign n5415 = n2833 & n5316;
  assign n5416 = ~n2764 & n5415;
  assign n5417 = n2855 & n5316;
  assign n5418 = ~P1_REG1_REG_18_ & n4056;
  assign n5419 = P1_REG1_REG_19_ & n2764;
  assign n5420 = ~P1_REG1_REG_19_ & ~n2764;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = P1_REG1_REG_16_ & ~n3914;
  assign n5423 = P1_REG1_REG_17_ & n5422;
  assign n5424 = ~P1_REG1_REG_17_ & ~n5422;
  assign n5425 = ~n3981 & ~n5424;
  assign n5426 = ~P1_REG1_REG_16_ & n3914;
  assign n5427 = ~P1_REG1_REG_17_ & n3981;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = P1_REG1_REG_15_ & ~n3857;
  assign n5430 = ~P1_REG1_REG_15_ & n3857;
  assign n5431 = P1_REG1_REG_14_ & ~n3795;
  assign n5432 = ~P1_REG1_REG_14_ & n3795;
  assign n5433 = ~P1_REG1_REG_13_ & n3712;
  assign n5434 = P1_REG1_REG_13_ & ~n3712;
  assign n5435 = P1_REG1_REG_12_ & ~n3645;
  assign n5436 = P1_REG1_REG_11_ & ~n3575;
  assign n5437 = ~P1_REG1_REG_12_ & n3645;
  assign n5438 = ~n5433 & ~n5437;
  assign n5439 = n5436 & n5438;
  assign n5440 = ~n5434 & ~n5435;
  assign n5441 = ~n5439 & n5440;
  assign n5442 = ~n5433 & ~n5441;
  assign n5443 = ~P1_REG1_REG_11_ & n3575;
  assign n5444 = ~P1_REG1_REG_10_ & n3522;
  assign n5445 = P1_REG1_REG_10_ & ~n3522;
  assign n5446 = P1_REG1_REG_9_ & ~n3455;
  assign n5447 = P1_REG1_REG_8_ & ~n3387;
  assign n5448 = ~P1_REG1_REG_9_ & n3455;
  assign n5449 = ~n5444 & ~n5448;
  assign n5450 = n5447 & n5449;
  assign n5451 = ~n5445 & ~n5446;
  assign n5452 = ~n5450 & n5451;
  assign n5453 = ~n5444 & ~n5452;
  assign n5454 = ~P1_REG1_REG_8_ & n3387;
  assign n5455 = P1_REG1_REG_6_ & ~n3244;
  assign n5456 = P1_REG1_REG_7_ & n5455;
  assign n5457 = ~P1_REG1_REG_7_ & ~n5455;
  assign n5458 = ~n3318 & ~n5457;
  assign n5459 = ~P1_REG1_REG_6_ & n3244;
  assign n5460 = ~P1_REG1_REG_7_ & n3318;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = P1_REG1_REG_4_ & ~n3111;
  assign n5463 = P1_REG1_REG_5_ & n5462;
  assign n5464 = ~P1_REG1_REG_5_ & ~n5462;
  assign n5465 = ~n3180 & ~n5464;
  assign n5466 = ~P1_REG1_REG_4_ & n3111;
  assign n5467 = ~P1_REG1_REG_5_ & n3180;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = P1_REG1_REG_3_ & ~n3045;
  assign n5470 = ~P1_REG1_REG_3_ & n3045;
  assign n5471 = P1_REG1_REG_2_ & ~n2981;
  assign n5472 = ~n5470 & n5471;
  assign n5473 = ~P1_REG1_REG_2_ & n2981;
  assign n5474 = ~n5470 & ~n5473;
  assign n5475 = P1_REG1_REG_0_ & ~n2859;
  assign n5476 = ~P1_REG1_REG_1_ & n2925;
  assign n5477 = n5475 & ~n5476;
  assign n5478 = P1_REG1_REG_1_ & ~n2925;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = n5474 & ~n5479;
  assign n5481 = ~n5469 & ~n5472;
  assign n5482 = ~n5480 & n5481;
  assign n5483 = n5468 & ~n5482;
  assign n5484 = ~n5463 & ~n5465;
  assign n5485 = ~n5483 & n5484;
  assign n5486 = n5461 & ~n5485;
  assign n5487 = ~n5456 & ~n5458;
  assign n5488 = ~n5486 & n5487;
  assign n5489 = n5449 & ~n5454;
  assign n5490 = ~n5488 & n5489;
  assign n5491 = ~n5453 & ~n5490;
  assign n5492 = n5438 & ~n5443;
  assign n5493 = ~n5491 & n5492;
  assign n5494 = ~n5442 & ~n5493;
  assign n5495 = ~n5432 & ~n5494;
  assign n5496 = ~n5431 & ~n5495;
  assign n5497 = ~n5430 & ~n5496;
  assign n5498 = ~n5429 & ~n5497;
  assign n5499 = n5428 & ~n5498;
  assign n5500 = ~n5423 & ~n5425;
  assign n5501 = ~n5499 & n5500;
  assign n5502 = P1_REG1_REG_18_ & ~n4056;
  assign n5503 = n5501 & ~n5502;
  assign n5504 = ~n5418 & ~n5421;
  assign n5505 = ~n5503 & n5504;
  assign n5506 = ~n5418 & ~n5501;
  assign n5507 = n5421 & ~n5502;
  assign n5508 = ~n5506 & n5507;
  assign n5509 = ~n5505 & ~n5508;
  assign n5510 = n5417 & n5509;
  assign n5511 = ~n5414 & ~n5416;
  assign n5512 = ~n5510 & n5511;
  assign n5513 = n2696 & ~n5315;
  assign n5514 = ~n2887 & ~n2896;
  assign n5515 = ~n2904 & n5514;
  assign n5516 = ~n2892 & ~n4912;
  assign n5517 = ~n2890 & n5516;
  assign n5518 = ~n2898 & ~n2901;
  assign n5519 = ~n4889 & n5518;
  assign n5520 = n5515 & n5517;
  assign n5521 = n5519 & n5520;
  assign n5522 = n4900 & n5521;
  assign n5523 = ~n4890 & n5522;
  assign n5524 = n2833 & ~n5523;
  assign n5525 = ~n2764 & n5524;
  assign n5526 = n5317 & ~n5523;
  assign n5527 = n5410 & n5526;
  assign n5528 = n2855 & ~n5523;
  assign n5529 = n5509 & n5528;
  assign n5530 = ~n5525 & ~n5527;
  assign n5531 = ~n5529 & n5530;
  assign n5532 = n5513 & ~n5531;
  assign n5533 = n5413 & n5512;
  assign n910 = n5532 | ~n5533;
  assign n5535 = P1_REG2_REG_18_ & n4056;
  assign n5536 = ~P1_REG2_REG_18_ & ~n4056;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = n5402 & ~n5537;
  assign n5539 = ~n5402 & n5537;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = n5318 & ~n5540;
  assign n5542 = P1_REG3_REG_18_ & ~P1_STATE_REG;
  assign n5543 = ~n5541 & ~n5542;
  assign n5544 = P1_ADDR_REG_18_ & n5315;
  assign n5545 = ~n4056 & n5415;
  assign n5546 = P1_REG1_REG_18_ & n4056;
  assign n5547 = ~P1_REG1_REG_18_ & ~n4056;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = n5501 & ~n5548;
  assign n5550 = ~n5501 & n5548;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = n5417 & ~n5551;
  assign n5553 = ~n5544 & ~n5545;
  assign n5554 = ~n5552 & n5553;
  assign n5555 = ~n4056 & n5524;
  assign n5556 = n5526 & ~n5540;
  assign n5557 = n5528 & ~n5551;
  assign n5558 = ~n5555 & ~n5556;
  assign n5559 = ~n5557 & n5558;
  assign n5560 = n5513 & ~n5559;
  assign n5561 = n5543 & n5554;
  assign n915 = n5560 | ~n5561;
  assign n5563 = P1_REG2_REG_17_ & ~n3981;
  assign n5564 = ~n5323 & n5399;
  assign n5565 = n5329 & ~n5563;
  assign n5566 = ~n5564 & n5565;
  assign n5567 = P1_REG2_REG_17_ & n3981;
  assign n5568 = ~P1_REG2_REG_17_ & ~n3981;
  assign n5569 = ~n5327 & ~n5399;
  assign n5570 = ~n5567 & ~n5568;
  assign n5571 = ~n5323 & n5570;
  assign n5572 = ~n5569 & n5571;
  assign n5573 = ~n5566 & ~n5572;
  assign n5574 = n5318 & n5573;
  assign n5575 = P1_REG3_REG_17_ & ~P1_STATE_REG;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = P1_ADDR_REG_17_ & n5315;
  assign n5578 = ~n3981 & n5415;
  assign n5579 = P1_REG1_REG_17_ & ~n3981;
  assign n5580 = ~n5422 & n5498;
  assign n5581 = n5428 & ~n5579;
  assign n5582 = ~n5580 & n5581;
  assign n5583 = P1_REG1_REG_17_ & n3981;
  assign n5584 = ~P1_REG1_REG_17_ & ~n3981;
  assign n5585 = ~n5426 & ~n5498;
  assign n5586 = ~n5583 & ~n5584;
  assign n5587 = ~n5422 & n5586;
  assign n5588 = ~n5585 & n5587;
  assign n5589 = ~n5582 & ~n5588;
  assign n5590 = n5417 & n5589;
  assign n5591 = ~n5577 & ~n5578;
  assign n5592 = ~n5590 & n5591;
  assign n5593 = ~n3981 & n5524;
  assign n5594 = n5526 & n5573;
  assign n5595 = n5528 & n5589;
  assign n5596 = ~n5593 & ~n5594;
  assign n5597 = ~n5595 & n5596;
  assign n5598 = n5513 & ~n5597;
  assign n5599 = n5576 & n5592;
  assign n920 = n5598 | ~n5599;
  assign n5601 = P1_REG2_REG_16_ & n3914;
  assign n5602 = ~P1_REG2_REG_16_ & ~n3914;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = n5399 & ~n5603;
  assign n5605 = ~n5323 & ~n5327;
  assign n5606 = ~n5399 & ~n5605;
  assign n5607 = ~n5604 & ~n5606;
  assign n5608 = n5318 & ~n5607;
  assign n5609 = P1_REG3_REG_16_ & ~P1_STATE_REG;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = P1_ADDR_REG_16_ & n5315;
  assign n5612 = ~n3914 & n5415;
  assign n5613 = P1_REG1_REG_16_ & n3914;
  assign n5614 = ~P1_REG1_REG_16_ & ~n3914;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = n5498 & ~n5615;
  assign n5617 = ~n5422 & ~n5426;
  assign n5618 = ~n5498 & ~n5617;
  assign n5619 = ~n5616 & ~n5618;
  assign n5620 = n5417 & ~n5619;
  assign n5621 = ~n5611 & ~n5612;
  assign n5622 = ~n5620 & n5621;
  assign n5623 = ~n3914 & n5524;
  assign n5624 = n5526 & ~n5607;
  assign n5625 = n5528 & ~n5619;
  assign n5626 = ~n5623 & ~n5624;
  assign n5627 = ~n5625 & n5626;
  assign n5628 = n5513 & ~n5627;
  assign n5629 = n5610 & n5622;
  assign n925 = n5628 | ~n5629;
  assign n5631 = P1_REG2_REG_15_ & n3857;
  assign n5632 = ~P1_REG2_REG_15_ & ~n3857;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = n5397 & ~n5633;
  assign n5635 = ~n5397 & n5633;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = n5318 & ~n5636;
  assign n5638 = P1_REG3_REG_15_ & ~P1_STATE_REG;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = P1_ADDR_REG_15_ & n5315;
  assign n5641 = ~n3857 & n5415;
  assign n5642 = P1_REG1_REG_15_ & n3857;
  assign n5643 = ~P1_REG1_REG_15_ & ~n3857;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = n5496 & ~n5644;
  assign n5646 = ~n5496 & n5644;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = n5417 & ~n5647;
  assign n5649 = ~n5640 & ~n5641;
  assign n5650 = ~n5648 & n5649;
  assign n5651 = ~n3857 & n5524;
  assign n5652 = n5526 & ~n5636;
  assign n5653 = n5528 & ~n5647;
  assign n5654 = ~n5651 & ~n5652;
  assign n5655 = ~n5653 & n5654;
  assign n5656 = n5513 & ~n5655;
  assign n5657 = n5639 & n5650;
  assign n930 = n5656 | ~n5657;
  assign n5659 = P1_REG2_REG_14_ & n3795;
  assign n5660 = ~P1_REG2_REG_14_ & ~n3795;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = n5395 & ~n5661;
  assign n5663 = ~n5395 & n5661;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = n5318 & ~n5664;
  assign n5666 = P1_REG3_REG_14_ & ~P1_STATE_REG;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = P1_ADDR_REG_14_ & n5315;
  assign n5669 = ~n3795 & n5415;
  assign n5670 = P1_REG1_REG_14_ & n3795;
  assign n5671 = ~P1_REG1_REG_14_ & ~n3795;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = n5494 & ~n5672;
  assign n5674 = ~n5494 & n5672;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = n5417 & ~n5675;
  assign n5677 = ~n5668 & ~n5669;
  assign n5678 = ~n5676 & n5677;
  assign n5679 = ~n3795 & n5524;
  assign n5680 = n5526 & ~n5664;
  assign n5681 = n5528 & ~n5675;
  assign n5682 = ~n5679 & ~n5680;
  assign n5683 = ~n5681 & n5682;
  assign n5684 = n5513 & ~n5683;
  assign n5685 = n5667 & n5678;
  assign n935 = n5684 | ~n5685;
  assign n5687 = ~n5344 & ~n5392;
  assign n5688 = ~n5337 & ~n5687;
  assign n5689 = ~n5336 & n5688;
  assign n5690 = ~n5335 & n5339;
  assign n5691 = ~n5689 & n5690;
  assign n5692 = P1_REG2_REG_13_ & n3712;
  assign n5693 = ~P1_REG2_REG_13_ & ~n3712;
  assign n5694 = ~n5338 & ~n5688;
  assign n5695 = ~n5692 & ~n5693;
  assign n5696 = ~n5336 & n5695;
  assign n5697 = ~n5694 & n5696;
  assign n5698 = ~n5691 & ~n5697;
  assign n5699 = n5318 & n5698;
  assign n5700 = P1_REG3_REG_13_ & ~P1_STATE_REG;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = P1_ADDR_REG_13_ & n5315;
  assign n5703 = ~n3712 & n5415;
  assign n5704 = ~n5443 & ~n5491;
  assign n5705 = ~n5436 & ~n5704;
  assign n5706 = ~n5435 & n5705;
  assign n5707 = ~n5434 & n5438;
  assign n5708 = ~n5706 & n5707;
  assign n5709 = P1_REG1_REG_13_ & n3712;
  assign n5710 = ~P1_REG1_REG_13_ & ~n3712;
  assign n5711 = ~n5437 & ~n5705;
  assign n5712 = ~n5709 & ~n5710;
  assign n5713 = ~n5435 & n5712;
  assign n5714 = ~n5711 & n5713;
  assign n5715 = ~n5708 & ~n5714;
  assign n5716 = n5417 & n5715;
  assign n5717 = ~n5702 & ~n5703;
  assign n5718 = ~n5716 & n5717;
  assign n5719 = ~n3712 & n5524;
  assign n5720 = n5526 & n5698;
  assign n5721 = n5528 & n5715;
  assign n5722 = ~n5719 & ~n5720;
  assign n5723 = ~n5721 & n5722;
  assign n5724 = n5513 & ~n5723;
  assign n5725 = n5701 & n5718;
  assign n940 = n5724 | ~n5725;
  assign n5727 = P1_REG2_REG_12_ & n3645;
  assign n5728 = ~P1_REG2_REG_12_ & ~n3645;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = n5688 & ~n5729;
  assign n5731 = ~n5336 & ~n5338;
  assign n5732 = ~n5688 & ~n5731;
  assign n5733 = ~n5730 & ~n5732;
  assign n5734 = n5318 & ~n5733;
  assign n5735 = P1_REG3_REG_12_ & ~P1_STATE_REG;
  assign n5736 = ~n5734 & ~n5735;
  assign n5737 = P1_ADDR_REG_12_ & n5315;
  assign n5738 = ~n3645 & n5415;
  assign n5739 = P1_REG1_REG_12_ & n3645;
  assign n5740 = ~P1_REG1_REG_12_ & ~n3645;
  assign n5741 = ~n5739 & ~n5740;
  assign n5742 = n5705 & ~n5741;
  assign n5743 = ~n5435 & ~n5437;
  assign n5744 = ~n5705 & ~n5743;
  assign n5745 = ~n5742 & ~n5744;
  assign n5746 = n5417 & ~n5745;
  assign n5747 = ~n5737 & ~n5738;
  assign n5748 = ~n5746 & n5747;
  assign n5749 = ~n3645 & n5524;
  assign n5750 = n5526 & ~n5733;
  assign n5751 = n5528 & ~n5745;
  assign n5752 = ~n5749 & ~n5750;
  assign n5753 = ~n5751 & n5752;
  assign n5754 = n5513 & ~n5753;
  assign n5755 = n5736 & n5748;
  assign n945 = n5754 | ~n5755;
  assign n5757 = P1_REG2_REG_11_ & n3575;
  assign n5758 = ~P1_REG2_REG_11_ & ~n3575;
  assign n5759 = ~n5757 & ~n5758;
  assign n5760 = n5392 & ~n5759;
  assign n5761 = ~n5337 & ~n5344;
  assign n5762 = ~n5392 & ~n5761;
  assign n5763 = ~n5760 & ~n5762;
  assign n5764 = n5318 & ~n5763;
  assign n5765 = P1_REG3_REG_11_ & ~P1_STATE_REG;
  assign n5766 = ~n5764 & ~n5765;
  assign n5767 = P1_ADDR_REG_11_ & n5315;
  assign n5768 = ~n3575 & n5415;
  assign n5769 = P1_REG1_REG_11_ & n3575;
  assign n5770 = ~P1_REG1_REG_11_ & ~n3575;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = n5491 & ~n5771;
  assign n5773 = ~n5436 & ~n5443;
  assign n5774 = ~n5491 & ~n5773;
  assign n5775 = ~n5772 & ~n5774;
  assign n5776 = n5417 & ~n5775;
  assign n5777 = ~n5767 & ~n5768;
  assign n5778 = ~n5776 & n5777;
  assign n5779 = ~n3575 & n5524;
  assign n5780 = n5526 & ~n5763;
  assign n5781 = n5528 & ~n5775;
  assign n5782 = ~n5779 & ~n5780;
  assign n5783 = ~n5781 & n5782;
  assign n5784 = n5513 & ~n5783;
  assign n5785 = n5766 & n5778;
  assign n950 = n5784 | ~n5785;
  assign n5787 = ~n5355 & ~n5389;
  assign n5788 = ~n5348 & ~n5787;
  assign n5789 = ~n5347 & n5788;
  assign n5790 = ~n5346 & n5350;
  assign n5791 = ~n5789 & n5790;
  assign n5792 = P1_REG2_REG_10_ & n3522;
  assign n5793 = ~P1_REG2_REG_10_ & ~n3522;
  assign n5794 = ~n5349 & ~n5788;
  assign n5795 = ~n5792 & ~n5793;
  assign n5796 = ~n5347 & n5795;
  assign n5797 = ~n5794 & n5796;
  assign n5798 = ~n5791 & ~n5797;
  assign n5799 = n5318 & n5798;
  assign n5800 = P1_REG3_REG_10_ & ~P1_STATE_REG;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = P1_ADDR_REG_10_ & n5315;
  assign n5803 = ~n3522 & n5415;
  assign n5804 = ~n5454 & ~n5488;
  assign n5805 = ~n5447 & ~n5804;
  assign n5806 = ~n5446 & n5805;
  assign n5807 = ~n5445 & n5449;
  assign n5808 = ~n5806 & n5807;
  assign n5809 = P1_REG1_REG_10_ & n3522;
  assign n5810 = ~P1_REG1_REG_10_ & ~n3522;
  assign n5811 = ~n5448 & ~n5805;
  assign n5812 = ~n5809 & ~n5810;
  assign n5813 = ~n5446 & n5812;
  assign n5814 = ~n5811 & n5813;
  assign n5815 = ~n5808 & ~n5814;
  assign n5816 = n5417 & n5815;
  assign n5817 = ~n5802 & ~n5803;
  assign n5818 = ~n5816 & n5817;
  assign n5819 = ~n3522 & n5524;
  assign n5820 = n5526 & n5798;
  assign n5821 = n5528 & n5815;
  assign n5822 = ~n5819 & ~n5820;
  assign n5823 = ~n5821 & n5822;
  assign n5824 = n5513 & ~n5823;
  assign n5825 = n5801 & n5818;
  assign n955 = n5824 | ~n5825;
  assign n5827 = P1_REG2_REG_9_ & n3455;
  assign n5828 = ~P1_REG2_REG_9_ & ~n3455;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = n5788 & ~n5829;
  assign n5831 = ~n5347 & ~n5349;
  assign n5832 = ~n5788 & ~n5831;
  assign n5833 = ~n5830 & ~n5832;
  assign n5834 = n5318 & ~n5833;
  assign n5835 = P1_REG3_REG_9_ & ~P1_STATE_REG;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = P1_ADDR_REG_9_ & n5315;
  assign n5838 = ~n3455 & n5415;
  assign n5839 = P1_REG1_REG_9_ & n3455;
  assign n5840 = ~P1_REG1_REG_9_ & ~n3455;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = n5805 & ~n5841;
  assign n5843 = ~n5446 & ~n5448;
  assign n5844 = ~n5805 & ~n5843;
  assign n5845 = ~n5842 & ~n5844;
  assign n5846 = n5417 & ~n5845;
  assign n5847 = ~n5837 & ~n5838;
  assign n5848 = ~n5846 & n5847;
  assign n5849 = ~n3455 & n5524;
  assign n5850 = n5526 & ~n5833;
  assign n5851 = n5528 & ~n5845;
  assign n5852 = ~n5849 & ~n5850;
  assign n5853 = ~n5851 & n5852;
  assign n5854 = n5513 & ~n5853;
  assign n5855 = n5836 & n5848;
  assign n960 = n5854 | ~n5855;
  assign n5857 = P1_REG2_REG_8_ & n3387;
  assign n5858 = ~P1_REG2_REG_8_ & ~n3387;
  assign n5859 = ~n5857 & ~n5858;
  assign n5860 = n5389 & ~n5859;
  assign n5861 = ~n5348 & ~n5355;
  assign n5862 = ~n5389 & ~n5861;
  assign n5863 = ~n5860 & ~n5862;
  assign n5864 = n5318 & ~n5863;
  assign n5865 = P1_REG3_REG_8_ & ~P1_STATE_REG;
  assign n5866 = ~n5864 & ~n5865;
  assign n5867 = P1_ADDR_REG_8_ & n5315;
  assign n5868 = ~n3387 & n5415;
  assign n5869 = P1_REG1_REG_8_ & n3387;
  assign n5870 = ~P1_REG1_REG_8_ & ~n3387;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = n5488 & ~n5871;
  assign n5873 = ~n5447 & ~n5454;
  assign n5874 = ~n5488 & ~n5873;
  assign n5875 = ~n5872 & ~n5874;
  assign n5876 = n5417 & ~n5875;
  assign n5877 = ~n5867 & ~n5868;
  assign n5878 = ~n5876 & n5877;
  assign n5879 = ~n3387 & n5524;
  assign n5880 = n5526 & ~n5863;
  assign n5881 = n5528 & ~n5875;
  assign n5882 = ~n5879 & ~n5880;
  assign n5883 = ~n5881 & n5882;
  assign n5884 = n5513 & ~n5883;
  assign n5885 = n5866 & n5878;
  assign n965 = n5884 | ~n5885;
  assign n5887 = P1_REG2_REG_7_ & ~n3318;
  assign n5888 = ~n5356 & n5386;
  assign n5889 = n5362 & ~n5887;
  assign n5890 = ~n5888 & n5889;
  assign n5891 = P1_REG2_REG_7_ & n3318;
  assign n5892 = ~P1_REG2_REG_7_ & ~n3318;
  assign n5893 = ~n5360 & ~n5386;
  assign n5894 = ~n5891 & ~n5892;
  assign n5895 = ~n5356 & n5894;
  assign n5896 = ~n5893 & n5895;
  assign n5897 = ~n5890 & ~n5896;
  assign n5898 = n5318 & n5897;
  assign n5899 = P1_REG3_REG_7_ & ~P1_STATE_REG;
  assign n5900 = ~n5898 & ~n5899;
  assign n5901 = P1_REG1_REG_7_ & ~n3318;
  assign n5902 = ~n5455 & n5485;
  assign n5903 = n5461 & ~n5901;
  assign n5904 = ~n5902 & n5903;
  assign n5905 = P1_REG1_REG_7_ & n3318;
  assign n5906 = ~P1_REG1_REG_7_ & ~n3318;
  assign n5907 = ~n5459 & ~n5485;
  assign n5908 = ~n5905 & ~n5906;
  assign n5909 = ~n5455 & n5908;
  assign n5910 = ~n5907 & n5909;
  assign n5911 = ~n5904 & ~n5910;
  assign n5912 = n5417 & n5911;
  assign n5913 = ~n3318 & n5415;
  assign n5914 = P1_ADDR_REG_7_ & n5315;
  assign n5915 = ~n5912 & ~n5913;
  assign n5916 = ~n5914 & n5915;
  assign n5917 = ~n3318 & n5524;
  assign n5918 = n5526 & n5897;
  assign n5919 = n5528 & n5911;
  assign n5920 = ~n5917 & ~n5918;
  assign n5921 = ~n5919 & n5920;
  assign n5922 = n5513 & ~n5921;
  assign n5923 = n5900 & n5916;
  assign n970 = n5922 | ~n5923;
  assign n5925 = P1_REG1_REG_6_ & n3244;
  assign n5926 = ~P1_REG1_REG_6_ & ~n3244;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = n5485 & ~n5927;
  assign n5929 = ~n5455 & ~n5459;
  assign n5930 = ~n5485 & ~n5929;
  assign n5931 = ~n5928 & ~n5930;
  assign n5932 = n5417 & ~n5931;
  assign n5933 = ~n3244 & n5415;
  assign n5934 = P1_ADDR_REG_6_ & n5315;
  assign n5935 = ~n5932 & ~n5933;
  assign n5936 = ~n5934 & n5935;
  assign n5937 = P1_REG2_REG_6_ & n3244;
  assign n5938 = ~P1_REG2_REG_6_ & ~n3244;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = n5386 & ~n5939;
  assign n5941 = ~n5356 & ~n5360;
  assign n5942 = ~n5386 & ~n5941;
  assign n5943 = ~n5940 & ~n5942;
  assign n5944 = n5318 & ~n5943;
  assign n5945 = P1_REG3_REG_6_ & ~P1_STATE_REG;
  assign n5946 = ~n3244 & n5524;
  assign n5947 = n5526 & ~n5943;
  assign n5948 = n5528 & ~n5931;
  assign n5949 = ~n5946 & ~n5947;
  assign n5950 = ~n5948 & n5949;
  assign n5951 = n5513 & ~n5950;
  assign n5952 = ~n5944 & ~n5945;
  assign n5953 = ~n5951 & n5952;
  assign n975 = ~n5936 | ~n5953;
  assign n5955 = P1_REG1_REG_5_ & ~n3180;
  assign n5956 = n5474 & n5477;
  assign n5957 = ~n5473 & n5478;
  assign n5958 = ~n5471 & ~n5957;
  assign n5959 = ~n5470 & ~n5958;
  assign n5960 = ~n5469 & ~n5956;
  assign n5961 = ~n5959 & n5960;
  assign n5962 = ~n5462 & n5961;
  assign n5963 = n5468 & ~n5955;
  assign n5964 = ~n5962 & n5963;
  assign n5965 = P1_REG1_REG_5_ & n3180;
  assign n5966 = ~P1_REG1_REG_5_ & ~n3180;
  assign n5967 = ~n5466 & ~n5961;
  assign n5968 = ~n5965 & ~n5966;
  assign n5969 = ~n5462 & n5968;
  assign n5970 = ~n5967 & n5969;
  assign n5971 = ~n5964 & ~n5970;
  assign n5972 = n5417 & n5971;
  assign n5973 = ~n3180 & n5415;
  assign n5974 = P1_ADDR_REG_5_ & n5315;
  assign n5975 = ~n5972 & ~n5973;
  assign n5976 = ~n5974 & n5975;
  assign n5977 = P1_REG2_REG_5_ & ~n3180;
  assign n5978 = n5375 & n5378;
  assign n5979 = ~n5374 & n5379;
  assign n5980 = ~n5372 & ~n5979;
  assign n5981 = ~n5371 & ~n5980;
  assign n5982 = ~n5370 & ~n5978;
  assign n5983 = ~n5981 & n5982;
  assign n5984 = ~n5363 & n5983;
  assign n5985 = n5369 & ~n5977;
  assign n5986 = ~n5984 & n5985;
  assign n5987 = P1_REG2_REG_5_ & n3180;
  assign n5988 = ~P1_REG2_REG_5_ & ~n3180;
  assign n5989 = ~n5367 & ~n5983;
  assign n5990 = ~n5987 & ~n5988;
  assign n5991 = ~n5363 & n5990;
  assign n5992 = ~n5989 & n5991;
  assign n5993 = ~n5986 & ~n5992;
  assign n5994 = n5318 & n5993;
  assign n5995 = P1_REG3_REG_5_ & ~P1_STATE_REG;
  assign n5996 = ~n3180 & n5524;
  assign n5997 = n5526 & n5993;
  assign n5998 = n5528 & n5971;
  assign n5999 = ~n5996 & ~n5997;
  assign n6000 = ~n5998 & n5999;
  assign n6001 = n5513 & ~n6000;
  assign n6002 = ~n5994 & ~n5995;
  assign n6003 = ~n6001 & n6002;
  assign n980 = ~n5976 | ~n6003;
  assign n6005 = P1_REG1_REG_4_ & n3111;
  assign n6006 = ~P1_REG1_REG_4_ & ~n3111;
  assign n6007 = ~n6005 & ~n6006;
  assign n6008 = n5961 & ~n6007;
  assign n6009 = ~n5462 & ~n5466;
  assign n6010 = ~n5961 & ~n6009;
  assign n6011 = ~n6008 & ~n6010;
  assign n6012 = n5417 & ~n6011;
  assign n6013 = ~n3111 & n5415;
  assign n6014 = P1_ADDR_REG_4_ & n5315;
  assign n6015 = ~n6012 & ~n6013;
  assign n6016 = ~n6014 & n6015;
  assign n6017 = P1_REG3_REG_4_ & ~P1_STATE_REG;
  assign n6018 = P1_REG2_REG_4_ & n3111;
  assign n6019 = ~P1_REG2_REG_4_ & ~n3111;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n5983 & ~n6020;
  assign n6022 = ~n5363 & ~n5367;
  assign n6023 = ~n5983 & ~n6022;
  assign n6024 = ~n6021 & ~n6023;
  assign n6025 = n5318 & ~n6024;
  assign n6026 = ~n3111 & n5524;
  assign n6027 = n5526 & ~n6024;
  assign n6028 = n5528 & ~n6011;
  assign n6029 = ~n6026 & ~n6027;
  assign n6030 = ~n6028 & n6029;
  assign n6031 = n5513 & ~n6030;
  assign n1330 = P1_STATE_REG & n5310;
  assign n6033 = P1_REG2_REG_0_ & n5317;
  assign n6034 = n2859 & n6033;
  assign n6035 = ~P1_REG2_REG_0_ & ~n2855;
  assign n6036 = ~n2833 & ~n6035;
  assign n6037 = ~n2859 & ~n6036;
  assign n6038 = n2758 & ~n2764;
  assign n6039 = ~n2755 & ~n2758;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n2694 & n2863;
  assign n6042 = n6040 & ~n6041;
  assign n6043 = ~n2694 & ~n6042;
  assign n6044 = ~n2866 & ~n2887;
  assign n6045 = ~n2896 & n6044;
  assign n6046 = ~n2694 & ~n6045;
  assign n6047 = ~n2694 & n6038;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = ~n2878 & ~n6048;
  assign n6050 = n2694 & ~n2859;
  assign n6051 = ~n2694 & ~n5516;
  assign n6052 = ~n2862 & n6051;
  assign n6053 = ~n6049 & ~n6050;
  assign n6054 = ~n6052 & n6053;
  assign n6055 = n6043 & n6054;
  assign n6056 = ~n6043 & ~n6054;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n2878 & n6051;
  assign n6059 = P1_REG1_REG_0_ & n2694;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = ~n6041 & n6048;
  assign n6062 = ~n2862 & ~n6061;
  assign n6063 = n6060 & ~n6062;
  assign n6064 = ~n6043 & ~n6063;
  assign n6065 = n6043 & n6063;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = ~n6057 & n6066;
  assign n6068 = n6057 & ~n6066;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n2833 & n2855;
  assign n6071 = ~n6069 & n6070;
  assign n6072 = ~n6034 & ~n6037;
  assign n6073 = ~n6071 & n6072;
  assign n6074 = n1330 & ~n6073;
  assign n6075 = ~n6031 & ~n6074;
  assign n6076 = ~n6017 & ~n6025;
  assign n6077 = n6075 & n6076;
  assign n985 = ~n6016 | ~n6077;
  assign n6079 = ~n5473 & n5477;
  assign n6080 = n5958 & ~n6079;
  assign n6081 = P1_REG1_REG_3_ & n3045;
  assign n6082 = ~P1_REG1_REG_3_ & ~n3045;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = n6080 & ~n6083;
  assign n6085 = ~n5469 & ~n5470;
  assign n6086 = ~n6080 & ~n6085;
  assign n6087 = ~n6084 & ~n6086;
  assign n6088 = n5417 & ~n6087;
  assign n6089 = ~n3045 & n5415;
  assign n6090 = P1_ADDR_REG_3_ & n5315;
  assign n6091 = ~n6088 & ~n6089;
  assign n6092 = ~n6090 & n6091;
  assign n6093 = ~n5374 & n5378;
  assign n6094 = n5980 & ~n6093;
  assign n6095 = P1_REG2_REG_3_ & n3045;
  assign n6096 = ~P1_REG2_REG_3_ & ~n3045;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = n6094 & ~n6097;
  assign n6099 = ~n5370 & ~n5371;
  assign n6100 = ~n6094 & ~n6099;
  assign n6101 = ~n6098 & ~n6100;
  assign n6102 = n5318 & ~n6101;
  assign n6103 = P1_REG3_REG_3_ & ~P1_STATE_REG;
  assign n6104 = ~n3045 & n5524;
  assign n6105 = n5526 & ~n6101;
  assign n6106 = n5528 & ~n6087;
  assign n6107 = ~n6104 & ~n6105;
  assign n6108 = ~n6106 & n6107;
  assign n6109 = n5513 & ~n6108;
  assign n6110 = ~n6102 & ~n6103;
  assign n6111 = ~n6109 & n6110;
  assign n990 = ~n6092 | ~n6111;
  assign n6113 = ~n5471 & ~n5473;
  assign n6114 = ~n5479 & n6113;
  assign n6115 = P1_REG1_REG_2_ & n2981;
  assign n6116 = ~P1_REG1_REG_2_ & ~n2981;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = ~n5478 & n6117;
  assign n6119 = ~n5477 & n6118;
  assign n6120 = ~n6114 & ~n6119;
  assign n6121 = n5417 & n6120;
  assign n6122 = ~n2981 & n5415;
  assign n6123 = P1_ADDR_REG_2_ & n5315;
  assign n6124 = ~n6121 & ~n6122;
  assign n6125 = ~n6123 & n6124;
  assign n6126 = P1_REG3_REG_2_ & ~P1_STATE_REG;
  assign n6127 = ~n5372 & ~n5374;
  assign n6128 = ~n5380 & n6127;
  assign n6129 = P1_REG2_REG_2_ & n2981;
  assign n6130 = ~P1_REG2_REG_2_ & ~n2981;
  assign n6131 = n5380 & ~n6129;
  assign n6132 = ~n6130 & n6131;
  assign n6133 = ~n6128 & ~n6132;
  assign n6134 = n5318 & n6133;
  assign n6135 = ~n2981 & n5524;
  assign n6136 = n5526 & n6133;
  assign n6137 = n5528 & n6120;
  assign n6138 = ~n6135 & ~n6136;
  assign n6139 = ~n6137 & n6138;
  assign n6140 = n5513 & ~n6139;
  assign n6141 = ~n6074 & ~n6140;
  assign n6142 = ~n6126 & ~n6134;
  assign n6143 = n6141 & n6142;
  assign n995 = ~n6125 | ~n6143;
  assign n6145 = ~n5476 & ~n5478;
  assign n6146 = ~n5475 & n6145;
  assign n6147 = n5475 & ~n6145;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = n5417 & ~n6148;
  assign n6150 = ~n2925 & n5415;
  assign n6151 = P1_ADDR_REG_1_ & n5315;
  assign n6152 = ~n6149 & ~n6150;
  assign n6153 = ~n6151 & n6152;
  assign n6154 = ~n5377 & ~n5379;
  assign n6155 = ~n5376 & n6154;
  assign n6156 = n5376 & ~n6154;
  assign n6157 = ~n6155 & ~n6156;
  assign n6158 = n5318 & ~n6157;
  assign n6159 = P1_REG3_REG_1_ & ~P1_STATE_REG;
  assign n6160 = ~n2925 & n5524;
  assign n6161 = n5526 & ~n6157;
  assign n6162 = n5528 & ~n6148;
  assign n6163 = ~n6160 & ~n6161;
  assign n6164 = ~n6162 & n6163;
  assign n6165 = n5513 & ~n6164;
  assign n6166 = ~n6158 & ~n6159;
  assign n6167 = ~n6165 & n6166;
  assign n1000 = ~n6153 | ~n6167;
  assign n6169 = P1_REG1_REG_0_ & n2859;
  assign n6170 = ~P1_REG1_REG_0_ & ~n2859;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = n5417 & ~n6171;
  assign n6173 = ~n2859 & n5415;
  assign n6174 = P1_ADDR_REG_0_ & n5315;
  assign n6175 = ~n6172 & ~n6173;
  assign n6176 = ~n6174 & n6175;
  assign n6177 = P1_REG2_REG_0_ & n2859;
  assign n6178 = ~P1_REG2_REG_0_ & ~n2859;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = n5318 & ~n6179;
  assign n6181 = P1_REG3_REG_0_ & ~P1_STATE_REG;
  assign n6182 = ~n2859 & n5524;
  assign n6183 = n5526 & ~n6179;
  assign n6184 = n5528 & ~n6171;
  assign n6185 = ~n6182 & ~n6183;
  assign n6186 = ~n6184 & n6185;
  assign n6187 = n5513 & ~n6186;
  assign n6188 = ~n6180 & ~n6181;
  assign n6189 = ~n6187 & n6188;
  assign n1005 = ~n6176 | ~n6189;
  assign n6191 = ~n2878 & n1330;
  assign n6192 = P1_DATAO_REG_0_ & ~n1330;
  assign n1010 = n6191 | n6192;
  assign n6194 = ~n2851 & n1330;
  assign n6195 = P1_DATAO_REG_1_ & ~n1330;
  assign n1015 = n6194 | n6195;
  assign n6197 = ~n2921 & n1330;
  assign n6198 = P1_DATAO_REG_2_ & ~n1330;
  assign n1020 = n6197 | n6198;
  assign n6200 = ~n2977 & n1330;
  assign n6201 = P1_DATAO_REG_3_ & ~n1330;
  assign n1025 = n6200 | n6201;
  assign n6203 = ~n3041 & n1330;
  assign n6204 = P1_DATAO_REG_4_ & ~n1330;
  assign n1030 = n6203 | n6204;
  assign n6206 = ~n3107 & n1330;
  assign n6207 = P1_DATAO_REG_5_ & ~n1330;
  assign n1035 = n6206 | n6207;
  assign n6209 = ~n3176 & n1330;
  assign n6210 = P1_DATAO_REG_6_ & ~n1330;
  assign n1040 = n6209 | n6210;
  assign n6212 = ~n3240 & n1330;
  assign n6213 = P1_DATAO_REG_7_ & ~n1330;
  assign n1045 = n6212 | n6213;
  assign n6215 = ~n3314 & n1330;
  assign n6216 = P1_DATAO_REG_8_ & ~n1330;
  assign n1050 = n6215 | n6216;
  assign n6218 = ~n3383 & n1330;
  assign n6219 = P1_DATAO_REG_9_ & ~n1330;
  assign n1055 = n6218 | n6219;
  assign n6221 = ~n3451 & n1330;
  assign n6222 = P1_DATAO_REG_10_ & ~n1330;
  assign n1060 = n6221 | n6222;
  assign n6224 = ~n3518 & n1330;
  assign n6225 = P1_DATAO_REG_11_ & ~n1330;
  assign n1065 = n6224 | n6225;
  assign n6227 = ~n3607 & n1330;
  assign n6228 = P1_DATAO_REG_12_ & ~n1330;
  assign n1070 = n6227 | n6228;
  assign n6230 = ~n3672 & n1330;
  assign n6231 = P1_DATAO_REG_13_ & ~n1330;
  assign n1075 = n6230 | n6231;
  assign n6233 = ~n3731 & n1330;
  assign n6234 = P1_DATAO_REG_14_ & ~n1330;
  assign n1080 = n6233 | n6234;
  assign n6236 = ~n3784 & n1330;
  assign n6237 = P1_DATAO_REG_15_ & ~n1330;
  assign n1085 = n6236 | n6237;
  assign n6239 = ~n3849 & n1330;
  assign n6240 = P1_DATAO_REG_16_ & ~n1330;
  assign n1090 = n6239 | n6240;
  assign n6242 = ~n3910 & n1330;
  assign n6243 = P1_DATAO_REG_17_ & ~n1330;
  assign n1095 = n6242 | n6243;
  assign n6245 = ~n3977 & n1330;
  assign n6246 = P1_DATAO_REG_18_ & ~n1330;
  assign n1100 = n6245 | n6246;
  assign n6248 = ~n4046 & n1330;
  assign n6249 = P1_DATAO_REG_19_ & ~n1330;
  assign n1105 = n6248 | n6249;
  assign n6251 = ~n4113 & n1330;
  assign n6252 = P1_DATAO_REG_20_ & ~n1330;
  assign n1110 = n6251 | n6252;
  assign n6254 = ~n4180 & n1330;
  assign n6255 = P1_DATAO_REG_21_ & ~n1330;
  assign n1115 = n6254 | n6255;
  assign n6257 = ~n4233 & n1330;
  assign n6258 = P1_DATAO_REG_22_ & ~n1330;
  assign n1120 = n6257 | n6258;
  assign n6260 = ~n4298 & n1330;
  assign n6261 = P1_DATAO_REG_23_ & ~n1330;
  assign n1125 = n6260 | n6261;
  assign n6263 = ~n4367 & n1330;
  assign n6264 = P1_DATAO_REG_24_ & ~n1330;
  assign n1130 = n6263 | n6264;
  assign n6266 = ~n4413 & n1330;
  assign n6267 = P1_DATAO_REG_25_ & ~n1330;
  assign n1135 = n6266 | n6267;
  assign n6269 = ~n4477 & n1330;
  assign n6270 = P1_DATAO_REG_26_ & ~n1330;
  assign n1140 = n6269 | n6270;
  assign n6272 = ~n4534 & n1330;
  assign n6273 = P1_DATAO_REG_27_ & ~n1330;
  assign n1145 = n6272 | n6273;
  assign n6275 = ~n4594 & n1330;
  assign n6276 = P1_DATAO_REG_28_ & ~n1330;
  assign n1150 = n6275 | n6276;
  assign n6278 = ~n4651 & n1330;
  assign n6279 = P1_DATAO_REG_29_ & ~n1330;
  assign n1155 = n6278 | n6279;
  assign n6281 = ~n4737 & n1330;
  assign n6282 = P1_DATAO_REG_30_ & ~n1330;
  assign n1160 = n6281 | n6282;
  assign n6284 = ~n4769 & n1330;
  assign n6285 = P1_DATAO_REG_31_ & ~n1330;
  assign n1165 = n6284 | n6285;
  assign n6287 = ~n2683 & ~n2752;
  assign n6288 = P1_STATE_REG & ~n6287;
  assign n6289 = ~n5310 & n6288;
  assign n6290 = ~n2752 & n2892;
  assign n6291 = n5317 & n6290;
  assign n6292 = n2683 & ~n6291;
  assign n6293 = n6289 & ~n6292;
  assign n6294 = P1_B_REG & ~n6293;
  assign n6295 = ~P1_STATE_REG & ~n6294;
  assign n6296 = n2868 & n4780;
  assign n6297 = ~n4737 & n4769;
  assign n6298 = ~n4769 & ~n6297;
  assign n6299 = n4737 & ~n4769;
  assign n6300 = ~n6297 & ~n6299;
  assign n6301 = n6297 & n6300;
  assign n6302 = ~n6298 & ~n6301;
  assign n6303 = ~n2683 & n2764;
  assign n6304 = ~n6287 & ~n6303;
  assign n6305 = ~n6302 & ~n6304;
  assign n6306 = ~n6296 & ~n6305;
  assign n6307 = n2868 & ~n6302;
  assign n6308 = n4780 & ~n6304;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = ~n6306 & n6309;
  assign n6311 = n6306 & ~n6309;
  assign n6312 = ~n6310 & ~n6311;
  assign n6313 = n2868 & n4479;
  assign n6314 = ~n2683 & ~n6313;
  assign n6315 = ~n4413 & ~n6297;
  assign n6316 = ~n4413 & n6297;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~n6304 & ~n6317;
  assign n6319 = n6314 & ~n6318;
  assign n6320 = n2683 & ~n4367;
  assign n6321 = n4479 & ~n6304;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = n2868 & ~n6317;
  assign n6324 = n6322 & ~n6323;
  assign n6325 = ~n6319 & n6324;
  assign n6326 = n2868 & n4536;
  assign n6327 = ~n2683 & ~n6326;
  assign n6328 = ~n4477 & ~n6297;
  assign n6329 = ~n4477 & n6297;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = ~n6304 & ~n6330;
  assign n6332 = n6327 & ~n6331;
  assign n6333 = n2683 & ~n4413;
  assign n6334 = n4536 & ~n6304;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = n2868 & ~n6330;
  assign n6337 = n6335 & ~n6336;
  assign n6338 = ~n6332 & n6337;
  assign n6339 = ~n6325 & ~n6338;
  assign n6340 = n6332 & ~n6337;
  assign n6341 = n2683 & ~n4477;
  assign n6342 = n4596 & ~n6304;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = ~n4534 & ~n6297;
  assign n6345 = ~n4534 & n6297;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = n2868 & ~n6346;
  assign n6348 = n6343 & ~n6347;
  assign n6349 = n2868 & n4596;
  assign n6350 = ~n2683 & ~n6349;
  assign n6351 = ~n6304 & ~n6346;
  assign n6352 = n6350 & ~n6351;
  assign n6353 = ~n6348 & n6352;
  assign n6354 = n2683 & ~n4534;
  assign n6355 = n4653 & ~n6304;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n4594 & ~n6297;
  assign n6358 = ~n4594 & n6297;
  assign n6359 = ~n6357 & ~n6358;
  assign n6360 = n2868 & ~n6359;
  assign n6361 = n6356 & ~n6360;
  assign n6362 = n2868 & n4653;
  assign n6363 = ~n2683 & ~n6362;
  assign n6364 = ~n6304 & ~n6359;
  assign n6365 = n6363 & ~n6364;
  assign n6366 = ~n6361 & n6365;
  assign n6367 = ~n4651 & ~n6297;
  assign n6368 = ~n4651 & n6297;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = n2868 & ~n6369;
  assign n6371 = n2683 & ~n4594;
  assign n6372 = n4707 & ~n6304;
  assign n6373 = ~n6370 & ~n6371;
  assign n6374 = ~n6372 & n6373;
  assign n6375 = ~n6304 & ~n6369;
  assign n6376 = n2868 & n4707;
  assign n6377 = ~n2683 & ~n6375;
  assign n6378 = ~n6376 & n6377;
  assign n6379 = ~n6374 & n6378;
  assign n6380 = ~n6339 & ~n6340;
  assign n6381 = ~n6353 & n6380;
  assign n6382 = ~n6366 & n6381;
  assign n6383 = ~n6379 & n6382;
  assign n6384 = ~n4737 & ~n6297;
  assign n6385 = n4737 & n6297;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = n2868 & ~n6386;
  assign n6388 = n4763 & ~n6304;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = n2868 & n4763;
  assign n6391 = ~n6304 & ~n6386;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = ~n6389 & n6392;
  assign n6394 = n6312 & n6383;
  assign n6395 = ~n6393 & n6394;
  assign n6396 = n2683 & ~n2868;
  assign n6397 = n6309 & n6396;
  assign n6398 = ~n6306 & n6397;
  assign n6399 = ~n6309 & ~n6396;
  assign n6400 = n6306 & n6399;
  assign n6401 = ~n6398 & ~n6400;
  assign n6402 = ~n6395 & n6401;
  assign n6403 = n2868 & n4235;
  assign n6404 = ~n2683 & ~n6403;
  assign n6405 = ~n4180 & ~n6297;
  assign n6406 = ~n4180 & n6297;
  assign n6407 = ~n6405 & ~n6406;
  assign n6408 = ~n6304 & ~n6407;
  assign n6409 = n6404 & ~n6408;
  assign n6410 = n2683 & ~n4113;
  assign n6411 = n4235 & ~n6304;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = n2868 & ~n6407;
  assign n6414 = n6412 & ~n6413;
  assign n6415 = ~n6409 & n6414;
  assign n6416 = n2868 & n4282;
  assign n6417 = ~n2683 & ~n6416;
  assign n6418 = ~n4233 & ~n6297;
  assign n6419 = ~n4233 & n6297;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = ~n6304 & ~n6420;
  assign n6422 = n6417 & ~n6421;
  assign n6423 = n2683 & ~n4180;
  assign n6424 = n4282 & ~n6304;
  assign n6425 = ~n6423 & ~n6424;
  assign n6426 = n2868 & ~n6420;
  assign n6427 = n6425 & ~n6426;
  assign n6428 = ~n6422 & n6427;
  assign n6429 = ~n6415 & ~n6428;
  assign n6430 = n2868 & n4164;
  assign n6431 = ~n2683 & ~n6430;
  assign n6432 = ~n4113 & ~n6297;
  assign n6433 = ~n4113 & n6297;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = ~n6304 & ~n6434;
  assign n6436 = n6431 & ~n6435;
  assign n6437 = n2683 & ~n4046;
  assign n6438 = n4164 & ~n6304;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = n2868 & ~n6434;
  assign n6441 = n6439 & ~n6440;
  assign n6442 = ~n6436 & n6441;
  assign n6443 = n2868 & ~n4117;
  assign n6444 = ~n2683 & ~n6443;
  assign n6445 = ~n4046 & ~n6297;
  assign n6446 = ~n4046 & n6297;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = ~n6304 & ~n6447;
  assign n6449 = n6444 & ~n6448;
  assign n6450 = n2683 & ~n3977;
  assign n6451 = ~n4117 & ~n6304;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = n2868 & ~n6447;
  assign n6454 = n6452 & ~n6453;
  assign n6455 = ~n6449 & n6454;
  assign n6456 = n2868 & ~n3798;
  assign n6457 = ~n2683 & ~n6456;
  assign n6458 = ~n3731 & ~n6297;
  assign n6459 = ~n3731 & n6297;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = ~n6304 & ~n6460;
  assign n6462 = n6457 & ~n6461;
  assign n6463 = n2683 & ~n3672;
  assign n6464 = ~n3798 & ~n6304;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = n2868 & ~n6460;
  assign n6467 = n6465 & ~n6466;
  assign n6468 = ~n6462 & n6467;
  assign n6469 = ~n3672 & ~n6297;
  assign n6470 = ~n3672 & n6297;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n6304 & ~n6471;
  assign n6473 = n2868 & ~n3715;
  assign n6474 = ~n2683 & ~n6472;
  assign n6475 = ~n6473 & n6474;
  assign n6476 = n2868 & ~n6471;
  assign n6477 = n2683 & ~n3607;
  assign n6478 = ~n3715 & ~n6304;
  assign n6479 = ~n6476 & ~n6477;
  assign n6480 = ~n6478 & n6479;
  assign n6481 = ~n6475 & n6480;
  assign n6482 = ~n3383 & ~n6297;
  assign n6483 = ~n3383 & n6297;
  assign n6484 = ~n6482 & ~n6483;
  assign n6485 = n2868 & ~n6484;
  assign n6486 = n2683 & ~n3314;
  assign n6487 = ~n3458 & ~n6304;
  assign n6488 = ~n6485 & ~n6486;
  assign n6489 = ~n6487 & n6488;
  assign n6490 = ~n6304 & ~n6484;
  assign n6491 = n2868 & ~n3458;
  assign n6492 = ~n2683 & ~n6490;
  assign n6493 = ~n6491 & n6492;
  assign n6494 = ~n6489 & n6493;
  assign n6495 = ~n3314 & ~n6297;
  assign n6496 = ~n3314 & n6297;
  assign n6497 = ~n6495 & ~n6496;
  assign n6498 = n2868 & ~n6497;
  assign n6499 = n2683 & ~n3240;
  assign n6500 = ~n3390 & ~n6304;
  assign n6501 = ~n6498 & ~n6499;
  assign n6502 = ~n6500 & n6501;
  assign n6503 = ~n6304 & ~n6497;
  assign n6504 = n2868 & ~n3390;
  assign n6505 = ~n2683 & ~n6503;
  assign n6506 = ~n6504 & n6505;
  assign n6507 = ~n6502 & n6506;
  assign n6508 = ~n6494 & ~n6507;
  assign n6509 = ~n3240 & ~n6297;
  assign n6510 = ~n3240 & n6297;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = n2868 & ~n6511;
  assign n6513 = n2683 & ~n3176;
  assign n6514 = ~n3321 & ~n6304;
  assign n6515 = ~n6512 & ~n6513;
  assign n6516 = ~n6514 & n6515;
  assign n6517 = ~n6304 & ~n6511;
  assign n6518 = n2868 & ~n3321;
  assign n6519 = ~n2683 & ~n6517;
  assign n6520 = ~n6518 & n6519;
  assign n6521 = ~n6516 & n6520;
  assign n6522 = ~n3176 & ~n6297;
  assign n6523 = ~n3176 & n6297;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = n2868 & ~n6524;
  assign n6526 = n2683 & ~n3107;
  assign n6527 = ~n3247 & ~n6304;
  assign n6528 = ~n6525 & ~n6526;
  assign n6529 = ~n6527 & n6528;
  assign n6530 = ~n6304 & ~n6524;
  assign n6531 = n2868 & ~n3247;
  assign n6532 = ~n2683 & ~n6530;
  assign n6533 = ~n6531 & n6532;
  assign n6534 = ~n6529 & n6533;
  assign n6535 = ~n6521 & ~n6534;
  assign n6536 = n6508 & n6535;
  assign n6537 = ~n3041 & ~n6297;
  assign n6538 = ~n3041 & n6297;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = ~n6304 & ~n6539;
  assign n6541 = n2868 & ~n3114;
  assign n6542 = ~n2683 & ~n6540;
  assign n6543 = ~n6541 & n6542;
  assign n6544 = n2868 & ~n6539;
  assign n6545 = n2683 & ~n2977;
  assign n6546 = ~n3114 & ~n6304;
  assign n6547 = ~n6544 & ~n6545;
  assign n6548 = ~n6546 & n6547;
  assign n6549 = ~n6543 & n6548;
  assign n6550 = ~n2977 & ~n6297;
  assign n6551 = ~n2977 & n6297;
  assign n6552 = ~n6550 & ~n6551;
  assign n6553 = ~n6304 & ~n6552;
  assign n6554 = n2868 & ~n3048;
  assign n6555 = ~n2683 & ~n6553;
  assign n6556 = ~n6554 & n6555;
  assign n6557 = n2868 & ~n6552;
  assign n6558 = n2683 & ~n2921;
  assign n6559 = ~n3048 & ~n6304;
  assign n6560 = ~n6557 & ~n6558;
  assign n6561 = ~n6559 & n6560;
  assign n6562 = ~n6556 & n6561;
  assign n6563 = ~n2921 & ~n6297;
  assign n6564 = ~n2921 & n6297;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = ~n6304 & ~n6565;
  assign n6567 = n2868 & ~n2984;
  assign n6568 = ~n2683 & ~n6566;
  assign n6569 = ~n6567 & n6568;
  assign n6570 = n2868 & ~n6565;
  assign n6571 = n2683 & ~n2851;
  assign n6572 = ~n2984 & ~n6304;
  assign n6573 = ~n6570 & ~n6571;
  assign n6574 = ~n6572 & n6573;
  assign n6575 = ~n6569 & n6574;
  assign n6576 = ~n2851 & ~n6297;
  assign n6577 = ~n2851 & n6297;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = ~n6304 & ~n6578;
  assign n6580 = n2868 & ~n2928;
  assign n6581 = ~n2683 & ~n6579;
  assign n6582 = ~n6580 & n6581;
  assign n6583 = n2868 & ~n6578;
  assign n6584 = n2683 & ~n2878;
  assign n6585 = ~n2928 & ~n6304;
  assign n6586 = ~n6583 & ~n6584;
  assign n6587 = ~n6585 & n6586;
  assign n6588 = ~n6582 & n6587;
  assign n6589 = n6569 & ~n6574;
  assign n6590 = n6588 & ~n6589;
  assign n6591 = ~n6575 & ~n6590;
  assign n6592 = n6556 & ~n6561;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = ~n6562 & ~n6593;
  assign n6595 = n6543 & ~n6548;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = ~n6549 & ~n6596;
  assign n6598 = ~n3107 & ~n6297;
  assign n6599 = ~n3107 & n6297;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = n2868 & ~n6600;
  assign n6602 = n2683 & ~n3041;
  assign n6603 = ~n3183 & ~n6304;
  assign n6604 = ~n6601 & ~n6602;
  assign n6605 = ~n6603 & n6604;
  assign n6606 = ~n6304 & ~n6600;
  assign n6607 = n2868 & ~n3183;
  assign n6608 = ~n2683 & ~n6606;
  assign n6609 = ~n6607 & n6608;
  assign n6610 = ~n6605 & n6609;
  assign n6611 = ~n6597 & ~n6610;
  assign n6612 = n6529 & ~n6533;
  assign n6613 = n6605 & ~n6609;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n2862 & n2868;
  assign n6616 = ~n2683 & ~n6615;
  assign n6617 = ~n2878 & ~n6297;
  assign n6618 = ~n2878 & n6297;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = ~n6304 & ~n6619;
  assign n6621 = n6616 & ~n6620;
  assign n6622 = ~n2683 & n2868;
  assign n6623 = n6621 & n6622;
  assign n6624 = n6582 & ~n6587;
  assign n6625 = n2868 & ~n6619;
  assign n6626 = ~n2862 & ~n6304;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = ~n6621 & ~n6622;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = ~n6623 & ~n6624;
  assign n6631 = ~n6629 & n6630;
  assign n6632 = ~n6589 & ~n6592;
  assign n6633 = ~n6610 & n6632;
  assign n6634 = ~n6595 & n6633;
  assign n6635 = n6631 & n6634;
  assign n6636 = n6614 & ~n6635;
  assign n6637 = ~n6611 & n6636;
  assign n6638 = n6536 & ~n6637;
  assign n6639 = n6516 & ~n6520;
  assign n6640 = n6508 & n6639;
  assign n6641 = n6502 & ~n6506;
  assign n6642 = ~n6494 & n6641;
  assign n6643 = ~n3451 & ~n6297;
  assign n6644 = ~n3451 & n6297;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = ~n6304 & ~n6645;
  assign n6647 = n2868 & ~n3525;
  assign n6648 = ~n2683 & ~n6646;
  assign n6649 = ~n6647 & n6648;
  assign n6650 = n2868 & ~n6645;
  assign n6651 = n2683 & ~n3383;
  assign n6652 = ~n3525 & ~n6304;
  assign n6653 = ~n6650 & ~n6651;
  assign n6654 = ~n6652 & n6653;
  assign n6655 = ~n6649 & n6654;
  assign n6656 = n6489 & ~n6493;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n3607 & ~n6297;
  assign n6659 = ~n3607 & n6297;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = ~n6304 & ~n6660;
  assign n6662 = n2868 & ~n3648;
  assign n6663 = ~n2683 & ~n6661;
  assign n6664 = ~n6662 & n6663;
  assign n6665 = n2868 & ~n6660;
  assign n6666 = n2683 & ~n3518;
  assign n6667 = ~n3648 & ~n6304;
  assign n6668 = ~n6665 & ~n6666;
  assign n6669 = ~n6667 & n6668;
  assign n6670 = ~n6664 & n6669;
  assign n6671 = ~n3518 & ~n6297;
  assign n6672 = ~n3518 & n6297;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = ~n6304 & ~n6673;
  assign n6675 = n2868 & ~n3578;
  assign n6676 = ~n2683 & ~n6674;
  assign n6677 = ~n6675 & n6676;
  assign n6678 = n2868 & ~n6673;
  assign n6679 = n2683 & ~n3451;
  assign n6680 = ~n3578 & ~n6304;
  assign n6681 = ~n6678 & ~n6679;
  assign n6682 = ~n6680 & n6681;
  assign n6683 = ~n6677 & n6682;
  assign n6684 = ~n6670 & ~n6683;
  assign n6685 = n6657 & n6684;
  assign n6686 = ~n6640 & ~n6642;
  assign n6687 = n6685 & n6686;
  assign n6688 = ~n6638 & n6687;
  assign n6689 = n6649 & ~n6654;
  assign n6690 = n6684 & n6689;
  assign n6691 = n6664 & ~n6669;
  assign n6692 = n6475 & ~n6480;
  assign n6693 = n6677 & ~n6682;
  assign n6694 = ~n6670 & n6693;
  assign n6695 = ~n6692 & ~n6694;
  assign n6696 = ~n6690 & ~n6691;
  assign n6697 = n6695 & n6696;
  assign n6698 = ~n6688 & n6697;
  assign n6699 = ~n6481 & ~n6698;
  assign n6700 = n6462 & ~n6467;
  assign n6701 = ~n6699 & ~n6700;
  assign n6702 = ~n6468 & ~n6701;
  assign n6703 = n2683 & ~n3731;
  assign n6704 = ~n3860 & ~n6304;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = ~n3784 & ~n6297;
  assign n6707 = ~n3784 & n6297;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = n2868 & ~n6708;
  assign n6710 = n6705 & ~n6709;
  assign n6711 = n2868 & ~n3860;
  assign n6712 = ~n2683 & ~n6711;
  assign n6713 = ~n6304 & ~n6708;
  assign n6714 = n6712 & ~n6713;
  assign n6715 = ~n6710 & n6714;
  assign n6716 = ~n6702 & ~n6715;
  assign n6717 = n2868 & ~n4059;
  assign n6718 = ~n2683 & ~n6717;
  assign n6719 = ~n3977 & ~n6297;
  assign n6720 = ~n3977 & n6297;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n6304 & ~n6721;
  assign n6723 = n6718 & ~n6722;
  assign n6724 = n2683 & ~n3910;
  assign n6725 = ~n4059 & ~n6304;
  assign n6726 = ~n6724 & ~n6725;
  assign n6727 = n2868 & ~n6721;
  assign n6728 = n6726 & ~n6727;
  assign n6729 = ~n6723 & n6728;
  assign n6730 = n2868 & ~n3984;
  assign n6731 = ~n2683 & ~n6730;
  assign n6732 = ~n3910 & ~n6297;
  assign n6733 = ~n3910 & n6297;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = ~n6304 & ~n6734;
  assign n6736 = n6731 & ~n6735;
  assign n6737 = n2683 & ~n3849;
  assign n6738 = ~n3984 & ~n6304;
  assign n6739 = ~n6737 & ~n6738;
  assign n6740 = n2868 & ~n6734;
  assign n6741 = n6739 & ~n6740;
  assign n6742 = ~n6736 & n6741;
  assign n6743 = ~n6729 & ~n6742;
  assign n6744 = n6710 & ~n6714;
  assign n6745 = n2868 & ~n3917;
  assign n6746 = ~n2683 & ~n6745;
  assign n6747 = ~n3849 & ~n6297;
  assign n6748 = ~n3849 & n6297;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = ~n6304 & ~n6749;
  assign n6751 = n6746 & ~n6750;
  assign n6752 = n2683 & ~n3784;
  assign n6753 = ~n3917 & ~n6304;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = n2868 & ~n6749;
  assign n6756 = n6754 & ~n6755;
  assign n6757 = ~n6751 & n6756;
  assign n6758 = ~n6744 & ~n6757;
  assign n6759 = n6743 & n6758;
  assign n6760 = ~n6716 & n6759;
  assign n6761 = n6751 & ~n6756;
  assign n6762 = n6743 & n6761;
  assign n6763 = n6736 & ~n6741;
  assign n6764 = ~n6729 & n6763;
  assign n6765 = n6449 & ~n6454;
  assign n6766 = n6723 & ~n6728;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n6762 & ~n6764;
  assign n6769 = n6767 & n6768;
  assign n6770 = ~n6760 & n6769;
  assign n6771 = ~n6455 & ~n6770;
  assign n6772 = n6436 & ~n6441;
  assign n6773 = ~n6771 & ~n6772;
  assign n6774 = ~n6442 & ~n6773;
  assign n6775 = n6409 & ~n6414;
  assign n6776 = ~n6774 & ~n6775;
  assign n6777 = n2868 & n4415;
  assign n6778 = ~n2683 & ~n6777;
  assign n6779 = ~n4367 & ~n6297;
  assign n6780 = ~n4367 & n6297;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = ~n6304 & ~n6781;
  assign n6783 = n6778 & ~n6782;
  assign n6784 = n2683 & ~n4298;
  assign n6785 = n4415 & ~n6304;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = n2868 & ~n6781;
  assign n6788 = n6786 & ~n6787;
  assign n6789 = ~n6783 & n6788;
  assign n6790 = n2868 & n4344;
  assign n6791 = ~n2683 & ~n6790;
  assign n6792 = ~n4298 & ~n6297;
  assign n6793 = ~n4298 & n6297;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = ~n6304 & ~n6794;
  assign n6796 = n6791 & ~n6795;
  assign n6797 = n2683 & ~n4233;
  assign n6798 = n4344 & ~n6304;
  assign n6799 = ~n6797 & ~n6798;
  assign n6800 = n2868 & ~n6794;
  assign n6801 = n6799 & ~n6800;
  assign n6802 = ~n6796 & n6801;
  assign n6803 = ~n6789 & ~n6802;
  assign n6804 = n6429 & ~n6776;
  assign n6805 = n6803 & n6804;
  assign n6806 = n6422 & ~n6427;
  assign n6807 = n6803 & n6806;
  assign n6808 = n6796 & ~n6801;
  assign n6809 = ~n6789 & n6808;
  assign n6810 = n6783 & ~n6788;
  assign n6811 = n6319 & ~n6324;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6807 & ~n6809;
  assign n6814 = n6812 & n6813;
  assign n6815 = ~n6340 & ~n6805;
  assign n6816 = ~n6353 & n6815;
  assign n6817 = n6814 & n6816;
  assign n6818 = ~n6366 & n6817;
  assign n6819 = ~n6379 & n6818;
  assign n6820 = n6312 & n6819;
  assign n6821 = ~n6393 & n6820;
  assign n6822 = n6312 & n6389;
  assign n6823 = ~n6392 & n6822;
  assign n6824 = n6374 & ~n6378;
  assign n6825 = n6312 & n6824;
  assign n6826 = ~n6393 & n6825;
  assign n6827 = n6361 & ~n6365;
  assign n6828 = n6348 & ~n6352;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = ~n6366 & ~n6379;
  assign n6831 = n6312 & ~n6829;
  assign n6832 = n6830 & n6831;
  assign n6833 = ~n6393 & n6832;
  assign n6834 = ~n6823 & ~n6826;
  assign n6835 = ~n6833 & n6834;
  assign n6836 = n6402 & ~n6821;
  assign n6837 = n6835 & n6836;
  assign n6838 = n2696 & n6291;
  assign n6839 = n6837 & n6838;
  assign n6840 = n4769 & n4780;
  assign n6841 = n4607 & ~n4670;
  assign n6842 = ~n6840 & n6841;
  assign n6843 = ~n4189 & ~n4237;
  assign n6844 = n2998 & ~n3059;
  assign n6845 = ~n3058 & ~n6844;
  assign n6846 = ~n3121 & ~n6845;
  assign n6847 = ~n3195 & n3347;
  assign n6848 = ~n6846 & n6847;
  assign n6849 = n3196 & ~n3254;
  assign n6850 = ~n3255 & ~n3334;
  assign n6851 = ~n3403 & n6850;
  assign n6852 = ~n3465 & n6851;
  assign n6853 = ~n6848 & ~n6849;
  assign n6854 = n6852 & n6853;
  assign n6855 = n3333 & ~n3403;
  assign n6856 = ~n3402 & ~n6855;
  assign n6857 = ~n3465 & ~n6856;
  assign n6858 = ~n3464 & ~n3538;
  assign n6859 = ~n3587 & ~n3650;
  assign n6860 = n6858 & n6859;
  assign n6861 = ~n3059 & ~n3121;
  assign n6862 = ~n6849 & n6861;
  assign n6863 = n2758 & ~n2879;
  assign n6864 = ~n2880 & ~n6863;
  assign n6865 = ~n2928 & n6864;
  assign n6866 = ~n2851 & ~n6865;
  assign n6867 = n2928 & ~n6864;
  assign n6868 = ~n2999 & ~n6867;
  assign n6869 = n6852 & n6868;
  assign n6870 = n6862 & ~n6866;
  assign n6871 = n6869 & n6870;
  assign n6872 = ~n6854 & ~n6857;
  assign n6873 = n6860 & n6872;
  assign n6874 = ~n6871 & n6873;
  assign n6875 = n3539 & n6859;
  assign n6876 = n3588 & ~n3650;
  assign n6877 = ~n3740 & ~n6876;
  assign n6878 = ~n3651 & ~n6875;
  assign n6879 = n6877 & n6878;
  assign n6880 = ~n6874 & n6879;
  assign n6881 = ~n3739 & ~n6880;
  assign n6882 = ~n3800 & ~n6881;
  assign n6883 = ~n3799 & ~n6882;
  assign n6884 = ~n3862 & ~n6883;
  assign n6885 = ~n3991 & ~n4060;
  assign n6886 = ~n3861 & ~n3918;
  assign n6887 = n6885 & n6886;
  assign n6888 = ~n6884 & n6887;
  assign n6889 = n3919 & n6885;
  assign n6890 = n3992 & ~n4060;
  assign n6891 = ~n4061 & ~n4119;
  assign n6892 = ~n6889 & ~n6890;
  assign n6893 = n6891 & n6892;
  assign n6894 = ~n6888 & n6893;
  assign n6895 = ~n4118 & ~n6894;
  assign n6896 = n6843 & ~n6895;
  assign n6897 = ~n4737 & ~n4763;
  assign n6898 = n4718 & ~n6897;
  assign n6899 = n4737 & ~n6840;
  assign n6900 = n4763 & n6899;
  assign n6901 = n4620 & ~n4670;
  assign n6902 = n4485 & n6901;
  assign n6903 = ~n6840 & n6902;
  assign n6904 = ~n6900 & ~n6903;
  assign n6905 = n4188 & ~n4237;
  assign n6906 = ~n4350 & ~n4425;
  assign n6907 = ~n4236 & ~n6905;
  assign n6908 = ~n4310 & n6907;
  assign n6909 = n6906 & n6908;
  assign n6910 = ~n4769 & ~n4780;
  assign n6911 = n4669 & ~n6840;
  assign n6912 = n4550 & n6901;
  assign n6913 = ~n6840 & n6912;
  assign n6914 = n6909 & ~n6910;
  assign n6915 = ~n6911 & n6914;
  assign n6916 = ~n6913 & n6915;
  assign n6917 = ~n6842 & ~n6896;
  assign n6918 = ~n6898 & n6917;
  assign n6919 = n6904 & n6918;
  assign n6920 = n6916 & n6919;
  assign n6921 = ~n6898 & ~n6910;
  assign n6922 = ~n6900 & n6921;
  assign n6923 = n4311 & n6906;
  assign n6924 = n4351 & ~n4425;
  assign n6925 = ~n4486 & ~n6924;
  assign n6926 = ~n4426 & ~n6923;
  assign n6927 = n6925 & n6926;
  assign n6928 = n6901 & n6927;
  assign n6929 = ~n6842 & ~n6911;
  assign n6930 = ~n6913 & ~n6928;
  assign n6931 = n6929 & n6930;
  assign n6932 = ~n6903 & n6931;
  assign n6933 = ~n4719 & n4737;
  assign n6934 = ~n4719 & n4763;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = ~n6932 & ~n6935;
  assign n6937 = n6922 & ~n6936;
  assign n6938 = ~n6840 & ~n6920;
  assign n6939 = ~n6937 & n6938;
  assign n6940 = n2755 & n6303;
  assign n6941 = n6939 & n6940;
  assign n6942 = ~n2683 & n2903;
  assign n6943 = ~n6939 & n6942;
  assign n6944 = ~n6941 & ~n6943;
  assign n6945 = n2755 & n6944;
  assign n6946 = ~n6294 & ~n6839;
  assign n6947 = n6945 & n6946;
  assign n6948 = ~n6295 & ~n6947;
  assign n6949 = ~n3189 & ~n3190;
  assign n6950 = ~n2994 & ~n3064;
  assign n6951 = ~n6949 & n6950;
  assign n6952 = ~n3327 & ~n3328;
  assign n6953 = ~n3270 & ~n6952;
  assign n6954 = ~n3658 & n6953;
  assign n6955 = n6951 & n6954;
  assign n6956 = ~n3928 & n6955;
  assign n6957 = n2862 & n2878;
  assign n6958 = ~n2937 & ~n6957;
  assign n6959 = ~n3851 & ~n3852;
  assign n6960 = ~n2936 & ~n6958;
  assign n6961 = ~n6959 & n6960;
  assign n6962 = ~n3733 & ~n3734;
  assign n6963 = ~n3408 & ~n3472;
  assign n6964 = ~n6962 & n6963;
  assign n6965 = ~n3921 & ~n3922;
  assign n6966 = n6961 & n6964;
  assign n6967 = ~n6965 & n6966;
  assign n6968 = ~n3985 & ~n3986;
  assign n6969 = ~n3532 & ~n3533;
  assign n6970 = ~n4182 & ~n4184;
  assign n6971 = ~n3593 & ~n6969;
  assign n6972 = ~n3131 & n6971;
  assign n6973 = ~n4126 & n6972;
  assign n6974 = ~n6970 & n6973;
  assign n6975 = n6956 & n6967;
  assign n6976 = ~n6968 & n6975;
  assign n6977 = ~n4066 & n6976;
  assign n6978 = n6974 & n6977;
  assign n6979 = n4769 & ~n4780;
  assign n6980 = ~n4769 & n4780;
  assign n6981 = ~n6979 & ~n6980;
  assign n6982 = n4737 & ~n4763;
  assign n6983 = ~n4737 & n4763;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = n4477 & ~n4536;
  assign n6986 = ~n4543 & ~n6985;
  assign n6987 = ~n4493 & ~n6986;
  assign n6988 = ~n4346 & ~n4347;
  assign n6989 = ~n4300 & ~n4304;
  assign n6990 = ~n4421 & ~n4422;
  assign n6991 = ~n6988 & ~n6989;
  assign n6992 = ~n6990 & n6991;
  assign n6993 = ~n4431 & n6992;
  assign n6994 = ~n4659 & ~n4665;
  assign n6995 = n4594 & ~n4653;
  assign n6996 = ~n4715 & ~n6995;
  assign n6997 = n4651 & ~n4707;
  assign n6998 = ~n4651 & n4707;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = n6987 & n6993;
  assign n7001 = ~n6994 & n7000;
  assign n7002 = ~n6996 & n7001;
  assign n7003 = ~n6999 & n7002;
  assign n7004 = ~n6984 & n7003;
  assign n7005 = n6978 & ~n6981;
  assign n7006 = n7004 & n7005;
  assign n7007 = ~n6303 & n7006;
  assign n7008 = ~n2683 & ~n2764;
  assign n7009 = ~n7006 & ~n7008;
  assign n7010 = ~n7007 & ~n7009;
  assign n7011 = n2758 & n7010;
  assign n7012 = n2896 & n6287;
  assign n7013 = ~n6837 & n7012;
  assign n7014 = n2752 & ~n2758;
  assign n7015 = ~n2683 & n7014;
  assign n7016 = n6837 & n7015;
  assign n7017 = ~n7013 & ~n7016;
  assign n7018 = n4763 & n6386;
  assign n7019 = ~n4707 & ~n6369;
  assign n7020 = ~n4780 & ~n6302;
  assign n7021 = n7019 & ~n7020;
  assign n7022 = ~n6386 & ~n7020;
  assign n7023 = ~n4763 & n7022;
  assign n7024 = ~n7021 & ~n7023;
  assign n7025 = n4596 & n6346;
  assign n7026 = ~n4536 & ~n6330;
  assign n7027 = n4536 & n6330;
  assign n7028 = n4479 & n6317;
  assign n7029 = ~n7027 & ~n7028;
  assign n7030 = ~n4344 & ~n6794;
  assign n7031 = n4415 & n6781;
  assign n7032 = n7030 & ~n7031;
  assign n7033 = n4282 & n6420;
  assign n7034 = n4344 & n6794;
  assign n7035 = ~n7033 & ~n7034;
  assign n7036 = ~n3860 & n6708;
  assign n7037 = ~n3798 & n6460;
  assign n7038 = ~n3458 & n6484;
  assign n7039 = ~n3390 & n6497;
  assign n7040 = n3321 & ~n6511;
  assign n7041 = n3247 & ~n6524;
  assign n7042 = ~n3321 & n6511;
  assign n7043 = n7041 & ~n7042;
  assign n7044 = n3390 & ~n6497;
  assign n7045 = ~n7040 & ~n7043;
  assign n7046 = ~n7044 & n7045;
  assign n7047 = ~n3183 & n6600;
  assign n7048 = ~n3114 & n6539;
  assign n7049 = ~n3048 & n6552;
  assign n7050 = n3114 & ~n6539;
  assign n7051 = n7049 & ~n7050;
  assign n7052 = ~n3247 & n6524;
  assign n7053 = ~n7042 & ~n7052;
  assign n7054 = ~n7048 & ~n7051;
  assign n7055 = n7053 & n7054;
  assign n7056 = n3183 & ~n6600;
  assign n7057 = n7053 & n7056;
  assign n7058 = ~n7055 & ~n7057;
  assign n7059 = ~n7047 & ~n7058;
  assign n7060 = n7046 & ~n7059;
  assign n7061 = ~n7039 & ~n7060;
  assign n7062 = n3458 & ~n6484;
  assign n7063 = ~n7061 & ~n7062;
  assign n7064 = ~n7038 & ~n7063;
  assign n7065 = n3525 & ~n6645;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = ~n2984 & n6565;
  assign n7068 = ~n7062 & ~n7065;
  assign n7069 = n3048 & ~n6552;
  assign n7070 = ~n7050 & ~n7069;
  assign n7071 = ~n7040 & n7070;
  assign n7072 = ~n7044 & n7071;
  assign n7073 = ~n7043 & ~n7057;
  assign n7074 = n7068 & n7073;
  assign n7075 = n7072 & n7074;
  assign n7076 = n7067 & n7075;
  assign n7077 = ~n2862 & n6619;
  assign n7078 = n2928 & ~n7077;
  assign n7079 = n2984 & ~n6565;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = ~n2928 & n7077;
  assign n7082 = ~n6578 & ~n7081;
  assign n7083 = n7080 & ~n7082;
  assign n7084 = n7075 & n7083;
  assign n7085 = ~n3578 & n6673;
  assign n7086 = ~n3525 & n6645;
  assign n7087 = ~n7085 & ~n7086;
  assign n7088 = ~n3715 & n6471;
  assign n7089 = ~n3648 & n6660;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = n7087 & n7090;
  assign n7092 = ~n7076 & ~n7084;
  assign n7093 = n7091 & n7092;
  assign n7094 = ~n7066 & n7093;
  assign n7095 = n3648 & ~n6660;
  assign n7096 = ~n7088 & n7095;
  assign n7097 = n3715 & ~n6471;
  assign n7098 = n3798 & ~n6460;
  assign n7099 = ~n7097 & ~n7098;
  assign n7100 = ~n7096 & n7099;
  assign n7101 = n3578 & ~n6673;
  assign n7102 = n7090 & n7101;
  assign n7103 = n7100 & ~n7102;
  assign n7104 = ~n7094 & n7103;
  assign n7105 = ~n7037 & ~n7104;
  assign n7106 = n3860 & ~n6708;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = ~n7036 & ~n7107;
  assign n7109 = n3917 & ~n6749;
  assign n7110 = n4117 & ~n6447;
  assign n7111 = n4059 & ~n6721;
  assign n7112 = ~n4117 & n6447;
  assign n7113 = n7111 & ~n7112;
  assign n7114 = ~n7110 & ~n7113;
  assign n7115 = n3984 & ~n6734;
  assign n7116 = ~n4059 & n6721;
  assign n7117 = ~n7112 & ~n7116;
  assign n7118 = n7115 & n7117;
  assign n7119 = ~n4164 & ~n6434;
  assign n7120 = ~n4282 & ~n6420;
  assign n7121 = ~n4235 & ~n6407;
  assign n7122 = ~n7120 & ~n7121;
  assign n7123 = n7114 & ~n7118;
  assign n7124 = ~n7119 & n7123;
  assign n7125 = n7122 & n7124;
  assign n7126 = ~n7108 & ~n7109;
  assign n7127 = n7125 & n7126;
  assign n7128 = ~n3917 & n6749;
  assign n7129 = ~n3984 & n6734;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = n7117 & n7130;
  assign n7132 = n7125 & ~n7131;
  assign n7133 = n4164 & n6434;
  assign n7134 = n7122 & n7133;
  assign n7135 = ~n7132 & ~n7134;
  assign n7136 = n4235 & n6407;
  assign n7137 = ~n7120 & n7136;
  assign n7138 = ~n7031 & ~n7137;
  assign n7139 = n7035 & ~n7127;
  assign n7140 = n7135 & n7139;
  assign n7141 = n7138 & n7140;
  assign n7142 = ~n4479 & ~n6317;
  assign n7143 = ~n4415 & ~n6781;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = ~n7032 & ~n7141;
  assign n7146 = n7144 & n7145;
  assign n7147 = n7029 & ~n7146;
  assign n7148 = ~n4596 & ~n6346;
  assign n7149 = ~n7026 & ~n7147;
  assign n7150 = ~n7148 & n7149;
  assign n7151 = ~n7025 & ~n7150;
  assign n7152 = ~n4653 & n7151;
  assign n7153 = n6359 & ~n7152;
  assign n7154 = n4707 & n6369;
  assign n7155 = n4653 & ~n7151;
  assign n7156 = ~n7154 & ~n7155;
  assign n7157 = ~n7020 & ~n7153;
  assign n7158 = n7156 & n7157;
  assign n7159 = n7024 & ~n7158;
  assign n7160 = ~n7018 & ~n7159;
  assign n7161 = n4780 & n6302;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = n2830 & n6303;
  assign n7164 = n7162 & n7163;
  assign n7165 = n6946 & ~n7164;
  assign n7166 = ~n7011 & n7017;
  assign n7167 = n6944 & n7166;
  assign n7168 = n7165 & n7167;
  assign n1170 = n6948 & ~n7168;
  assign n7170 = n2696 & ~n4900;
  assign n7171 = ~n2745 & ~n2749;
  assign n7172 = n2827 & n7171;
  assign n7173 = n7170 & ~n7172;
  assign n7174 = n2683 & ~n4891;
  assign n7175 = ~n5310 & n7174;
  assign n7176 = ~n2898 & ~n2904;
  assign n7177 = ~n2901 & n7176;
  assign n7178 = n2758 & ~n7177;
  assign n7179 = ~n2890 & ~n4912;
  assign n7180 = ~n2896 & n7179;
  assign n7181 = n2752 & ~n7180;
  assign n7182 = ~n2888 & ~n2893;
  assign n7183 = ~n4889 & n7182;
  assign n7184 = ~n7178 & ~n7181;
  assign n7185 = n7183 & n7184;
  assign n7186 = ~n7172 & ~n7185;
  assign n7187 = n7175 & ~n7186;
  assign n7188 = P1_STATE_REG & ~n7187;
  assign n7189 = ~n7173 & ~n7188;
  assign n7190 = ~n3780 & ~n7189;
  assign n7191 = n7170 & n7172;
  assign n7192 = n2696 & n4890;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 = ~n3860 & ~n7193;
  assign n7195 = n2696 & n6290;
  assign n7196 = ~n3780 & ~n7172;
  assign n7197 = ~n2833 & n7172;
  assign n7198 = ~n3731 & n7197;
  assign n7199 = n2833 & n7172;
  assign n7200 = ~n3849 & n7199;
  assign n7201 = ~n7196 & ~n7198;
  assign n7202 = ~n7200 & n7201;
  assign n7203 = n7195 & ~n7202;
  assign n7204 = ~n3731 & ~n6048;
  assign n7205 = ~n3798 & n6051;
  assign n7206 = ~n7204 & ~n7205;
  assign n7207 = ~n3731 & n6051;
  assign n7208 = ~n3798 & ~n6061;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = ~n6043 & ~n7209;
  assign n7211 = n6043 & n7209;
  assign n7212 = ~n7210 & ~n7211;
  assign n7213 = ~n7206 & ~n7212;
  assign n7214 = n7206 & n7212;
  assign n7215 = ~n3672 & n6051;
  assign n7216 = ~n3715 & ~n6061;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = ~n6043 & ~n7217;
  assign n7219 = n6043 & n7217;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = ~n3672 & ~n6048;
  assign n7222 = ~n3715 & n6051;
  assign n7223 = ~n7221 & ~n7222;
  assign n7224 = n7220 & n7223;
  assign n7225 = ~n7220 & ~n7223;
  assign n7226 = ~n3607 & ~n6048;
  assign n7227 = ~n3648 & n6051;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = ~n3607 & n6051;
  assign n7230 = ~n3648 & ~n6061;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = ~n6043 & ~n7231;
  assign n7233 = n6043 & n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = ~n7228 & ~n7234;
  assign n7236 = ~n7225 & ~n7235;
  assign n7237 = ~n3518 & ~n6048;
  assign n7238 = ~n3578 & n6051;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = ~n3518 & n6051;
  assign n7241 = ~n3578 & ~n6061;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = ~n6043 & ~n7242;
  assign n7244 = n6043 & n7242;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n7239 & ~n7245;
  assign n7247 = n7228 & n7234;
  assign n7248 = ~n7224 & ~n7247;
  assign n7249 = n7246 & n7248;
  assign n7250 = n7236 & ~n7249;
  assign n7251 = ~n7224 & ~n7250;
  assign n7252 = n7239 & n7245;
  assign n7253 = n7248 & ~n7252;
  assign n7254 = ~n3451 & ~n6048;
  assign n7255 = ~n3525 & n6051;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = ~n3451 & n6051;
  assign n7258 = ~n3525 & ~n6061;
  assign n7259 = ~n7257 & ~n7258;
  assign n7260 = ~n6043 & ~n7259;
  assign n7261 = n6043 & n7259;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7256 & ~n7262;
  assign n7264 = n7256 & n7262;
  assign n7265 = ~n3383 & n6051;
  assign n7266 = ~n3458 & ~n6061;
  assign n7267 = ~n7265 & ~n7266;
  assign n7268 = ~n6043 & ~n7267;
  assign n7269 = n6043 & n7267;
  assign n7270 = ~n7268 & ~n7269;
  assign n7271 = ~n3383 & ~n6048;
  assign n7272 = ~n3458 & n6051;
  assign n7273 = ~n7271 & ~n7272;
  assign n7274 = n7270 & n7273;
  assign n7275 = ~n3314 & ~n6048;
  assign n7276 = ~n3390 & n6051;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = ~n3314 & n6051;
  assign n7279 = ~n3390 & ~n6061;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = ~n6043 & ~n7280;
  assign n7282 = n6043 & n7280;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 = ~n7277 & ~n7283;
  assign n7285 = n7277 & n7283;
  assign n7286 = ~n3240 & ~n6048;
  assign n7287 = ~n3321 & n6051;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = ~n3176 & ~n6048;
  assign n7290 = ~n3247 & n6051;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n3176 & n6051;
  assign n7293 = ~n3247 & ~n6061;
  assign n7294 = ~n7292 & ~n7293;
  assign n7295 = ~n6043 & ~n7294;
  assign n7296 = n6043 & n7294;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = ~n7291 & ~n7297;
  assign n7299 = ~n7288 & n7298;
  assign n7300 = ~n3240 & n6051;
  assign n7301 = ~n3321 & ~n6061;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = ~n6043 & ~n7302;
  assign n7304 = n6043 & n7302;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = n7288 & ~n7298;
  assign n7307 = ~n7305 & ~n7306;
  assign n7308 = ~n7299 & ~n7307;
  assign n7309 = n7291 & n7297;
  assign n7310 = n7288 & n7305;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~n3107 & ~n6048;
  assign n7313 = ~n3183 & n6051;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n3107 & n6051;
  assign n7316 = ~n3183 & ~n6061;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = ~n6043 & ~n7317;
  assign n7319 = n6043 & n7317;
  assign n7320 = ~n7318 & ~n7319;
  assign n7321 = ~n7314 & ~n7320;
  assign n7322 = n7314 & n7320;
  assign n7323 = ~n3041 & n6051;
  assign n7324 = ~n3114 & ~n6061;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~n6043 & ~n7325;
  assign n7327 = n6043 & n7325;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~n3041 & ~n6048;
  assign n7330 = ~n3114 & n6051;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = n7328 & n7331;
  assign n7333 = ~n2977 & ~n6048;
  assign n7334 = ~n3048 & n6051;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n2921 & ~n6048;
  assign n7337 = ~n2984 & n6051;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~n2921 & n6051;
  assign n7340 = ~n2984 & ~n6061;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = ~n6043 & ~n7341;
  assign n7343 = n6043 & n7341;
  assign n7344 = ~n7342 & ~n7343;
  assign n7345 = ~n7338 & ~n7344;
  assign n7346 = ~n7335 & n7345;
  assign n7347 = ~n2977 & n6051;
  assign n7348 = ~n3048 & ~n6061;
  assign n7349 = ~n7347 & ~n7348;
  assign n7350 = ~n6043 & ~n7349;
  assign n7351 = n6043 & n7349;
  assign n7352 = ~n7350 & ~n7351;
  assign n7353 = n7335 & ~n7345;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n7346 & ~n7354;
  assign n7356 = n7338 & n7344;
  assign n7357 = n7335 & n7352;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = ~n2851 & ~n6048;
  assign n7360 = ~n2928 & n6051;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = ~n2851 & n6051;
  assign n7363 = ~n2928 & ~n6061;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = ~n6043 & ~n7364;
  assign n7366 = n6043 & n7364;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = ~n7361 & ~n7367;
  assign n7369 = n7361 & n7367;
  assign n7370 = n6043 & ~n6054;
  assign n7371 = ~n6043 & n6054;
  assign n7372 = ~n6066 & ~n7371;
  assign n7373 = ~n7370 & ~n7372;
  assign n7374 = ~n7369 & ~n7373;
  assign n7375 = ~n7368 & ~n7374;
  assign n7376 = n7358 & ~n7375;
  assign n7377 = n7355 & ~n7376;
  assign n7378 = ~n7332 & ~n7377;
  assign n7379 = ~n7328 & ~n7331;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = ~n7322 & ~n7380;
  assign n7382 = ~n7321 & ~n7381;
  assign n7383 = n7311 & ~n7382;
  assign n7384 = n7308 & ~n7383;
  assign n7385 = ~n7285 & ~n7384;
  assign n7386 = ~n7284 & ~n7385;
  assign n7387 = ~n7274 & ~n7386;
  assign n7388 = ~n7270 & ~n7273;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = ~n7264 & ~n7389;
  assign n7391 = ~n7263 & ~n7390;
  assign n7392 = n7253 & ~n7391;
  assign n7393 = ~n7251 & ~n7392;
  assign n7394 = ~n7214 & ~n7393;
  assign n7395 = ~n7213 & ~n7394;
  assign n7396 = ~n3784 & n6051;
  assign n7397 = ~n3860 & ~n6061;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = ~n6043 & ~n7398;
  assign n7400 = n6043 & n7398;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = ~n3784 & ~n6048;
  assign n7403 = ~n3860 & n6051;
  assign n7404 = ~n7402 & ~n7403;
  assign n7405 = ~n7401 & n7404;
  assign n7406 = n7401 & ~n7404;
  assign n7407 = ~n7405 & ~n7406;
  assign n7408 = n7395 & ~n7407;
  assign n7409 = ~n7395 & n7407;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = n2696 & ~n7185;
  assign n7412 = n7172 & n7411;
  assign n7413 = ~n7410 & n7412;
  assign n7414 = ~n7190 & ~n7194;
  assign n7415 = ~n5638 & n7414;
  assign n7416 = ~n7203 & n7415;
  assign n1175 = n7413 | ~n7416;
  assign n7418 = ~n4900 & ~n7172;
  assign n7419 = n7187 & ~n7418;
  assign n7420 = P1_STATE_REG & ~n7419;
  assign n7421 = ~n4473 & n7420;
  assign n7422 = ~n4900 & n7172;
  assign n7423 = ~n4890 & ~n7422;
  assign n7424 = n2696 & ~n7423;
  assign n7425 = n4536 & n7424;
  assign n7426 = P1_REG3_REG_26_ & ~P1_STATE_REG;
  assign n7427 = ~n4473 & ~n7172;
  assign n7428 = ~n4413 & n7197;
  assign n7429 = ~n4534 & n7199;
  assign n7430 = ~n7427 & ~n7428;
  assign n7431 = ~n7429 & n7430;
  assign n7432 = n7195 & ~n7431;
  assign n7433 = ~n4477 & n6051;
  assign n7434 = n4536 & ~n6061;
  assign n7435 = ~n7433 & ~n7434;
  assign n7436 = ~n6043 & ~n7435;
  assign n7437 = n6043 & n7435;
  assign n7438 = ~n7436 & ~n7437;
  assign n7439 = ~n4477 & ~n6048;
  assign n7440 = n4536 & n6051;
  assign n7441 = ~n7439 & ~n7440;
  assign n7442 = ~n7438 & n7441;
  assign n7443 = n7438 & ~n7441;
  assign n7444 = ~n7442 & ~n7443;
  assign n7445 = ~n4413 & ~n6048;
  assign n7446 = n4479 & n6051;
  assign n7447 = ~n7445 & ~n7446;
  assign n7448 = ~n4413 & n6051;
  assign n7449 = n4479 & ~n6061;
  assign n7450 = ~n7448 & ~n7449;
  assign n7451 = ~n6043 & ~n7450;
  assign n7452 = n6043 & n7450;
  assign n7453 = ~n7451 & ~n7452;
  assign n7454 = ~n7447 & ~n7453;
  assign n7455 = n7444 & ~n7454;
  assign n7456 = ~n4367 & ~n6048;
  assign n7457 = n4415 & n6051;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = ~n4367 & n6051;
  assign n7460 = n4415 & ~n6061;
  assign n7461 = ~n7459 & ~n7460;
  assign n7462 = ~n6043 & ~n7461;
  assign n7463 = n6043 & n7461;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = ~n7458 & ~n7464;
  assign n7466 = n7458 & n7464;
  assign n7467 = ~n4298 & ~n6048;
  assign n7468 = n4344 & n6051;
  assign n7469 = ~n7467 & ~n7468;
  assign n7470 = ~n4298 & n6051;
  assign n7471 = n4344 & ~n6061;
  assign n7472 = ~n7470 & ~n7471;
  assign n7473 = ~n6043 & ~n7472;
  assign n7474 = n6043 & n7472;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = ~n7469 & ~n7475;
  assign n7477 = n7469 & n7475;
  assign n7478 = ~n4233 & ~n6048;
  assign n7479 = n4282 & n6051;
  assign n7480 = ~n7478 & ~n7479;
  assign n7481 = ~n4233 & n6051;
  assign n7482 = n4282 & ~n6061;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n6043 & ~n7483;
  assign n7485 = n6043 & n7483;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = ~n7480 & ~n7486;
  assign n7488 = n7480 & n7486;
  assign n7489 = ~n4180 & n6051;
  assign n7490 = n4235 & ~n6061;
  assign n7491 = ~n7489 & ~n7490;
  assign n7492 = ~n6043 & ~n7491;
  assign n7493 = n6043 & n7491;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~n4180 & ~n6048;
  assign n7496 = n4235 & n6051;
  assign n7497 = ~n7495 & ~n7496;
  assign n7498 = n7494 & n7497;
  assign n7499 = ~n7494 & ~n7497;
  assign n7500 = ~n4113 & ~n6048;
  assign n7501 = n4164 & n6051;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = ~n4113 & n6051;
  assign n7504 = n4164 & ~n6061;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n6043 & ~n7505;
  assign n7507 = n6043 & n7505;
  assign n7508 = ~n7506 & ~n7507;
  assign n7509 = ~n7502 & ~n7508;
  assign n7510 = ~n7499 & ~n7509;
  assign n7511 = ~n4046 & ~n6048;
  assign n7512 = ~n4117 & n6051;
  assign n7513 = ~n7511 & ~n7512;
  assign n7514 = ~n4046 & n6051;
  assign n7515 = ~n4117 & ~n6061;
  assign n7516 = ~n7514 & ~n7515;
  assign n7517 = ~n6043 & ~n7516;
  assign n7518 = n6043 & n7516;
  assign n7519 = ~n7517 & ~n7518;
  assign n7520 = ~n7513 & ~n7519;
  assign n7521 = n7502 & n7508;
  assign n7522 = ~n7498 & ~n7521;
  assign n7523 = n7520 & n7522;
  assign n7524 = n7510 & ~n7523;
  assign n7525 = ~n7498 & ~n7524;
  assign n7526 = n7513 & n7519;
  assign n7527 = n7522 & ~n7526;
  assign n7528 = ~n3977 & ~n6048;
  assign n7529 = ~n4059 & n6051;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = ~n3977 & n6051;
  assign n7532 = ~n4059 & ~n6061;
  assign n7533 = ~n7531 & ~n7532;
  assign n7534 = ~n6043 & ~n7533;
  assign n7535 = n6043 & n7533;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = ~n7530 & ~n7536;
  assign n7538 = n7530 & n7536;
  assign n7539 = ~n3910 & ~n6048;
  assign n7540 = ~n3984 & n6051;
  assign n7541 = ~n7539 & ~n7540;
  assign n7542 = ~n3849 & ~n6048;
  assign n7543 = ~n3917 & n6051;
  assign n7544 = ~n7542 & ~n7543;
  assign n7545 = ~n3849 & n6051;
  assign n7546 = ~n3917 & ~n6061;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = ~n6043 & ~n7547;
  assign n7549 = n6043 & n7547;
  assign n7550 = ~n7548 & ~n7549;
  assign n7551 = ~n7544 & ~n7550;
  assign n7552 = ~n7541 & n7551;
  assign n7553 = ~n3910 & n6051;
  assign n7554 = ~n3984 & ~n6061;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = ~n6043 & ~n7555;
  assign n7557 = n6043 & n7555;
  assign n7558 = ~n7556 & ~n7557;
  assign n7559 = n7541 & ~n7551;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~n7552 & ~n7560;
  assign n7562 = n7544 & n7550;
  assign n7563 = n7541 & n7558;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = ~n7401 & ~n7404;
  assign n7566 = n7401 & n7404;
  assign n7567 = ~n7395 & ~n7566;
  assign n7568 = ~n7565 & ~n7567;
  assign n7569 = n7564 & ~n7568;
  assign n7570 = n7561 & ~n7569;
  assign n7571 = ~n7538 & ~n7570;
  assign n7572 = ~n7537 & ~n7571;
  assign n7573 = n7527 & ~n7572;
  assign n7574 = ~n7525 & ~n7573;
  assign n7575 = ~n7488 & ~n7574;
  assign n7576 = ~n7487 & ~n7575;
  assign n7577 = ~n7477 & ~n7576;
  assign n7578 = ~n7476 & ~n7577;
  assign n7579 = ~n7466 & ~n7578;
  assign n7580 = ~n7465 & ~n7579;
  assign n7581 = n7455 & n7580;
  assign n7582 = n7447 & n7453;
  assign n7583 = n7444 & n7582;
  assign n7584 = ~n7438 & ~n7441;
  assign n7585 = ~n7441 & ~n7582;
  assign n7586 = ~n7438 & ~n7582;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = ~n7584 & ~n7587;
  assign n7589 = ~n7454 & ~n7465;
  assign n7590 = ~n7579 & n7589;
  assign n7591 = n7588 & ~n7590;
  assign n7592 = ~n7581 & ~n7583;
  assign n7593 = ~n7591 & n7592;
  assign n7594 = n7412 & n7593;
  assign n7595 = ~n7421 & ~n7425;
  assign n7596 = ~n7426 & n7595;
  assign n7597 = ~n7432 & n7596;
  assign n1180 = n7594 | ~n7597;
  assign n7599 = ~n3169 & ~n7189;
  assign n7600 = ~n3247 & ~n7193;
  assign n7601 = ~n3240 & n7199;
  assign n7602 = ~n3107 & n7197;
  assign n7603 = ~n3169 & ~n7172;
  assign n7604 = ~n7601 & ~n7602;
  assign n7605 = ~n7603 & n7604;
  assign n7606 = n7195 & ~n7605;
  assign n7607 = n7291 & ~n7297;
  assign n7608 = ~n7291 & n7297;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = n7382 & ~n7609;
  assign n7611 = ~n7298 & ~n7309;
  assign n7612 = ~n7382 & ~n7611;
  assign n7613 = ~n7610 & ~n7612;
  assign n7614 = n7412 & ~n7613;
  assign n7615 = ~n7599 & ~n7600;
  assign n7616 = ~n5945 & n7615;
  assign n7617 = ~n7606 & n7616;
  assign n1185 = n7614 | ~n7617;
  assign n7619 = ~n3973 & ~n7189;
  assign n7620 = ~n4059 & ~n7193;
  assign n7621 = ~n3973 & ~n7172;
  assign n7622 = ~n3910 & n7197;
  assign n7623 = ~n4046 & n7199;
  assign n7624 = ~n7621 & ~n7622;
  assign n7625 = ~n7623 & n7624;
  assign n7626 = n7195 & ~n7625;
  assign n7627 = n7530 & ~n7536;
  assign n7628 = ~n7530 & n7536;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = n7570 & ~n7629;
  assign n7631 = ~n7570 & n7629;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = n7412 & ~n7632;
  assign n7634 = ~n7619 & ~n7620;
  assign n7635 = ~n5542 & n7634;
  assign n7636 = ~n7626 & n7635;
  assign n1190 = n7633 | ~n7636;
  assign n7638 = P1_REG3_REG_2_ & ~n7189;
  assign n7639 = ~n2984 & ~n7193;
  assign n7640 = ~n2977 & n7199;
  assign n7641 = ~n2851 & n7197;
  assign n7642 = P1_REG3_REG_2_ & ~n7172;
  assign n7643 = ~n7640 & ~n7641;
  assign n7644 = ~n7642 & n7643;
  assign n7645 = n7195 & ~n7644;
  assign n7646 = n7338 & ~n7344;
  assign n7647 = ~n7338 & n7344;
  assign n7648 = ~n7646 & ~n7647;
  assign n7649 = n7375 & ~n7648;
  assign n7650 = ~n7345 & ~n7356;
  assign n7651 = ~n7375 & ~n7650;
  assign n7652 = ~n7649 & ~n7651;
  assign n7653 = n7412 & ~n7652;
  assign n7654 = ~n6126 & ~n7653;
  assign n7655 = ~n7638 & ~n7639;
  assign n7656 = ~n7645 & n7655;
  assign n1195 = ~n7654 | ~n7656;
  assign n7658 = ~n3514 & ~n7189;
  assign n7659 = ~n3578 & ~n7193;
  assign n7660 = ~n3607 & n7199;
  assign n7661 = ~n3451 & n7197;
  assign n7662 = ~n3514 & ~n7172;
  assign n7663 = ~n7660 & ~n7661;
  assign n7664 = ~n7662 & n7663;
  assign n7665 = n7195 & ~n7664;
  assign n7666 = n7239 & ~n7245;
  assign n7667 = ~n7239 & n7245;
  assign n7668 = ~n7666 & ~n7667;
  assign n7669 = n7391 & ~n7668;
  assign n7670 = ~n7246 & ~n7252;
  assign n7671 = ~n7391 & ~n7670;
  assign n7672 = ~n7669 & ~n7671;
  assign n7673 = n7412 & ~n7672;
  assign n7674 = ~n7658 & ~n7659;
  assign n7675 = ~n5765 & n7674;
  assign n7676 = ~n7665 & n7675;
  assign n1200 = n7673 | ~n7676;
  assign n7678 = ~n4229 & n7420;
  assign n7679 = n4282 & n7424;
  assign n7680 = P1_REG3_REG_22_ & ~P1_STATE_REG;
  assign n7681 = ~n4229 & ~n7172;
  assign n7682 = ~n4180 & n7197;
  assign n7683 = ~n4298 & n7199;
  assign n7684 = ~n7681 & ~n7682;
  assign n7685 = ~n7683 & n7684;
  assign n7686 = n7195 & ~n7685;
  assign n7687 = n7480 & ~n7486;
  assign n7688 = ~n7480 & n7486;
  assign n7689 = ~n7687 & ~n7688;
  assign n7690 = n7574 & ~n7689;
  assign n7691 = ~n7574 & n7689;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = n7412 & ~n7692;
  assign n7694 = ~n7678 & ~n7679;
  assign n7695 = ~n7680 & n7694;
  assign n7696 = ~n7686 & n7695;
  assign n1205 = n7693 | ~n7696;
  assign n7698 = ~n3668 & ~n7189;
  assign n7699 = ~n3715 & ~n7193;
  assign n7700 = ~n3668 & ~n7172;
  assign n7701 = ~n3607 & n7197;
  assign n7702 = ~n3731 & n7199;
  assign n7703 = ~n7700 & ~n7701;
  assign n7704 = ~n7702 & n7703;
  assign n7705 = n7195 & ~n7704;
  assign n7706 = ~n7225 & n7248;
  assign n7707 = ~n7252 & ~n7391;
  assign n7708 = ~n7246 & ~n7707;
  assign n7709 = ~n7235 & n7708;
  assign n7710 = n7706 & ~n7709;
  assign n7711 = ~n7220 & n7223;
  assign n7712 = n7220 & ~n7223;
  assign n7713 = ~n7711 & ~n7712;
  assign n7714 = ~n7235 & n7713;
  assign n7715 = ~n7247 & ~n7708;
  assign n7716 = n7714 & ~n7715;
  assign n7717 = ~n7710 & ~n7716;
  assign n7718 = n7412 & n7717;
  assign n7719 = ~n7698 & ~n7699;
  assign n7720 = ~n5700 & n7719;
  assign n7721 = ~n7705 & n7720;
  assign n1210 = n7718 | ~n7721;
  assign n7723 = ~n4109 & n7420;
  assign n7724 = n4164 & n7424;
  assign n7725 = P1_REG3_REG_20_ & ~P1_STATE_REG;
  assign n7726 = ~n4109 & ~n7172;
  assign n7727 = ~n4046 & n7197;
  assign n7728 = ~n4180 & n7199;
  assign n7729 = ~n7726 & ~n7727;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = n7195 & ~n7730;
  assign n7732 = n7502 & ~n7508;
  assign n7733 = ~n7502 & n7508;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = ~n7526 & ~n7572;
  assign n7736 = ~n7520 & ~n7735;
  assign n7737 = ~n7734 & n7736;
  assign n7738 = ~n7509 & ~n7521;
  assign n7739 = ~n7736 & ~n7738;
  assign n7740 = ~n7737 & ~n7739;
  assign n7741 = n7412 & ~n7740;
  assign n7742 = ~n7723 & ~n7724;
  assign n7743 = ~n7725 & n7742;
  assign n7744 = ~n7731 & n7743;
  assign n1215 = n7741 | ~n7744;
  assign n7746 = ~n6069 & n7412;
  assign n7747 = ~n6181 & ~n7746;
  assign n7748 = ~n7170 & ~n7195;
  assign n7749 = ~n7172 & ~n7748;
  assign n7750 = ~n7188 & ~n7749;
  assign n7751 = P1_REG3_REG_0_ & ~n7750;
  assign n7752 = ~n2862 & ~n7193;
  assign n7753 = ~n2851 & n7195;
  assign n7754 = n7199 & n7753;
  assign n7755 = ~n7752 & ~n7754;
  assign n7756 = n7747 & ~n7751;
  assign n1220 = ~n7755 | ~n7756;
  assign n7758 = ~n3379 & ~n7189;
  assign n7759 = ~n3458 & ~n7193;
  assign n7760 = ~n3451 & n7199;
  assign n7761 = ~n3314 & n7197;
  assign n7762 = ~n3379 & ~n7172;
  assign n7763 = ~n7760 & ~n7761;
  assign n7764 = ~n7762 & n7763;
  assign n7765 = n7195 & ~n7764;
  assign n7766 = ~n7270 & n7273;
  assign n7767 = n7270 & ~n7273;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = n7386 & ~n7768;
  assign n7770 = ~n7386 & n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = n7412 & ~n7771;
  assign n7773 = ~n7758 & ~n7759;
  assign n7774 = ~n5835 & n7773;
  assign n7775 = ~n7765 & n7774;
  assign n1225 = n7772 | ~n7775;
  assign n7777 = ~n3034 & ~n7189;
  assign n7778 = ~n3114 & ~n7193;
  assign n7779 = ~n3107 & n7199;
  assign n7780 = ~n2977 & n7197;
  assign n7781 = ~n3034 & ~n7172;
  assign n7782 = ~n7779 & ~n7780;
  assign n7783 = ~n7781 & n7782;
  assign n7784 = n7195 & ~n7783;
  assign n7785 = ~n7328 & n7331;
  assign n7786 = n7328 & ~n7331;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = n7377 & ~n7787;
  assign n7789 = ~n7377 & n7787;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = n7412 & ~n7790;
  assign n7792 = ~n7777 & ~n7778;
  assign n7793 = ~n6017 & n7792;
  assign n7794 = ~n7784 & n7793;
  assign n1230 = n7791 | ~n7794;
  assign n7796 = ~n4363 & n7420;
  assign n7797 = n4415 & n7424;
  assign n7798 = P1_REG3_REG_24_ & ~P1_STATE_REG;
  assign n7799 = ~n4363 & ~n7172;
  assign n7800 = ~n4298 & n7197;
  assign n7801 = ~n4413 & n7199;
  assign n7802 = ~n7799 & ~n7800;
  assign n7803 = ~n7801 & n7802;
  assign n7804 = n7195 & ~n7803;
  assign n7805 = n7458 & ~n7464;
  assign n7806 = ~n7458 & n7464;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = n7578 & ~n7807;
  assign n7809 = ~n7465 & ~n7466;
  assign n7810 = ~n7578 & ~n7809;
  assign n7811 = ~n7808 & ~n7810;
  assign n7812 = n7412 & ~n7811;
  assign n7813 = ~n7796 & ~n7797;
  assign n7814 = ~n7798 & n7813;
  assign n7815 = ~n7804 & n7814;
  assign n1235 = n7812 | ~n7815;
  assign n7817 = ~n3906 & ~n7189;
  assign n7818 = ~n3984 & ~n7193;
  assign n7819 = ~n3906 & ~n7172;
  assign n7820 = ~n3849 & n7197;
  assign n7821 = ~n3977 & n7199;
  assign n7822 = ~n7819 & ~n7820;
  assign n7823 = ~n7821 & n7822;
  assign n7824 = n7195 & ~n7823;
  assign n7825 = ~n7541 & ~n7558;
  assign n7826 = n7564 & ~n7825;
  assign n7827 = ~n7551 & n7568;
  assign n7828 = n7826 & ~n7827;
  assign n7829 = n7541 & ~n7558;
  assign n7830 = ~n7541 & n7558;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = ~n7551 & n7831;
  assign n7833 = ~n7562 & ~n7568;
  assign n7834 = n7832 & ~n7833;
  assign n7835 = ~n7828 & ~n7834;
  assign n7836 = n7412 & n7835;
  assign n7837 = ~n7817 & ~n7818;
  assign n7838 = ~n5575 & n7837;
  assign n7839 = ~n7824 & n7838;
  assign n1240 = n7836 | ~n7839;
  assign n7841 = ~n3100 & ~n7189;
  assign n7842 = ~n3183 & ~n7193;
  assign n7843 = ~n3176 & n7199;
  assign n7844 = ~n3041 & n7197;
  assign n7845 = ~n3100 & ~n7172;
  assign n7846 = ~n7843 & ~n7844;
  assign n7847 = ~n7845 & n7846;
  assign n7848 = n7195 & ~n7847;
  assign n7849 = n7314 & ~n7320;
  assign n7850 = ~n7314 & n7320;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = n7380 & ~n7851;
  assign n7853 = ~n7380 & n7851;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = n7412 & ~n7854;
  assign n7856 = ~n7841 & ~n7842;
  assign n7857 = ~n5995 & n7856;
  assign n7858 = ~n7848 & n7857;
  assign n1245 = n7855 | ~n7858;
  assign n7860 = ~n3845 & ~n7189;
  assign n7861 = ~n3917 & ~n7193;
  assign n7862 = ~n3845 & ~n7172;
  assign n7863 = ~n3784 & n7197;
  assign n7864 = ~n3910 & n7199;
  assign n7865 = ~n7862 & ~n7863;
  assign n7866 = ~n7864 & n7865;
  assign n7867 = n7195 & ~n7866;
  assign n7868 = n7544 & ~n7550;
  assign n7869 = ~n7544 & n7550;
  assign n7870 = ~n7868 & ~n7869;
  assign n7871 = n7568 & ~n7870;
  assign n7872 = ~n7551 & ~n7562;
  assign n7873 = ~n7568 & ~n7872;
  assign n7874 = ~n7871 & ~n7873;
  assign n7875 = n7412 & ~n7874;
  assign n7876 = ~n7860 & ~n7861;
  assign n7877 = ~n5609 & n7876;
  assign n7878 = ~n7867 & n7877;
  assign n1250 = n7875 | ~n7878;
  assign n7880 = ~n4409 & n7420;
  assign n7881 = n4479 & n7424;
  assign n7882 = P1_REG3_REG_25_ & ~P1_STATE_REG;
  assign n7883 = ~n4409 & ~n7172;
  assign n7884 = ~n4367 & n7197;
  assign n7885 = ~n4477 & n7199;
  assign n7886 = ~n7883 & ~n7884;
  assign n7887 = ~n7885 & n7886;
  assign n7888 = n7195 & ~n7887;
  assign n7889 = n7447 & ~n7453;
  assign n7890 = ~n7447 & n7453;
  assign n7891 = ~n7889 & ~n7890;
  assign n7892 = n7580 & ~n7891;
  assign n7893 = ~n7454 & ~n7582;
  assign n7894 = ~n7580 & ~n7893;
  assign n7895 = ~n7892 & ~n7894;
  assign n7896 = n7412 & ~n7895;
  assign n7897 = ~n7880 & ~n7881;
  assign n7898 = ~n7882 & n7897;
  assign n7899 = ~n7888 & n7898;
  assign n1255 = n7896 | ~n7899;
  assign n7901 = ~n3603 & ~n7189;
  assign n7902 = ~n3648 & ~n7193;
  assign n7903 = ~n3603 & ~n7172;
  assign n7904 = ~n3518 & n7197;
  assign n7905 = ~n3672 & n7199;
  assign n7906 = ~n7903 & ~n7904;
  assign n7907 = ~n7905 & n7906;
  assign n7908 = n7195 & ~n7907;
  assign n7909 = n7228 & ~n7234;
  assign n7910 = ~n7228 & n7234;
  assign n7911 = ~n7909 & ~n7910;
  assign n7912 = n7708 & ~n7911;
  assign n7913 = ~n7235 & ~n7247;
  assign n7914 = ~n7708 & ~n7913;
  assign n7915 = ~n7912 & ~n7914;
  assign n7916 = n7412 & ~n7915;
  assign n7917 = ~n7901 & ~n7902;
  assign n7918 = ~n5735 & n7917;
  assign n7919 = ~n7908 & n7918;
  assign n1260 = n7916 | ~n7919;
  assign n7921 = ~n4176 & n7420;
  assign n7922 = n4235 & n7424;
  assign n7923 = P1_REG3_REG_21_ & ~P1_STATE_REG;
  assign n7924 = ~n4176 & ~n7172;
  assign n7925 = ~n4113 & n7197;
  assign n7926 = ~n4233 & n7199;
  assign n7927 = ~n7924 & ~n7925;
  assign n7928 = ~n7926 & n7927;
  assign n7929 = n7195 & ~n7928;
  assign n7930 = ~n7499 & n7522;
  assign n7931 = ~n7509 & n7736;
  assign n7932 = n7930 & ~n7931;
  assign n7933 = ~n7494 & n7497;
  assign n7934 = n7494 & ~n7497;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7509 & n7935;
  assign n7937 = ~n7521 & ~n7736;
  assign n7938 = n7936 & ~n7937;
  assign n7939 = ~n7932 & ~n7938;
  assign n7940 = n7412 & n7939;
  assign n7941 = ~n7921 & ~n7922;
  assign n7942 = ~n7923 & n7941;
  assign n7943 = ~n7929 & n7942;
  assign n1265 = n7940 | ~n7943;
  assign n7945 = P1_REG3_REG_1_ & ~n7189;
  assign n7946 = ~n2928 & ~n7193;
  assign n7947 = n7361 & ~n7367;
  assign n7948 = ~n7361 & n7367;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = n7373 & ~n7949;
  assign n7951 = ~n7373 & n7949;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = n7412 & ~n7952;
  assign n7954 = ~n6159 & ~n7953;
  assign n7955 = ~n2921 & n7199;
  assign n7956 = ~n2878 & n7197;
  assign n7957 = P1_REG3_REG_1_ & ~n7172;
  assign n7958 = ~n7955 & ~n7956;
  assign n7959 = ~n7957 & n7958;
  assign n7960 = n7195 & ~n7959;
  assign n7961 = ~n7945 & ~n7946;
  assign n7962 = n7954 & n7961;
  assign n1270 = n7960 | ~n7962;
  assign n7964 = ~n3307 & ~n7189;
  assign n7965 = ~n3390 & ~n7193;
  assign n7966 = ~n3383 & n7199;
  assign n7967 = ~n3240 & n7197;
  assign n7968 = ~n3307 & ~n7172;
  assign n7969 = ~n7966 & ~n7967;
  assign n7970 = ~n7968 & n7969;
  assign n7971 = n7195 & ~n7970;
  assign n7972 = n7277 & ~n7283;
  assign n7973 = ~n7277 & n7283;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = n7384 & ~n7974;
  assign n7976 = ~n7384 & n7974;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = n7412 & ~n7977;
  assign n7979 = ~n7964 & ~n7965;
  assign n7980 = ~n5865 & n7979;
  assign n7981 = ~n7971 & n7980;
  assign n1275 = n7978 | ~n7981;
  assign n7983 = ~n4590 & n7420;
  assign n7984 = n4653 & n7424;
  assign n7985 = P1_REG3_REG_28_ & ~P1_STATE_REG;
  assign n7986 = ~n4651 & n7199;
  assign n7987 = ~n4534 & n7197;
  assign n7988 = ~n4590 & ~n7172;
  assign n7989 = ~n7986 & ~n7987;
  assign n7990 = ~n7988 & n7989;
  assign n7991 = n7195 & ~n7990;
  assign n7992 = ~n4534 & n6051;
  assign n7993 = n4596 & ~n6061;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = ~n6043 & ~n7994;
  assign n7996 = n6043 & n7994;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = ~n4534 & ~n6048;
  assign n7999 = n4596 & n6051;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = n7997 & n8000;
  assign n8002 = n7584 & ~n8001;
  assign n8003 = ~n7466 & ~n8001;
  assign n8004 = ~n7578 & ~n7587;
  assign n8005 = n8003 & n8004;
  assign n8006 = ~n7587 & ~n7589;
  assign n8007 = ~n8001 & n8006;
  assign n8008 = ~n7997 & ~n8000;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~n4594 & ~n6048;
  assign n8011 = n4653 & n6051;
  assign n8012 = ~n8010 & ~n8011;
  assign n8013 = ~n6043 & ~n8012;
  assign n8014 = n6043 & n8012;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~n4594 & n6051;
  assign n8017 = n4653 & ~n6061;
  assign n8018 = ~n8016 & ~n8017;
  assign n8019 = ~n8015 & n8018;
  assign n8020 = n8015 & ~n8018;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = ~n8002 & ~n8005;
  assign n8023 = n8009 & n8022;
  assign n8024 = ~n8021 & n8023;
  assign n8025 = n7579 & ~n7587;
  assign n8026 = ~n7584 & ~n8008;
  assign n8027 = ~n8006 & ~n8025;
  assign n8028 = n8026 & n8027;
  assign n8029 = ~n8001 & ~n8028;
  assign n8030 = n8021 & n8029;
  assign n8031 = ~n8024 & ~n8030;
  assign n8032 = n7412 & ~n8031;
  assign n8033 = ~n7983 & ~n7984;
  assign n8034 = ~n7985 & n8033;
  assign n8035 = ~n7991 & n8034;
  assign n1280 = n8032 | ~n8035;
  assign n8037 = ~n4042 & ~n7189;
  assign n8038 = ~n4117 & ~n7193;
  assign n8039 = ~n4042 & ~n7172;
  assign n8040 = ~n3977 & n7197;
  assign n8041 = ~n4113 & n7199;
  assign n8042 = ~n8039 & ~n8040;
  assign n8043 = ~n8041 & n8042;
  assign n8044 = n7195 & ~n8043;
  assign n8045 = n7513 & ~n7519;
  assign n8046 = ~n7513 & n7519;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = n7572 & ~n8047;
  assign n8049 = ~n7520 & ~n7526;
  assign n8050 = ~n7572 & ~n8049;
  assign n8051 = ~n8048 & ~n8050;
  assign n8052 = n7412 & ~n8051;
  assign n8053 = ~n8037 & ~n8038;
  assign n8054 = ~n5412 & n8053;
  assign n8055 = ~n8044 & n8054;
  assign n1285 = n8052 | ~n8055;
  assign n8057 = ~P1_REG3_REG_3_ & ~n7189;
  assign n8058 = ~n3048 & ~n7193;
  assign n8059 = ~n3041 & n7199;
  assign n8060 = ~n2921 & n7197;
  assign n8061 = ~P1_REG3_REG_3_ & ~n7172;
  assign n8062 = ~n8059 & ~n8060;
  assign n8063 = ~n8061 & n8062;
  assign n8064 = n7195 & ~n8063;
  assign n8065 = ~n7335 & ~n7352;
  assign n8066 = n7358 & ~n8065;
  assign n8067 = ~n7345 & n7375;
  assign n8068 = n8066 & ~n8067;
  assign n8069 = n7335 & ~n7352;
  assign n8070 = ~n7335 & n7352;
  assign n8071 = ~n8069 & ~n8070;
  assign n8072 = ~n7345 & n8071;
  assign n8073 = ~n7356 & ~n7375;
  assign n8074 = n8072 & ~n8073;
  assign n8075 = ~n8068 & ~n8074;
  assign n8076 = n7412 & n8075;
  assign n8077 = ~n8057 & ~n8058;
  assign n8078 = ~n6103 & n8077;
  assign n8079 = ~n8064 & n8078;
  assign n1290 = n8076 | ~n8079;
  assign n8081 = ~n3447 & ~n7189;
  assign n8082 = ~n3525 & ~n7193;
  assign n8083 = ~n3518 & n7199;
  assign n8084 = ~n3383 & n7197;
  assign n8085 = ~n3447 & ~n7172;
  assign n8086 = ~n8083 & ~n8084;
  assign n8087 = ~n8085 & n8086;
  assign n8088 = n7195 & ~n8087;
  assign n8089 = n7256 & ~n7262;
  assign n8090 = ~n7256 & n7262;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = n7389 & ~n8091;
  assign n8093 = ~n7389 & n8091;
  assign n8094 = ~n8092 & ~n8093;
  assign n8095 = n7412 & ~n8094;
  assign n8096 = ~n8081 & ~n8082;
  assign n8097 = ~n5800 & n8096;
  assign n8098 = ~n8088 & n8097;
  assign n1295 = n8095 | ~n8098;
  assign n8100 = ~n4294 & n7420;
  assign n8101 = n4344 & n7424;
  assign n8102 = P1_REG3_REG_23_ & ~P1_STATE_REG;
  assign n8103 = ~n4294 & ~n7172;
  assign n8104 = ~n4233 & n7197;
  assign n8105 = ~n4367 & n7199;
  assign n8106 = ~n8103 & ~n8104;
  assign n8107 = ~n8105 & n8106;
  assign n8108 = n7195 & ~n8107;
  assign n8109 = n7469 & ~n7475;
  assign n8110 = ~n7469 & n7475;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = n7576 & ~n8111;
  assign n8113 = ~n7576 & n8111;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = n7412 & ~n8114;
  assign n8116 = ~n8100 & ~n8101;
  assign n8117 = ~n8102 & n8116;
  assign n8118 = ~n8108 & n8117;
  assign n1300 = n8115 | ~n8118;
  assign n8120 = ~n3727 & ~n7189;
  assign n8121 = ~n3798 & ~n7193;
  assign n8122 = ~n3727 & ~n7172;
  assign n8123 = ~n3672 & n7197;
  assign n8124 = ~n3784 & n7199;
  assign n8125 = ~n8122 & ~n8123;
  assign n8126 = ~n8124 & n8125;
  assign n8127 = n7195 & ~n8126;
  assign n8128 = n7206 & ~n7212;
  assign n8129 = ~n7206 & n7212;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = n7393 & ~n8130;
  assign n8132 = ~n7393 & n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = n7412 & ~n8133;
  assign n8135 = ~n8120 & ~n8121;
  assign n8136 = ~n5666 & n8135;
  assign n8137 = ~n8127 & n8136;
  assign n1305 = n8134 | ~n8137;
  assign n8139 = ~n4530 & n7420;
  assign n8140 = n4596 & n7424;
  assign n8141 = P1_REG3_REG_27_ & ~P1_STATE_REG;
  assign n8142 = ~n4530 & ~n7172;
  assign n8143 = ~n4477 & n7197;
  assign n8144 = ~n4594 & n7199;
  assign n8145 = ~n8142 & ~n8143;
  assign n8146 = ~n8144 & n8145;
  assign n8147 = n7195 & ~n8146;
  assign n8148 = ~n7584 & ~n8006;
  assign n8149 = ~n8025 & n8148;
  assign n8150 = ~n7997 & n8000;
  assign n8151 = n7997 & ~n8000;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = n8149 & ~n8152;
  assign n8154 = ~n8149 & n8152;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = n7412 & ~n8155;
  assign n8157 = ~n8139 & ~n8140;
  assign n8158 = ~n8141 & n8157;
  assign n8159 = ~n8147 & n8158;
  assign n1310 = n8156 | ~n8159;
  assign n8161 = ~n3233 & ~n7189;
  assign n8162 = ~n3321 & ~n7193;
  assign n8163 = ~n3314 & n7199;
  assign n8164 = ~n3176 & n7197;
  assign n8165 = ~n3233 & ~n7172;
  assign n8166 = ~n8163 & ~n8164;
  assign n8167 = ~n8165 & n8166;
  assign n8168 = n7195 & ~n8167;
  assign n8169 = ~n7288 & ~n7305;
  assign n8170 = n7311 & ~n8169;
  assign n8171 = ~n7298 & n7382;
  assign n8172 = n8170 & ~n8171;
  assign n8173 = n7288 & ~n7305;
  assign n8174 = ~n7288 & n7305;
  assign n8175 = ~n8173 & ~n8174;
  assign n8176 = ~n7298 & n8175;
  assign n8177 = ~n7309 & ~n7382;
  assign n8178 = n8176 & ~n8177;
  assign n8179 = ~n8172 & ~n8178;
  assign n8180 = n7412 & n8179;
  assign n8181 = ~n8161 & ~n8162;
  assign n8182 = ~n5899 & n8181;
  assign n8183 = ~n8168 & n8182;
  assign n1315 = n8180 | ~n8183;
  assign n8185 = ~P2_IR_REG_31_ & P2_STATE_REG;
  assign n8186 = P2_STATE_REG & ~n8185;
  assign n8187 = P2_IR_REG_0_ & n8186;
  assign n8188 = P2_IR_REG_0_ & n8185;
  assign n8189 = n1734 & ~n1741;
  assign n8190 = P1_DATAO_REG_0_ & ~n1734;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = ~P2_STATE_REG & ~n8191;
  assign n8193 = ~n8187 & ~n8188;
  assign n1335 = n8192 | ~n8193;
  assign n8195 = P2_IR_REG_0_ & ~P2_IR_REG_1_;
  assign n8196 = ~P2_IR_REG_0_ & P2_IR_REG_1_;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = n8186 & ~n8197;
  assign n8199 = P2_IR_REG_1_ & n8185;
  assign n8200 = n1734 & ~n1767;
  assign n8201 = P1_DATAO_REG_1_ & ~n1734;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = ~P2_STATE_REG & ~n8202;
  assign n8204 = ~n8198 & ~n8199;
  assign n1340 = n8203 | ~n8204;
  assign n8206 = ~P2_IR_REG_0_ & ~P2_IR_REG_1_;
  assign n8207 = P2_IR_REG_2_ & ~n8206;
  assign n8208 = ~P2_IR_REG_2_ & n8206;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = n8186 & n8209;
  assign n8211 = P2_IR_REG_2_ & n8185;
  assign n8212 = n1734 & ~n1792;
  assign n8213 = P1_DATAO_REG_2_ & ~n1734;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~P2_STATE_REG & ~n8214;
  assign n8216 = ~n8210 & ~n8211;
  assign n1345 = n8215 | ~n8216;
  assign n8218 = P2_IR_REG_3_ & ~n8208;
  assign n8219 = ~P2_IR_REG_3_ & n8208;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = n8186 & n8220;
  assign n8222 = P2_IR_REG_3_ & n8185;
  assign n8223 = n1734 & ~n1816;
  assign n8224 = P1_DATAO_REG_3_ & ~n1734;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = ~P2_STATE_REG & ~n8225;
  assign n8227 = ~n8221 & ~n8222;
  assign n1350 = n8226 | ~n8227;
  assign n8229 = P2_IR_REG_4_ & ~n8219;
  assign n8230 = ~P2_IR_REG_4_ & n8219;
  assign n8231 = ~n8229 & ~n8230;
  assign n8232 = n8186 & n8231;
  assign n8233 = P2_IR_REG_4_ & n8185;
  assign n8234 = n1734 & ~n1844;
  assign n8235 = P1_DATAO_REG_4_ & ~n1734;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = ~P2_STATE_REG & ~n8236;
  assign n8238 = ~n8232 & ~n8233;
  assign n1355 = n8237 | ~n8238;
  assign n8240 = ~P2_IR_REG_5_ & n8230;
  assign n8241 = P2_IR_REG_5_ & ~n8230;
  assign n8242 = ~n8240 & ~n8241;
  assign n8243 = n8186 & n8242;
  assign n8244 = P2_IR_REG_5_ & n8185;
  assign n8245 = n1734 & ~n1868;
  assign n8246 = P1_DATAO_REG_5_ & ~n1734;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = ~P2_STATE_REG & ~n8247;
  assign n8249 = ~n8243 & ~n8244;
  assign n1360 = n8248 | ~n8249;
  assign n8251 = P2_IR_REG_6_ & ~n8240;
  assign n8252 = ~P2_IR_REG_5_ & ~P2_IR_REG_6_;
  assign n8253 = n8230 & n8252;
  assign n8254 = ~n8251 & ~n8253;
  assign n8255 = n8186 & n8254;
  assign n8256 = P2_IR_REG_6_ & n8185;
  assign n8257 = n1734 & ~n1896;
  assign n8258 = P1_DATAO_REG_6_ & ~n1734;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~P2_STATE_REG & ~n8259;
  assign n8261 = ~n8255 & ~n8256;
  assign n1365 = n8260 | ~n8261;
  assign n8263 = P2_IR_REG_7_ & ~n8253;
  assign n8264 = ~P2_IR_REG_7_ & n8253;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = n8186 & n8265;
  assign n8267 = P2_IR_REG_7_ & n8185;
  assign n8268 = n1734 & ~n1923;
  assign n8269 = P1_DATAO_REG_7_ & ~n1734;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~P2_STATE_REG & ~n8270;
  assign n8272 = ~n8266 & ~n8267;
  assign n1370 = n8271 | ~n8272;
  assign n8274 = P2_IR_REG_8_ & ~n8264;
  assign n8275 = ~P2_IR_REG_7_ & n8252;
  assign n8276 = ~P2_IR_REG_8_ & n8275;
  assign n8277 = ~P2_IR_REG_3_ & ~P2_IR_REG_4_;
  assign n8278 = ~P2_IR_REG_2_ & n8277;
  assign n8279 = ~P2_IR_REG_1_ & n8278;
  assign n8280 = ~P2_IR_REG_0_ & n8279;
  assign n8281 = n8276 & n8280;
  assign n8282 = ~n8274 & ~n8281;
  assign n8283 = n8186 & n8282;
  assign n8284 = P2_IR_REG_8_ & n8185;
  assign n8285 = n1734 & ~n1951;
  assign n8286 = P1_DATAO_REG_8_ & ~n1734;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~P2_STATE_REG & ~n8287;
  assign n8289 = ~n8283 & ~n8284;
  assign n1375 = n8288 | ~n8289;
  assign n8291 = ~P2_IR_REG_9_ & n8281;
  assign n8292 = P2_IR_REG_9_ & ~n8281;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = n8186 & n8293;
  assign n8295 = P2_IR_REG_9_ & n8185;
  assign n8296 = n1734 & ~n1978;
  assign n8297 = P1_DATAO_REG_9_ & ~n1734;
  assign n8298 = ~n8296 & ~n8297;
  assign n8299 = ~P2_STATE_REG & ~n8298;
  assign n8300 = ~n8294 & ~n8295;
  assign n1380 = n8299 | ~n8300;
  assign n8302 = P2_IR_REG_10_ & ~n8291;
  assign n8303 = ~P2_IR_REG_9_ & ~P2_IR_REG_10_;
  assign n8304 = n8281 & n8303;
  assign n8305 = ~n8302 & ~n8304;
  assign n8306 = n8186 & n8305;
  assign n8307 = P2_IR_REG_10_ & n8185;
  assign n8308 = n1734 & ~n2006;
  assign n8309 = P1_DATAO_REG_10_ & ~n1734;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = ~P2_STATE_REG & ~n8310;
  assign n8312 = ~n8306 & ~n8307;
  assign n1385 = n8311 | ~n8312;
  assign n8314 = P2_IR_REG_11_ & ~n8304;
  assign n8315 = ~P2_IR_REG_11_ & n8304;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = n8186 & n8316;
  assign n8318 = P2_IR_REG_11_ & n8185;
  assign n8319 = n1734 & ~n2033;
  assign n8320 = P1_DATAO_REG_11_ & ~n1734;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = ~P2_STATE_REG & ~n8321;
  assign n8323 = ~n8317 & ~n8318;
  assign n1390 = n8322 | ~n8323;
  assign n8325 = P2_IR_REG_12_ & ~n8315;
  assign n8326 = ~P2_IR_REG_9_ & ~P2_IR_REG_12_;
  assign n8327 = ~P2_IR_REG_10_ & n8326;
  assign n8328 = ~P2_IR_REG_11_ & n8327;
  assign n8329 = n8281 & n8328;
  assign n8330 = ~n8325 & ~n8329;
  assign n8331 = n8186 & n8330;
  assign n8332 = P2_IR_REG_12_ & n8185;
  assign n8333 = n1734 & ~n2060_1;
  assign n8334 = P1_DATAO_REG_12_ & ~n1734;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = ~P2_STATE_REG & ~n8335;
  assign n8337 = ~n8331 & ~n8332;
  assign n1395 = n8336 | ~n8337;
  assign n8339 = ~P2_IR_REG_13_ & n8329;
  assign n8340 = P2_IR_REG_13_ & ~n8329;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8186 & n8341;
  assign n8343 = P2_IR_REG_13_ & n8185;
  assign n8344 = n1734 & ~n2087;
  assign n8345 = P1_DATAO_REG_13_ & ~n1734;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = ~P2_STATE_REG & ~n8346;
  assign n8348 = ~n8342 & ~n8343;
  assign n1400 = n8347 | ~n8348;
  assign n8350 = P2_IR_REG_14_ & ~n8339;
  assign n8351 = ~P2_IR_REG_13_ & ~P2_IR_REG_14_;
  assign n8352 = n8329 & n8351;
  assign n8353 = ~n8350 & ~n8352;
  assign n8354 = n8186 & n8353;
  assign n8355 = P2_IR_REG_14_ & n8185;
  assign n8356 = n1734 & ~n2115_1;
  assign n8357 = P1_DATAO_REG_14_ & ~n1734;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = ~P2_STATE_REG & ~n8358;
  assign n8360 = ~n8354 & ~n8355;
  assign n1405 = n8359 | ~n8360;
  assign n8362 = P2_IR_REG_15_ & ~n8352;
  assign n8363 = ~P2_IR_REG_15_ & n8352;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n8186 & n8364;
  assign n8366 = P2_IR_REG_15_ & n8185;
  assign n8367 = n1734 & ~n2142;
  assign n8368 = P1_DATAO_REG_15_ & ~n1734;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = ~P2_STATE_REG & ~n8369;
  assign n8371 = ~n8365 & ~n8366;
  assign n1410 = n8370 | ~n8371;
  assign n8373 = P2_IR_REG_16_ & ~n8363;
  assign n8374 = ~P2_IR_REG_13_ & ~P2_IR_REG_15_;
  assign n8375 = ~P2_IR_REG_14_ & n8374;
  assign n8376 = ~P2_IR_REG_16_ & n8328;
  assign n8377 = n8375 & n8376;
  assign n8378 = n8281 & n8377;
  assign n8379 = ~n8373 & ~n8378;
  assign n8380 = n8186 & n8379;
  assign n8381 = P2_IR_REG_16_ & n8185;
  assign n8382 = n1734 & ~n2180_1;
  assign n8383 = P1_DATAO_REG_16_ & ~n1734;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~P2_STATE_REG & ~n8384;
  assign n8386 = ~n8380 & ~n8381;
  assign n1415 = n8385 | ~n8386;
  assign n8388 = ~P2_IR_REG_17_ & n8378;
  assign n8389 = P2_IR_REG_17_ & ~n8378;
  assign n8390 = ~n8388 & ~n8389;
  assign n8391 = n8186 & n8390;
  assign n8392 = P2_IR_REG_17_ & n8185;
  assign n8393 = n1734 & ~n2204;
  assign n8394 = P1_DATAO_REG_17_ & ~n1734;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~P2_STATE_REG & ~n8395;
  assign n8397 = ~n8391 & ~n8392;
  assign n1420 = n8396 | ~n8397;
  assign n8399 = P2_IR_REG_18_ & ~n8388;
  assign n8400 = ~P2_IR_REG_17_ & ~P2_IR_REG_18_;
  assign n8401 = n8378 & n8400;
  assign n8402 = ~n8399 & ~n8401;
  assign n8403 = n8186 & n8402;
  assign n8404 = P2_IR_REG_18_ & n8185;
  assign n8405 = n1734 & ~n2238;
  assign n8406 = P1_DATAO_REG_18_ & ~n1734;
  assign n8407 = ~n8405 & ~n8406;
  assign n8408 = ~P2_STATE_REG & ~n8407;
  assign n8409 = ~n8403 & ~n8404;
  assign n1425 = n8408 | ~n8409;
  assign n8411 = P2_IR_REG_19_ & ~n8401;
  assign n8412 = ~P2_IR_REG_19_ & n8401;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = n8186 & n8413;
  assign n8415 = P2_IR_REG_19_ & n8185;
  assign n8416 = n1734 & ~n2275_1;
  assign n8417 = P1_DATAO_REG_19_ & ~n1734;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = ~P2_STATE_REG & ~n8418;
  assign n8420 = ~n8414 & ~n8415;
  assign n1430 = n8419 | ~n8420;
  assign n8422 = P2_IR_REG_20_ & ~n8412;
  assign n8423 = ~P2_IR_REG_19_ & ~P2_IR_REG_20_;
  assign n8424 = ~P2_IR_REG_17_ & n8423;
  assign n8425 = ~P2_IR_REG_18_ & n8424;
  assign n8426 = n8378 & n8425;
  assign n8427 = ~n8422 & ~n8426;
  assign n8428 = n8186 & n8427;
  assign n8429 = P2_IR_REG_20_ & n8185;
  assign n8430 = n1734 & ~n2312;
  assign n8431 = P1_DATAO_REG_20_ & ~n1734;
  assign n8432 = ~n8430 & ~n8431;
  assign n8433 = ~P2_STATE_REG & ~n8432;
  assign n8434 = ~n8428 & ~n8429;
  assign n1435 = n8433 | ~n8434;
  assign n8436 = ~P2_IR_REG_21_ & n8426;
  assign n8437 = P2_IR_REG_21_ & ~n8426;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = n8186 & n8438;
  assign n8440 = P2_IR_REG_21_ & n8185;
  assign n8441 = n1734 & ~n2336;
  assign n8442 = P1_DATAO_REG_21_ & ~n1734;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = ~P2_STATE_REG & ~n8443;
  assign n8445 = ~n8439 & ~n8440;
  assign n1440 = n8444 | ~n8445;
  assign n8447 = P2_IR_REG_22_ & ~n8436;
  assign n8448 = ~P2_IR_REG_21_ & ~P2_IR_REG_22_;
  assign n8449 = n8426 & n8448;
  assign n8450 = ~n8447 & ~n8449;
  assign n8451 = n8186 & n8450;
  assign n8452 = P2_IR_REG_22_ & n8185;
  assign n8453 = n1734 & ~n2373;
  assign n8454 = P1_DATAO_REG_22_ & ~n1734;
  assign n8455 = ~n8453 & ~n8454;
  assign n8456 = ~P2_STATE_REG & ~n8455;
  assign n8457 = ~n8451 & ~n8452;
  assign n1445 = n8456 | ~n8457;
  assign n8459 = P2_IR_REG_23_ & ~n8449;
  assign n8460 = ~P2_IR_REG_23_ & n8449;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = n8186 & n8461;
  assign n8463 = P2_IR_REG_23_ & n8185;
  assign n8464 = n1734 & ~n2415_1;
  assign n8465 = P1_DATAO_REG_23_ & ~n1734;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = ~P2_STATE_REG & ~n8466;
  assign n8468 = ~n8462 & ~n8463;
  assign n1450 = n8467 | ~n8468;
  assign n8470 = P2_IR_REG_24_ & ~n8460;
  assign n8471 = ~P2_IR_REG_21_ & ~P2_IR_REG_23_;
  assign n8472 = ~P2_IR_REG_22_ & n8471;
  assign n8473 = ~P2_IR_REG_24_ & n8425;
  assign n8474 = n8472 & n8473;
  assign n8475 = n8378 & n8474;
  assign n8476 = ~n8470 & ~n8475;
  assign n8477 = n8186 & n8476;
  assign n8478 = P2_IR_REG_24_ & n8185;
  assign n8479 = n1734 & ~n2455_1;
  assign n8480 = P1_DATAO_REG_24_ & ~n1734;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~P2_STATE_REG & ~n8481;
  assign n8483 = ~n8477 & ~n8478;
  assign n1455 = n8482 | ~n8483;
  assign n8485 = ~P2_IR_REG_25_ & n8475;
  assign n8486 = P2_IR_REG_25_ & ~n8475;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = n8186 & n8487;
  assign n8489 = P2_IR_REG_25_ & n8185;
  assign n8490 = n1734 & ~n2479;
  assign n8491 = P1_DATAO_REG_25_ & ~n1734;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = ~P2_STATE_REG & ~n8492;
  assign n8494 = ~n8488 & ~n8489;
  assign n1460 = n8493 | ~n8494;
  assign n8496 = P2_IR_REG_26_ & ~n8485;
  assign n8497 = ~P2_IR_REG_25_ & ~P2_IR_REG_26_;
  assign n8498 = n8475 & n8497;
  assign n8499 = ~n8496 & ~n8498;
  assign n8500 = n8186 & n8499;
  assign n8501 = P2_IR_REG_26_ & n8185;
  assign n8502 = n1734 & ~n2522;
  assign n8503 = P1_DATAO_REG_26_ & ~n1734;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = ~P2_STATE_REG & ~n8504;
  assign n8506 = ~n8500 & ~n8501;
  assign n1465 = n8505 | ~n8506;
  assign n8508 = ~P2_IR_REG_27_ & n8498;
  assign n8509 = P2_IR_REG_27_ & ~n8498;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = n8186 & n8510;
  assign n8512 = P2_IR_REG_27_ & n8185;
  assign n8513 = n1734 & ~n2546;
  assign n8514 = P1_DATAO_REG_27_ & ~n1734;
  assign n8515 = ~n8513 & ~n8514;
  assign n8516 = ~P2_STATE_REG & ~n8515;
  assign n8517 = ~n8511 & ~n8512;
  assign n1470 = n8516 | ~n8517;
  assign n8519 = P2_IR_REG_27_ & P2_IR_REG_28_;
  assign n8520 = ~P2_IR_REG_27_ & n8497;
  assign n8521 = ~P2_IR_REG_28_ & n8520;
  assign n8522 = n8475 & n8521;
  assign n8523 = ~n8519 & ~n8522;
  assign n8524 = P2_IR_REG_28_ & ~n8498;
  assign n8525 = n8523 & ~n8524;
  assign n8526 = n8186 & n8525;
  assign n8527 = P2_IR_REG_28_ & n8185;
  assign n8528 = n1734 & ~n2591;
  assign n8529 = P1_DATAO_REG_28_ & ~n1734;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = ~P2_STATE_REG & ~n8530;
  assign n8532 = ~n8526 & ~n8527;
  assign n1475 = n8531 | ~n8532;
  assign n8534 = P2_IR_REG_29_ & ~n8522;
  assign n8535 = ~P2_IR_REG_29_ & n8522;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = n8186 & n8536;
  assign n8538 = P2_IR_REG_29_ & n8185;
  assign n8539 = n1734 & ~n2620;
  assign n8540 = P1_DATAO_REG_29_ & ~n1734;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = ~P2_STATE_REG & ~n8541;
  assign n8543 = ~n8537 & ~n8538;
  assign n1480 = n8542 | ~n8543;
  assign n8545 = ~P2_IR_REG_30_ & n8535;
  assign n8546 = P2_IR_REG_30_ & ~n8535;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n8186 & n8547;
  assign n8549 = P2_IR_REG_30_ & n8185;
  assign n8550 = n1734 & ~n2644;
  assign n8551 = P1_DATAO_REG_30_ & ~n1734;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = ~P2_STATE_REG & ~n8552;
  assign n8554 = ~n8548 & ~n8549;
  assign n1485 = n8553 | ~n8554;
  assign n8556 = P2_IR_REG_31_ & n8545;
  assign n8557 = ~P2_IR_REG_31_ & ~n8545;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = n8186 & ~n8558;
  assign n8560 = P2_IR_REG_31_ & n8185;
  assign n8561 = n1734 & n2675;
  assign n8562 = P1_DATAO_REG_31_ & ~n1734;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = ~P2_STATE_REG & ~n8563;
  assign n8565 = ~n8559 & ~n8560;
  assign n1490 = n8564 | ~n8565;
  assign n8567 = P2_IR_REG_31_ & n8461;
  assign n8568 = P2_IR_REG_23_ & ~P2_IR_REG_31_;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = P2_IR_REG_31_ & n8487;
  assign n8571 = P2_IR_REG_25_ & ~P2_IR_REG_31_;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = P2_IR_REG_31_ & n8499;
  assign n8574 = P2_IR_REG_26_ & ~P2_IR_REG_31_;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = P2_IR_REG_31_ & n8476;
  assign n8577 = P2_IR_REG_24_ & ~P2_IR_REG_31_;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n8572 & ~n8575;
  assign n8580 = ~n8578 & n8579;
  assign n8581 = n8569 & ~n8580;
  assign n8582 = P2_STATE_REG & n8581;
  assign n8583 = n8572 & ~n8575;
  assign n8584 = ~P2_B_REG & ~n8578;
  assign n8585 = P2_B_REG & n8578;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = n8583 & ~n8586;
  assign n8588 = ~n8575 & ~n8587;
  assign n8589 = n8582 & ~n8588;
  assign n8590 = n8578 & ~n8583;
  assign n8591 = n8589 & ~n8590;
  assign n8592 = P2_D_REG_0_ & ~n8589;
  assign n1495 = n8591 | n8592;
  assign n8594 = n8572 & ~n8583;
  assign n8595 = n8589 & ~n8594;
  assign n8596 = P2_D_REG_1_ & ~n8589;
  assign n1500 = n8595 | n8596;
  assign n1505 = P2_D_REG_2_ & ~n8589;
  assign n1510 = P2_D_REG_3_ & ~n8589;
  assign n1515 = P2_D_REG_4_ & ~n8589;
  assign n1520 = P2_D_REG_5_ & ~n8589;
  assign n1525 = P2_D_REG_6_ & ~n8589;
  assign n1530 = P2_D_REG_7_ & ~n8589;
  assign n1535 = P2_D_REG_8_ & ~n8589;
  assign n1540 = P2_D_REG_9_ & ~n8589;
  assign n1545 = P2_D_REG_10_ & ~n8589;
  assign n1550 = P2_D_REG_11_ & ~n8589;
  assign n1555 = P2_D_REG_12_ & ~n8589;
  assign n1560 = P2_D_REG_13_ & ~n8589;
  assign n1565 = P2_D_REG_14_ & ~n8589;
  assign n1570 = P2_D_REG_15_ & ~n8589;
  assign n1575 = P2_D_REG_16_ & ~n8589;
  assign n1580 = P2_D_REG_17_ & ~n8589;
  assign n1585 = P2_D_REG_18_ & ~n8589;
  assign n1590 = P2_D_REG_19_ & ~n8589;
  assign n1595 = P2_D_REG_20_ & ~n8589;
  assign n1600 = P2_D_REG_21_ & ~n8589;
  assign n1605 = P2_D_REG_22_ & ~n8589;
  assign n1610 = P2_D_REG_23_ & ~n8589;
  assign n1615 = P2_D_REG_24_ & ~n8589;
  assign n1620 = P2_D_REG_25_ & ~n8589;
  assign n1625 = P2_D_REG_26_ & ~n8589;
  assign n1630 = P2_D_REG_27_ & ~n8589;
  assign n1635 = P2_D_REG_28_ & ~n8589;
  assign n1640 = P2_D_REG_29_ & ~n8589;
  assign n1645 = P2_D_REG_30_ & ~n8589;
  assign n1650 = P2_D_REG_31_ & ~n8589;
  assign n8628 = ~n8588 & ~n8594;
  assign n8629 = P2_D_REG_1_ & n8588;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = P2_D_REG_0_ & n8588;
  assign n8632 = n8575 & n8578;
  assign n8633 = ~n8588 & ~n8632;
  assign n8634 = ~n8631 & ~n8633;
  assign n8635 = n8630 & n8634;
  assign n8636 = P2_D_REG_8_ & n8588;
  assign n8637 = P2_D_REG_7_ & n8588;
  assign n8638 = P2_D_REG_9_ & n8588;
  assign n8639 = ~n8636 & ~n8637;
  assign n8640 = ~n8638 & n8639;
  assign n8641 = P2_D_REG_6_ & n8588;
  assign n8642 = P2_D_REG_5_ & n8588;
  assign n8643 = P2_D_REG_4_ & n8588;
  assign n8644 = P2_D_REG_3_ & n8588;
  assign n8645 = ~n8641 & ~n8642;
  assign n8646 = ~n8643 & n8645;
  assign n8647 = ~n8644 & n8646;
  assign n8648 = P2_D_REG_31_ & n8588;
  assign n8649 = P2_D_REG_30_ & n8588;
  assign n8650 = P2_D_REG_2_ & n8588;
  assign n8651 = P2_D_REG_29_ & n8588;
  assign n8652 = ~n8648 & ~n8649;
  assign n8653 = ~n8650 & n8652;
  assign n8654 = ~n8651 & n8653;
  assign n8655 = P2_D_REG_28_ & n8588;
  assign n8656 = P2_D_REG_27_ & n8588;
  assign n8657 = P2_D_REG_26_ & n8588;
  assign n8658 = P2_D_REG_25_ & n8588;
  assign n8659 = ~n8655 & ~n8656;
  assign n8660 = ~n8657 & n8659;
  assign n8661 = ~n8658 & n8660;
  assign n8662 = n8640 & n8647;
  assign n8663 = n8654 & n8662;
  assign n8664 = n8661 & n8663;
  assign n8665 = P2_D_REG_23_ & n8588;
  assign n8666 = P2_D_REG_22_ & n8588;
  assign n8667 = P2_D_REG_24_ & n8588;
  assign n8668 = ~n8665 & ~n8666;
  assign n8669 = ~n8667 & n8668;
  assign n8670 = P2_D_REG_21_ & n8588;
  assign n8671 = P2_D_REG_20_ & n8588;
  assign n8672 = P2_D_REG_19_ & n8588;
  assign n8673 = P2_D_REG_18_ & n8588;
  assign n8674 = ~n8670 & ~n8671;
  assign n8675 = ~n8672 & n8674;
  assign n8676 = ~n8673 & n8675;
  assign n8677 = P2_D_REG_17_ & n8588;
  assign n8678 = P2_D_REG_16_ & n8588;
  assign n8679 = P2_D_REG_15_ & n8588;
  assign n8680 = P2_D_REG_14_ & n8588;
  assign n8681 = ~n8677 & ~n8678;
  assign n8682 = ~n8679 & n8681;
  assign n8683 = ~n8680 & n8682;
  assign n8684 = P2_D_REG_13_ & n8588;
  assign n8685 = P2_D_REG_12_ & n8588;
  assign n8686 = P2_D_REG_11_ & n8588;
  assign n8687 = P2_D_REG_10_ & n8588;
  assign n8688 = ~n8684 & ~n8685;
  assign n8689 = ~n8686 & n8688;
  assign n8690 = ~n8687 & n8689;
  assign n8691 = n8669 & n8676;
  assign n8692 = n8683 & n8691;
  assign n8693 = n8690 & n8692;
  assign n8694 = n8664 & n8693;
  assign n8695 = n8635 & n8694;
  assign n8696 = P2_IR_REG_31_ & n8450;
  assign n8697 = P2_IR_REG_22_ & ~P2_IR_REG_31_;
  assign n8698 = ~n8696 & ~n8697;
  assign n8699 = P2_IR_REG_31_ & n8438;
  assign n8700 = P2_IR_REG_21_ & ~P2_IR_REG_31_;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = P2_IR_REG_31_ & n8427;
  assign n8703 = P2_IR_REG_20_ & ~P2_IR_REG_31_;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8701 & n8704;
  assign n8706 = ~n8698 & ~n8705;
  assign n8707 = n8698 & n8705;
  assign n8708 = ~n8706 & ~n8707;
  assign n8709 = P2_IR_REG_31_ & n8413;
  assign n8710 = P2_IR_REG_19_ & ~P2_IR_REG_31_;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = n8701 & n8711;
  assign n8713 = ~n8708 & ~n8712;
  assign n8714 = n8695 & ~n8713;
  assign n8715 = ~n8630 & ~n8634;
  assign n8716 = n8694 & n8715;
  assign n8717 = ~n8698 & ~n8711;
  assign n8718 = n8701 & n8717;
  assign n8719 = ~n8704 & n8718;
  assign n8720 = ~n8698 & n8711;
  assign n8721 = n8704 & n8720;
  assign n8722 = ~n8701 & n8721;
  assign n8723 = ~n8719 & ~n8722;
  assign n8724 = n8716 & ~n8723;
  assign n8725 = ~n8714 & ~n8724;
  assign n8726 = n8582 & ~n8725;
  assign n8727 = P2_IR_REG_31_ & n8510;
  assign n8728 = P2_IR_REG_27_ & ~P2_IR_REG_31_;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = P2_IR_REG_31_ & n8525;
  assign n8731 = P2_IR_REG_28_ & ~P2_IR_REG_31_;
  assign n8732 = ~n8730 & ~n8731;
  assign n8733 = n8729 & n8732;
  assign n8734 = P2_IR_REG_0_ & P2_IR_REG_31_;
  assign n8735 = P2_IR_REG_0_ & ~P2_IR_REG_31_;
  assign n8736 = ~n8734 & ~n8735;
  assign n8737 = n8733 & ~n8736;
  assign n8738 = ~n8191 & ~n8733;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = n8698 & n8711;
  assign n8741 = n8701 & n8740;
  assign n8742 = n8698 & ~n8711;
  assign n8743 = n8701 & n8742;
  assign n8744 = ~n8741 & ~n8743;
  assign n8745 = ~n8739 & ~n8744;
  assign n8746 = P2_IR_REG_31_ & n8547;
  assign n8747 = P2_IR_REG_30_ & ~P2_IR_REG_31_;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = P2_IR_REG_31_ & n8536;
  assign n8750 = P2_IR_REG_29_ & ~P2_IR_REG_31_;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8748 & ~n8751;
  assign n8753 = P2_REG3_REG_0_ & n8752;
  assign n8754 = ~n8748 & n8751;
  assign n8755 = P2_REG2_REG_0_ & n8754;
  assign n8756 = n8748 & ~n8751;
  assign n8757 = P2_REG1_REG_0_ & n8756;
  assign n8758 = n8748 & n8751;
  assign n8759 = P2_REG0_REG_0_ & n8758;
  assign n8760 = ~n8753 & ~n8755;
  assign n8761 = ~n8757 & n8760;
  assign n8762 = ~n8759 & n8761;
  assign n8763 = ~n8739 & n8762;
  assign n8764 = n8739 & ~n8762;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = n8704 & n8742;
  assign n8767 = ~n8765 & n8766;
  assign n8768 = ~n8698 & ~n8701;
  assign n8769 = ~n8729 & ~n8732;
  assign n8770 = ~n8733 & ~n8769;
  assign n8771 = n8768 & ~n8770;
  assign n8772 = P2_REG3_REG_1_ & n8752;
  assign n8773 = P2_REG2_REG_1_ & n8754;
  assign n8774 = P2_REG1_REG_1_ & n8756;
  assign n8775 = P2_REG0_REG_1_ & n8758;
  assign n8776 = ~n8772 & ~n8773;
  assign n8777 = ~n8774 & n8776;
  assign n8778 = ~n8775 & n8777;
  assign n8779 = n8771 & ~n8778;
  assign n8780 = ~n8745 & ~n8767;
  assign n8781 = ~n8779 & n8780;
  assign n8782 = n8701 & n8720;
  assign n8783 = n8704 & n8782;
  assign n8784 = ~n8765 & n8783;
  assign n8785 = ~n8701 & n8711;
  assign n8786 = ~n8704 & n8785;
  assign n8787 = ~n8765 & n8786;
  assign n8788 = ~n8701 & n8740;
  assign n8789 = n8704 & n8788;
  assign n8790 = ~n8765 & n8789;
  assign n8791 = ~n8701 & ~n8711;
  assign n8792 = ~n8704 & n8791;
  assign n8793 = ~n8765 & n8792;
  assign n8794 = ~n8704 & n8720;
  assign n8795 = ~n8765 & n8794;
  assign n8796 = ~n8793 & ~n8795;
  assign n8797 = ~n8704 & n8717;
  assign n8798 = ~n8765 & n8797;
  assign n8799 = n8704 & n8717;
  assign n8800 = ~n8765 & n8799;
  assign n8801 = ~n8798 & ~n8800;
  assign n8802 = ~n8784 & ~n8787;
  assign n8803 = ~n8790 & n8802;
  assign n8804 = n8796 & n8803;
  assign n8805 = n8801 & n8804;
  assign n8806 = n8781 & n8805;
  assign n8807 = n8726 & ~n8806;
  assign n8808 = P2_REG0_REG_0_ & ~n8726;
  assign n1655 = n8807 | n8808;
  assign n8810 = P2_REG3_REG_2_ & n8752;
  assign n8811 = P2_REG2_REG_2_ & n8754;
  assign n8812 = P2_REG1_REG_2_ & n8756;
  assign n8813 = P2_REG0_REG_2_ & n8758;
  assign n8814 = ~n8810 & ~n8811;
  assign n8815 = ~n8812 & n8814;
  assign n8816 = ~n8813 & n8815;
  assign n8817 = n8771 & ~n8816;
  assign n8818 = P2_IR_REG_31_ & ~n8197;
  assign n8819 = P2_IR_REG_1_ & ~P2_IR_REG_31_;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = n8733 & ~n8820;
  assign n8822 = ~n8202 & ~n8733;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = ~n8744 & ~n8823;
  assign n8825 = ~n8778 & n8823;
  assign n8826 = n8778 & ~n8823;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = ~n8763 & ~n8827;
  assign n8829 = n8763 & n8827;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = n8766 & ~n8830;
  assign n8832 = ~n8817 & ~n8824;
  assign n8833 = ~n8831 & n8832;
  assign n8834 = ~n8778 & ~n8823;
  assign n8835 = n8778 & n8823;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = ~n8739 & ~n8762;
  assign n8838 = n8836 & ~n8837;
  assign n8839 = ~n8836 & n8837;
  assign n8840 = ~n8838 & ~n8839;
  assign n8841 = n8799 & ~n8840;
  assign n8842 = ~n8729 & n8732;
  assign n8843 = n8729 & ~n8732;
  assign n8844 = ~n8842 & ~n8843;
  assign n8845 = n8768 & ~n8844;
  assign n8846 = ~n8762 & n8845;
  assign n8847 = n8794 & ~n8830;
  assign n8848 = n8797 & ~n8840;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = n8789 & ~n8830;
  assign n8851 = n8783 & ~n8830;
  assign n8852 = n8786 & ~n8840;
  assign n8853 = n8792 & ~n8840;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = ~n8850 & ~n8851;
  assign n8856 = n8854 & n8855;
  assign n8857 = ~n8841 & ~n8846;
  assign n8858 = n8849 & n8857;
  assign n8859 = n8856 & n8858;
  assign n8860 = n8833 & n8859;
  assign n8861 = n8726 & ~n8860;
  assign n8862 = P2_REG0_REG_1_ & ~n8726;
  assign n1660 = n8861 | n8862;
  assign n8864 = ~P2_REG3_REG_3_ & n8752;
  assign n8865 = P2_REG2_REG_3_ & n8754;
  assign n8866 = P2_REG1_REG_3_ & n8756;
  assign n8867 = P2_REG0_REG_3_ & n8758;
  assign n8868 = ~n8864 & ~n8865;
  assign n8869 = ~n8866 & n8868;
  assign n8870 = ~n8867 & n8869;
  assign n8871 = n8771 & ~n8870;
  assign n8872 = P2_IR_REG_31_ & n8209;
  assign n8873 = P2_IR_REG_2_ & ~P2_IR_REG_31_;
  assign n8874 = ~n8872 & ~n8873;
  assign n8875 = n8733 & ~n8874;
  assign n8876 = ~n8214 & ~n8733;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~n8744 & ~n8877;
  assign n8879 = ~n8816 & n8877;
  assign n8880 = n8816 & ~n8877;
  assign n8881 = ~n8879 & ~n8880;
  assign n8882 = ~n8763 & ~n8778;
  assign n8883 = ~n8763 & n8823;
  assign n8884 = ~n8882 & ~n8883;
  assign n8885 = ~n8825 & n8884;
  assign n8886 = n8881 & n8885;
  assign n8887 = ~n8881 & ~n8885;
  assign n8888 = ~n8886 & ~n8887;
  assign n8889 = n8766 & ~n8888;
  assign n8890 = ~n8871 & ~n8878;
  assign n8891 = ~n8889 & n8890;
  assign n8892 = ~n8816 & ~n8877;
  assign n8893 = n8816 & n8877;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 = ~n8835 & n8837;
  assign n8896 = ~n8834 & ~n8895;
  assign n8897 = n8894 & ~n8896;
  assign n8898 = ~n8834 & n8881;
  assign n8899 = ~n8895 & n8898;
  assign n8900 = ~n8897 & ~n8899;
  assign n8901 = n8799 & n8900;
  assign n8902 = ~n8778 & n8845;
  assign n8903 = n8794 & ~n8888;
  assign n8904 = n8797 & n8900;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = n8789 & ~n8888;
  assign n8907 = n8783 & ~n8888;
  assign n8908 = n8786 & n8900;
  assign n8909 = n8792 & n8900;
  assign n8910 = ~n8908 & ~n8909;
  assign n8911 = ~n8906 & ~n8907;
  assign n8912 = n8910 & n8911;
  assign n8913 = ~n8901 & ~n8902;
  assign n8914 = n8905 & n8913;
  assign n8915 = n8912 & n8914;
  assign n8916 = n8891 & n8915;
  assign n8917 = n8726 & ~n8916;
  assign n8918 = P2_REG0_REG_2_ & ~n8726;
  assign n1665 = n8917 | n8918;
  assign n8920 = ~P2_REG3_REG_4_ & ~P2_REG3_REG_3_;
  assign n8921 = P2_REG3_REG_4_ & P2_REG3_REG_3_;
  assign n8922 = ~n8920 & ~n8921;
  assign n8923 = n8752 & ~n8922;
  assign n8924 = P2_REG2_REG_4_ & n8754;
  assign n8925 = P2_REG1_REG_4_ & n8756;
  assign n8926 = P2_REG0_REG_4_ & n8758;
  assign n8927 = ~n8923 & ~n8924;
  assign n8928 = ~n8925 & n8927;
  assign n8929 = ~n8926 & n8928;
  assign n8930 = n8771 & ~n8929;
  assign n8931 = P2_IR_REG_31_ & n8220;
  assign n8932 = P2_IR_REG_3_ & ~P2_IR_REG_31_;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = n8733 & ~n8933;
  assign n8935 = ~n8225 & ~n8733;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8744 & ~n8936;
  assign n8938 = ~n8870 & n8936;
  assign n8939 = n8870 & ~n8936;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = ~n8880 & ~n8940;
  assign n8942 = ~n8879 & n8885;
  assign n8943 = n8941 & ~n8942;
  assign n8944 = ~n8879 & n8940;
  assign n8945 = ~n8880 & ~n8885;
  assign n8946 = n8944 & ~n8945;
  assign n8947 = ~n8943 & ~n8946;
  assign n8948 = n8766 & ~n8947;
  assign n8949 = ~n8930 & ~n8937;
  assign n8950 = ~n8948 & n8949;
  assign n8951 = n8834 & ~n8893;
  assign n8952 = ~n8892 & ~n8951;
  assign n8953 = ~n8893 & n8895;
  assign n8954 = n8952 & ~n8953;
  assign n8955 = ~n8940 & n8954;
  assign n8956 = ~n8870 & ~n8936;
  assign n8957 = n8870 & n8936;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n8954 & ~n8958;
  assign n8960 = ~n8955 & ~n8959;
  assign n8961 = n8799 & ~n8960;
  assign n8962 = ~n8816 & n8845;
  assign n8963 = n8794 & ~n8947;
  assign n8964 = n8797 & ~n8960;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = n8789 & ~n8947;
  assign n8967 = n8783 & ~n8947;
  assign n8968 = n8786 & ~n8960;
  assign n8969 = n8792 & ~n8960;
  assign n8970 = ~n8968 & ~n8969;
  assign n8971 = ~n8966 & ~n8967;
  assign n8972 = n8970 & n8971;
  assign n8973 = ~n8961 & ~n8962;
  assign n8974 = n8965 & n8973;
  assign n8975 = n8972 & n8974;
  assign n8976 = n8950 & n8975;
  assign n8977 = n8726 & ~n8976;
  assign n8978 = P2_REG0_REG_3_ & ~n8726;
  assign n1670 = n8977 | n8978;
  assign n8980 = ~P2_REG3_REG_5_ & n8920;
  assign n8981 = P2_REG3_REG_5_ & ~n8920;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = n8752 & ~n8982;
  assign n8984 = P2_REG2_REG_5_ & n8754;
  assign n8985 = P2_REG1_REG_5_ & n8756;
  assign n8986 = P2_REG0_REG_5_ & n8758;
  assign n8987 = ~n8983 & ~n8984;
  assign n8988 = ~n8985 & n8987;
  assign n8989 = ~n8986 & n8988;
  assign n8990 = n8771 & ~n8989;
  assign n8991 = P2_IR_REG_31_ & n8231;
  assign n8992 = P2_IR_REG_4_ & ~P2_IR_REG_31_;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = n8733 & ~n8993;
  assign n8995 = ~n8236 & ~n8733;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = ~n8744 & ~n8996;
  assign n8998 = ~n8870 & n8879;
  assign n8999 = n8870 & ~n8879;
  assign n9000 = n8936 & ~n8999;
  assign n9001 = ~n8998 & ~n9000;
  assign n9002 = ~n8880 & ~n8939;
  assign n9003 = ~n8885 & n9002;
  assign n9004 = n9001 & ~n9003;
  assign n9005 = ~n8929 & n8996;
  assign n9006 = n8929 & ~n8996;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = n9004 & n9007;
  assign n9009 = ~n9004 & ~n9007;
  assign n9010 = ~n9008 & ~n9009;
  assign n9011 = n8766 & ~n9010;
  assign n9012 = ~n8990 & ~n8997;
  assign n9013 = ~n9011 & n9012;
  assign n9014 = ~n8893 & ~n8957;
  assign n9015 = n8895 & n9014;
  assign n9016 = ~n8956 & ~n9015;
  assign n9017 = ~n8952 & ~n8957;
  assign n9018 = n9016 & ~n9017;
  assign n9019 = ~n9007 & n9018;
  assign n9020 = n8929 & n8996;
  assign n9021 = ~n8929 & ~n8996;
  assign n9022 = ~n9020 & ~n9021;
  assign n9023 = ~n9018 & ~n9022;
  assign n9024 = ~n9019 & ~n9023;
  assign n9025 = n8799 & ~n9024;
  assign n9026 = n8845 & ~n8870;
  assign n9027 = n8794 & ~n9010;
  assign n9028 = n8797 & ~n9024;
  assign n9029 = ~n9027 & ~n9028;
  assign n9030 = n8789 & ~n9010;
  assign n9031 = n8783 & ~n9010;
  assign n9032 = n8786 & ~n9024;
  assign n9033 = n8792 & ~n9024;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = ~n9030 & ~n9031;
  assign n9036 = n9034 & n9035;
  assign n9037 = ~n9025 & ~n9026;
  assign n9038 = n9029 & n9037;
  assign n9039 = n9036 & n9038;
  assign n9040 = n9013 & n9039;
  assign n9041 = n8726 & ~n9040;
  assign n9042 = P2_REG0_REG_4_ & ~n8726;
  assign n1675 = n9041 | n9042;
  assign n9044 = ~P2_REG3_REG_6_ & ~P2_REG3_REG_5_;
  assign n9045 = ~P2_REG3_REG_4_ & n9044;
  assign n9046 = ~P2_REG3_REG_3_ & n9045;
  assign n9047 = P2_REG3_REG_6_ & ~n8980;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 = n8752 & ~n9048;
  assign n9050 = P2_REG2_REG_6_ & n8754;
  assign n9051 = P2_REG1_REG_6_ & n8756;
  assign n9052 = P2_REG0_REG_6_ & n8758;
  assign n9053 = ~n9049 & ~n9050;
  assign n9054 = ~n9051 & n9053;
  assign n9055 = ~n9052 & n9054;
  assign n9056 = n8771 & ~n9055;
  assign n9057 = P2_IR_REG_31_ & n8242;
  assign n9058 = P2_IR_REG_5_ & ~P2_IR_REG_31_;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = n8733 & ~n9059;
  assign n9061 = ~n8247 & ~n8733;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~n8744 & ~n9062;
  assign n9064 = ~n8989 & n9062;
  assign n9065 = n8989 & ~n9062;
  assign n9066 = ~n9064 & ~n9065;
  assign n9067 = ~n9004 & ~n9006;
  assign n9068 = ~n9005 & ~n9067;
  assign n9069 = n9066 & n9068;
  assign n9070 = ~n9066 & ~n9068;
  assign n9071 = ~n9069 & ~n9070;
  assign n9072 = n8766 & ~n9071;
  assign n9073 = ~n9056 & ~n9063;
  assign n9074 = ~n9072 & n9073;
  assign n9075 = ~n8989 & ~n9062;
  assign n9076 = n8989 & n9062;
  assign n9077 = ~n9020 & ~n9076;
  assign n9078 = ~n9075 & n9077;
  assign n9079 = n9018 & ~n9021;
  assign n9080 = n9078 & ~n9079;
  assign n9081 = ~n9021 & n9066;
  assign n9082 = ~n9018 & ~n9020;
  assign n9083 = n9081 & ~n9082;
  assign n9084 = ~n9080 & ~n9083;
  assign n9085 = n8799 & n9084;
  assign n9086 = n8845 & ~n8929;
  assign n9087 = n8794 & ~n9071;
  assign n9088 = n8797 & n9084;
  assign n9089 = ~n9087 & ~n9088;
  assign n9090 = n8789 & ~n9071;
  assign n9091 = n8783 & ~n9071;
  assign n9092 = n8786 & n9084;
  assign n9093 = n8792 & n9084;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = ~n9090 & ~n9091;
  assign n9096 = n9094 & n9095;
  assign n9097 = ~n9085 & ~n9086;
  assign n9098 = n9089 & n9097;
  assign n9099 = n9096 & n9098;
  assign n9100 = n9074 & n9099;
  assign n9101 = n8726 & ~n9100;
  assign n9102 = P2_REG0_REG_5_ & ~n8726;
  assign n1680 = n9101 | n9102;
  assign n9104 = ~P2_REG3_REG_6_ & n8980;
  assign n9105 = ~P2_REG3_REG_7_ & n9104;
  assign n9106 = P2_REG3_REG_7_ & ~n9046;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = n8752 & ~n9107;
  assign n9109 = P2_REG2_REG_7_ & n8754;
  assign n9110 = P2_REG1_REG_7_ & n8756;
  assign n9111 = P2_REG0_REG_7_ & n8758;
  assign n9112 = ~n9108 & ~n9109;
  assign n9113 = ~n9110 & n9112;
  assign n9114 = ~n9111 & n9113;
  assign n9115 = n8771 & ~n9114;
  assign n9116 = P2_IR_REG_31_ & n8254;
  assign n9117 = P2_IR_REG_6_ & ~P2_IR_REG_31_;
  assign n9118 = ~n9116 & ~n9117;
  assign n9119 = n8733 & ~n9118;
  assign n9120 = ~n8259 & ~n8733;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = ~n8744 & ~n9121;
  assign n9123 = ~n9055 & n9121;
  assign n9124 = n9055 & ~n9121;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = ~n9065 & ~n9125;
  assign n9127 = ~n9064 & n9068;
  assign n9128 = n9126 & ~n9127;
  assign n9129 = ~n9064 & ~n9123;
  assign n9130 = ~n9124 & n9129;
  assign n9131 = ~n9065 & ~n9068;
  assign n9132 = n9130 & ~n9131;
  assign n9133 = ~n9128 & ~n9132;
  assign n9134 = n8766 & ~n9133;
  assign n9135 = ~n9115 & ~n9122;
  assign n9136 = ~n9134 & n9135;
  assign n9137 = n9021 & ~n9062;
  assign n9138 = ~n9021 & n9062;
  assign n9139 = ~n8989 & ~n9138;
  assign n9140 = ~n9137 & ~n9139;
  assign n9141 = ~n8957 & n9077;
  assign n9142 = ~n8892 & ~n8956;
  assign n9143 = ~n8893 & ~n8896;
  assign n9144 = n9142 & ~n9143;
  assign n9145 = n9141 & ~n9144;
  assign n9146 = n9140 & ~n9145;
  assign n9147 = ~n9125 & n9146;
  assign n9148 = n9055 & n9121;
  assign n9149 = ~n9055 & ~n9121;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = ~n9146 & ~n9150;
  assign n9152 = ~n9147 & ~n9151;
  assign n9153 = n8799 & ~n9152;
  assign n9154 = n8845 & ~n8989;
  assign n9155 = n8794 & ~n9133;
  assign n9156 = n8797 & ~n9152;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = n8789 & ~n9133;
  assign n9159 = n8783 & ~n9133;
  assign n9160 = n8786 & ~n9152;
  assign n9161 = n8792 & ~n9152;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = ~n9158 & ~n9159;
  assign n9164 = n9162 & n9163;
  assign n9165 = ~n9153 & ~n9154;
  assign n9166 = n9157 & n9165;
  assign n9167 = n9164 & n9166;
  assign n9168 = n9136 & n9167;
  assign n9169 = n8726 & ~n9168;
  assign n9170 = P2_REG0_REG_6_ & ~n8726;
  assign n1685 = n9169 | n9170;
  assign n9172 = ~P2_REG3_REG_8_ & n9105;
  assign n9173 = P2_REG3_REG_8_ & ~n9105;
  assign n9174 = ~n9172 & ~n9173;
  assign n9175 = n8752 & ~n9174;
  assign n9176 = P2_REG2_REG_8_ & n8754;
  assign n9177 = P2_REG1_REG_8_ & n8756;
  assign n9178 = P2_REG0_REG_8_ & n8758;
  assign n9179 = ~n9175 & ~n9176;
  assign n9180 = ~n9177 & n9179;
  assign n9181 = ~n9178 & n9180;
  assign n9182 = n8771 & ~n9181;
  assign n9183 = P2_IR_REG_31_ & n8265;
  assign n9184 = P2_IR_REG_7_ & ~P2_IR_REG_31_;
  assign n9185 = ~n9183 & ~n9184;
  assign n9186 = n8733 & ~n9185;
  assign n9187 = ~n8270 & ~n8733;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = ~n8744 & ~n9188;
  assign n9190 = ~n9114 & n9188;
  assign n9191 = n9114 & ~n9188;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = n9005 & ~n9065;
  assign n9194 = n9129 & ~n9193;
  assign n9195 = ~n9124 & ~n9194;
  assign n9196 = ~n9065 & ~n9124;
  assign n9197 = ~n9006 & n9196;
  assign n9198 = ~n9004 & n9197;
  assign n9199 = ~n9195 & ~n9198;
  assign n9200 = n9192 & n9199;
  assign n9201 = ~n9192 & ~n9199;
  assign n9202 = ~n9200 & ~n9201;
  assign n9203 = n8766 & ~n9202;
  assign n9204 = ~n9182 & ~n9189;
  assign n9205 = ~n9203 & n9204;
  assign n9206 = ~n9114 & ~n9188;
  assign n9207 = n9114 & n9188;
  assign n9208 = ~n9148 & ~n9207;
  assign n9209 = ~n9206 & n9208;
  assign n9210 = n9146 & ~n9149;
  assign n9211 = n9209 & ~n9210;
  assign n9212 = ~n9149 & n9192;
  assign n9213 = ~n9146 & ~n9148;
  assign n9214 = n9212 & ~n9213;
  assign n9215 = ~n9211 & ~n9214;
  assign n9216 = n8799 & n9215;
  assign n9217 = n8845 & ~n9055;
  assign n9218 = n8794 & ~n9202;
  assign n9219 = n8797 & n9215;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = n8789 & ~n9202;
  assign n9222 = n8783 & ~n9202;
  assign n9223 = n8786 & n9215;
  assign n9224 = n8792 & n9215;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n9221 & ~n9222;
  assign n9227 = n9225 & n9226;
  assign n9228 = ~n9216 & ~n9217;
  assign n9229 = n9220 & n9228;
  assign n9230 = n9227 & n9229;
  assign n9231 = n9205 & n9230;
  assign n9232 = n8726 & ~n9231;
  assign n9233 = P2_REG0_REG_7_ & ~n8726;
  assign n1690 = n9232 | n9233;
  assign n9235 = ~P2_REG3_REG_9_ & ~P2_REG3_REG_8_;
  assign n9236 = n9105 & n9235;
  assign n9237 = P2_REG3_REG_9_ & ~n9172;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = n8752 & ~n9238;
  assign n9240 = P2_REG2_REG_9_ & n8754;
  assign n9241 = P2_REG1_REG_9_ & n8756;
  assign n9242 = P2_REG0_REG_9_ & n8758;
  assign n9243 = ~n9239 & ~n9240;
  assign n9244 = ~n9241 & n9243;
  assign n9245 = ~n9242 & n9244;
  assign n9246 = n8771 & ~n9245;
  assign n9247 = P2_IR_REG_31_ & n8282;
  assign n9248 = P2_IR_REG_8_ & ~P2_IR_REG_31_;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = n8733 & ~n9249;
  assign n9251 = ~n8287 & ~n8733;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = ~n8744 & ~n9252;
  assign n9254 = ~n9181 & n9252;
  assign n9255 = n9181 & ~n9252;
  assign n9256 = ~n9254 & ~n9255;
  assign n9257 = ~n9191 & ~n9256;
  assign n9258 = ~n9190 & n9199;
  assign n9259 = n9257 & ~n9258;
  assign n9260 = ~n9190 & n9256;
  assign n9261 = ~n9191 & ~n9199;
  assign n9262 = n9260 & ~n9261;
  assign n9263 = ~n9259 & ~n9262;
  assign n9264 = n8766 & ~n9263;
  assign n9265 = ~n9246 & ~n9253;
  assign n9266 = ~n9264 & n9265;
  assign n9267 = n9149 & ~n9188;
  assign n9268 = ~n9149 & n9188;
  assign n9269 = ~n9114 & ~n9268;
  assign n9270 = ~n9267 & ~n9269;
  assign n9271 = ~n9146 & n9208;
  assign n9272 = n9270 & ~n9271;
  assign n9273 = ~n9256 & n9272;
  assign n9274 = n9181 & n9252;
  assign n9275 = ~n9181 & ~n9252;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = ~n9272 & ~n9276;
  assign n9278 = ~n9273 & ~n9277;
  assign n9279 = n8799 & ~n9278;
  assign n9280 = n8845 & ~n9114;
  assign n9281 = n8797 & ~n9278;
  assign n9282 = n8794 & ~n9263;
  assign n9283 = n8789 & ~n9263;
  assign n9284 = n8783 & ~n9263;
  assign n9285 = n8786 & ~n9278;
  assign n9286 = n8792 & ~n9278;
  assign n9287 = ~n9285 & ~n9286;
  assign n9288 = ~n9283 & ~n9284;
  assign n9289 = n9287 & n9288;
  assign n9290 = ~n9279 & ~n9280;
  assign n9291 = ~n9281 & n9290;
  assign n9292 = ~n9282 & n9291;
  assign n9293 = n9289 & n9292;
  assign n9294 = n9266 & n9293;
  assign n9295 = n8726 & ~n9294;
  assign n9296 = P2_REG0_REG_8_ & ~n8726;
  assign n1695 = n9295 | n9296;
  assign n9298 = ~P2_REG3_REG_9_ & ~P2_REG3_REG_10_;
  assign n9299 = ~P2_REG3_REG_8_ & n9298;
  assign n9300 = n9105 & n9299;
  assign n9301 = P2_REG3_REG_10_ & ~n9236;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = n8752 & ~n9302;
  assign n9304 = P2_REG2_REG_10_ & n8754;
  assign n9305 = P2_REG1_REG_10_ & n8756;
  assign n9306 = P2_REG0_REG_10_ & n8758;
  assign n9307 = ~n9303 & ~n9304;
  assign n9308 = ~n9305 & n9307;
  assign n9309 = ~n9306 & n9308;
  assign n9310 = n8771 & ~n9309;
  assign n9311 = P2_IR_REG_31_ & n8293;
  assign n9312 = P2_IR_REG_9_ & ~P2_IR_REG_31_;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = n8733 & ~n9313;
  assign n9315 = ~n8298 & ~n8733;
  assign n9316 = ~n9314 & ~n9315;
  assign n9317 = ~n8744 & ~n9316;
  assign n9318 = ~n9191 & ~n9255;
  assign n9319 = n9195 & n9318;
  assign n9320 = n9181 & ~n9190;
  assign n9321 = n9252 & ~n9320;
  assign n9322 = ~n9181 & n9190;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = ~n9319 & n9323;
  assign n9325 = n9197 & n9318;
  assign n9326 = ~n9004 & n9325;
  assign n9327 = n9324 & ~n9326;
  assign n9328 = ~n9245 & n9316;
  assign n9329 = n9245 & ~n9316;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = n9327 & n9330;
  assign n9332 = ~n9327 & ~n9330;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = n8766 & ~n9333;
  assign n9335 = ~n9310 & ~n9317;
  assign n9336 = ~n9334 & n9335;
  assign n9337 = ~n9272 & ~n9274;
  assign n9338 = ~n9275 & ~n9337;
  assign n9339 = ~n9330 & n9338;
  assign n9340 = n9245 & n9316;
  assign n9341 = ~n9245 & ~n9316;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = ~n9338 & ~n9342;
  assign n9344 = ~n9339 & ~n9343;
  assign n9345 = n8799 & ~n9344;
  assign n9346 = n8845 & ~n9181;
  assign n9347 = n8797 & ~n9344;
  assign n9348 = n8794 & ~n9333;
  assign n9349 = n8789 & ~n9333;
  assign n9350 = n8783 & ~n9333;
  assign n9351 = n8786 & ~n9344;
  assign n9352 = n8792 & ~n9344;
  assign n9353 = ~n9351 & ~n9352;
  assign n9354 = ~n9349 & ~n9350;
  assign n9355 = n9353 & n9354;
  assign n9356 = ~n9345 & ~n9346;
  assign n9357 = ~n9347 & n9356;
  assign n9358 = ~n9348 & n9357;
  assign n9359 = n9355 & n9358;
  assign n9360 = n9336 & n9359;
  assign n9361 = n8726 & ~n9360;
  assign n9362 = P2_REG0_REG_9_ & ~n8726;
  assign n1700 = n9361 | n9362;
  assign n9364 = ~P2_REG3_REG_11_ & ~P2_REG3_REG_10_;
  assign n9365 = ~P2_REG3_REG_8_ & n9364;
  assign n9366 = ~P2_REG3_REG_9_ & n9365;
  assign n9367 = n9105 & n9366;
  assign n9368 = P2_REG3_REG_11_ & ~n9300;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = n8752 & ~n9369;
  assign n9371 = P2_REG2_REG_11_ & n8754;
  assign n9372 = P2_REG1_REG_11_ & n8756;
  assign n9373 = P2_REG0_REG_11_ & n8758;
  assign n9374 = ~n9370 & ~n9371;
  assign n9375 = ~n9372 & n9374;
  assign n9376 = ~n9373 & n9375;
  assign n9377 = n8771 & ~n9376;
  assign n9378 = P2_IR_REG_31_ & n8305;
  assign n9379 = P2_IR_REG_10_ & ~P2_IR_REG_31_;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = n8733 & ~n9380;
  assign n9382 = ~n8310 & ~n8733;
  assign n9383 = ~n9381 & ~n9382;
  assign n9384 = ~n8744 & ~n9383;
  assign n9385 = ~n9309 & n9383;
  assign n9386 = n9309 & ~n9383;
  assign n9387 = ~n9385 & ~n9386;
  assign n9388 = ~n9327 & ~n9329;
  assign n9389 = ~n9328 & ~n9388;
  assign n9390 = n9387 & n9389;
  assign n9391 = ~n9387 & ~n9389;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = n8766 & ~n9392;
  assign n9394 = ~n9377 & ~n9384;
  assign n9395 = ~n9393 & n9394;
  assign n9396 = ~n9309 & ~n9383;
  assign n9397 = n9309 & n9383;
  assign n9398 = ~n9340 & ~n9397;
  assign n9399 = ~n9396 & n9398;
  assign n9400 = n9338 & ~n9341;
  assign n9401 = n9399 & ~n9400;
  assign n9402 = ~n9341 & n9387;
  assign n9403 = ~n9338 & ~n9340;
  assign n9404 = n9402 & ~n9403;
  assign n9405 = ~n9401 & ~n9404;
  assign n9406 = n8799 & n9405;
  assign n9407 = n8845 & ~n9245;
  assign n9408 = n8797 & n9405;
  assign n9409 = n8794 & ~n9392;
  assign n9410 = n8789 & ~n9392;
  assign n9411 = n8783 & ~n9392;
  assign n9412 = n8786 & n9405;
  assign n9413 = n8792 & n9405;
  assign n9414 = ~n9412 & ~n9413;
  assign n9415 = ~n9410 & ~n9411;
  assign n9416 = n9414 & n9415;
  assign n9417 = ~n9406 & ~n9407;
  assign n9418 = ~n9408 & n9417;
  assign n9419 = ~n9409 & n9418;
  assign n9420 = n9416 & n9419;
  assign n9421 = n9395 & n9420;
  assign n9422 = n8726 & ~n9421;
  assign n9423 = P2_REG0_REG_10_ & ~n8726;
  assign n1705 = n9422 | n9423;
  assign n9425 = ~P2_REG3_REG_12_ & n9367;
  assign n9426 = P2_REG3_REG_12_ & ~n9367;
  assign n9427 = ~n9425 & ~n9426;
  assign n9428 = n8752 & ~n9427;
  assign n9429 = P2_REG2_REG_12_ & n8754;
  assign n9430 = P2_REG1_REG_12_ & n8756;
  assign n9431 = P2_REG0_REG_12_ & n8758;
  assign n9432 = ~n9428 & ~n9429;
  assign n9433 = ~n9430 & n9432;
  assign n9434 = ~n9431 & n9433;
  assign n9435 = n8771 & ~n9434;
  assign n9436 = P2_IR_REG_31_ & n8316;
  assign n9437 = P2_IR_REG_11_ & ~P2_IR_REG_31_;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = n8733 & ~n9438;
  assign n9440 = ~n8321 & ~n8733;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = ~n8744 & ~n9441;
  assign n9443 = ~n9376 & n9441;
  assign n9444 = n9376 & ~n9441;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n9386 & ~n9445;
  assign n9447 = ~n9385 & n9389;
  assign n9448 = n9446 & ~n9447;
  assign n9449 = ~n9385 & ~n9443;
  assign n9450 = ~n9444 & n9449;
  assign n9451 = ~n9386 & ~n9389;
  assign n9452 = n9450 & ~n9451;
  assign n9453 = ~n9448 & ~n9452;
  assign n9454 = n8766 & ~n9453;
  assign n9455 = ~n9435 & ~n9442;
  assign n9456 = ~n9454 & n9455;
  assign n9457 = n9275 & n9398;
  assign n9458 = ~n9341 & ~n9457;
  assign n9459 = ~n9397 & ~n9458;
  assign n9460 = ~n9396 & ~n9459;
  assign n9461 = ~n9274 & n9398;
  assign n9462 = ~n9272 & n9461;
  assign n9463 = n9460 & ~n9462;
  assign n9464 = ~n9445 & n9463;
  assign n9465 = n9376 & n9441;
  assign n9466 = ~n9376 & ~n9441;
  assign n9467 = ~n9465 & ~n9466;
  assign n9468 = ~n9463 & ~n9467;
  assign n9469 = ~n9464 & ~n9468;
  assign n9470 = n8799 & ~n9469;
  assign n9471 = n8845 & ~n9309;
  assign n9472 = n8797 & ~n9469;
  assign n9473 = n8794 & ~n9453;
  assign n9474 = n8789 & ~n9453;
  assign n9475 = n8783 & ~n9453;
  assign n9476 = n8786 & ~n9469;
  assign n9477 = n8792 & ~n9469;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = ~n9474 & ~n9475;
  assign n9480 = n9478 & n9479;
  assign n9481 = ~n9470 & ~n9471;
  assign n9482 = ~n9472 & n9481;
  assign n9483 = ~n9473 & n9482;
  assign n9484 = n9480 & n9483;
  assign n9485 = n9456 & n9484;
  assign n9486 = n8726 & ~n9485;
  assign n9487 = P2_REG0_REG_11_ & ~n8726;
  assign n1710 = n9486 | n9487;
  assign n9489 = ~P2_REG3_REG_13_ & ~P2_REG3_REG_12_;
  assign n9490 = n9367 & n9489;
  assign n9491 = P2_REG3_REG_13_ & ~n9425;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = n8752 & ~n9492;
  assign n9494 = P2_REG2_REG_13_ & n8754;
  assign n9495 = P2_REG1_REG_13_ & n8756;
  assign n9496 = P2_REG0_REG_13_ & n8758;
  assign n9497 = ~n9493 & ~n9494;
  assign n9498 = ~n9495 & n9497;
  assign n9499 = ~n9496 & n9498;
  assign n9500 = n8771 & ~n9499;
  assign n9501 = P2_IR_REG_31_ & n8330;
  assign n9502 = P2_IR_REG_12_ & ~P2_IR_REG_31_;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = n8733 & ~n9503;
  assign n9505 = ~n8335 & ~n8733;
  assign n9506 = ~n9504 & ~n9505;
  assign n9507 = ~n8744 & ~n9506;
  assign n9508 = ~n9434 & n9506;
  assign n9509 = n9434 & ~n9506;
  assign n9510 = ~n9508 & ~n9509;
  assign n9511 = ~n9329 & ~n9386;
  assign n9512 = ~n9444 & n9511;
  assign n9513 = ~n9327 & n9512;
  assign n9514 = n9328 & ~n9386;
  assign n9515 = n9449 & ~n9514;
  assign n9516 = ~n9444 & ~n9515;
  assign n9517 = ~n9513 & ~n9516;
  assign n9518 = ~n9510 & ~n9517;
  assign n9519 = n9510 & n9517;
  assign n9520 = ~n9518 & ~n9519;
  assign n9521 = n8766 & ~n9520;
  assign n9522 = ~n9500 & ~n9507;
  assign n9523 = ~n9521 & n9522;
  assign n9524 = ~n9463 & ~n9465;
  assign n9525 = ~n9466 & ~n9524;
  assign n9526 = ~n9510 & n9525;
  assign n9527 = n9434 & n9506;
  assign n9528 = ~n9434 & ~n9506;
  assign n9529 = ~n9527 & ~n9528;
  assign n9530 = ~n9525 & ~n9529;
  assign n9531 = ~n9526 & ~n9530;
  assign n9532 = n8799 & ~n9531;
  assign n9533 = n8845 & ~n9376;
  assign n9534 = n8794 & ~n9520;
  assign n9535 = n8797 & ~n9531;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = n8789 & ~n9520;
  assign n9538 = n8783 & ~n9520;
  assign n9539 = n8786 & ~n9531;
  assign n9540 = n8792 & ~n9531;
  assign n9541 = ~n9539 & ~n9540;
  assign n9542 = ~n9537 & ~n9538;
  assign n9543 = n9541 & n9542;
  assign n9544 = ~n9532 & ~n9533;
  assign n9545 = n9536 & n9544;
  assign n9546 = n9543 & n9545;
  assign n9547 = n9523 & n9546;
  assign n9548 = n8726 & ~n9547;
  assign n9549 = P2_REG0_REG_12_ & ~n8726;
  assign n1715 = n9548 | n9549;
  assign n9551 = ~P2_REG3_REG_14_ & n9490;
  assign n9552 = P2_REG3_REG_14_ & ~n9490;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = n8752 & ~n9553;
  assign n9555 = P2_REG2_REG_14_ & n8754;
  assign n9556 = P2_REG1_REG_14_ & n8756;
  assign n9557 = P2_REG0_REG_14_ & n8758;
  assign n9558 = ~n9554 & ~n9555;
  assign n9559 = ~n9556 & n9558;
  assign n9560 = ~n9557 & n9559;
  assign n9561 = n8771 & ~n9560;
  assign n9562 = P2_IR_REG_31_ & n8341;
  assign n9563 = P2_IR_REG_13_ & ~P2_IR_REG_31_;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = n8733 & ~n9564;
  assign n9566 = ~n8346 & ~n8733;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = ~n8744 & ~n9567;
  assign n9569 = ~n9499 & n9567;
  assign n9570 = n9499 & ~n9567;
  assign n9571 = ~n9569 & ~n9570;
  assign n9572 = ~n9509 & n9516;
  assign n9573 = ~n9508 & ~n9572;
  assign n9574 = ~n9509 & n9512;
  assign n9575 = ~n9327 & n9574;
  assign n9576 = n9573 & ~n9575;
  assign n9577 = ~n9571 & ~n9576;
  assign n9578 = n9571 & n9576;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = n8766 & ~n9579;
  assign n9581 = ~n9561 & ~n9568;
  assign n9582 = ~n9580 & n9581;
  assign n9583 = ~n9499 & ~n9567;
  assign n9584 = n9499 & n9567;
  assign n9585 = ~n9527 & ~n9584;
  assign n9586 = ~n9583 & n9585;
  assign n9587 = n9525 & ~n9528;
  assign n9588 = n9586 & ~n9587;
  assign n9589 = ~n9528 & n9571;
  assign n9590 = ~n9525 & ~n9527;
  assign n9591 = n9589 & ~n9590;
  assign n9592 = ~n9588 & ~n9591;
  assign n9593 = n8799 & n9592;
  assign n9594 = n8845 & ~n9434;
  assign n9595 = n8794 & ~n9579;
  assign n9596 = n8797 & n9592;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = n8789 & ~n9579;
  assign n9599 = n8783 & ~n9579;
  assign n9600 = n8786 & n9592;
  assign n9601 = n8792 & n9592;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = ~n9598 & ~n9599;
  assign n9604 = n9602 & n9603;
  assign n9605 = ~n9593 & ~n9594;
  assign n9606 = n9597 & n9605;
  assign n9607 = n9604 & n9606;
  assign n9608 = n9582 & n9607;
  assign n9609 = n8726 & ~n9608;
  assign n9610 = P2_REG0_REG_13_ & ~n8726;
  assign n1720 = n9609 | n9610;
  assign n9612 = ~P2_REG3_REG_14_ & n9489;
  assign n9613 = ~P2_REG3_REG_15_ & n9612;
  assign n9614 = n9367 & n9613;
  assign n9615 = P2_REG3_REG_15_ & ~n9551;
  assign n9616 = ~n9614 & ~n9615;
  assign n9617 = n8752 & ~n9616;
  assign n9618 = P2_REG2_REG_15_ & n8754;
  assign n9619 = P2_REG1_REG_15_ & n8756;
  assign n9620 = P2_REG0_REG_15_ & n8758;
  assign n9621 = ~n9617 & ~n9618;
  assign n9622 = ~n9619 & n9621;
  assign n9623 = ~n9620 & n9622;
  assign n9624 = n8771 & ~n9623;
  assign n9625 = P2_IR_REG_31_ & n8353;
  assign n9626 = P2_IR_REG_14_ & ~P2_IR_REG_31_;
  assign n9627 = ~n9625 & ~n9626;
  assign n9628 = n8733 & ~n9627;
  assign n9629 = ~n8358 & ~n8733;
  assign n9630 = ~n9628 & ~n9629;
  assign n9631 = ~n8744 & ~n9630;
  assign n9632 = ~n9570 & ~n9576;
  assign n9633 = ~n9569 & ~n9632;
  assign n9634 = ~n9560 & n9630;
  assign n9635 = n9560 & ~n9630;
  assign n9636 = ~n9634 & ~n9635;
  assign n9637 = n9633 & n9636;
  assign n9638 = ~n9633 & ~n9636;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = n8766 & ~n9639;
  assign n9641 = ~n9624 & ~n9631;
  assign n9642 = ~n9640 & n9641;
  assign n9643 = n9466 & n9585;
  assign n9644 = ~n9528 & ~n9643;
  assign n9645 = ~n9584 & ~n9644;
  assign n9646 = ~n9583 & ~n9645;
  assign n9647 = ~n9465 & n9585;
  assign n9648 = ~n9463 & n9647;
  assign n9649 = n9646 & ~n9648;
  assign n9650 = ~n9636 & n9649;
  assign n9651 = n9636 & ~n9649;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = n8799 & ~n9652;
  assign n9654 = n8845 & ~n9499;
  assign n9655 = n8797 & ~n9652;
  assign n9656 = n8794 & ~n9639;
  assign n9657 = n8789 & ~n9639;
  assign n9658 = n8783 & ~n9639;
  assign n9659 = n8786 & ~n9652;
  assign n9660 = n8792 & ~n9652;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = ~n9657 & ~n9658;
  assign n9663 = n9661 & n9662;
  assign n9664 = ~n9653 & ~n9654;
  assign n9665 = ~n9655 & n9664;
  assign n9666 = ~n9656 & n9665;
  assign n9667 = n9663 & n9666;
  assign n9668 = n9642 & n9667;
  assign n9669 = n8726 & ~n9668;
  assign n9670 = P2_REG0_REG_14_ & ~n8726;
  assign n1725 = n9669 | n9670;
  assign n9672 = ~P2_REG3_REG_16_ & n9614;
  assign n9673 = P2_REG3_REG_16_ & ~n9614;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = n8752 & ~n9674;
  assign n9676 = P2_REG2_REG_16_ & n8754;
  assign n9677 = P2_REG1_REG_16_ & n8756;
  assign n9678 = P2_REG0_REG_16_ & n8758;
  assign n9679 = ~n9675 & ~n9676;
  assign n9680 = ~n9677 & n9679;
  assign n9681 = ~n9678 & n9680;
  assign n9682 = n8771 & ~n9681;
  assign n9683 = P2_IR_REG_31_ & n8364;
  assign n9684 = P2_IR_REG_15_ & ~P2_IR_REG_31_;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = n8733 & ~n9685;
  assign n9687 = ~n8369 & ~n8733;
  assign n9688 = ~n9686 & ~n9687;
  assign n9689 = ~n8744 & ~n9688;
  assign n9690 = ~n9623 & n9688;
  assign n9691 = n9623 & ~n9688;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = ~n9633 & ~n9635;
  assign n9694 = ~n9634 & ~n9693;
  assign n9695 = n9692 & n9694;
  assign n9696 = ~n9692 & ~n9694;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = n8766 & ~n9697;
  assign n9699 = ~n9682 & ~n9689;
  assign n9700 = ~n9698 & n9699;
  assign n9701 = ~n9560 & ~n9630;
  assign n9702 = n9560 & n9630;
  assign n9703 = ~n9649 & ~n9702;
  assign n9704 = ~n9701 & ~n9703;
  assign n9705 = ~n9692 & n9704;
  assign n9706 = n9692 & ~n9704;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = n8799 & ~n9707;
  assign n9709 = n8845 & ~n9560;
  assign n9710 = n8797 & ~n9707;
  assign n9711 = n8794 & ~n9697;
  assign n9712 = n8789 & ~n9697;
  assign n9713 = n8783 & ~n9697;
  assign n9714 = n8786 & ~n9707;
  assign n9715 = n8792 & ~n9707;
  assign n9716 = ~n9714 & ~n9715;
  assign n9717 = ~n9712 & ~n9713;
  assign n9718 = n9716 & n9717;
  assign n9719 = ~n9708 & ~n9709;
  assign n9720 = ~n9710 & n9719;
  assign n9721 = ~n9711 & n9720;
  assign n9722 = n9718 & n9721;
  assign n9723 = n9700 & n9722;
  assign n9724 = n8726 & ~n9723;
  assign n9725 = P2_REG0_REG_15_ & ~n8726;
  assign n1730 = n9724 | n9725;
  assign n9727 = ~P2_REG3_REG_17_ & ~P2_REG3_REG_16_;
  assign n9728 = n9614 & n9727;
  assign n9729 = P2_REG3_REG_17_ & ~n9672;
  assign n9730 = ~n9728 & ~n9729;
  assign n9731 = n8752 & ~n9730;
  assign n9732 = P2_REG2_REG_17_ & n8754;
  assign n9733 = P2_REG1_REG_17_ & n8756;
  assign n9734 = P2_REG0_REG_17_ & n8758;
  assign n9735 = ~n9731 & ~n9732;
  assign n9736 = ~n9733 & n9735;
  assign n9737 = ~n9734 & n9736;
  assign n9738 = n8771 & ~n9737;
  assign n9739 = P2_IR_REG_31_ & n8379;
  assign n9740 = P2_IR_REG_16_ & ~P2_IR_REG_31_;
  assign n9741 = ~n9739 & ~n9740;
  assign n9742 = n8733 & ~n9741;
  assign n9743 = ~n8384 & ~n8733;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = ~n8744 & ~n9744;
  assign n9746 = ~n9681 & n9744;
  assign n9747 = n9681 & ~n9744;
  assign n9748 = ~n9746 & ~n9747;
  assign n9749 = ~n9691 & ~n9748;
  assign n9750 = ~n9690 & n9694;
  assign n9751 = n9749 & ~n9750;
  assign n9752 = ~n9690 & ~n9746;
  assign n9753 = ~n9747 & n9752;
  assign n9754 = ~n9691 & ~n9694;
  assign n9755 = n9753 & ~n9754;
  assign n9756 = ~n9751 & ~n9755;
  assign n9757 = n8766 & ~n9756;
  assign n9758 = ~n9738 & ~n9745;
  assign n9759 = ~n9757 & n9758;
  assign n9760 = ~n9623 & ~n9688;
  assign n9761 = n9623 & n9688;
  assign n9762 = ~n9704 & ~n9761;
  assign n9763 = ~n9760 & ~n9762;
  assign n9764 = ~n9748 & n9763;
  assign n9765 = n9681 & n9744;
  assign n9766 = ~n9681 & ~n9744;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = ~n9763 & ~n9767;
  assign n9769 = ~n9764 & ~n9768;
  assign n9770 = n8799 & ~n9769;
  assign n9771 = n8845 & ~n9623;
  assign n9772 = n8797 & ~n9769;
  assign n9773 = n8794 & ~n9756;
  assign n9774 = n8789 & ~n9756;
  assign n9775 = n8783 & ~n9756;
  assign n9776 = n8786 & ~n9769;
  assign n9777 = n8792 & ~n9769;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~n9774 & ~n9775;
  assign n9780 = n9778 & n9779;
  assign n9781 = ~n9770 & ~n9771;
  assign n9782 = ~n9772 & n9781;
  assign n9783 = ~n9773 & n9782;
  assign n9784 = n9780 & n9783;
  assign n9785 = n9759 & n9784;
  assign n9786 = n8726 & ~n9785;
  assign n9787 = P2_REG0_REG_16_ & ~n8726;
  assign n1735 = n9786 | n9787;
  assign n9789 = ~P2_REG3_REG_18_ & n9728;
  assign n9790 = P2_REG3_REG_18_ & ~n9728;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = n8752 & ~n9791;
  assign n9793 = P2_REG2_REG_18_ & n8754;
  assign n9794 = P2_REG1_REG_18_ & n8756;
  assign n9795 = P2_REG0_REG_18_ & n8758;
  assign n9796 = ~n9792 & ~n9793;
  assign n9797 = ~n9794 & n9796;
  assign n9798 = ~n9795 & n9797;
  assign n9799 = n8771 & ~n9798;
  assign n9800 = P2_IR_REG_31_ & n8390;
  assign n9801 = P2_IR_REG_17_ & ~P2_IR_REG_31_;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = n8733 & ~n9802;
  assign n9804 = ~n8395 & ~n8733;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~n8744 & ~n9805;
  assign n9807 = ~n9737 & n9805;
  assign n9808 = n9737 & ~n9805;
  assign n9809 = ~n9807 & ~n9808;
  assign n9810 = ~n9691 & ~n9747;
  assign n9811 = n9634 & n9810;
  assign n9812 = n9752 & ~n9811;
  assign n9813 = ~n9747 & ~n9812;
  assign n9814 = ~n9635 & n9810;
  assign n9815 = ~n9633 & n9814;
  assign n9816 = ~n9813 & ~n9815;
  assign n9817 = ~n9809 & ~n9816;
  assign n9818 = n9809 & n9816;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = n8766 & ~n9819;
  assign n9821 = ~n9799 & ~n9806;
  assign n9822 = ~n9820 & n9821;
  assign n9823 = ~n9737 & ~n9805;
  assign n9824 = n9737 & n9805;
  assign n9825 = ~n9765 & ~n9824;
  assign n9826 = ~n9823 & n9825;
  assign n9827 = n9763 & ~n9766;
  assign n9828 = n9826 & ~n9827;
  assign n9829 = ~n9766 & n9809;
  assign n9830 = ~n9763 & ~n9765;
  assign n9831 = n9829 & ~n9830;
  assign n9832 = ~n9828 & ~n9831;
  assign n9833 = n8799 & n9832;
  assign n9834 = n8845 & ~n9681;
  assign n9835 = n8794 & ~n9819;
  assign n9836 = n8797 & n9832;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = n8789 & ~n9819;
  assign n9839 = n8783 & ~n9819;
  assign n9840 = n8786 & n9832;
  assign n9841 = n8792 & n9832;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = ~n9838 & ~n9839;
  assign n9844 = n9842 & n9843;
  assign n9845 = ~n9833 & ~n9834;
  assign n9846 = n9837 & n9845;
  assign n9847 = n9844 & n9846;
  assign n9848 = n9822 & n9847;
  assign n9849 = n8726 & ~n9848;
  assign n9850 = P2_REG0_REG_17_ & ~n8726;
  assign n1740 = n9849 | n9850;
  assign n9852 = ~P2_REG3_REG_18_ & ~P2_REG3_REG_19_;
  assign n9853 = n9728 & n9852;
  assign n9854 = P2_REG3_REG_19_ & ~n9789;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = n8752 & ~n9855;
  assign n9857 = P2_REG2_REG_19_ & n8754;
  assign n9858 = P2_REG1_REG_19_ & n8756;
  assign n9859 = P2_REG0_REG_19_ & n8758;
  assign n9860 = ~n9856 & ~n9857;
  assign n9861 = ~n9858 & n9860;
  assign n9862 = ~n9859 & n9861;
  assign n9863 = n8771 & ~n9862;
  assign n9864 = P2_IR_REG_31_ & n8402;
  assign n9865 = P2_IR_REG_18_ & ~P2_IR_REG_31_;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n8733 & ~n9866;
  assign n9868 = ~n8407 & ~n8733;
  assign n9869 = ~n9867 & ~n9868;
  assign n9870 = ~n8744 & ~n9869;
  assign n9871 = ~n9798 & n9869;
  assign n9872 = n9798 & ~n9869;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9808 & ~n9816;
  assign n9875 = ~n9807 & ~n9874;
  assign n9876 = ~n9873 & ~n9875;
  assign n9877 = n9873 & n9875;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = n8766 & ~n9878;
  assign n9880 = ~n9863 & ~n9870;
  assign n9881 = ~n9879 & n9880;
  assign n9882 = n9766 & ~n9805;
  assign n9883 = ~n9766 & n9805;
  assign n9884 = ~n9737 & ~n9883;
  assign n9885 = ~n9882 & ~n9884;
  assign n9886 = ~n9763 & n9825;
  assign n9887 = n9885 & ~n9886;
  assign n9888 = ~n9873 & n9887;
  assign n9889 = n9798 & n9869;
  assign n9890 = ~n9798 & ~n9869;
  assign n9891 = ~n9889 & ~n9890;
  assign n9892 = ~n9887 & ~n9891;
  assign n9893 = ~n9888 & ~n9892;
  assign n9894 = n8799 & ~n9893;
  assign n9895 = n8845 & ~n9737;
  assign n9896 = n8794 & ~n9878;
  assign n9897 = n8797 & ~n9893;
  assign n9898 = ~n9896 & ~n9897;
  assign n9899 = n8789 & ~n9878;
  assign n9900 = n8783 & ~n9878;
  assign n9901 = n8786 & ~n9893;
  assign n9902 = n8792 & ~n9893;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = ~n9899 & ~n9900;
  assign n9905 = n9903 & n9904;
  assign n9906 = ~n9894 & ~n9895;
  assign n9907 = n9898 & n9906;
  assign n9908 = n9905 & n9907;
  assign n9909 = n9881 & n9908;
  assign n9910 = n8726 & ~n9909;
  assign n9911 = P2_REG0_REG_18_ & ~n8726;
  assign n1745 = n9910 | n9911;
  assign n9913 = ~P2_REG3_REG_20_ & n9853;
  assign n9914 = P2_REG3_REG_20_ & ~n9853;
  assign n9915 = ~n9913 & ~n9914;
  assign n9916 = n8752 & ~n9915;
  assign n9917 = P2_REG0_REG_20_ & n8758;
  assign n9918 = P2_REG1_REG_20_ & n8756;
  assign n9919 = P2_REG2_REG_20_ & n8754;
  assign n9920 = ~n9916 & ~n9917;
  assign n9921 = ~n9918 & n9920;
  assign n9922 = ~n9919 & n9921;
  assign n9923 = n8771 & ~n9922;
  assign n9924 = ~n8711 & n8733;
  assign n9925 = ~n8418 & ~n8733;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = ~n8744 & ~n9926;
  assign n9928 = ~n9862 & n9926;
  assign n9929 = n9862 & ~n9926;
  assign n9930 = ~n9928 & ~n9929;
  assign n9931 = ~n9798 & ~n9875;
  assign n9932 = n9869 & ~n9875;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = ~n9871 & n9933;
  assign n9935 = ~n9930 & ~n9934;
  assign n9936 = n9930 & n9934;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = n8766 & ~n9937;
  assign n9939 = ~n9923 & ~n9927;
  assign n9940 = ~n9938 & n9939;
  assign n9941 = ~n9887 & ~n9889;
  assign n9942 = ~n9890 & ~n9941;
  assign n9943 = ~n9930 & n9942;
  assign n9944 = n9862 & n9926;
  assign n9945 = ~n9862 & ~n9926;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9942 & ~n9946;
  assign n9948 = ~n9943 & ~n9947;
  assign n9949 = n8799 & ~n9948;
  assign n9950 = n8845 & ~n9798;
  assign n9951 = n8794 & ~n9937;
  assign n9952 = n8797 & ~n9948;
  assign n9953 = ~n9951 & ~n9952;
  assign n9954 = n8789 & ~n9937;
  assign n9955 = n8783 & ~n9937;
  assign n9956 = n8786 & ~n9948;
  assign n9957 = n8792 & ~n9948;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = ~n9954 & ~n9955;
  assign n9960 = n9958 & n9959;
  assign n9961 = ~n9949 & ~n9950;
  assign n9962 = n9953 & n9961;
  assign n9963 = n9960 & n9962;
  assign n9964 = n9940 & n9963;
  assign n9965 = n8726 & ~n9964;
  assign n9966 = P2_REG0_REG_19_ & ~n8726;
  assign n1750 = n9965 | n9966;
  assign n9968 = ~P2_REG3_REG_20_ & ~P2_REG3_REG_21_;
  assign n9969 = n9853 & n9968;
  assign n9970 = P2_REG3_REG_21_ & ~n9913;
  assign n9971 = ~n9969 & ~n9970;
  assign n9972 = n8752 & ~n9971;
  assign n9973 = P2_REG0_REG_21_ & n8758;
  assign n9974 = P2_REG1_REG_21_ & n8756;
  assign n9975 = P2_REG2_REG_21_ & n8754;
  assign n9976 = ~n9972 & ~n9973;
  assign n9977 = ~n9974 & n9976;
  assign n9978 = ~n9975 & n9977;
  assign n9979 = n8771 & ~n9978;
  assign n9980 = ~n8432 & ~n8733;
  assign n9981 = ~n8744 & n9980;
  assign n9982 = ~n9922 & ~n9980;
  assign n9983 = n9922 & n9980;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9929 & ~n9934;
  assign n9986 = ~n9928 & ~n9985;
  assign n9987 = ~n9984 & ~n9986;
  assign n9988 = n9984 & n9986;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = n8766 & ~n9989;
  assign n9991 = ~n9979 & ~n9981;
  assign n9992 = ~n9990 & n9991;
  assign n9993 = ~n9922 & n9980;
  assign n9994 = n9922 & ~n9980;
  assign n9995 = ~n9944 & ~n9994;
  assign n9996 = ~n9993 & n9995;
  assign n9997 = n9942 & ~n9945;
  assign n9998 = n9996 & ~n9997;
  assign n9999 = ~n9945 & n9984;
  assign n10000 = ~n9942 & ~n9944;
  assign n10001 = n9999 & ~n10000;
  assign n10002 = ~n9998 & ~n10001;
  assign n10003 = n8799 & n10002;
  assign n10004 = n8845 & ~n9862;
  assign n10005 = n8794 & ~n9989;
  assign n10006 = n8797 & n10002;
  assign n10007 = ~n10005 & ~n10006;
  assign n10008 = n8789 & ~n9989;
  assign n10009 = n8783 & ~n9989;
  assign n10010 = n8786 & n10002;
  assign n10011 = n8792 & n10002;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = ~n10008 & ~n10009;
  assign n10014 = n10012 & n10013;
  assign n10015 = ~n10003 & ~n10004;
  assign n10016 = n10007 & n10015;
  assign n10017 = n10014 & n10016;
  assign n10018 = n9992 & n10017;
  assign n10019 = n8726 & ~n10018;
  assign n10020 = P2_REG0_REG_20_ & ~n8726;
  assign n1755 = n10019 | n10020;
  assign n10022 = ~P2_REG3_REG_22_ & n9969;
  assign n10023 = P2_REG3_REG_22_ & ~n9969;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n8752 & ~n10024;
  assign n10026 = P2_REG0_REG_22_ & n8758;
  assign n10027 = P2_REG1_REG_22_ & n8756;
  assign n10028 = P2_REG2_REG_22_ & n8754;
  assign n10029 = ~n10025 & ~n10026;
  assign n10030 = ~n10027 & n10029;
  assign n10031 = ~n10028 & n10030;
  assign n10032 = n8771 & ~n10031;
  assign n10033 = ~n8443 & ~n8733;
  assign n10034 = ~n8744 & n10033;
  assign n10035 = ~n9983 & ~n9986;
  assign n10036 = ~n9982 & ~n10035;
  assign n10037 = ~n9978 & ~n10033;
  assign n10038 = n9978 & n10033;
  assign n10039 = ~n10037 & ~n10038;
  assign n10040 = n10036 & n10039;
  assign n10041 = ~n10036 & ~n10039;
  assign n10042 = ~n10040 & ~n10041;
  assign n10043 = n8766 & ~n10042;
  assign n10044 = ~n10032 & ~n10034;
  assign n10045 = ~n10043 & n10044;
  assign n10046 = ~n9942 & n9995;
  assign n10047 = ~n9945 & ~n9980;
  assign n10048 = n9945 & n9980;
  assign n10049 = n9922 & ~n10048;
  assign n10050 = ~n10047 & ~n10049;
  assign n10051 = ~n10046 & ~n10050;
  assign n10052 = ~n10039 & ~n10051;
  assign n10053 = n10039 & ~n10050;
  assign n10054 = ~n10046 & n10053;
  assign n10055 = ~n10052 & ~n10054;
  assign n10056 = n8799 & n10055;
  assign n10057 = n8845 & ~n9922;
  assign n10058 = n8797 & n10055;
  assign n10059 = n8794 & ~n10042;
  assign n10060 = n8789 & ~n10042;
  assign n10061 = n8783 & ~n10042;
  assign n10062 = n8786 & n10055;
  assign n10063 = n8792 & n10055;
  assign n10064 = ~n10062 & ~n10063;
  assign n10065 = ~n10060 & ~n10061;
  assign n10066 = n10064 & n10065;
  assign n10067 = ~n10056 & ~n10057;
  assign n10068 = ~n10058 & n10067;
  assign n10069 = ~n10059 & n10068;
  assign n10070 = n10066 & n10069;
  assign n10071 = n10045 & n10070;
  assign n10072 = n8726 & ~n10071;
  assign n10073 = P2_REG0_REG_21_ & ~n8726;
  assign n1760 = n10072 | n10073;
  assign n10075 = ~P2_REG3_REG_22_ & ~P2_REG3_REG_23_;
  assign n10076 = n9969 & n10075;
  assign n10077 = P2_REG3_REG_23_ & ~n10022;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = n8752 & ~n10078;
  assign n10080 = P2_REG0_REG_23_ & n8758;
  assign n10081 = P2_REG1_REG_23_ & n8756;
  assign n10082 = P2_REG2_REG_23_ & n8754;
  assign n10083 = ~n10079 & ~n10080;
  assign n10084 = ~n10081 & n10083;
  assign n10085 = ~n10082 & n10084;
  assign n10086 = n8771 & ~n10085;
  assign n10087 = ~n8455 & ~n8733;
  assign n10088 = ~n8744 & n10087;
  assign n10089 = ~n10031 & ~n10087;
  assign n10090 = n10031 & n10087;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = ~n10036 & ~n10038;
  assign n10093 = ~n10037 & ~n10092;
  assign n10094 = n10091 & n10093;
  assign n10095 = ~n10091 & ~n10093;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = n8766 & ~n10096;
  assign n10098 = ~n10086 & ~n10088;
  assign n10099 = ~n10097 & n10098;
  assign n10100 = n9978 & ~n10033;
  assign n10101 = n9890 & n9995;
  assign n10102 = ~n10050 & ~n10101;
  assign n10103 = ~n10100 & ~n10102;
  assign n10104 = ~n9978 & n10033;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = ~n9889 & n9995;
  assign n10107 = ~n9887 & ~n10100;
  assign n10108 = n10106 & n10107;
  assign n10109 = n10105 & ~n10108;
  assign n10110 = ~n10091 & n10109;
  assign n10111 = n10091 & ~n10109;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = n8799 & ~n10112;
  assign n10114 = n8845 & ~n9978;
  assign n10115 = n8797 & ~n10112;
  assign n10116 = n8794 & ~n10096;
  assign n10117 = n8789 & ~n10096;
  assign n10118 = n8783 & ~n10096;
  assign n10119 = n8786 & ~n10112;
  assign n10120 = n8792 & ~n10112;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 = ~n10117 & ~n10118;
  assign n10123 = n10121 & n10122;
  assign n10124 = ~n10113 & ~n10114;
  assign n10125 = ~n10115 & n10124;
  assign n10126 = ~n10116 & n10125;
  assign n10127 = n10123 & n10126;
  assign n10128 = n10099 & n10127;
  assign n10129 = n8726 & ~n10128;
  assign n10130 = P2_REG0_REG_22_ & ~n8726;
  assign n1765 = n10129 | n10130;
  assign n10132 = ~P2_REG3_REG_24_ & n10076;
  assign n10133 = P2_REG3_REG_24_ & ~n10076;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = n8752 & ~n10134;
  assign n10136 = P2_REG0_REG_24_ & n8758;
  assign n10137 = P2_REG1_REG_24_ & n8756;
  assign n10138 = P2_REG2_REG_24_ & n8754;
  assign n10139 = ~n10135 & ~n10136;
  assign n10140 = ~n10137 & n10139;
  assign n10141 = ~n10138 & n10140;
  assign n10142 = n8771 & ~n10141;
  assign n10143 = ~n8466 & ~n8733;
  assign n10144 = ~n8744 & n10143;
  assign n10145 = ~n10085 & ~n10143;
  assign n10146 = n10085 & n10143;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = ~n10090 & ~n10147;
  assign n10149 = ~n10089 & n10093;
  assign n10150 = n10148 & ~n10149;
  assign n10151 = ~n10089 & ~n10145;
  assign n10152 = ~n10146 & n10151;
  assign n10153 = ~n10090 & ~n10093;
  assign n10154 = n10152 & ~n10153;
  assign n10155 = ~n10150 & ~n10154;
  assign n10156 = n8766 & ~n10155;
  assign n10157 = ~n10142 & ~n10144;
  assign n10158 = ~n10156 & n10157;
  assign n10159 = ~n10031 & n10087;
  assign n10160 = n10031 & ~n10087;
  assign n10161 = ~n10109 & ~n10160;
  assign n10162 = ~n10159 & ~n10161;
  assign n10163 = ~n10147 & n10162;
  assign n10164 = n10147 & ~n10162;
  assign n10165 = ~n10163 & ~n10164;
  assign n10166 = n8799 & ~n10165;
  assign n10167 = n8845 & ~n10031;
  assign n10168 = n8797 & ~n10165;
  assign n10169 = n8794 & ~n10155;
  assign n10170 = n8789 & ~n10155;
  assign n10171 = n8783 & ~n10155;
  assign n10172 = n8786 & ~n10165;
  assign n10173 = n8792 & ~n10165;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = ~n10170 & ~n10171;
  assign n10176 = n10174 & n10175;
  assign n10177 = ~n10166 & ~n10167;
  assign n10178 = ~n10168 & n10177;
  assign n10179 = ~n10169 & n10178;
  assign n10180 = n10176 & n10179;
  assign n10181 = n10158 & n10180;
  assign n10182 = n8726 & ~n10181;
  assign n10183 = P2_REG0_REG_23_ & ~n8726;
  assign n1770 = n10182 | n10183;
  assign n10185 = ~P2_REG3_REG_24_ & ~P2_REG3_REG_25_;
  assign n10186 = n10076 & n10185;
  assign n10187 = P2_REG3_REG_25_ & ~n10132;
  assign n10188 = ~n10186 & ~n10187;
  assign n10189 = n8752 & ~n10188;
  assign n10190 = P2_REG0_REG_25_ & n8758;
  assign n10191 = P2_REG1_REG_25_ & n8756;
  assign n10192 = P2_REG2_REG_25_ & n8754;
  assign n10193 = ~n10189 & ~n10190;
  assign n10194 = ~n10191 & n10193;
  assign n10195 = ~n10192 & n10194;
  assign n10196 = n8771 & ~n10195;
  assign n10197 = ~n8481 & ~n8733;
  assign n10198 = ~n8744 & n10197;
  assign n10199 = ~n10141 & ~n10197;
  assign n10200 = n10141 & n10197;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = ~n10090 & ~n10146;
  assign n10203 = n10037 & n10202;
  assign n10204 = n10151 & ~n10203;
  assign n10205 = ~n10146 & ~n10204;
  assign n10206 = ~n10038 & n10202;
  assign n10207 = ~n10036 & n10206;
  assign n10208 = ~n10205 & ~n10207;
  assign n10209 = ~n10201 & ~n10208;
  assign n10210 = n10201 & n10208;
  assign n10211 = ~n10209 & ~n10210;
  assign n10212 = n8766 & ~n10211;
  assign n10213 = ~n10196 & ~n10198;
  assign n10214 = ~n10212 & n10213;
  assign n10215 = ~n10085 & n10143;
  assign n10216 = n10085 & ~n10143;
  assign n10217 = ~n10162 & ~n10216;
  assign n10218 = ~n10215 & ~n10217;
  assign n10219 = ~n10201 & n10218;
  assign n10220 = n10141 & ~n10197;
  assign n10221 = ~n10141 & n10197;
  assign n10222 = ~n10220 & ~n10221;
  assign n10223 = ~n10218 & ~n10222;
  assign n10224 = ~n10219 & ~n10223;
  assign n10225 = n8799 & ~n10224;
  assign n10226 = n8845 & ~n10085;
  assign n10227 = n8794 & ~n10211;
  assign n10228 = n8797 & ~n10224;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = n8789 & ~n10211;
  assign n10231 = n8783 & ~n10211;
  assign n10232 = n8786 & ~n10224;
  assign n10233 = n8792 & ~n10224;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = ~n10230 & ~n10231;
  assign n10236 = n10234 & n10235;
  assign n10237 = ~n10225 & ~n10226;
  assign n10238 = n10229 & n10237;
  assign n10239 = n10236 & n10238;
  assign n10240 = n10214 & n10239;
  assign n10241 = n8726 & ~n10240;
  assign n10242 = P2_REG0_REG_24_ & ~n8726;
  assign n1775 = n10241 | n10242;
  assign n10244 = ~P2_REG3_REG_26_ & n10186;
  assign n10245 = P2_REG3_REG_26_ & ~n10186;
  assign n10246 = ~n10244 & ~n10245;
  assign n10247 = n8752 & ~n10246;
  assign n10248 = P2_REG0_REG_26_ & n8758;
  assign n10249 = P2_REG1_REG_26_ & n8756;
  assign n10250 = P2_REG2_REG_26_ & n8754;
  assign n10251 = ~n10247 & ~n10248;
  assign n10252 = ~n10249 & n10251;
  assign n10253 = ~n10250 & n10252;
  assign n10254 = n8771 & ~n10253;
  assign n10255 = ~n8492 & ~n8733;
  assign n10256 = ~n8744 & n10255;
  assign n10257 = ~n10195 & ~n10255;
  assign n10258 = n10195 & n10255;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = ~n10200 & ~n10208;
  assign n10261 = ~n10199 & ~n10260;
  assign n10262 = ~n10259 & ~n10261;
  assign n10263 = n10259 & n10261;
  assign n10264 = ~n10262 & ~n10263;
  assign n10265 = n8766 & ~n10264;
  assign n10266 = ~n10254 & ~n10256;
  assign n10267 = ~n10265 & n10266;
  assign n10268 = ~n10218 & ~n10220;
  assign n10269 = ~n10221 & ~n10268;
  assign n10270 = ~n10259 & n10269;
  assign n10271 = n10195 & ~n10255;
  assign n10272 = ~n10195 & n10255;
  assign n10273 = ~n10271 & ~n10272;
  assign n10274 = ~n10269 & ~n10273;
  assign n10275 = ~n10270 & ~n10274;
  assign n10276 = n8799 & ~n10275;
  assign n10277 = n8845 & ~n10141;
  assign n10278 = n8794 & ~n10264;
  assign n10279 = n8797 & ~n10275;
  assign n10280 = ~n10278 & ~n10279;
  assign n10281 = n8789 & ~n10264;
  assign n10282 = n8783 & ~n10264;
  assign n10283 = n8786 & ~n10275;
  assign n10284 = n8792 & ~n10275;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = ~n10281 & ~n10282;
  assign n10287 = n10285 & n10286;
  assign n10288 = ~n10276 & ~n10277;
  assign n10289 = n10280 & n10288;
  assign n10290 = n10287 & n10289;
  assign n10291 = n10267 & n10290;
  assign n10292 = n8726 & ~n10291;
  assign n10293 = P2_REG0_REG_25_ & ~n8726;
  assign n1780 = n10292 | n10293;
  assign n10295 = ~P2_REG3_REG_26_ & ~P2_REG3_REG_27_;
  assign n10296 = n10186 & n10295;
  assign n10297 = P2_REG3_REG_27_ & ~n10244;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = n8752 & ~n10298;
  assign n10300 = P2_REG0_REG_27_ & n8758;
  assign n10301 = P2_REG1_REG_27_ & n8756;
  assign n10302 = P2_REG2_REG_27_ & n8754;
  assign n10303 = ~n10299 & ~n10300;
  assign n10304 = ~n10301 & n10303;
  assign n10305 = ~n10302 & n10304;
  assign n10306 = n8771 & ~n10305;
  assign n10307 = ~n8504 & ~n8733;
  assign n10308 = ~n8744 & n10307;
  assign n10309 = ~n10253 & ~n10307;
  assign n10310 = n10253 & n10307;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = ~n10258 & ~n10261;
  assign n10313 = ~n10257 & ~n10312;
  assign n10314 = n10311 & n10313;
  assign n10315 = ~n10311 & ~n10313;
  assign n10316 = ~n10314 & ~n10315;
  assign n10317 = n8766 & ~n10316;
  assign n10318 = ~n10306 & ~n10308;
  assign n10319 = ~n10317 & n10318;
  assign n10320 = n10269 & ~n10272;
  assign n10321 = ~n10253 & n10307;
  assign n10322 = ~n10271 & n10307;
  assign n10323 = ~n10253 & ~n10271;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = ~n10320 & ~n10321;
  assign n10326 = ~n10324 & n10325;
  assign n10327 = ~n10269 & ~n10271;
  assign n10328 = ~n10272 & ~n10327;
  assign n10329 = n10311 & n10328;
  assign n10330 = ~n10326 & ~n10329;
  assign n10331 = n8799 & n10330;
  assign n10332 = n8845 & ~n10195;
  assign n10333 = n8794 & ~n10316;
  assign n10334 = n8797 & n10330;
  assign n10335 = ~n10333 & ~n10334;
  assign n10336 = n8789 & ~n10316;
  assign n10337 = n8783 & ~n10316;
  assign n10338 = n8786 & n10330;
  assign n10339 = n8792 & n10330;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = ~n10336 & ~n10337;
  assign n10342 = n10340 & n10341;
  assign n10343 = ~n10331 & ~n10332;
  assign n10344 = n10335 & n10343;
  assign n10345 = n10342 & n10344;
  assign n10346 = n10319 & n10345;
  assign n10347 = n8726 & ~n10346;
  assign n10348 = P2_REG0_REG_26_ & ~n8726;
  assign n1785 = n10347 | n10348;
  assign n10350 = ~P2_REG3_REG_28_ & n10296;
  assign n10351 = P2_REG3_REG_28_ & ~n10296;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = n8752 & ~n10352;
  assign n10354 = P2_REG0_REG_28_ & n8758;
  assign n10355 = P2_REG1_REG_28_ & n8756;
  assign n10356 = P2_REG2_REG_28_ & n8754;
  assign n10357 = ~n10353 & ~n10354;
  assign n10358 = ~n10355 & n10357;
  assign n10359 = ~n10356 & n10358;
  assign n10360 = n8771 & ~n10359;
  assign n10361 = ~n8515 & ~n8733;
  assign n10362 = ~n8744 & n10361;
  assign n10363 = ~n10305 & ~n10361;
  assign n10364 = n10305 & n10361;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = ~n10310 & ~n10365;
  assign n10367 = ~n10309 & n10313;
  assign n10368 = n10366 & ~n10367;
  assign n10369 = ~n10309 & n10365;
  assign n10370 = ~n10310 & ~n10313;
  assign n10371 = n10369 & ~n10370;
  assign n10372 = ~n10368 & ~n10371;
  assign n10373 = n8766 & ~n10372;
  assign n10374 = ~n10360 & ~n10362;
  assign n10375 = ~n10373 & n10374;
  assign n10376 = ~n10221 & ~n10272;
  assign n10377 = ~n10324 & ~n10376;
  assign n10378 = n10268 & ~n10324;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = ~n10321 & n10379;
  assign n10381 = ~n10365 & n10380;
  assign n10382 = n10365 & ~n10380;
  assign n10383 = ~n10381 & ~n10382;
  assign n10384 = n8799 & ~n10383;
  assign n10385 = n8845 & ~n10253;
  assign n10386 = n8794 & ~n10372;
  assign n10387 = n8797 & ~n10383;
  assign n10388 = ~n10386 & ~n10387;
  assign n10389 = n8789 & ~n10372;
  assign n10390 = n8783 & ~n10372;
  assign n10391 = n8786 & ~n10383;
  assign n10392 = n8792 & ~n10383;
  assign n10393 = ~n10391 & ~n10392;
  assign n10394 = ~n10389 & ~n10390;
  assign n10395 = n10393 & n10394;
  assign n10396 = ~n10384 & ~n10385;
  assign n10397 = n10388 & n10396;
  assign n10398 = n10395 & n10397;
  assign n10399 = n10375 & n10398;
  assign n10400 = n8726 & ~n10399;
  assign n10401 = P2_REG0_REG_27_ & ~n8726;
  assign n1790 = n10400 | n10401;
  assign n10403 = P2_REG0_REG_29_ & n8758;
  assign n10404 = P2_REG1_REG_29_ & n8756;
  assign n10405 = P2_REG2_REG_29_ & n8754;
  assign n10406 = n8752 & n10350;
  assign n10407 = ~n10403 & ~n10404;
  assign n10408 = ~n10405 & n10407;
  assign n10409 = ~n10406 & n10408;
  assign n10410 = n8771 & ~n10409;
  assign n10411 = ~n8530 & ~n8733;
  assign n10412 = ~n8744 & n10411;
  assign n10413 = ~n10359 & ~n10411;
  assign n10414 = n10359 & n10411;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416 = ~n10305 & n10309;
  assign n10417 = n10305 & ~n10309;
  assign n10418 = ~n10361 & ~n10417;
  assign n10419 = ~n10416 & ~n10418;
  assign n10420 = ~n10310 & ~n10364;
  assign n10421 = ~n10313 & n10420;
  assign n10422 = n10419 & ~n10421;
  assign n10423 = ~n10415 & ~n10422;
  assign n10424 = n10415 & n10422;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = n8766 & ~n10425;
  assign n10427 = ~n10410 & ~n10412;
  assign n10428 = ~n10426 & n10427;
  assign n10429 = n10305 & ~n10361;
  assign n10430 = n10321 & ~n10429;
  assign n10431 = ~n10220 & ~n10429;
  assign n10432 = ~n10218 & ~n10324;
  assign n10433 = n10431 & n10432;
  assign n10434 = n10377 & ~n10429;
  assign n10435 = ~n10305 & n10361;
  assign n10436 = ~n10434 & ~n10435;
  assign n10437 = ~n10430 & ~n10433;
  assign n10438 = n10436 & n10437;
  assign n10439 = ~n10415 & n10438;
  assign n10440 = n10415 & ~n10438;
  assign n10441 = ~n10439 & ~n10440;
  assign n10442 = n8799 & ~n10441;
  assign n10443 = n8845 & ~n10305;
  assign n10444 = n8794 & ~n10425;
  assign n10445 = n8797 & ~n10441;
  assign n10446 = ~n10444 & ~n10445;
  assign n10447 = n8789 & ~n10425;
  assign n10448 = n8783 & ~n10425;
  assign n10449 = n8786 & ~n10441;
  assign n10450 = n8792 & ~n10441;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = ~n10447 & ~n10448;
  assign n10453 = n10451 & n10452;
  assign n10454 = ~n10442 & ~n10443;
  assign n10455 = n10446 & n10454;
  assign n10456 = n10453 & n10455;
  assign n10457 = n10428 & n10456;
  assign n10458 = n8726 & ~n10457;
  assign n10459 = P2_REG0_REG_28_ & ~n8726;
  assign n1795 = n10458 | n10459;
  assign n10461 = ~n8541 & ~n8733;
  assign n10462 = ~n8744 & n10461;
  assign n10463 = ~n10409 & ~n10461;
  assign n10464 = n10409 & n10461;
  assign n10465 = ~n10463 & ~n10464;
  assign n10466 = ~n10413 & n10419;
  assign n10467 = n10465 & n10466;
  assign n10468 = ~n10421 & n10467;
  assign n10469 = n10359 & n10465;
  assign n10470 = n10411 & n10469;
  assign n10471 = ~n10359 & ~n10465;
  assign n10472 = ~n10411 & n10471;
  assign n10473 = ~n10470 & ~n10472;
  assign n10474 = ~n10468 & n10473;
  assign n10475 = ~n10414 & ~n10465;
  assign n10476 = ~n10422 & n10475;
  assign n10477 = n10474 & ~n10476;
  assign n10478 = n8766 & ~n10477;
  assign n10479 = ~n10462 & ~n10478;
  assign n10480 = n8789 & ~n10477;
  assign n10481 = n8783 & ~n10477;
  assign n10482 = n10411 & ~n10438;
  assign n10483 = ~n10359 & ~n10438;
  assign n10484 = ~n10359 & n10411;
  assign n10485 = ~n10482 & ~n10483;
  assign n10486 = ~n10484 & n10485;
  assign n10487 = ~n10465 & n10486;
  assign n10488 = n10465 & ~n10486;
  assign n10489 = ~n10487 & ~n10488;
  assign n10490 = n8786 & ~n10489;
  assign n10491 = n8792 & ~n10489;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = ~n10480 & ~n10481;
  assign n10494 = n10492 & n10493;
  assign n10495 = n8845 & ~n10359;
  assign n10496 = ~P2_B_REG & n8769;
  assign n10497 = ~n8733 & ~n10496;
  assign n10498 = P2_REG0_REG_30_ & n8758;
  assign n10499 = P2_REG1_REG_30_ & n8756;
  assign n10500 = P2_REG2_REG_30_ & n8754;
  assign n10501 = ~n10406 & ~n10498;
  assign n10502 = ~n10499 & n10501;
  assign n10503 = ~n10500 & n10502;
  assign n10504 = n8768 & ~n10497;
  assign n10505 = ~n10503 & n10504;
  assign n10506 = n8799 & ~n10489;
  assign n10507 = n8797 & ~n10489;
  assign n10508 = n8794 & ~n10477;
  assign n10509 = ~n10495 & ~n10505;
  assign n10510 = ~n10506 & n10509;
  assign n10511 = ~n10507 & n10510;
  assign n10512 = ~n10508 & n10511;
  assign n10513 = n10494 & n10512;
  assign n10514 = n10479 & n10513;
  assign n10515 = n8726 & ~n10514;
  assign n10516 = P2_REG0_REG_29_ & ~n8726;
  assign n1800 = n10515 | n10516;
  assign n10518 = P2_REG0_REG_31_ & n8758;
  assign n10519 = P2_REG1_REG_31_ & n8756;
  assign n10520 = P2_REG2_REG_31_ & n8754;
  assign n10521 = ~n10518 & ~n10519;
  assign n10522 = ~n10520 & n10521;
  assign n10523 = ~n10406 & n10522;
  assign n10524 = n10504 & ~n10523;
  assign n10525 = ~n8552 & ~n8733;
  assign n10526 = ~n8744 & n10525;
  assign n10527 = ~n10524 & ~n10526;
  assign n10528 = n8726 & ~n10527;
  assign n10529 = P2_REG0_REG_30_ & ~n8726;
  assign n1805 = n10528 | n10529;
  assign n10531 = ~n8563 & ~n8733;
  assign n10532 = ~n8744 & n10531;
  assign n10533 = ~n10524 & ~n10532;
  assign n10534 = n8726 & ~n10533;
  assign n10535 = P2_REG0_REG_31_ & ~n8726;
  assign n1810 = n10534 | n10535;
  assign n10537 = n8630 & ~n8634;
  assign n10538 = n8694 & n10537;
  assign n10539 = n8705 & n8711;
  assign n10540 = n8698 & ~n8705;
  assign n10541 = ~n10539 & ~n10540;
  assign n10542 = ~n8718 & n10541;
  assign n10543 = n10538 & ~n10542;
  assign n10544 = ~n8630 & n8634;
  assign n10545 = n8694 & n10544;
  assign n10546 = ~n8704 & n8782;
  assign n10547 = ~n8722 & ~n10546;
  assign n10548 = n10545 & ~n10547;
  assign n10549 = ~n10543 & ~n10548;
  assign n10550 = n8582 & ~n10549;
  assign n10551 = ~n8806 & n10550;
  assign n10552 = P2_REG1_REG_0_ & ~n10550;
  assign n1815 = n10551 | n10552;
  assign n10554 = ~n8860 & n10550;
  assign n10555 = P2_REG1_REG_1_ & ~n10550;
  assign n1820 = n10554 | n10555;
  assign n10557 = ~n8916 & n10550;
  assign n10558 = P2_REG1_REG_2_ & ~n10550;
  assign n1825 = n10557 | n10558;
  assign n10560 = ~n8976 & n10550;
  assign n10561 = P2_REG1_REG_3_ & ~n10550;
  assign n1830 = n10560 | n10561;
  assign n10563 = ~n9040 & n10550;
  assign n10564 = P2_REG1_REG_4_ & ~n10550;
  assign n1835 = n10563 | n10564;
  assign n10566 = ~n9100 & n10550;
  assign n10567 = P2_REG1_REG_5_ & ~n10550;
  assign n1840 = n10566 | n10567;
  assign n10569 = ~n9168 & n10550;
  assign n10570 = P2_REG1_REG_6_ & ~n10550;
  assign n1845 = n10569 | n10570;
  assign n10572 = ~n9231 & n10550;
  assign n10573 = P2_REG1_REG_7_ & ~n10550;
  assign n1850 = n10572 | n10573;
  assign n10575 = ~n9294 & n10550;
  assign n10576 = P2_REG1_REG_8_ & ~n10550;
  assign n1855 = n10575 | n10576;
  assign n10578 = ~n9360 & n10550;
  assign n10579 = P2_REG1_REG_9_ & ~n10550;
  assign n1860 = n10578 | n10579;
  assign n10581 = ~n9421 & n10550;
  assign n10582 = P2_REG1_REG_10_ & ~n10550;
  assign n1865 = n10581 | n10582;
  assign n10584 = ~n9485 & n10550;
  assign n10585 = P2_REG1_REG_11_ & ~n10550;
  assign n1870 = n10584 | n10585;
  assign n10587 = ~n9547 & n10550;
  assign n10588 = P2_REG1_REG_12_ & ~n10550;
  assign n1875 = n10587 | n10588;
  assign n10590 = ~n9608 & n10550;
  assign n10591 = P2_REG1_REG_13_ & ~n10550;
  assign n1880 = n10590 | n10591;
  assign n10593 = ~n9668 & n10550;
  assign n10594 = P2_REG1_REG_14_ & ~n10550;
  assign n1885 = n10593 | n10594;
  assign n10596 = ~n9723 & n10550;
  assign n10597 = P2_REG1_REG_15_ & ~n10550;
  assign n1890 = n10596 | n10597;
  assign n10599 = ~n9785 & n10550;
  assign n10600 = P2_REG1_REG_16_ & ~n10550;
  assign n1895 = n10599 | n10600;
  assign n10602 = ~n9848 & n10550;
  assign n10603 = P2_REG1_REG_17_ & ~n10550;
  assign n1900 = n10602 | n10603;
  assign n10605 = ~n9909 & n10550;
  assign n10606 = P2_REG1_REG_18_ & ~n10550;
  assign n1905 = n10605 | n10606;
  assign n10608 = ~n9964 & n10550;
  assign n10609 = P2_REG1_REG_19_ & ~n10550;
  assign n1910 = n10608 | n10609;
  assign n10611 = ~n10018 & n10550;
  assign n10612 = P2_REG1_REG_20_ & ~n10550;
  assign n1915 = n10611 | n10612;
  assign n10614 = ~n10071 & n10550;
  assign n10615 = P2_REG1_REG_21_ & ~n10550;
  assign n1920 = n10614 | n10615;
  assign n10617 = ~n10128 & n10550;
  assign n10618 = P2_REG1_REG_22_ & ~n10550;
  assign n1925 = n10617 | n10618;
  assign n10620 = ~n10181 & n10550;
  assign n10621 = P2_REG1_REG_23_ & ~n10550;
  assign n1930 = n10620 | n10621;
  assign n10623 = ~n10240 & n10550;
  assign n10624 = P2_REG1_REG_24_ & ~n10550;
  assign n1935 = n10623 | n10624;
  assign n10626 = ~n10291 & n10550;
  assign n10627 = P2_REG1_REG_25_ & ~n10550;
  assign n1940 = n10626 | n10627;
  assign n10629 = ~n10346 & n10550;
  assign n10630 = P2_REG1_REG_26_ & ~n10550;
  assign n1945 = n10629 | n10630;
  assign n10632 = ~n10399 & n10550;
  assign n10633 = P2_REG1_REG_27_ & ~n10550;
  assign n1950 = n10632 | n10633;
  assign n10635 = ~n10457 & n10550;
  assign n10636 = P2_REG1_REG_28_ & ~n10550;
  assign n1955 = n10635 | n10636;
  assign n10638 = ~n10514 & n10550;
  assign n10639 = P2_REG1_REG_29_ & ~n10550;
  assign n1960 = n10638 | n10639;
  assign n10641 = ~n10527 & n10550;
  assign n10642 = P2_REG1_REG_30_ & ~n10550;
  assign n1965 = n10641 | n10642;
  assign n10644 = ~n10533 & n10550;
  assign n10645 = P2_REG1_REG_31_ & ~n10550;
  assign n1970 = n10644 | n10645;
  assign n10647 = ~n8701 & n8704;
  assign n10648 = ~n8711 & n10647;
  assign n10649 = n8701 & ~n8711;
  assign n10650 = ~n8698 & ~n10649;
  assign n10651 = ~n8705 & n10650;
  assign n10652 = n10545 & ~n10651;
  assign n10653 = n8704 & n8743;
  assign n10654 = n10538 & ~n10547;
  assign n10655 = ~n10652 & ~n10653;
  assign n10656 = ~n10654 & n10655;
  assign n10657 = n8582 & ~n10656;
  assign n10658 = n10648 & n10657;
  assign n10659 = ~n8765 & n10658;
  assign n10660 = n8771 & n10657;
  assign n10661 = ~n8778 & n10660;
  assign n10662 = ~n8704 & n8743;
  assign n10663 = ~n8741 & ~n10662;
  assign n10664 = n10657 & ~n10663;
  assign n10665 = ~n8739 & n10664;
  assign n10666 = ~n8805 & n10657;
  assign n10667 = P2_REG2_REG_0_ & ~n10657;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = n10653 & n10657;
  assign n10670 = P2_REG3_REG_0_ & n10669;
  assign n10671 = ~n10659 & ~n10661;
  assign n10672 = ~n10665 & n10671;
  assign n10673 = n10668 & n10672;
  assign n1975 = n10670 | ~n10673;
  assign n10675 = ~n8830 & n10658;
  assign n10676 = ~n8816 & n10660;
  assign n10677 = ~n8823 & n10664;
  assign n10678 = ~n8859 & n10657;
  assign n10679 = P2_REG2_REG_1_ & ~n10657;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = P2_REG3_REG_1_ & n10669;
  assign n10682 = ~n10675 & ~n10676;
  assign n10683 = ~n10677 & n10682;
  assign n10684 = n10680 & n10683;
  assign n1980 = n10681 | ~n10684;
  assign n10686 = ~n8888 & n10658;
  assign n10687 = ~n8870 & n10660;
  assign n10688 = ~n8877 & n10664;
  assign n10689 = ~n8915 & n10657;
  assign n10690 = P2_REG2_REG_2_ & ~n10657;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = P2_REG3_REG_2_ & n10669;
  assign n10693 = ~n10686 & ~n10687;
  assign n10694 = ~n10688 & n10693;
  assign n10695 = n10691 & n10694;
  assign n1985 = n10692 | ~n10695;
  assign n10697 = ~n8947 & n10658;
  assign n10698 = ~n8929 & n10660;
  assign n10699 = ~n8936 & n10664;
  assign n10700 = ~n8975 & n10657;
  assign n10701 = P2_REG2_REG_3_ & ~n10657;
  assign n10702 = ~n10700 & ~n10701;
  assign n10703 = ~P2_REG3_REG_3_ & n10669;
  assign n10704 = ~n10697 & ~n10698;
  assign n10705 = ~n10699 & n10704;
  assign n10706 = n10702 & n10705;
  assign n1990 = n10703 | ~n10706;
  assign n10708 = ~n9010 & n10658;
  assign n10709 = ~n8989 & n10660;
  assign n10710 = ~n8996 & n10664;
  assign n10711 = ~n9039 & n10657;
  assign n10712 = P2_REG2_REG_4_ & ~n10657;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~n8922 & n10669;
  assign n10715 = ~n10708 & ~n10709;
  assign n10716 = ~n10710 & n10715;
  assign n10717 = n10713 & n10716;
  assign n1995 = n10714 | ~n10717;
  assign n10719 = ~n9071 & n10658;
  assign n10720 = ~n9055 & n10660;
  assign n10721 = ~n9062 & n10664;
  assign n10722 = ~n9099 & n10657;
  assign n10723 = P2_REG2_REG_5_ & ~n10657;
  assign n10724 = ~n10722 & ~n10723;
  assign n10725 = ~n8982 & n10669;
  assign n10726 = ~n10719 & ~n10720;
  assign n10727 = ~n10721 & n10726;
  assign n10728 = n10724 & n10727;
  assign n2000 = n10725 | ~n10728;
  assign n10730 = ~n9133 & n10658;
  assign n10731 = ~n9114 & n10660;
  assign n10732 = ~n9121 & n10664;
  assign n10733 = ~n9167 & n10657;
  assign n10734 = P2_REG2_REG_6_ & ~n10657;
  assign n10735 = ~n10733 & ~n10734;
  assign n10736 = ~n9048 & n10669;
  assign n10737 = ~n10730 & ~n10731;
  assign n10738 = ~n10732 & n10737;
  assign n10739 = n10735 & n10738;
  assign n2005 = n10736 | ~n10739;
  assign n10741 = ~n9107 & n10669;
  assign n10742 = ~n9188 & n10664;
  assign n10743 = ~n9202 & n10658;
  assign n10744 = ~n9181 & n10660;
  assign n10745 = ~n9230 & n10657;
  assign n10746 = P2_REG2_REG_7_ & ~n10657;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = ~n10741 & ~n10742;
  assign n10749 = ~n10743 & n10748;
  assign n10750 = ~n10744 & n10749;
  assign n2010 = ~n10747 | ~n10750;
  assign n10752 = ~n9174 & n10669;
  assign n10753 = ~n9252 & n10664;
  assign n10754 = ~n9263 & n10658;
  assign n10755 = ~n9245 & n10660;
  assign n10756 = ~n9293 & n10657;
  assign n10757 = P2_REG2_REG_8_ & ~n10657;
  assign n10758 = ~n10756 & ~n10757;
  assign n10759 = ~n10752 & ~n10753;
  assign n10760 = ~n10754 & n10759;
  assign n10761 = ~n10755 & n10760;
  assign n2015 = ~n10758 | ~n10761;
  assign n10763 = ~n9316 & n10664;
  assign n10764 = ~n9309 & n10660;
  assign n10765 = ~n9238 & n10669;
  assign n10766 = ~n9333 & n10658;
  assign n10767 = ~n9359 & n10657;
  assign n10768 = P2_REG2_REG_9_ & ~n10657;
  assign n10769 = ~n10767 & ~n10768;
  assign n10770 = ~n10763 & ~n10764;
  assign n10771 = ~n10765 & n10770;
  assign n10772 = ~n10766 & n10771;
  assign n2020 = ~n10769 | ~n10772;
  assign n10774 = ~n9383 & n10664;
  assign n10775 = ~n9376 & n10660;
  assign n10776 = ~n9302 & n10669;
  assign n10777 = ~n9392 & n10658;
  assign n10778 = ~n9420 & n10657;
  assign n10779 = P2_REG2_REG_10_ & ~n10657;
  assign n10780 = ~n10778 & ~n10779;
  assign n10781 = ~n10774 & ~n10775;
  assign n10782 = ~n10776 & n10781;
  assign n10783 = ~n10777 & n10782;
  assign n2025 = ~n10780 | ~n10783;
  assign n10785 = ~n9441 & n10664;
  assign n10786 = ~n9434 & n10660;
  assign n10787 = ~n9369 & n10669;
  assign n10788 = ~n9453 & n10658;
  assign n10789 = ~n9484 & n10657;
  assign n10790 = P2_REG2_REG_11_ & ~n10657;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = ~n10785 & ~n10786;
  assign n10793 = ~n10787 & n10792;
  assign n10794 = ~n10788 & n10793;
  assign n2030 = ~n10791 | ~n10794;
  assign n10796 = ~n9506 & n10664;
  assign n10797 = ~n9499 & n10660;
  assign n10798 = ~n9427 & n10669;
  assign n10799 = ~n9520 & n10658;
  assign n10800 = ~n9546 & n10657;
  assign n10801 = P2_REG2_REG_12_ & ~n10657;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~n10796 & ~n10797;
  assign n10804 = ~n10798 & n10803;
  assign n10805 = ~n10799 & n10804;
  assign n2035 = ~n10802 | ~n10805;
  assign n10807 = ~n9567 & n10664;
  assign n10808 = ~n9560 & n10660;
  assign n10809 = ~n9492 & n10669;
  assign n10810 = ~n9579 & n10658;
  assign n10811 = ~n9607 & n10657;
  assign n10812 = P2_REG2_REG_13_ & ~n10657;
  assign n10813 = ~n10811 & ~n10812;
  assign n10814 = ~n10807 & ~n10808;
  assign n10815 = ~n10809 & n10814;
  assign n10816 = ~n10810 & n10815;
  assign n2040 = ~n10813 | ~n10816;
  assign n10818 = ~n9630 & n10664;
  assign n10819 = ~n9623 & n10660;
  assign n10820 = ~n9553 & n10669;
  assign n10821 = ~n9639 & n10658;
  assign n10822 = ~n9667 & n10657;
  assign n10823 = P2_REG2_REG_14_ & ~n10657;
  assign n10824 = ~n10822 & ~n10823;
  assign n10825 = ~n10818 & ~n10819;
  assign n10826 = ~n10820 & n10825;
  assign n10827 = ~n10821 & n10826;
  assign n2045 = ~n10824 | ~n10827;
  assign n10829 = ~n9688 & n10664;
  assign n10830 = ~n9681 & n10660;
  assign n10831 = ~n9616 & n10669;
  assign n10832 = ~n9697 & n10658;
  assign n10833 = ~n9722 & n10657;
  assign n10834 = P2_REG2_REG_15_ & ~n10657;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = ~n10829 & ~n10830;
  assign n10837 = ~n10831 & n10836;
  assign n10838 = ~n10832 & n10837;
  assign n2050 = ~n10835 | ~n10838;
  assign n10840 = ~n9744 & n10664;
  assign n10841 = ~n9737 & n10660;
  assign n10842 = ~n9674 & n10669;
  assign n10843 = ~n9756 & n10658;
  assign n10844 = ~n9784 & n10657;
  assign n10845 = P2_REG2_REG_16_ & ~n10657;
  assign n10846 = ~n10844 & ~n10845;
  assign n10847 = ~n10840 & ~n10841;
  assign n10848 = ~n10842 & n10847;
  assign n10849 = ~n10843 & n10848;
  assign n2055 = ~n10846 | ~n10849;
  assign n10851 = ~n9805 & n10664;
  assign n10852 = ~n9798 & n10660;
  assign n10853 = ~n9730 & n10669;
  assign n10854 = ~n9819 & n10658;
  assign n10855 = ~n9847 & n10657;
  assign n10856 = P2_REG2_REG_17_ & ~n10657;
  assign n10857 = ~n10855 & ~n10856;
  assign n10858 = ~n10851 & ~n10852;
  assign n10859 = ~n10853 & n10858;
  assign n10860 = ~n10854 & n10859;
  assign n2060 = ~n10857 | ~n10860;
  assign n10862 = ~n9869 & n10664;
  assign n10863 = ~n9862 & n10660;
  assign n10864 = ~n9791 & n10669;
  assign n10865 = ~n9878 & n10658;
  assign n10866 = ~n9908 & n10657;
  assign n10867 = P2_REG2_REG_18_ & ~n10657;
  assign n10868 = ~n10866 & ~n10867;
  assign n10869 = ~n10862 & ~n10863;
  assign n10870 = ~n10864 & n10869;
  assign n10871 = ~n10865 & n10870;
  assign n2065 = ~n10868 | ~n10871;
  assign n10873 = ~n9926 & n10664;
  assign n10874 = ~n9922 & n10660;
  assign n10875 = ~n9855 & n10669;
  assign n10876 = ~n9937 & n10658;
  assign n10877 = ~n9963 & n10657;
  assign n10878 = P2_REG2_REG_19_ & ~n10657;
  assign n10879 = ~n10877 & ~n10878;
  assign n10880 = ~n10873 & ~n10874;
  assign n10881 = ~n10875 & n10880;
  assign n10882 = ~n10876 & n10881;
  assign n2070 = ~n10879 | ~n10882;
  assign n10884 = n9980 & n10664;
  assign n10885 = ~n9978 & n10660;
  assign n10886 = ~n9915 & n10669;
  assign n10887 = ~n9989 & n10658;
  assign n10888 = ~n10017 & n10657;
  assign n10889 = P2_REG2_REG_20_ & ~n10657;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = ~n10884 & ~n10885;
  assign n10892 = ~n10886 & n10891;
  assign n10893 = ~n10887 & n10892;
  assign n2075 = ~n10890 | ~n10893;
  assign n10895 = n10033 & n10664;
  assign n10896 = ~n10031 & n10660;
  assign n10897 = ~n9971 & n10669;
  assign n10898 = ~n10042 & n10658;
  assign n10899 = ~n10070 & n10657;
  assign n10900 = P2_REG2_REG_21_ & ~n10657;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 = ~n10895 & ~n10896;
  assign n10903 = ~n10897 & n10902;
  assign n10904 = ~n10898 & n10903;
  assign n2080 = ~n10901 | ~n10904;
  assign n10906 = n10087 & n10664;
  assign n10907 = ~n10085 & n10660;
  assign n10908 = ~n10024 & n10669;
  assign n10909 = ~n10096 & n10658;
  assign n10910 = ~n10127 & n10657;
  assign n10911 = P2_REG2_REG_22_ & ~n10657;
  assign n10912 = ~n10910 & ~n10911;
  assign n10913 = ~n10906 & ~n10907;
  assign n10914 = ~n10908 & n10913;
  assign n10915 = ~n10909 & n10914;
  assign n2085 = ~n10912 | ~n10915;
  assign n10917 = n10143 & n10664;
  assign n10918 = ~n10141 & n10660;
  assign n10919 = ~n10078 & n10669;
  assign n10920 = ~n10155 & n10658;
  assign n10921 = ~n10180 & n10657;
  assign n10922 = P2_REG2_REG_23_ & ~n10657;
  assign n10923 = ~n10921 & ~n10922;
  assign n10924 = ~n10917 & ~n10918;
  assign n10925 = ~n10919 & n10924;
  assign n10926 = ~n10920 & n10925;
  assign n2090 = ~n10923 | ~n10926;
  assign n10928 = n10197 & n10664;
  assign n10929 = ~n10195 & n10660;
  assign n10930 = ~n10134 & n10669;
  assign n10931 = ~n10211 & n10658;
  assign n10932 = ~n10239 & n10657;
  assign n10933 = P2_REG2_REG_24_ & ~n10657;
  assign n10934 = ~n10932 & ~n10933;
  assign n10935 = ~n10928 & ~n10929;
  assign n10936 = ~n10930 & n10935;
  assign n10937 = ~n10931 & n10936;
  assign n2095 = ~n10934 | ~n10937;
  assign n10939 = n10255 & n10664;
  assign n10940 = ~n10253 & n10660;
  assign n10941 = ~n10188 & n10669;
  assign n10942 = ~n10264 & n10658;
  assign n10943 = ~n10290 & n10657;
  assign n10944 = P2_REG2_REG_25_ & ~n10657;
  assign n10945 = ~n10943 & ~n10944;
  assign n10946 = ~n10939 & ~n10940;
  assign n10947 = ~n10941 & n10946;
  assign n10948 = ~n10942 & n10947;
  assign n2100 = ~n10945 | ~n10948;
  assign n10950 = n10307 & n10664;
  assign n10951 = ~n10305 & n10660;
  assign n10952 = ~n10246 & n10669;
  assign n10953 = ~n10316 & n10658;
  assign n10954 = ~n10345 & n10657;
  assign n10955 = P2_REG2_REG_26_ & ~n10657;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = ~n10950 & ~n10951;
  assign n10958 = ~n10952 & n10957;
  assign n10959 = ~n10953 & n10958;
  assign n2105 = ~n10956 | ~n10959;
  assign n10961 = n10361 & n10664;
  assign n10962 = ~n10359 & n10660;
  assign n10963 = ~n10298 & n10669;
  assign n10964 = ~n10372 & n10658;
  assign n10965 = ~n10398 & n10657;
  assign n10966 = P2_REG2_REG_27_ & ~n10657;
  assign n10967 = ~n10965 & ~n10966;
  assign n10968 = ~n10961 & ~n10962;
  assign n10969 = ~n10963 & n10968;
  assign n10970 = ~n10964 & n10969;
  assign n2110 = ~n10967 | ~n10970;
  assign n10972 = n10411 & n10664;
  assign n10973 = ~n10409 & n10660;
  assign n10974 = ~n10352 & n10669;
  assign n10975 = ~n10425 & n10658;
  assign n10976 = ~n10456 & n10657;
  assign n10977 = P2_REG2_REG_28_ & ~n10657;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~n10972 & ~n10973;
  assign n10980 = ~n10974 & n10979;
  assign n10981 = ~n10975 & n10980;
  assign n2115 = ~n10978 | ~n10981;
  assign n10983 = n10461 & n10664;
  assign n10984 = n10350 & n10669;
  assign n10985 = ~n10477 & n10658;
  assign n10986 = ~n10513 & n10657;
  assign n10987 = P2_REG2_REG_29_ & ~n10657;
  assign n10988 = ~n10986 & ~n10987;
  assign n10989 = ~n10983 & ~n10984;
  assign n10990 = ~n10985 & n10989;
  assign n2120 = ~n10988 | ~n10990;
  assign n10992 = P2_REG2_REG_30_ & ~n10657;
  assign n10993 = n10524 & n10657;
  assign n10994 = ~n10984 & ~n10993;
  assign n10995 = n10525 & n10664;
  assign n10996 = ~n10992 & n10994;
  assign n2125 = n10995 | ~n10996;
  assign n10998 = P2_REG2_REG_31_ & ~n10657;
  assign n10999 = n10531 & n10664;
  assign n11000 = n10994 & ~n10998;
  assign n2130 = n10999 | ~n11000;
  assign n11002 = ~n8569 & ~n8733;
  assign n11003 = ~n8733 & ~n8768;
  assign n11004 = ~n11002 & ~n11003;
  assign n11005 = n8569 & n8580;
  assign n11006 = P2_STATE_REG & ~n11005;
  assign n11007 = n11004 & n11006;
  assign n11008 = n8582 & ~n11007;
  assign n11009 = ~n8786 & ~n10653;
  assign n11010 = ~n8721 & ~n8792;
  assign n11011 = ~n8799 & n11010;
  assign n11012 = ~n8797 & n11011;
  assign n11013 = ~n8794 & n11012;
  assign n11014 = ~n10647 & n10663;
  assign n11015 = n11009 & n11014;
  assign n11016 = n11013 & n11015;
  assign n11017 = n8732 & ~n11016;
  assign n11018 = ~n8711 & n11017;
  assign n11019 = P2_REG2_REG_18_ & n9866;
  assign n11020 = ~P2_REG2_REG_19_ & ~n8711;
  assign n11021 = P2_REG2_REG_19_ & n8711;
  assign n11022 = ~n11020 & ~n11021;
  assign n11023 = ~n11019 & ~n11022;
  assign n11024 = ~P2_REG2_REG_17_ & ~n9802;
  assign n11025 = P2_REG2_REG_17_ & n9802;
  assign n11026 = ~P2_REG2_REG_16_ & ~n9741;
  assign n11027 = P2_REG2_REG_16_ & n9741;
  assign n11028 = ~P2_REG2_REG_14_ & ~n9627;
  assign n11029 = P2_REG2_REG_14_ & n9627;
  assign n11030 = ~P2_REG2_REG_13_ & ~n9564;
  assign n11031 = P2_REG2_REG_13_ & n9564;
  assign n11032 = ~P2_REG2_REG_12_ & ~n9503;
  assign n11033 = P2_REG2_REG_12_ & n9503;
  assign n11034 = ~P2_REG2_REG_11_ & ~n9438;
  assign n11035 = P2_REG2_REG_11_ & n9438;
  assign n11036 = ~P2_REG2_REG_10_ & ~n9380;
  assign n11037 = P2_REG2_REG_10_ & n9380;
  assign n11038 = ~P2_REG2_REG_9_ & ~n9313;
  assign n11039 = P2_REG2_REG_9_ & n9313;
  assign n11040 = ~P2_REG2_REG_8_ & ~n9249;
  assign n11041 = P2_REG2_REG_8_ & n9249;
  assign n11042 = ~P2_REG2_REG_7_ & ~n9185;
  assign n11043 = P2_REG2_REG_7_ & n9185;
  assign n11044 = ~P2_REG2_REG_6_ & ~n9118;
  assign n11045 = P2_REG2_REG_6_ & n9118;
  assign n11046 = ~P2_REG2_REG_5_ & ~n9059;
  assign n11047 = P2_REG2_REG_5_ & n9059;
  assign n11048 = ~P2_REG2_REG_4_ & ~n8993;
  assign n11049 = P2_REG2_REG_4_ & n8993;
  assign n11050 = ~P2_REG2_REG_3_ & ~n8933;
  assign n11051 = P2_REG2_REG_3_ & n8933;
  assign n11052 = ~P2_REG2_REG_2_ & ~n8874;
  assign n11053 = P2_REG2_REG_2_ & n8874;
  assign n11054 = P2_REG2_REG_0_ & n8736;
  assign n11055 = ~P2_REG2_REG_1_ & ~n11054;
  assign n11056 = P2_REG2_REG_1_ & n11054;
  assign n11057 = ~n8820 & ~n11056;
  assign n11058 = ~n11055 & ~n11057;
  assign n11059 = ~n11053 & ~n11058;
  assign n11060 = ~n11052 & ~n11059;
  assign n11061 = ~n11051 & ~n11060;
  assign n11062 = ~n11050 & ~n11061;
  assign n11063 = ~n11049 & ~n11062;
  assign n11064 = ~n11048 & ~n11063;
  assign n11065 = ~n11047 & ~n11064;
  assign n11066 = ~n11046 & ~n11065;
  assign n11067 = ~n11045 & ~n11066;
  assign n11068 = ~n11044 & ~n11067;
  assign n11069 = ~n11043 & ~n11068;
  assign n11070 = ~n11042 & ~n11069;
  assign n11071 = ~n11041 & ~n11070;
  assign n11072 = ~n11040 & ~n11071;
  assign n11073 = ~n11039 & ~n11072;
  assign n11074 = ~n11038 & ~n11073;
  assign n11075 = ~n11037 & ~n11074;
  assign n11076 = ~n11036 & ~n11075;
  assign n11077 = ~n11035 & ~n11076;
  assign n11078 = ~n11034 & ~n11077;
  assign n11079 = ~n11033 & ~n11078;
  assign n11080 = ~n11032 & ~n11079;
  assign n11081 = ~n11031 & ~n11080;
  assign n11082 = ~n11030 & ~n11081;
  assign n11083 = ~n11029 & ~n11082;
  assign n11084 = ~n11028 & ~n11083;
  assign n11085 = ~P2_REG2_REG_15_ & ~n11084;
  assign n11086 = P2_REG2_REG_15_ & n11084;
  assign n11087 = ~n9685 & ~n11086;
  assign n11088 = ~n11085 & ~n11087;
  assign n11089 = ~n11027 & ~n11088;
  assign n11090 = ~n11026 & ~n11089;
  assign n11091 = ~n11025 & ~n11090;
  assign n11092 = ~n11024 & ~n11091;
  assign n11093 = ~P2_REG2_REG_18_ & ~n9866;
  assign n11094 = n11092 & ~n11093;
  assign n11095 = n11023 & ~n11094;
  assign n11096 = n11022 & ~n11093;
  assign n11097 = ~n11019 & ~n11092;
  assign n11098 = n11096 & ~n11097;
  assign n11099 = ~n11095 & ~n11098;
  assign n11100 = n8769 & ~n11016;
  assign n11101 = ~n11099 & n11100;
  assign n11102 = P2_REG1_REG_18_ & n9866;
  assign n11103 = ~P2_REG1_REG_19_ & ~n8711;
  assign n11104 = P2_REG1_REG_19_ & n8711;
  assign n11105 = ~n11103 & ~n11104;
  assign n11106 = ~n11102 & ~n11105;
  assign n11107 = ~P2_REG1_REG_17_ & ~n9802;
  assign n11108 = P2_REG1_REG_17_ & n9802;
  assign n11109 = ~P2_REG1_REG_16_ & ~n9741;
  assign n11110 = P2_REG1_REG_16_ & n9741;
  assign n11111 = ~P2_REG1_REG_14_ & ~n9627;
  assign n11112 = P2_REG1_REG_14_ & n9627;
  assign n11113 = ~P2_REG1_REG_13_ & ~n9564;
  assign n11114 = P2_REG1_REG_13_ & n9564;
  assign n11115 = ~P2_REG1_REG_12_ & ~n9503;
  assign n11116 = P2_REG1_REG_12_ & n9503;
  assign n11117 = ~P2_REG1_REG_11_ & ~n9438;
  assign n11118 = P2_REG1_REG_11_ & n9438;
  assign n11119 = ~P2_REG1_REG_10_ & ~n9380;
  assign n11120 = P2_REG1_REG_10_ & n9380;
  assign n11121 = ~P2_REG1_REG_9_ & ~n9313;
  assign n11122 = P2_REG1_REG_9_ & n9313;
  assign n11123 = ~P2_REG1_REG_8_ & ~n9249;
  assign n11124 = P2_REG1_REG_8_ & n9249;
  assign n11125 = ~P2_REG1_REG_7_ & ~n9185;
  assign n11126 = P2_REG1_REG_7_ & n9185;
  assign n11127 = ~P2_REG1_REG_6_ & ~n9118;
  assign n11128 = P2_REG1_REG_6_ & n9118;
  assign n11129 = ~P2_REG1_REG_5_ & ~n9059;
  assign n11130 = P2_REG1_REG_5_ & n9059;
  assign n11131 = ~P2_REG1_REG_4_ & ~n8993;
  assign n11132 = P2_REG1_REG_4_ & n8993;
  assign n11133 = ~P2_REG1_REG_3_ & ~n8933;
  assign n11134 = P2_REG1_REG_3_ & n8933;
  assign n11135 = ~P2_REG1_REG_2_ & ~n8874;
  assign n11136 = P2_REG1_REG_2_ & n8874;
  assign n11137 = P2_REG1_REG_0_ & n8736;
  assign n11138 = ~P2_REG1_REG_1_ & ~n11137;
  assign n11139 = P2_REG1_REG_1_ & n11137;
  assign n11140 = ~n8820 & ~n11139;
  assign n11141 = ~n11138 & ~n11140;
  assign n11142 = ~n11136 & ~n11141;
  assign n11143 = ~n11135 & ~n11142;
  assign n11144 = ~n11134 & ~n11143;
  assign n11145 = ~n11133 & ~n11144;
  assign n11146 = ~n11132 & ~n11145;
  assign n11147 = ~n11131 & ~n11146;
  assign n11148 = ~n11130 & ~n11147;
  assign n11149 = ~n11129 & ~n11148;
  assign n11150 = ~n11128 & ~n11149;
  assign n11151 = ~n11127 & ~n11150;
  assign n11152 = ~n11126 & ~n11151;
  assign n11153 = ~n11125 & ~n11152;
  assign n11154 = ~n11124 & ~n11153;
  assign n11155 = ~n11123 & ~n11154;
  assign n11156 = ~n11122 & ~n11155;
  assign n11157 = ~n11121 & ~n11156;
  assign n11158 = ~n11120 & ~n11157;
  assign n11159 = ~n11119 & ~n11158;
  assign n11160 = ~n11118 & ~n11159;
  assign n11161 = ~n11117 & ~n11160;
  assign n11162 = ~n11116 & ~n11161;
  assign n11163 = ~n11115 & ~n11162;
  assign n11164 = ~n11114 & ~n11163;
  assign n11165 = ~n11113 & ~n11164;
  assign n11166 = ~n11112 & ~n11165;
  assign n11167 = ~n11111 & ~n11166;
  assign n11168 = ~P2_REG1_REG_15_ & ~n11167;
  assign n11169 = P2_REG1_REG_15_ & n11167;
  assign n11170 = ~n9685 & ~n11169;
  assign n11171 = ~n11168 & ~n11170;
  assign n11172 = ~n11110 & ~n11171;
  assign n11173 = ~n11109 & ~n11172;
  assign n11174 = ~n11108 & ~n11173;
  assign n11175 = ~n11107 & ~n11174;
  assign n11176 = ~P2_REG1_REG_18_ & ~n9866;
  assign n11177 = n11175 & ~n11176;
  assign n11178 = n11106 & ~n11177;
  assign n11179 = n11105 & ~n11176;
  assign n11180 = ~n11102 & ~n11175;
  assign n11181 = n11179 & ~n11180;
  assign n11182 = ~n11178 & ~n11181;
  assign n11183 = n8729 & ~n11016;
  assign n11184 = ~n11182 & n11183;
  assign n11185 = ~n11018 & ~n11101;
  assign n11186 = ~n11184 & n11185;
  assign n11187 = n11008 & ~n11186;
  assign n11188 = P2_STATE_REG & n8569;
  assign n2555 = n8580 & n11188;
  assign n11190 = ~n8732 & n2555;
  assign n11191 = P2_STATE_REG & ~n8569;
  assign n11192 = ~n11007 & n11191;
  assign n11193 = n8732 & n11192;
  assign n11194 = ~n11190 & ~n11193;
  assign n11195 = ~n8711 & ~n11194;
  assign n11196 = P2_REG2_REG_19_ & ~n8729;
  assign n11197 = P2_REG1_REG_19_ & n8729;
  assign n11198 = ~n11196 & ~n11197;
  assign n11199 = n8711 & ~n11198;
  assign n11200 = ~n8711 & n11198;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = P2_REG2_REG_18_ & ~n8729;
  assign n11203 = P2_REG1_REG_18_ & n8729;
  assign n11204 = ~n11202 & ~n11203;
  assign n11205 = P2_REG2_REG_17_ & ~n8729;
  assign n11206 = P2_REG1_REG_17_ & n8729;
  assign n11207 = ~n11205 & ~n11206;
  assign n11208 = n9802 & ~n11207;
  assign n11209 = ~n9802 & n11207;
  assign n11210 = P2_REG2_REG_16_ & ~n8729;
  assign n11211 = P2_REG1_REG_16_ & n8729;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n9741 & n11212;
  assign n11214 = P2_REG2_REG_15_ & ~n8729;
  assign n11215 = P2_REG1_REG_15_ & n8729;
  assign n11216 = ~n11214 & ~n11215;
  assign n11217 = n9685 & ~n11216;
  assign n11218 = n9741 & ~n11212;
  assign n11219 = ~n11217 & ~n11218;
  assign n11220 = P2_REG2_REG_14_ & ~n8729;
  assign n11221 = P2_REG1_REG_14_ & n8729;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = n9627 & ~n11222;
  assign n11224 = ~n9685 & n11216;
  assign n11225 = ~n11213 & ~n11224;
  assign n11226 = n11223 & n11225;
  assign n11227 = n11219 & ~n11226;
  assign n11228 = ~n11213 & ~n11227;
  assign n11229 = ~n9627 & n11222;
  assign n11230 = P2_REG2_REG_13_ & ~n8729;
  assign n11231 = P2_REG1_REG_13_ & n8729;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = n9564 & ~n11232;
  assign n11234 = ~n9564 & n11232;
  assign n11235 = P2_REG2_REG_12_ & ~n8729;
  assign n11236 = P2_REG1_REG_12_ & n8729;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = n9503 & ~n11237;
  assign n11239 = ~n9503 & n11237;
  assign n11240 = P2_REG2_REG_11_ & ~n8729;
  assign n11241 = P2_REG1_REG_11_ & n8729;
  assign n11242 = ~n11240 & ~n11241;
  assign n11243 = ~n9438 & n11242;
  assign n11244 = P2_REG2_REG_10_ & ~n8729;
  assign n11245 = P2_REG1_REG_10_ & n8729;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = n9380 & ~n11246;
  assign n11248 = n9438 & ~n11242;
  assign n11249 = ~n11247 & ~n11248;
  assign n11250 = P2_REG2_REG_9_ & ~n8729;
  assign n11251 = P2_REG1_REG_9_ & n8729;
  assign n11252 = ~n11250 & ~n11251;
  assign n11253 = n9313 & ~n11252;
  assign n11254 = ~n9380 & n11246;
  assign n11255 = ~n11243 & ~n11254;
  assign n11256 = n11253 & n11255;
  assign n11257 = n11249 & ~n11256;
  assign n11258 = ~n11243 & ~n11257;
  assign n11259 = ~n9313 & n11252;
  assign n11260 = P2_REG2_REG_8_ & ~n8729;
  assign n11261 = P2_REG1_REG_8_ & n8729;
  assign n11262 = ~n11260 & ~n11261;
  assign n11263 = P2_REG2_REG_7_ & ~n8729;
  assign n11264 = P2_REG1_REG_7_ & n8729;
  assign n11265 = ~n11263 & ~n11264;
  assign n11266 = n9185 & ~n11265;
  assign n11267 = n11262 & ~n11266;
  assign n11268 = n9249 & ~n11267;
  assign n11269 = ~n11262 & n11266;
  assign n11270 = ~n9249 & n11262;
  assign n11271 = ~n9185 & n11265;
  assign n11272 = P2_REG2_REG_6_ & ~n8729;
  assign n11273 = P2_REG1_REG_6_ & n8729;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~n9118 & n11274;
  assign n11276 = P2_REG2_REG_5_ & ~n8729;
  assign n11277 = P2_REG1_REG_5_ & n8729;
  assign n11278 = ~n11276 & ~n11277;
  assign n11279 = n9059 & ~n11278;
  assign n11280 = n9118 & ~n11274;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = P2_REG2_REG_4_ & ~n8729;
  assign n11283 = P2_REG1_REG_4_ & n8729;
  assign n11284 = ~n11282 & ~n11283;
  assign n11285 = n8993 & ~n11284;
  assign n11286 = ~n9059 & n11278;
  assign n11287 = ~n11275 & ~n11286;
  assign n11288 = n11285 & n11287;
  assign n11289 = n11281 & ~n11288;
  assign n11290 = ~n11275 & ~n11289;
  assign n11291 = ~n8993 & n11284;
  assign n11292 = P2_REG2_REG_3_ & ~n8729;
  assign n11293 = P2_REG1_REG_3_ & n8729;
  assign n11294 = ~n11292 & ~n11293;
  assign n11295 = P2_REG2_REG_2_ & ~n8729;
  assign n11296 = P2_REG1_REG_2_ & n8729;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = n8874 & ~n11297;
  assign n11299 = n11294 & ~n11298;
  assign n11300 = n8933 & ~n11299;
  assign n11301 = ~n11294 & n11298;
  assign n11302 = ~n8933 & n11294;
  assign n11303 = ~n8874 & n11297;
  assign n11304 = P2_REG2_REG_1_ & ~n8729;
  assign n11305 = P2_REG1_REG_1_ & n8729;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = P2_REG2_REG_0_ & ~n8729;
  assign n11308 = P2_REG1_REG_0_ & n8729;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = ~n8736 & n11309;
  assign n11311 = ~n11306 & ~n11310;
  assign n11312 = n11306 & n11310;
  assign n11313 = n8820 & ~n11312;
  assign n11314 = ~n11311 & ~n11313;
  assign n11315 = ~n11302 & ~n11303;
  assign n11316 = ~n11314 & n11315;
  assign n11317 = ~n11300 & ~n11301;
  assign n11318 = ~n11316 & n11317;
  assign n11319 = n11287 & ~n11291;
  assign n11320 = ~n11318 & n11319;
  assign n11321 = ~n11290 & ~n11320;
  assign n11322 = ~n11270 & ~n11271;
  assign n11323 = ~n11321 & n11322;
  assign n11324 = ~n11268 & ~n11269;
  assign n11325 = ~n11323 & n11324;
  assign n11326 = n11255 & ~n11259;
  assign n11327 = ~n11325 & n11326;
  assign n11328 = ~n11258 & ~n11327;
  assign n11329 = ~n11239 & ~n11328;
  assign n11330 = ~n11238 & ~n11329;
  assign n11331 = ~n11234 & ~n11330;
  assign n11332 = ~n11233 & ~n11331;
  assign n11333 = n11225 & ~n11229;
  assign n11334 = ~n11332 & n11333;
  assign n11335 = ~n11228 & ~n11334;
  assign n11336 = ~n11209 & ~n11335;
  assign n11337 = ~n11208 & ~n11336;
  assign n11338 = ~n11204 & ~n11337;
  assign n11339 = n11204 & n11337;
  assign n11340 = n9866 & ~n11339;
  assign n11341 = ~n11338 & ~n11340;
  assign n11342 = ~n11201 & ~n11341;
  assign n11343 = n11201 & n11341;
  assign n11344 = ~n11342 & ~n11343;
  assign n11345 = ~n8733 & ~n8842;
  assign n11346 = n2555 & ~n11345;
  assign n11347 = ~n11344 & n11346;
  assign n11348 = n8769 & n11192;
  assign n11349 = ~n11099 & n11348;
  assign n11350 = P2_ADDR_REG_19_ & n11007;
  assign n11351 = P2_REG3_REG_19_ & ~P2_STATE_REG;
  assign n11352 = ~n11350 & ~n11351;
  assign n11353 = n8729 & n11192;
  assign n11354 = ~n11182 & n11353;
  assign n11355 = n11352 & ~n11354;
  assign n11356 = ~n11195 & ~n11347;
  assign n11357 = ~n11349 & n11356;
  assign n11358 = n11355 & n11357;
  assign n2135 = n11187 | ~n11358;
  assign n11360 = ~n9866 & n11017;
  assign n11361 = ~n11019 & ~n11093;
  assign n11362 = ~n11092 & ~n11361;
  assign n11363 = n11092 & n11361;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = n11100 & ~n11364;
  assign n11366 = ~n11102 & ~n11176;
  assign n11367 = ~n11175 & ~n11366;
  assign n11368 = n11175 & n11366;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = n11183 & ~n11369;
  assign n11371 = ~n11360 & ~n11365;
  assign n11372 = ~n11370 & n11371;
  assign n11373 = n11008 & ~n11372;
  assign n11374 = ~n9866 & ~n11194;
  assign n11375 = n9866 & ~n11204;
  assign n11376 = ~n9866 & n11204;
  assign n11377 = ~n11375 & ~n11376;
  assign n11378 = ~n11337 & ~n11377;
  assign n11379 = n11337 & n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = n11346 & ~n11380;
  assign n11382 = n11348 & ~n11364;
  assign n11383 = P2_ADDR_REG_18_ & n11007;
  assign n11384 = P2_REG3_REG_18_ & ~P2_STATE_REG;
  assign n11385 = ~n11383 & ~n11384;
  assign n11386 = n11353 & ~n11369;
  assign n11387 = n11385 & ~n11386;
  assign n11388 = ~n11374 & ~n11381;
  assign n11389 = ~n11382 & n11388;
  assign n11390 = n11387 & n11389;
  assign n2140 = n11373 | ~n11390;
  assign n11392 = ~n9802 & n11017;
  assign n11393 = ~n11024 & ~n11025;
  assign n11394 = ~n11090 & ~n11393;
  assign n11395 = n11090 & n11393;
  assign n11396 = ~n11394 & ~n11395;
  assign n11397 = n11100 & ~n11396;
  assign n11398 = ~n11107 & ~n11108;
  assign n11399 = ~n11173 & ~n11398;
  assign n11400 = n11173 & n11398;
  assign n11401 = ~n11399 & ~n11400;
  assign n11402 = n11183 & ~n11401;
  assign n11403 = ~n11392 & ~n11397;
  assign n11404 = ~n11402 & n11403;
  assign n11405 = n11008 & ~n11404;
  assign n11406 = ~n9802 & ~n11194;
  assign n11407 = ~n11208 & ~n11209;
  assign n11408 = ~n11335 & ~n11407;
  assign n11409 = n11335 & n11407;
  assign n11410 = ~n11408 & ~n11409;
  assign n11411 = n11346 & ~n11410;
  assign n11412 = n11348 & ~n11396;
  assign n11413 = P2_ADDR_REG_17_ & n11007;
  assign n11414 = P2_REG3_REG_17_ & ~P2_STATE_REG;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = n11353 & ~n11401;
  assign n11417 = n11415 & ~n11416;
  assign n11418 = ~n11406 & ~n11411;
  assign n11419 = ~n11412 & n11418;
  assign n11420 = n11417 & n11419;
  assign n2145 = n11405 | ~n11420;
  assign n11422 = ~n9741 & n11017;
  assign n11423 = ~n11026 & ~n11027;
  assign n11424 = ~n11088 & ~n11423;
  assign n11425 = n11088 & n11423;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = n11100 & ~n11426;
  assign n11428 = ~n11109 & ~n11110;
  assign n11429 = ~n11171 & ~n11428;
  assign n11430 = n11171 & n11428;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = n11183 & ~n11431;
  assign n11433 = ~n11422 & ~n11427;
  assign n11434 = ~n11432 & n11433;
  assign n11435 = n11008 & ~n11434;
  assign n11436 = ~n9741 & ~n11194;
  assign n11437 = ~n11213 & ~n11218;
  assign n11438 = ~n11229 & ~n11332;
  assign n11439 = ~n11223 & ~n11438;
  assign n11440 = ~n11217 & n11439;
  assign n11441 = ~n11224 & ~n11437;
  assign n11442 = ~n11440 & n11441;
  assign n11443 = ~n11224 & ~n11439;
  assign n11444 = ~n11213 & n11219;
  assign n11445 = ~n11443 & n11444;
  assign n11446 = ~n11442 & ~n11445;
  assign n11447 = n11346 & ~n11446;
  assign n11448 = n11348 & ~n11426;
  assign n11449 = P2_ADDR_REG_16_ & n11007;
  assign n11450 = P2_REG3_REG_16_ & ~P2_STATE_REG;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = n11353 & ~n11431;
  assign n11453 = n11451 & ~n11452;
  assign n11454 = ~n11436 & ~n11447;
  assign n11455 = ~n11448 & n11454;
  assign n11456 = n11453 & n11455;
  assign n2150 = n11435 | ~n11456;
  assign n11458 = ~n9685 & n11017;
  assign n11459 = P2_REG2_REG_15_ & n9685;
  assign n11460 = ~P2_REG2_REG_15_ & ~n9685;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = ~n11084 & ~n11461;
  assign n11463 = n11084 & n11461;
  assign n11464 = ~n11462 & ~n11463;
  assign n11465 = n11100 & ~n11464;
  assign n11466 = P2_REG1_REG_15_ & n9685;
  assign n11467 = ~P2_REG1_REG_15_ & ~n9685;
  assign n11468 = ~n11466 & ~n11467;
  assign n11469 = ~n11167 & ~n11468;
  assign n11470 = n11167 & n11468;
  assign n11471 = ~n11469 & ~n11470;
  assign n11472 = n11183 & ~n11471;
  assign n11473 = ~n11458 & ~n11465;
  assign n11474 = ~n11472 & n11473;
  assign n11475 = n11008 & ~n11474;
  assign n11476 = ~n9685 & ~n11194;
  assign n11477 = ~n11217 & ~n11224;
  assign n11478 = n11439 & n11477;
  assign n11479 = ~n11439 & ~n11477;
  assign n11480 = ~n11478 & ~n11479;
  assign n11481 = n11346 & ~n11480;
  assign n11482 = n11348 & ~n11464;
  assign n11483 = P2_ADDR_REG_15_ & n11007;
  assign n11484 = P2_REG3_REG_15_ & ~P2_STATE_REG;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = n11353 & ~n11471;
  assign n11487 = n11485 & ~n11486;
  assign n11488 = ~n11476 & ~n11481;
  assign n11489 = ~n11482 & n11488;
  assign n11490 = n11487 & n11489;
  assign n2155 = n11475 | ~n11490;
  assign n11492 = ~n9627 & n11017;
  assign n11493 = ~n11028 & ~n11029;
  assign n11494 = ~n11082 & ~n11493;
  assign n11495 = n11082 & n11493;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = n11100 & ~n11496;
  assign n11498 = ~n11111 & ~n11112;
  assign n11499 = ~n11165 & ~n11498;
  assign n11500 = n11165 & n11498;
  assign n11501 = ~n11499 & ~n11500;
  assign n11502 = n11183 & ~n11501;
  assign n11503 = ~n11492 & ~n11497;
  assign n11504 = ~n11502 & n11503;
  assign n11505 = n11008 & ~n11504;
  assign n11506 = ~n9627 & ~n11194;
  assign n11507 = ~n11223 & ~n11229;
  assign n11508 = n11332 & n11507;
  assign n11509 = ~n11332 & ~n11507;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = n11346 & ~n11510;
  assign n11512 = n11348 & ~n11496;
  assign n11513 = P2_ADDR_REG_14_ & n11007;
  assign n11514 = P2_REG3_REG_14_ & ~P2_STATE_REG;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = n11353 & ~n11501;
  assign n11517 = n11515 & ~n11516;
  assign n11518 = ~n11506 & ~n11511;
  assign n11519 = ~n11512 & n11518;
  assign n11520 = n11517 & n11519;
  assign n2160 = n11505 | ~n11520;
  assign n11522 = ~n9564 & n11017;
  assign n11523 = ~n11030 & ~n11031;
  assign n11524 = ~n11080 & ~n11523;
  assign n11525 = n11080 & n11523;
  assign n11526 = ~n11524 & ~n11525;
  assign n11527 = n11100 & ~n11526;
  assign n11528 = ~n11113 & ~n11114;
  assign n11529 = ~n11163 & ~n11528;
  assign n11530 = n11163 & n11528;
  assign n11531 = ~n11529 & ~n11530;
  assign n11532 = n11183 & ~n11531;
  assign n11533 = ~n11522 & ~n11527;
  assign n11534 = ~n11532 & n11533;
  assign n11535 = n11008 & ~n11534;
  assign n11536 = ~n9564 & ~n11194;
  assign n11537 = ~n11233 & ~n11234;
  assign n11538 = ~n11330 & ~n11537;
  assign n11539 = n11330 & n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = n11346 & ~n11540;
  assign n11542 = n11348 & ~n11526;
  assign n11543 = P2_ADDR_REG_13_ & n11007;
  assign n11544 = P2_REG3_REG_13_ & ~P2_STATE_REG;
  assign n11545 = ~n11543 & ~n11544;
  assign n11546 = n11353 & ~n11531;
  assign n11547 = n11545 & ~n11546;
  assign n11548 = ~n11536 & ~n11541;
  assign n11549 = ~n11542 & n11548;
  assign n11550 = n11547 & n11549;
  assign n2165 = n11535 | ~n11550;
  assign n11552 = ~n9503 & n11017;
  assign n11553 = ~n11032 & ~n11033;
  assign n11554 = ~n11078 & ~n11553;
  assign n11555 = n11078 & n11553;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = n11100 & ~n11556;
  assign n11558 = ~n11115 & ~n11116;
  assign n11559 = ~n11161 & ~n11558;
  assign n11560 = n11161 & n11558;
  assign n11561 = ~n11559 & ~n11560;
  assign n11562 = n11183 & ~n11561;
  assign n11563 = ~n11552 & ~n11557;
  assign n11564 = ~n11562 & n11563;
  assign n11565 = n11008 & ~n11564;
  assign n11566 = ~n9503 & ~n11194;
  assign n11567 = ~n11238 & ~n11239;
  assign n11568 = ~n11328 & ~n11567;
  assign n11569 = n11328 & n11567;
  assign n11570 = ~n11568 & ~n11569;
  assign n11571 = n11346 & ~n11570;
  assign n11572 = n11348 & ~n11556;
  assign n11573 = P2_ADDR_REG_12_ & n11007;
  assign n11574 = P2_REG3_REG_12_ & ~P2_STATE_REG;
  assign n11575 = ~n11573 & ~n11574;
  assign n11576 = n11353 & ~n11561;
  assign n11577 = n11575 & ~n11576;
  assign n11578 = ~n11566 & ~n11571;
  assign n11579 = ~n11572 & n11578;
  assign n11580 = n11577 & n11579;
  assign n2170 = n11565 | ~n11580;
  assign n11582 = ~n9438 & n11017;
  assign n11583 = ~n11034 & ~n11035;
  assign n11584 = ~n11076 & ~n11583;
  assign n11585 = n11076 & n11583;
  assign n11586 = ~n11584 & ~n11585;
  assign n11587 = n11100 & ~n11586;
  assign n11588 = ~n11117 & ~n11118;
  assign n11589 = ~n11159 & ~n11588;
  assign n11590 = n11159 & n11588;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = n11183 & ~n11591;
  assign n11593 = ~n11582 & ~n11587;
  assign n11594 = ~n11592 & n11593;
  assign n11595 = n11008 & ~n11594;
  assign n11596 = ~n9438 & ~n11194;
  assign n11597 = n11348 & ~n11586;
  assign n11598 = ~n11243 & ~n11248;
  assign n11599 = ~n11259 & ~n11325;
  assign n11600 = ~n11253 & ~n11599;
  assign n11601 = ~n11247 & n11600;
  assign n11602 = ~n11254 & ~n11598;
  assign n11603 = ~n11601 & n11602;
  assign n11604 = ~n11254 & ~n11600;
  assign n11605 = ~n11243 & n11249;
  assign n11606 = ~n11604 & n11605;
  assign n11607 = ~n11603 & ~n11606;
  assign n11608 = n11346 & ~n11607;
  assign n11609 = P2_ADDR_REG_11_ & n11007;
  assign n11610 = P2_REG3_REG_11_ & ~P2_STATE_REG;
  assign n11611 = ~n11609 & ~n11610;
  assign n11612 = n11353 & ~n11591;
  assign n11613 = n11611 & ~n11612;
  assign n11614 = ~n11596 & ~n11597;
  assign n11615 = ~n11608 & n11614;
  assign n11616 = n11613 & n11615;
  assign n2175 = n11595 | ~n11616;
  assign n11618 = ~n9380 & n11017;
  assign n11619 = ~n11036 & ~n11037;
  assign n11620 = ~n11074 & ~n11619;
  assign n11621 = n11074 & n11619;
  assign n11622 = ~n11620 & ~n11621;
  assign n11623 = n11100 & ~n11622;
  assign n11624 = ~n11119 & ~n11120;
  assign n11625 = ~n11157 & ~n11624;
  assign n11626 = n11157 & n11624;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = n11183 & ~n11627;
  assign n11629 = ~n11618 & ~n11623;
  assign n11630 = ~n11628 & n11629;
  assign n11631 = n11008 & ~n11630;
  assign n11632 = ~n9380 & ~n11194;
  assign n11633 = n11348 & ~n11622;
  assign n11634 = ~n11247 & ~n11254;
  assign n11635 = n11600 & n11634;
  assign n11636 = ~n11600 & ~n11634;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = n11346 & ~n11637;
  assign n11639 = P2_ADDR_REG_10_ & n11007;
  assign n11640 = P2_REG3_REG_10_ & ~P2_STATE_REG;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = n11353 & ~n11627;
  assign n11643 = n11641 & ~n11642;
  assign n11644 = ~n11632 & ~n11633;
  assign n11645 = ~n11638 & n11644;
  assign n11646 = n11643 & n11645;
  assign n2180 = n11631 | ~n11646;
  assign n11648 = ~n9313 & n11017;
  assign n11649 = ~n11038 & ~n11039;
  assign n11650 = ~n11072 & ~n11649;
  assign n11651 = n11072 & n11649;
  assign n11652 = ~n11650 & ~n11651;
  assign n11653 = n11100 & ~n11652;
  assign n11654 = ~n11121 & ~n11122;
  assign n11655 = ~n11155 & ~n11654;
  assign n11656 = n11155 & n11654;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = n11183 & ~n11657;
  assign n11659 = ~n11648 & ~n11653;
  assign n11660 = ~n11658 & n11659;
  assign n11661 = n11008 & ~n11660;
  assign n11662 = ~n9313 & ~n11194;
  assign n11663 = n11348 & ~n11652;
  assign n11664 = ~n11253 & ~n11259;
  assign n11665 = n11325 & n11664;
  assign n11666 = ~n11325 & ~n11664;
  assign n11667 = ~n11665 & ~n11666;
  assign n11668 = n11346 & ~n11667;
  assign n11669 = P2_ADDR_REG_9_ & n11007;
  assign n11670 = P2_REG3_REG_9_ & ~P2_STATE_REG;
  assign n11671 = ~n11669 & ~n11670;
  assign n11672 = n11353 & ~n11657;
  assign n11673 = n11671 & ~n11672;
  assign n11674 = ~n11662 & ~n11663;
  assign n11675 = ~n11668 & n11674;
  assign n11676 = n11673 & n11675;
  assign n2185 = n11661 | ~n11676;
  assign n11678 = P2_ADDR_REG_8_ & n11007;
  assign n11679 = P2_REG3_REG_8_ & ~P2_STATE_REG;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11123 & ~n11124;
  assign n11682 = ~n11153 & ~n11681;
  assign n11683 = n11153 & n11681;
  assign n11684 = ~n11682 & ~n11683;
  assign n11685 = n11353 & ~n11684;
  assign n11686 = ~n11040 & ~n11041;
  assign n11687 = ~n11070 & ~n11686;
  assign n11688 = n11070 & n11686;
  assign n11689 = ~n11687 & ~n11688;
  assign n11690 = n11348 & ~n11689;
  assign n11691 = n11680 & ~n11685;
  assign n11692 = ~n11690 & n11691;
  assign n11693 = ~n9249 & n11017;
  assign n11694 = n11100 & ~n11689;
  assign n11695 = n11183 & ~n11684;
  assign n11696 = ~n11693 & ~n11694;
  assign n11697 = ~n11695 & n11696;
  assign n11698 = n11008 & ~n11697;
  assign n11699 = ~n9249 & ~n11194;
  assign n11700 = n9249 & ~n11262;
  assign n11701 = ~n11270 & ~n11700;
  assign n11702 = ~n11266 & n11321;
  assign n11703 = ~n11271 & ~n11701;
  assign n11704 = ~n11702 & n11703;
  assign n11705 = ~n11271 & ~n11321;
  assign n11706 = ~n11266 & n11701;
  assign n11707 = ~n11705 & n11706;
  assign n11708 = ~n11704 & ~n11707;
  assign n11709 = n11346 & ~n11708;
  assign n11710 = ~n11699 & ~n11709;
  assign n11711 = n11692 & ~n11698;
  assign n2190 = ~n11710 | ~n11711;
  assign n11713 = P2_ADDR_REG_7_ & n11007;
  assign n11714 = P2_REG3_REG_7_ & ~P2_STATE_REG;
  assign n11715 = ~n11713 & ~n11714;
  assign n11716 = ~n11125 & ~n11126;
  assign n11717 = ~n11151 & ~n11716;
  assign n11718 = n11151 & n11716;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = n11353 & ~n11719;
  assign n11721 = ~n11042 & ~n11043;
  assign n11722 = ~n11068 & ~n11721;
  assign n11723 = n11068 & n11721;
  assign n11724 = ~n11722 & ~n11723;
  assign n11725 = n11348 & ~n11724;
  assign n11726 = n11715 & ~n11720;
  assign n11727 = ~n11725 & n11726;
  assign n11728 = ~n9185 & n11017;
  assign n11729 = n11100 & ~n11724;
  assign n11730 = n11183 & ~n11719;
  assign n11731 = ~n11728 & ~n11729;
  assign n11732 = ~n11730 & n11731;
  assign n11733 = n11008 & ~n11732;
  assign n11734 = ~n9185 & ~n11194;
  assign n11735 = ~n11266 & ~n11271;
  assign n11736 = n11321 & n11735;
  assign n11737 = ~n11321 & ~n11735;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = n11346 & ~n11738;
  assign n11740 = ~n11734 & ~n11739;
  assign n11741 = n11727 & ~n11733;
  assign n2195 = ~n11740 | ~n11741;
  assign n11743 = ~n9118 & n11017;
  assign n11744 = ~n11044 & ~n11045;
  assign n11745 = ~n11066 & ~n11744;
  assign n11746 = n11066 & n11744;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = n11100 & ~n11747;
  assign n11749 = ~n11127 & ~n11128;
  assign n11750 = ~n11149 & ~n11749;
  assign n11751 = n11149 & n11749;
  assign n11752 = ~n11750 & ~n11751;
  assign n11753 = n11183 & ~n11752;
  assign n11754 = ~n11743 & ~n11748;
  assign n11755 = ~n11753 & n11754;
  assign n11756 = n11008 & ~n11755;
  assign n11757 = n11348 & ~n11747;
  assign n11758 = ~n9118 & ~n11194;
  assign n11759 = P2_ADDR_REG_6_ & n11007;
  assign n11760 = P2_REG3_REG_6_ & ~P2_STATE_REG;
  assign n11761 = ~n11759 & ~n11760;
  assign n11762 = n11353 & ~n11752;
  assign n11763 = n11761 & ~n11762;
  assign n11764 = ~n11757 & ~n11758;
  assign n11765 = n11763 & n11764;
  assign n11766 = ~n11275 & ~n11280;
  assign n11767 = ~n11291 & ~n11318;
  assign n11768 = ~n11285 & ~n11767;
  assign n11769 = ~n11279 & n11768;
  assign n11770 = ~n11286 & ~n11766;
  assign n11771 = ~n11769 & n11770;
  assign n11772 = ~n11286 & ~n11768;
  assign n11773 = ~n11275 & n11281;
  assign n11774 = ~n11772 & n11773;
  assign n11775 = ~n11771 & ~n11774;
  assign n11776 = n11346 & ~n11775;
  assign n11777 = ~n11756 & n11765;
  assign n2200 = n11776 | ~n11777;
  assign n11779 = ~n9059 & n11017;
  assign n11780 = ~n11046 & ~n11047;
  assign n11781 = ~n11064 & ~n11780;
  assign n11782 = n11064 & n11780;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = n11100 & ~n11783;
  assign n11785 = ~n11129 & ~n11130;
  assign n11786 = ~n11147 & ~n11785;
  assign n11787 = n11147 & n11785;
  assign n11788 = ~n11786 & ~n11787;
  assign n11789 = n11183 & ~n11788;
  assign n11790 = ~n11779 & ~n11784;
  assign n11791 = ~n11789 & n11790;
  assign n11792 = n11008 & ~n11791;
  assign n11793 = n11348 & ~n11783;
  assign n11794 = ~n9059 & ~n11194;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = P2_ADDR_REG_5_ & n11007;
  assign n11797 = P2_REG3_REG_5_ & ~P2_STATE_REG;
  assign n11798 = ~n11796 & ~n11797;
  assign n11799 = n11353 & ~n11788;
  assign n11800 = n11798 & ~n11799;
  assign n11801 = ~n11279 & ~n11286;
  assign n11802 = n11768 & n11801;
  assign n11803 = ~n11768 & ~n11801;
  assign n11804 = ~n11802 & ~n11803;
  assign n11805 = n11346 & ~n11804;
  assign n11806 = ~n11792 & n11795;
  assign n11807 = n11800 & n11806;
  assign n2205 = n11805 | ~n11807;
  assign n11809 = ~n11048 & ~n11049;
  assign n11810 = ~n11062 & ~n11809;
  assign n11811 = n11062 & n11809;
  assign n11812 = ~n11810 & ~n11811;
  assign n11813 = n11348 & ~n11812;
  assign n11814 = ~n8993 & n11017;
  assign n11815 = n11100 & ~n11812;
  assign n11816 = ~n11131 & ~n11132;
  assign n11817 = ~n11145 & ~n11816;
  assign n11818 = n11145 & n11816;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = n11183 & ~n11819;
  assign n11821 = ~n11814 & ~n11815;
  assign n11822 = ~n11820 & n11821;
  assign n11823 = n11008 & ~n11822;
  assign n11824 = ~n8993 & ~n11194;
  assign n11825 = P2_ADDR_REG_4_ & n11007;
  assign n11826 = P2_REG3_REG_4_ & ~P2_STATE_REG;
  assign n11827 = ~n11825 & ~n11826;
  assign n11828 = n11353 & ~n11819;
  assign n11829 = n11827 & ~n11828;
  assign n11830 = ~n11285 & ~n11291;
  assign n11831 = n11318 & n11830;
  assign n11832 = ~n11318 & ~n11830;
  assign n11833 = ~n11831 & ~n11832;
  assign n11834 = n11346 & ~n11833;
  assign n11835 = ~n11824 & n11829;
  assign n11836 = ~n11834 & n11835;
  assign n11837 = ~n11813 & ~n11823;
  assign n2210 = ~n11836 | ~n11837;
  assign n11839 = ~n11050 & ~n11051;
  assign n11840 = ~n11060 & ~n11839;
  assign n11841 = n11060 & n11839;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = n11348 & ~n11842;
  assign n11844 = ~n8933 & n11017;
  assign n11845 = n11100 & ~n11842;
  assign n11846 = ~n11133 & ~n11134;
  assign n11847 = ~n11143 & ~n11846;
  assign n11848 = n11143 & n11846;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = n11183 & ~n11849;
  assign n11851 = ~n11844 & ~n11845;
  assign n11852 = ~n11850 & n11851;
  assign n11853 = n11008 & ~n11852;
  assign n11854 = ~n8933 & ~n11194;
  assign n11855 = P2_ADDR_REG_3_ & n11007;
  assign n11856 = P2_REG3_REG_3_ & ~P2_STATE_REG;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = n11353 & ~n11849;
  assign n11859 = n11857 & ~n11858;
  assign n11860 = n8933 & ~n11294;
  assign n11861 = ~n11302 & ~n11860;
  assign n11862 = ~n11298 & n11314;
  assign n11863 = ~n11303 & ~n11861;
  assign n11864 = ~n11862 & n11863;
  assign n11865 = ~n11303 & ~n11314;
  assign n11866 = ~n11298 & n11861;
  assign n11867 = ~n11865 & n11866;
  assign n11868 = ~n11864 & ~n11867;
  assign n11869 = n11346 & ~n11868;
  assign n11870 = ~n11854 & n11859;
  assign n11871 = ~n11869 & n11870;
  assign n11872 = ~n11843 & ~n11853;
  assign n2215 = ~n11871 | ~n11872;
  assign n11874 = ~n8874 & n11017;
  assign n11875 = ~n11052 & ~n11053;
  assign n11876 = ~n11058 & ~n11875;
  assign n11877 = n11058 & n11875;
  assign n11878 = ~n11876 & ~n11877;
  assign n11879 = n11100 & ~n11878;
  assign n11880 = ~n11135 & ~n11136;
  assign n11881 = ~n11141 & ~n11880;
  assign n11882 = n11141 & n11880;
  assign n11883 = ~n11881 & ~n11882;
  assign n11884 = n11183 & ~n11883;
  assign n11885 = ~n11874 & ~n11879;
  assign n11886 = ~n11884 & n11885;
  assign n11887 = n11008 & ~n11886;
  assign n11888 = ~n8874 & ~n11194;
  assign n11889 = n11348 & ~n11878;
  assign n11890 = ~n11298 & ~n11303;
  assign n11891 = n11314 & n11890;
  assign n11892 = ~n11314 & ~n11890;
  assign n11893 = ~n11891 & ~n11892;
  assign n11894 = n11346 & ~n11893;
  assign n11895 = P2_ADDR_REG_2_ & n11007;
  assign n11896 = P2_REG3_REG_2_ & ~P2_STATE_REG;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = n11353 & ~n11883;
  assign n11899 = n11897 & ~n11898;
  assign n11900 = ~n11888 & ~n11889;
  assign n11901 = ~n11894 & n11900;
  assign n11902 = n11899 & n11901;
  assign n2220 = n11887 | ~n11902;
  assign n11904 = ~n8820 & n11017;
  assign n11905 = P2_REG2_REG_1_ & ~n11054;
  assign n11906 = ~P2_REG2_REG_1_ & n11054;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = n8820 & ~n11907;
  assign n11909 = ~n8820 & n11907;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = n11100 & ~n11910;
  assign n11912 = P2_REG1_REG_1_ & ~n11137;
  assign n11913 = ~P2_REG1_REG_1_ & n11137;
  assign n11914 = ~n11912 & ~n11913;
  assign n11915 = n8820 & ~n11914;
  assign n11916 = ~n8820 & n11914;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = n11183 & ~n11917;
  assign n11919 = ~n11904 & ~n11911;
  assign n11920 = ~n11918 & n11919;
  assign n11921 = n11008 & ~n11920;
  assign n11922 = ~n8820 & ~n11194;
  assign n11923 = n8820 & ~n11306;
  assign n11924 = ~n8820 & n11306;
  assign n11925 = ~n11923 & ~n11924;
  assign n11926 = ~n11310 & ~n11925;
  assign n11927 = n11310 & n11925;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = n11346 & ~n11928;
  assign n11930 = n11348 & ~n11910;
  assign n11931 = P2_ADDR_REG_1_ & n11007;
  assign n11932 = P2_REG3_REG_1_ & ~P2_STATE_REG;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = n11353 & ~n11917;
  assign n11935 = n11933 & ~n11934;
  assign n11936 = ~n11922 & ~n11929;
  assign n11937 = ~n11930 & n11936;
  assign n11938 = n11935 & n11937;
  assign n2225 = n11921 | ~n11938;
  assign n11940 = ~n8736 & n11017;
  assign n11941 = ~P2_REG2_REG_0_ & ~n8736;
  assign n11942 = ~n11054 & ~n11941;
  assign n11943 = n11100 & ~n11942;
  assign n11944 = ~P2_REG1_REG_0_ & ~n8736;
  assign n11945 = ~n11137 & ~n11944;
  assign n11946 = n11183 & ~n11945;
  assign n11947 = ~n11940 & ~n11943;
  assign n11948 = ~n11946 & n11947;
  assign n11949 = n11008 & ~n11948;
  assign n11950 = ~n8736 & ~n11194;
  assign n11951 = n8736 & ~n11309;
  assign n11952 = ~n11310 & ~n11951;
  assign n11953 = n11346 & ~n11952;
  assign n11954 = n11348 & ~n11942;
  assign n11955 = P2_ADDR_REG_0_ & n11007;
  assign n11956 = P2_REG3_REG_0_ & ~P2_STATE_REG;
  assign n11957 = ~n11955 & ~n11956;
  assign n11958 = n11353 & ~n11945;
  assign n11959 = n11957 & ~n11958;
  assign n11960 = ~n11950 & ~n11953;
  assign n11961 = ~n11954 & n11960;
  assign n11962 = n11959 & n11961;
  assign n2230 = n11949 | ~n11962;
  assign n11964 = ~n8762 & n2555;
  assign n11965 = P2_DATAO_REG_0_ & ~n2555;
  assign n2235 = n11964 | n11965;
  assign n11967 = ~n8778 & n2555;
  assign n11968 = P2_DATAO_REG_1_ & ~n2555;
  assign n2240 = n11967 | n11968;
  assign n11970 = ~n8816 & n2555;
  assign n11971 = P2_DATAO_REG_2_ & ~n2555;
  assign n2245 = n11970 | n11971;
  assign n11973 = ~n8870 & n2555;
  assign n11974 = P2_DATAO_REG_3_ & ~n2555;
  assign n2250 = n11973 | n11974;
  assign n11976 = ~n8929 & n2555;
  assign n11977 = P2_DATAO_REG_4_ & ~n2555;
  assign n2255 = n11976 | n11977;
  assign n11979 = ~n8989 & n2555;
  assign n11980 = P2_DATAO_REG_5_ & ~n2555;
  assign n2260 = n11979 | n11980;
  assign n11982 = ~n9055 & n2555;
  assign n11983 = P2_DATAO_REG_6_ & ~n2555;
  assign n2265 = n11982 | n11983;
  assign n11985 = ~n9114 & n2555;
  assign n11986 = P2_DATAO_REG_7_ & ~n2555;
  assign n2270 = n11985 | n11986;
  assign n11988 = ~n9181 & n2555;
  assign n11989 = P2_DATAO_REG_8_ & ~n2555;
  assign n2275 = n11988 | n11989;
  assign n11991 = ~n9245 & n2555;
  assign n11992 = P2_DATAO_REG_9_ & ~n2555;
  assign n2280 = n11991 | n11992;
  assign n11994 = ~n9309 & n2555;
  assign n11995 = P2_DATAO_REG_10_ & ~n2555;
  assign n2285 = n11994 | n11995;
  assign n11997 = ~n9376 & n2555;
  assign n11998 = P2_DATAO_REG_11_ & ~n2555;
  assign n2290 = n11997 | n11998;
  assign n12000 = ~n9434 & n2555;
  assign n12001 = P2_DATAO_REG_12_ & ~n2555;
  assign n2295 = n12000 | n12001;
  assign n12003 = ~n9499 & n2555;
  assign n12004 = P2_DATAO_REG_13_ & ~n2555;
  assign n2300 = n12003 | n12004;
  assign n12006 = ~n9560 & n2555;
  assign n12007 = P2_DATAO_REG_14_ & ~n2555;
  assign n2305 = n12006 | n12007;
  assign n12009 = ~n9623 & n2555;
  assign n12010 = P2_DATAO_REG_15_ & ~n2555;
  assign n2310 = n12009 | n12010;
  assign n12012 = ~n9681 & n2555;
  assign n12013 = P2_DATAO_REG_16_ & ~n2555;
  assign n2315 = n12012 | n12013;
  assign n12015 = ~n9737 & n2555;
  assign n12016 = P2_DATAO_REG_17_ & ~n2555;
  assign n2320 = n12015 | n12016;
  assign n12018 = ~n9798 & n2555;
  assign n12019 = P2_DATAO_REG_18_ & ~n2555;
  assign n2325 = n12018 | n12019;
  assign n12021 = ~n9862 & n2555;
  assign n12022 = P2_DATAO_REG_19_ & ~n2555;
  assign n2330 = n12021 | n12022;
  assign n12024 = ~n9922 & n2555;
  assign n12025 = P2_DATAO_REG_20_ & ~n2555;
  assign n2335 = n12024 | n12025;
  assign n12027 = ~n9978 & n2555;
  assign n12028 = P2_DATAO_REG_21_ & ~n2555;
  assign n2340 = n12027 | n12028;
  assign n12030 = ~n10031 & n2555;
  assign n12031 = P2_DATAO_REG_22_ & ~n2555;
  assign n2345 = n12030 | n12031;
  assign n12033 = ~n10085 & n2555;
  assign n12034 = P2_DATAO_REG_23_ & ~n2555;
  assign n2350 = n12033 | n12034;
  assign n12036 = ~n10141 & n2555;
  assign n12037 = P2_DATAO_REG_24_ & ~n2555;
  assign n2355 = n12036 | n12037;
  assign n12039 = ~n10195 & n2555;
  assign n12040 = P2_DATAO_REG_25_ & ~n2555;
  assign n2360 = n12039 | n12040;
  assign n12042 = ~n10253 & n2555;
  assign n12043 = P2_DATAO_REG_26_ & ~n2555;
  assign n2365 = n12042 | n12043;
  assign n12045 = ~n10305 & n2555;
  assign n12046 = P2_DATAO_REG_27_ & ~n2555;
  assign n2370 = n12045 | n12046;
  assign n12048 = ~n10359 & n2555;
  assign n12049 = P2_DATAO_REG_28_ & ~n2555;
  assign n2375 = n12048 | n12049;
  assign n12051 = ~n10409 & n2555;
  assign n12052 = P2_DATAO_REG_29_ & ~n2555;
  assign n2380 = n12051 | n12052;
  assign n12054 = ~n10503 & n2555;
  assign n12055 = P2_DATAO_REG_30_ & ~n2555;
  assign n2385 = n12054 | n12055;
  assign n12057 = ~n10523 & n2555;
  assign n12058 = P2_DATAO_REG_31_ & ~n2555;
  assign n2390 = n12057 | n12058;
  assign n12060 = ~n8569 & ~n8698;
  assign n12061 = n8722 & n8843;
  assign n12062 = n8569 & ~n12061;
  assign n12063 = ~n12060 & ~n12062;
  assign n12064 = n11006 & n12063;
  assign n12065 = P2_B_REG & ~n12064;
  assign n12066 = n8569 & ~n10031;
  assign n12067 = ~n8701 & n8717;
  assign n12068 = ~n8569 & ~n8701;
  assign n12069 = n8720 & n12068;
  assign n12070 = ~n12067 & ~n12069;
  assign n12071 = ~n10085 & ~n12070;
  assign n12072 = n8744 & ~n8782;
  assign n12073 = ~n8701 & n8742;
  assign n12074 = ~n8788 & ~n12073;
  assign n12075 = ~n8718 & n12074;
  assign n12076 = n12072 & n12075;
  assign n12077 = n10143 & ~n12076;
  assign n12078 = ~n12066 & ~n12071;
  assign n12079 = ~n12077 & n12078;
  assign n12080 = ~n10085 & ~n12076;
  assign n12081 = n10143 & ~n12070;
  assign n12082 = ~n8569 & ~n12080;
  assign n12083 = ~n12081 & n12082;
  assign n12084 = ~n12079 & n12083;
  assign n12085 = n8569 & ~n9978;
  assign n12086 = ~n10031 & ~n12070;
  assign n12087 = n10087 & ~n12076;
  assign n12088 = ~n12085 & ~n12086;
  assign n12089 = ~n12087 & n12088;
  assign n12090 = ~n10031 & ~n12076;
  assign n12091 = n10087 & ~n12070;
  assign n12092 = ~n8569 & ~n12090;
  assign n12093 = ~n12091 & n12092;
  assign n12094 = ~n12089 & n12093;
  assign n12095 = n12079 & ~n12083;
  assign n12096 = n12094 & ~n12095;
  assign n12097 = ~n12084 & ~n12096;
  assign n12098 = ~n10141 & ~n12076;
  assign n12099 = n10197 & ~n12070;
  assign n12100 = ~n8569 & ~n12098;
  assign n12101 = ~n12099 & n12100;
  assign n12102 = n8569 & ~n10085;
  assign n12103 = ~n10141 & ~n12070;
  assign n12104 = n10197 & ~n12076;
  assign n12105 = ~n12102 & ~n12103;
  assign n12106 = ~n12104 & n12105;
  assign n12107 = ~n12101 & n12106;
  assign n12108 = ~n12097 & ~n12107;
  assign n12109 = ~n9560 & ~n12076;
  assign n12110 = ~n9630 & ~n12070;
  assign n12111 = ~n8569 & ~n12109;
  assign n12112 = ~n12110 & n12111;
  assign n12113 = ~n9560 & ~n12070;
  assign n12114 = n8569 & ~n9499;
  assign n12115 = ~n9630 & ~n12076;
  assign n12116 = ~n12113 & ~n12114;
  assign n12117 = ~n12115 & n12116;
  assign n12118 = ~n12112 & n12117;
  assign n12119 = ~n9499 & ~n12076;
  assign n12120 = ~n9567 & ~n12070;
  assign n12121 = ~n8569 & ~n12119;
  assign n12122 = ~n12120 & n12121;
  assign n12123 = ~n9499 & ~n12070;
  assign n12124 = n8569 & ~n9434;
  assign n12125 = ~n9567 & ~n12076;
  assign n12126 = ~n12123 & ~n12124;
  assign n12127 = ~n12125 & n12126;
  assign n12128 = ~n12122 & n12127;
  assign n12129 = ~n8823 & ~n12070;
  assign n12130 = ~n8569 & ~n12129;
  assign n12131 = ~n8778 & ~n12076;
  assign n12132 = n12130 & ~n12131;
  assign n12133 = ~n8778 & ~n12070;
  assign n12134 = ~n8823 & ~n12076;
  assign n12135 = n8569 & ~n8762;
  assign n12136 = ~n12133 & ~n12134;
  assign n12137 = ~n12135 & n12136;
  assign n12138 = ~n12132 & n12137;
  assign n12139 = ~n8816 & ~n12070;
  assign n12140 = ~n8877 & ~n12076;
  assign n12141 = n8569 & ~n8778;
  assign n12142 = ~n12139 & ~n12140;
  assign n12143 = ~n12141 & n12142;
  assign n12144 = ~n8877 & ~n12070;
  assign n12145 = ~n8569 & ~n12144;
  assign n12146 = ~n8816 & ~n12076;
  assign n12147 = n12145 & ~n12146;
  assign n12148 = ~n12143 & n12147;
  assign n12149 = ~n8870 & ~n12070;
  assign n12150 = ~n8936 & ~n12076;
  assign n12151 = n8569 & ~n8816;
  assign n12152 = ~n12149 & ~n12150;
  assign n12153 = ~n12151 & n12152;
  assign n12154 = ~n8936 & ~n12070;
  assign n12155 = ~n8569 & ~n12154;
  assign n12156 = ~n8870 & ~n12076;
  assign n12157 = n12155 & ~n12156;
  assign n12158 = ~n12153 & n12157;
  assign n12159 = ~n12148 & ~n12158;
  assign n12160 = ~n9055 & ~n12070;
  assign n12161 = n8569 & ~n8989;
  assign n12162 = ~n9121 & ~n12076;
  assign n12163 = ~n12160 & ~n12161;
  assign n12164 = ~n12162 & n12163;
  assign n12165 = ~n9055 & ~n12076;
  assign n12166 = ~n9121 & ~n12070;
  assign n12167 = ~n8569 & ~n12165;
  assign n12168 = ~n12166 & n12167;
  assign n12169 = ~n12164 & n12168;
  assign n12170 = ~n8989 & ~n12070;
  assign n12171 = n8569 & ~n8929;
  assign n12172 = ~n9062 & ~n12076;
  assign n12173 = ~n12170 & ~n12171;
  assign n12174 = ~n12172 & n12173;
  assign n12175 = ~n8989 & ~n12076;
  assign n12176 = ~n9062 & ~n12070;
  assign n12177 = ~n8569 & ~n12175;
  assign n12178 = ~n12176 & n12177;
  assign n12179 = ~n12174 & n12178;
  assign n12180 = n12164 & ~n12168;
  assign n12181 = n12179 & ~n12180;
  assign n12182 = ~n12169 & ~n12181;
  assign n12183 = ~n8929 & ~n12070;
  assign n12184 = ~n8996 & ~n12076;
  assign n12185 = n8569 & ~n8870;
  assign n12186 = ~n12183 & ~n12184;
  assign n12187 = ~n12185 & n12186;
  assign n12188 = ~n8996 & ~n12070;
  assign n12189 = ~n8569 & ~n12188;
  assign n12190 = ~n8929 & ~n12076;
  assign n12191 = n12189 & ~n12190;
  assign n12192 = ~n12187 & n12191;
  assign n12193 = n12174 & ~n12178;
  assign n12194 = ~n12180 & ~n12193;
  assign n12195 = n12192 & n12194;
  assign n12196 = ~n9245 & ~n12070;
  assign n12197 = n8569 & ~n9181;
  assign n12198 = ~n9316 & ~n12076;
  assign n12199 = ~n12196 & ~n12197;
  assign n12200 = ~n12198 & n12199;
  assign n12201 = ~n9245 & ~n12076;
  assign n12202 = ~n9316 & ~n12070;
  assign n12203 = ~n8569 & ~n12201;
  assign n12204 = ~n12202 & n12203;
  assign n12205 = ~n12200 & n12204;
  assign n12206 = ~n9181 & ~n12070;
  assign n12207 = n8569 & ~n9114;
  assign n12208 = ~n9252 & ~n12076;
  assign n12209 = ~n12206 & ~n12207;
  assign n12210 = ~n12208 & n12209;
  assign n12211 = ~n9181 & ~n12076;
  assign n12212 = ~n9252 & ~n12070;
  assign n12213 = ~n8569 & ~n12211;
  assign n12214 = ~n12212 & n12213;
  assign n12215 = ~n12210 & n12214;
  assign n12216 = ~n12205 & ~n12215;
  assign n12217 = ~n9114 & ~n12070;
  assign n12218 = n8569 & ~n9055;
  assign n12219 = ~n9188 & ~n12076;
  assign n12220 = ~n12217 & ~n12218;
  assign n12221 = ~n12219 & n12220;
  assign n12222 = ~n9114 & ~n12076;
  assign n12223 = ~n9188 & ~n12070;
  assign n12224 = ~n8569 & ~n12222;
  assign n12225 = ~n12223 & n12224;
  assign n12226 = ~n12221 & n12225;
  assign n12227 = n12216 & ~n12226;
  assign n12228 = n12182 & ~n12195;
  assign n12229 = n12227 & n12228;
  assign n12230 = n12159 & n12229;
  assign n12231 = n12138 & n12230;
  assign n12232 = n12221 & ~n12225;
  assign n12233 = n12216 & n12232;
  assign n12234 = n12210 & ~n12214;
  assign n12235 = ~n12205 & n12234;
  assign n12236 = ~n8739 & ~n12070;
  assign n12237 = ~n8569 & ~n12236;
  assign n12238 = ~n8762 & ~n12076;
  assign n12239 = n12237 & ~n12238;
  assign n12240 = n8698 & ~n8701;
  assign n12241 = ~n8569 & n12240;
  assign n12242 = n12239 & n12241;
  assign n12243 = n12132 & ~n12137;
  assign n12244 = ~n8762 & ~n12070;
  assign n12245 = ~n8739 & ~n12076;
  assign n12246 = ~n12244 & ~n12245;
  assign n12247 = ~n12239 & ~n12241;
  assign n12248 = ~n12246 & ~n12247;
  assign n12249 = ~n12242 & ~n12243;
  assign n12250 = ~n12248 & n12249;
  assign n12251 = n12230 & n12250;
  assign n12252 = n12153 & ~n12157;
  assign n12253 = n12187 & ~n12191;
  assign n12254 = n12143 & ~n12147;
  assign n12255 = ~n12158 & n12254;
  assign n12256 = n12194 & ~n12252;
  assign n12257 = ~n12253 & n12256;
  assign n12258 = ~n12255 & n12257;
  assign n12259 = n12229 & ~n12258;
  assign n12260 = ~n9434 & ~n12076;
  assign n12261 = ~n9506 & ~n12070;
  assign n12262 = ~n8569 & ~n12260;
  assign n12263 = ~n12261 & n12262;
  assign n12264 = ~n9434 & ~n12070;
  assign n12265 = n8569 & ~n9376;
  assign n12266 = ~n9506 & ~n12076;
  assign n12267 = ~n12264 & ~n12265;
  assign n12268 = ~n12266 & n12267;
  assign n12269 = ~n12263 & n12268;
  assign n12270 = ~n9376 & ~n12076;
  assign n12271 = ~n9441 & ~n12070;
  assign n12272 = ~n8569 & ~n12270;
  assign n12273 = ~n12271 & n12272;
  assign n12274 = ~n9376 & ~n12070;
  assign n12275 = n8569 & ~n9309;
  assign n12276 = ~n9441 & ~n12076;
  assign n12277 = ~n12274 & ~n12275;
  assign n12278 = ~n12276 & n12277;
  assign n12279 = ~n12273 & n12278;
  assign n12280 = ~n12269 & ~n12279;
  assign n12281 = n12200 & ~n12204;
  assign n12282 = ~n9309 & ~n12076;
  assign n12283 = ~n9383 & ~n12070;
  assign n12284 = ~n8569 & ~n12282;
  assign n12285 = ~n12283 & n12284;
  assign n12286 = ~n9309 & ~n12070;
  assign n12287 = n8569 & ~n9245;
  assign n12288 = ~n9383 & ~n12076;
  assign n12289 = ~n12286 & ~n12287;
  assign n12290 = ~n12288 & n12289;
  assign n12291 = ~n12285 & n12290;
  assign n12292 = ~n12281 & ~n12291;
  assign n12293 = n12280 & n12292;
  assign n12294 = ~n12259 & n12293;
  assign n12295 = ~n12231 & ~n12233;
  assign n12296 = ~n12235 & n12295;
  assign n12297 = ~n12251 & n12296;
  assign n12298 = n12294 & n12297;
  assign n12299 = n12273 & ~n12278;
  assign n12300 = ~n12269 & n12299;
  assign n12301 = n12263 & ~n12268;
  assign n12302 = n12122 & ~n12127;
  assign n12303 = ~n12301 & ~n12302;
  assign n12304 = ~n12300 & n12303;
  assign n12305 = n12285 & ~n12290;
  assign n12306 = n12280 & n12305;
  assign n12307 = n12304 & ~n12306;
  assign n12308 = ~n12298 & n12307;
  assign n12309 = ~n12128 & ~n12308;
  assign n12310 = n12112 & ~n12117;
  assign n12311 = ~n12309 & ~n12310;
  assign n12312 = ~n12118 & ~n12311;
  assign n12313 = ~n9623 & ~n12070;
  assign n12314 = n8569 & ~n9560;
  assign n12315 = ~n9688 & ~n12076;
  assign n12316 = ~n12313 & ~n12314;
  assign n12317 = ~n12315 & n12316;
  assign n12318 = ~n9623 & ~n12076;
  assign n12319 = ~n9688 & ~n12070;
  assign n12320 = ~n8569 & ~n12318;
  assign n12321 = ~n12319 & n12320;
  assign n12322 = ~n12317 & n12321;
  assign n12323 = ~n9798 & ~n12070;
  assign n12324 = n8569 & ~n9737;
  assign n12325 = ~n9869 & ~n12076;
  assign n12326 = ~n12323 & ~n12324;
  assign n12327 = ~n12325 & n12326;
  assign n12328 = ~n9798 & ~n12076;
  assign n12329 = ~n9869 & ~n12070;
  assign n12330 = ~n8569 & ~n12328;
  assign n12331 = ~n12329 & n12330;
  assign n12332 = ~n12327 & n12331;
  assign n12333 = ~n9737 & ~n12070;
  assign n12334 = n8569 & ~n9681;
  assign n12335 = ~n9805 & ~n12076;
  assign n12336 = ~n12333 & ~n12334;
  assign n12337 = ~n12335 & n12336;
  assign n12338 = ~n9737 & ~n12076;
  assign n12339 = ~n9805 & ~n12070;
  assign n12340 = ~n8569 & ~n12338;
  assign n12341 = ~n12339 & n12340;
  assign n12342 = ~n12337 & n12341;
  assign n12343 = n12327 & ~n12331;
  assign n12344 = n12342 & ~n12343;
  assign n12345 = ~n12332 & ~n12344;
  assign n12346 = ~n9681 & ~n12070;
  assign n12347 = n8569 & ~n9623;
  assign n12348 = ~n9744 & ~n12076;
  assign n12349 = ~n12346 & ~n12347;
  assign n12350 = ~n12348 & n12349;
  assign n12351 = ~n9681 & ~n12076;
  assign n12352 = ~n9744 & ~n12070;
  assign n12353 = ~n8569 & ~n12351;
  assign n12354 = ~n12352 & n12353;
  assign n12355 = ~n12350 & n12354;
  assign n12356 = n12337 & ~n12341;
  assign n12357 = ~n12343 & ~n12356;
  assign n12358 = n12355 & n12357;
  assign n12359 = ~n9862 & ~n12070;
  assign n12360 = n8569 & ~n9798;
  assign n12361 = ~n9926 & ~n12076;
  assign n12362 = ~n12359 & ~n12360;
  assign n12363 = ~n12361 & n12362;
  assign n12364 = ~n9862 & ~n12076;
  assign n12365 = ~n9926 & ~n12070;
  assign n12366 = ~n8569 & ~n12364;
  assign n12367 = ~n12365 & n12366;
  assign n12368 = ~n12363 & n12367;
  assign n12369 = n8569 & ~n9922;
  assign n12370 = ~n9978 & ~n12070;
  assign n12371 = n10033 & ~n12076;
  assign n12372 = ~n12369 & ~n12370;
  assign n12373 = ~n12371 & n12372;
  assign n12374 = ~n9978 & ~n12076;
  assign n12375 = n10033 & ~n12070;
  assign n12376 = ~n8569 & ~n12374;
  assign n12377 = ~n12375 & n12376;
  assign n12378 = ~n12373 & n12377;
  assign n12379 = n8569 & ~n9862;
  assign n12380 = ~n9922 & ~n12070;
  assign n12381 = n9980 & ~n12076;
  assign n12382 = ~n12379 & ~n12380;
  assign n12383 = ~n12381 & n12382;
  assign n12384 = ~n9922 & ~n12076;
  assign n12385 = n9980 & ~n12070;
  assign n12386 = ~n8569 & ~n12384;
  assign n12387 = ~n12385 & n12386;
  assign n12388 = ~n12383 & n12387;
  assign n12389 = ~n12378 & ~n12388;
  assign n12390 = n12345 & ~n12358;
  assign n12391 = ~n12368 & n12390;
  assign n12392 = n12389 & n12391;
  assign n12393 = ~n12312 & ~n12322;
  assign n12394 = n12392 & n12393;
  assign n12395 = n12317 & ~n12321;
  assign n12396 = n12350 & ~n12354;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = n12357 & n12397;
  assign n12399 = n12392 & ~n12398;
  assign n12400 = n12089 & ~n12093;
  assign n12401 = n12373 & ~n12377;
  assign n12402 = ~n12400 & ~n12401;
  assign n12403 = n12363 & ~n12367;
  assign n12404 = n12389 & n12403;
  assign n12405 = n12383 & ~n12387;
  assign n12406 = ~n12378 & n12405;
  assign n12407 = ~n12404 & ~n12406;
  assign n12408 = ~n12095 & n12407;
  assign n12409 = ~n12394 & ~n12399;
  assign n12410 = n12402 & n12409;
  assign n12411 = n12408 & n12410;
  assign n12412 = ~n12107 & n12411;
  assign n12413 = n12101 & ~n12106;
  assign n12414 = n8569 & ~n10141;
  assign n12415 = ~n10195 & ~n12070;
  assign n12416 = n10255 & ~n12076;
  assign n12417 = ~n12414 & ~n12415;
  assign n12418 = ~n12416 & n12417;
  assign n12419 = ~n10195 & ~n12076;
  assign n12420 = n10255 & ~n12070;
  assign n12421 = ~n8569 & ~n12419;
  assign n12422 = ~n12420 & n12421;
  assign n12423 = ~n12418 & n12422;
  assign n12424 = ~n12413 & ~n12423;
  assign n12425 = n8569 & ~n10195;
  assign n12426 = ~n10253 & ~n12070;
  assign n12427 = n10307 & ~n12076;
  assign n12428 = ~n12425 & ~n12426;
  assign n12429 = ~n12427 & n12428;
  assign n12430 = ~n10253 & ~n12076;
  assign n12431 = n10307 & ~n12070;
  assign n12432 = ~n8569 & ~n12430;
  assign n12433 = ~n12431 & n12432;
  assign n12434 = ~n12429 & n12433;
  assign n12435 = n8569 & ~n10253;
  assign n12436 = ~n10305 & ~n12070;
  assign n12437 = n10361 & ~n12076;
  assign n12438 = ~n12435 & ~n12436;
  assign n12439 = ~n12437 & n12438;
  assign n12440 = ~n10305 & ~n12076;
  assign n12441 = n10361 & ~n12070;
  assign n12442 = ~n8569 & ~n12440;
  assign n12443 = ~n12441 & n12442;
  assign n12444 = ~n12439 & n12443;
  assign n12445 = n8569 & ~n10305;
  assign n12446 = ~n10359 & ~n12070;
  assign n12447 = n10411 & ~n12076;
  assign n12448 = ~n12445 & ~n12446;
  assign n12449 = ~n12447 & n12448;
  assign n12450 = ~n10359 & ~n12076;
  assign n12451 = n10411 & ~n12070;
  assign n12452 = ~n8569 & ~n12450;
  assign n12453 = ~n12451 & n12452;
  assign n12454 = ~n12449 & n12453;
  assign n12455 = ~n12434 & ~n12444;
  assign n12456 = ~n12454 & n12455;
  assign n12457 = ~n10523 & ~n12076;
  assign n12458 = n10531 & ~n12070;
  assign n12459 = ~n12457 & ~n12458;
  assign n12460 = n10531 & ~n12076;
  assign n12461 = ~n10523 & ~n12070;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~n12459 & n12462;
  assign n12464 = n12459 & ~n12462;
  assign n12465 = ~n12463 & ~n12464;
  assign n12466 = ~n12108 & ~n12412;
  assign n12467 = n12424 & n12466;
  assign n12468 = n12456 & n12467;
  assign n12469 = n12465 & n12468;
  assign n12470 = n8569 & ~n10359;
  assign n12471 = ~n10409 & ~n12070;
  assign n12472 = n10461 & ~n12076;
  assign n12473 = ~n12470 & ~n12471;
  assign n12474 = ~n12472 & n12473;
  assign n12475 = ~n10409 & ~n12076;
  assign n12476 = n10461 & ~n12070;
  assign n12477 = ~n8569 & ~n12475;
  assign n12478 = ~n12476 & n12477;
  assign n12479 = ~n12474 & n12478;
  assign n12480 = n10525 & ~n12076;
  assign n12481 = ~n10503 & ~n12070;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = ~n12479 & n12482;
  assign n12484 = ~n10503 & ~n12076;
  assign n12485 = n10525 & ~n12070;
  assign n12486 = ~n12484 & ~n12485;
  assign n12487 = ~n12479 & ~n12486;
  assign n12488 = ~n12483 & ~n12487;
  assign n12489 = n12469 & ~n12488;
  assign n12490 = n12474 & ~n12478;
  assign n12491 = ~n12482 & n12486;
  assign n12492 = n12465 & n12490;
  assign n12493 = ~n12491 & n12492;
  assign n12494 = n12429 & ~n12433;
  assign n12495 = n12456 & n12494;
  assign n12496 = n12465 & n12495;
  assign n12497 = ~n12488 & n12496;
  assign n12498 = n12418 & ~n12422;
  assign n12499 = n12456 & n12498;
  assign n12500 = n12465 & n12499;
  assign n12501 = ~n12488 & n12500;
  assign n12502 = ~n12497 & ~n12501;
  assign n12503 = n12449 & ~n12453;
  assign n12504 = n12465 & n12503;
  assign n12505 = ~n12488 & n12504;
  assign n12506 = n12439 & ~n12443;
  assign n12507 = ~n12454 & n12506;
  assign n12508 = n12465 & n12507;
  assign n12509 = ~n12488 & n12508;
  assign n12510 = n12465 & n12482;
  assign n12511 = ~n12486 & n12510;
  assign n12512 = n8569 & ~n8701;
  assign n12513 = n8720 & n12512;
  assign n12514 = n12462 & ~n12513;
  assign n12515 = n12459 & n12513;
  assign n12516 = ~n12459 & ~n12462;
  assign n12517 = ~n12514 & ~n12515;
  assign n12518 = ~n12516 & n12517;
  assign n12519 = ~n12511 & ~n12518;
  assign n12520 = ~n12505 & ~n12509;
  assign n12521 = n12519 & n12520;
  assign n12522 = ~n12489 & ~n12493;
  assign n12523 = n12502 & n12522;
  assign n12524 = n12521 & n12523;
  assign n12525 = n8582 & n12061;
  assign n12526 = n12524 & n12525;
  assign n12527 = n8569 & ~n12065;
  assign n12528 = ~n12526 & n12527;
  assign n12529 = ~P2_STATE_REG & ~n12065;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = n8739 & n8762;
  assign n12532 = ~n8837 & ~n12531;
  assign n12533 = ~n8836 & ~n12532;
  assign n12534 = ~n9701 & ~n9702;
  assign n12535 = ~n9583 & ~n9584;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = ~n9276 & ~n9342;
  assign n12538 = n12533 & n12536;
  assign n12539 = n12537 & n12538;
  assign n12540 = ~n9891 & n12539;
  assign n12541 = ~n9075 & ~n9076;
  assign n12542 = ~n9206 & ~n9207;
  assign n12543 = ~n8894 & ~n12541;
  assign n12544 = ~n12542 & n12543;
  assign n12545 = ~n9767 & n12544;
  assign n12546 = ~n9760 & ~n9761;
  assign n12547 = ~n9150 & ~n9529;
  assign n12548 = ~n12546 & n12547;
  assign n12549 = ~n9823 & ~n9824;
  assign n12550 = n12545 & n12548;
  assign n12551 = ~n12549 & n12550;
  assign n12552 = ~n10215 & ~n10216;
  assign n12553 = n10253 & ~n10307;
  assign n12554 = ~n10321 & ~n12553;
  assign n12555 = ~n10222 & ~n12552;
  assign n12556 = ~n10273 & n12555;
  assign n12557 = ~n12554 & n12556;
  assign n12558 = n10503 & ~n10525;
  assign n12559 = ~n10503 & n10525;
  assign n12560 = ~n12558 & ~n12559;
  assign n12561 = n12540 & n12551;
  assign n12562 = ~n9946 & n12561;
  assign n12563 = n12557 & n12562;
  assign n12564 = ~n12560 & n12563;
  assign n12565 = ~n9396 & ~n9397;
  assign n12566 = ~n9022 & ~n12565;
  assign n12567 = ~n9467 & n12566;
  assign n12568 = ~n8958 & n12567;
  assign n12569 = ~n9993 & ~n9994;
  assign n12570 = ~n10100 & ~n10104;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = ~n10159 & ~n10160;
  assign n12573 = n10409 & ~n10461;
  assign n12574 = ~n10409 & n10461;
  assign n12575 = ~n12573 & ~n12574;
  assign n12576 = n10359 & ~n10411;
  assign n12577 = ~n10484 & ~n12576;
  assign n12578 = ~n10429 & ~n10435;
  assign n12579 = n10523 & ~n10531;
  assign n12580 = ~n10523 & n10531;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = ~n12577 & ~n12578;
  assign n12583 = ~n12581 & n12582;
  assign n12584 = n12568 & n12571;
  assign n12585 = ~n12572 & n12584;
  assign n12586 = ~n12575 & n12585;
  assign n12587 = n12583 & n12586;
  assign n12588 = n12564 & n12587;
  assign n12589 = ~n8711 & ~n12588;
  assign n12590 = n8711 & n12588;
  assign n12591 = ~n12589 & ~n12590;
  assign n12592 = n8701 & ~n12591;
  assign n12593 = ~n8704 & n12592;
  assign n12594 = n8711 & n8768;
  assign n12595 = ~n8711 & ~n8768;
  assign n12596 = ~n12594 & ~n12595;
  assign n12597 = n12524 & ~n12596;
  assign n12598 = ~n12524 & n12596;
  assign n12599 = ~n12597 & ~n12598;
  assign n12600 = n8704 & n12599;
  assign n12601 = ~n10503 & n10523;
  assign n12602 = ~n10523 & ~n12601;
  assign n12603 = n10503 & ~n10523;
  assign n12604 = ~n12601 & ~n12603;
  assign n12605 = n12601 & n12604;
  assign n12606 = ~n12602 & ~n12605;
  assign n12607 = n10531 & n12606;
  assign n12608 = ~n10531 & ~n12606;
  assign n12609 = ~n10525 & ~n12608;
  assign n12610 = ~n10503 & ~n12601;
  assign n12611 = n10503 & n12601;
  assign n12612 = ~n12610 & ~n12611;
  assign n12613 = ~n12608 & ~n12612;
  assign n12614 = ~n12609 & ~n12613;
  assign n12615 = ~n10359 & ~n12601;
  assign n12616 = ~n10359 & n12601;
  assign n12617 = ~n12615 & ~n12616;
  assign n12618 = ~n10411 & ~n12617;
  assign n12619 = ~n10409 & ~n12601;
  assign n12620 = ~n10409 & n12601;
  assign n12621 = ~n12619 & ~n12620;
  assign n12622 = n10461 & n12621;
  assign n12623 = n12618 & ~n12622;
  assign n12624 = ~n12614 & n12623;
  assign n12625 = ~n12607 & ~n12624;
  assign n12626 = ~n9623 & ~n12601;
  assign n12627 = ~n9623 & n12601;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = n9688 & ~n12628;
  assign n12630 = ~n9560 & ~n12601;
  assign n12631 = ~n9560 & n12601;
  assign n12632 = ~n12630 & ~n12631;
  assign n12633 = n9630 & ~n12632;
  assign n12634 = ~n9181 & ~n12601;
  assign n12635 = ~n9181 & n12601;
  assign n12636 = ~n12634 & ~n12635;
  assign n12637 = ~n9252 & n12636;
  assign n12638 = ~n9114 & ~n12601;
  assign n12639 = ~n9114 & n12601;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n9188 & n12640;
  assign n12642 = ~n9245 & ~n12601;
  assign n12643 = ~n9245 & n12601;
  assign n12644 = ~n12642 & ~n12643;
  assign n12645 = ~n9316 & n12644;
  assign n12646 = ~n9309 & ~n12601;
  assign n12647 = ~n9309 & n12601;
  assign n12648 = ~n12646 & ~n12647;
  assign n12649 = ~n9383 & n12648;
  assign n12650 = ~n12637 & ~n12641;
  assign n12651 = ~n12645 & n12650;
  assign n12652 = ~n12649 & n12651;
  assign n12653 = ~n9055 & ~n12601;
  assign n12654 = ~n9055 & n12601;
  assign n12655 = ~n12653 & ~n12654;
  assign n12656 = n9121 & ~n12655;
  assign n12657 = n9188 & ~n12640;
  assign n12658 = ~n12656 & ~n12657;
  assign n12659 = ~n8989 & ~n12601;
  assign n12660 = ~n8989 & n12601;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = ~n9062 & n12661;
  assign n12663 = ~n9121 & n12655;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = n9062 & ~n12661;
  assign n12666 = ~n8929 & ~n12601;
  assign n12667 = ~n8929 & n12601;
  assign n12668 = ~n12666 & ~n12667;
  assign n12669 = n8996 & ~n12668;
  assign n12670 = ~n12665 & ~n12669;
  assign n12671 = n12664 & ~n12670;
  assign n12672 = n12658 & ~n12671;
  assign n12673 = n12652 & ~n12672;
  assign n12674 = ~n8870 & ~n12601;
  assign n12675 = ~n8870 & n12601;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = n8936 & ~n12676;
  assign n12678 = ~n8996 & n12668;
  assign n12679 = n12664 & ~n12678;
  assign n12680 = n12652 & n12679;
  assign n12681 = n12677 & n12680;
  assign n12682 = n9383 & ~n12648;
  assign n12683 = ~n12645 & ~n12649;
  assign n12684 = n9316 & ~n12644;
  assign n12685 = n9252 & ~n12636;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = n12683 & ~n12686;
  assign n12688 = ~n9499 & ~n12601;
  assign n12689 = ~n9499 & n12601;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = n9567 & ~n12690;
  assign n12692 = ~n9434 & ~n12601;
  assign n12693 = ~n9434 & n12601;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = n9506 & ~n12694;
  assign n12696 = ~n12691 & ~n12695;
  assign n12697 = ~n9376 & ~n12601;
  assign n12698 = ~n9376 & n12601;
  assign n12699 = ~n12697 & ~n12698;
  assign n12700 = n9441 & ~n12699;
  assign n12701 = n12696 & ~n12700;
  assign n12702 = ~n12682 & ~n12687;
  assign n12703 = n12701 & n12702;
  assign n12704 = ~n8816 & ~n12601;
  assign n12705 = ~n8816 & n12601;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = n8877 & ~n12706;
  assign n12708 = ~n8936 & n12676;
  assign n12709 = n12680 & ~n12708;
  assign n12710 = n12707 & n12709;
  assign n12711 = ~n8877 & n12706;
  assign n12712 = ~n8778 & ~n12601;
  assign n12713 = ~n8778 & n12601;
  assign n12714 = ~n12712 & ~n12713;
  assign n12715 = ~n8823 & n12714;
  assign n12716 = ~n12711 & ~n12715;
  assign n12717 = ~n8762 & ~n12601;
  assign n12718 = ~n8762 & n12601;
  assign n12719 = ~n12717 & ~n12718;
  assign n12720 = ~n8739 & n12719;
  assign n12721 = n8823 & ~n12714;
  assign n12722 = n12720 & ~n12721;
  assign n12723 = n12716 & ~n12722;
  assign n12724 = n12709 & n12723;
  assign n12725 = ~n12673 & ~n12681;
  assign n12726 = n12703 & n12725;
  assign n12727 = ~n12710 & n12726;
  assign n12728 = ~n12724 & n12727;
  assign n12729 = ~n9506 & n12694;
  assign n12730 = ~n12691 & n12729;
  assign n12731 = ~n9567 & n12690;
  assign n12732 = ~n9630 & n12632;
  assign n12733 = ~n12731 & ~n12732;
  assign n12734 = ~n12730 & n12733;
  assign n12735 = ~n9441 & n12699;
  assign n12736 = n12696 & n12735;
  assign n12737 = n12734 & ~n12736;
  assign n12738 = ~n12728 & n12737;
  assign n12739 = ~n12633 & ~n12738;
  assign n12740 = ~n9688 & n12628;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = ~n12629 & ~n12741;
  assign n12743 = ~n9681 & ~n12601;
  assign n12744 = ~n9681 & n12601;
  assign n12745 = ~n12743 & ~n12744;
  assign n12746 = ~n9744 & n12745;
  assign n12747 = ~n9862 & ~n12601;
  assign n12748 = ~n9862 & n12601;
  assign n12749 = ~n12747 & ~n12748;
  assign n12750 = ~n9926 & n12749;
  assign n12751 = ~n9798 & ~n12601;
  assign n12752 = ~n9798 & n12601;
  assign n12753 = ~n12751 & ~n12752;
  assign n12754 = ~n9869 & n12753;
  assign n12755 = n9926 & ~n12749;
  assign n12756 = n12754 & ~n12755;
  assign n12757 = ~n12750 & ~n12756;
  assign n12758 = ~n9737 & ~n12601;
  assign n12759 = ~n9737 & n12601;
  assign n12760 = ~n12758 & ~n12759;
  assign n12761 = ~n9805 & n12760;
  assign n12762 = n9869 & ~n12753;
  assign n12763 = ~n12755 & ~n12762;
  assign n12764 = n12761 & n12763;
  assign n12765 = ~n9922 & ~n12601;
  assign n12766 = ~n9922 & n12601;
  assign n12767 = ~n12765 & ~n12766;
  assign n12768 = n9980 & n12767;
  assign n12769 = ~n10031 & ~n12601;
  assign n12770 = ~n10031 & n12601;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = n10087 & n12771;
  assign n12773 = ~n9978 & ~n12601;
  assign n12774 = ~n9978 & n12601;
  assign n12775 = ~n12773 & ~n12774;
  assign n12776 = n10033 & n12775;
  assign n12777 = ~n12772 & ~n12776;
  assign n12778 = n12757 & ~n12764;
  assign n12779 = ~n12768 & n12778;
  assign n12780 = n12777 & n12779;
  assign n12781 = ~n12742 & ~n12746;
  assign n12782 = n12780 & n12781;
  assign n12783 = n9744 & ~n12745;
  assign n12784 = n9805 & ~n12760;
  assign n12785 = ~n12783 & ~n12784;
  assign n12786 = n12763 & n12785;
  assign n12787 = n12780 & ~n12786;
  assign n12788 = ~n10085 & ~n12601;
  assign n12789 = ~n10085 & n12601;
  assign n12790 = ~n12788 & ~n12789;
  assign n12791 = ~n10143 & ~n12790;
  assign n12792 = ~n10087 & ~n12771;
  assign n12793 = ~n12791 & ~n12792;
  assign n12794 = ~n9980 & ~n12767;
  assign n12795 = n12777 & n12794;
  assign n12796 = ~n10033 & ~n12775;
  assign n12797 = ~n12772 & n12796;
  assign n12798 = ~n10141 & ~n12601;
  assign n12799 = ~n10141 & n12601;
  assign n12800 = ~n12798 & ~n12799;
  assign n12801 = ~n10197 & ~n12800;
  assign n12802 = ~n10195 & ~n12601;
  assign n12803 = ~n10195 & n12601;
  assign n12804 = ~n12802 & ~n12803;
  assign n12805 = ~n10255 & ~n12804;
  assign n12806 = ~n12795 & ~n12797;
  assign n12807 = ~n12801 & n12806;
  assign n12808 = ~n12805 & n12807;
  assign n12809 = ~n12782 & ~n12787;
  assign n12810 = n12793 & n12809;
  assign n12811 = n12808 & n12810;
  assign n12812 = n10197 & n12800;
  assign n12813 = n10143 & n12790;
  assign n12814 = ~n12812 & ~n12813;
  assign n12815 = ~n12801 & ~n12814;
  assign n12816 = ~n12805 & n12815;
  assign n12817 = ~n10253 & ~n12601;
  assign n12818 = ~n10253 & n12601;
  assign n12819 = ~n12817 & ~n12818;
  assign n12820 = n10307 & n12819;
  assign n12821 = n10255 & n12804;
  assign n12822 = ~n12820 & ~n12821;
  assign n12823 = ~n10305 & ~n12601;
  assign n12824 = ~n10305 & n12601;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = n10361 & n12825;
  assign n12827 = n10411 & n12617;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = ~n12622 & n12828;
  assign n12830 = n12822 & n12829;
  assign n12831 = ~n12811 & ~n12816;
  assign n12832 = ~n12614 & n12831;
  assign n12833 = n12830 & n12832;
  assign n12834 = ~n12825 & n12829;
  assign n12835 = ~n12614 & n12834;
  assign n12836 = ~n10361 & n12835;
  assign n12837 = ~n10461 & ~n12621;
  assign n12838 = ~n12614 & n12837;
  assign n12839 = ~n10525 & n12613;
  assign n12840 = ~n12819 & n12829;
  assign n12841 = ~n12614 & n12840;
  assign n12842 = ~n10307 & n12841;
  assign n12843 = ~n12836 & ~n12838;
  assign n12844 = ~n12839 & n12843;
  assign n12845 = ~n12842 & n12844;
  assign n12846 = n12625 & ~n12833;
  assign n12847 = n12845 & n12846;
  assign n12848 = n8786 & n12847;
  assign n12849 = n8792 & ~n12847;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = ~n12065 & n12850;
  assign n12852 = ~n12526 & n12851;
  assign n12853 = ~n12593 & ~n12600;
  assign n12854 = n12852 & n12853;
  assign n2395 = n12530 & ~n12854;
  assign n12856 = n8582 & ~n10663;
  assign n12857 = ~n8716 & n12856;
  assign n12858 = n8704 & n8718;
  assign n12859 = ~n8783 & ~n12073;
  assign n12860 = ~n10546 & n12859;
  assign n12861 = ~n12858 & n12860;
  assign n12862 = ~n8788 & n12861;
  assign n12863 = ~n8716 & ~n12862;
  assign n12864 = ~n8695 & n8719;
  assign n12865 = ~n8704 & n8768;
  assign n12866 = n8581 & ~n12865;
  assign n12867 = ~n12067 & n12866;
  assign n12868 = ~n12863 & ~n12864;
  assign n12869 = n12867 & n12868;
  assign n12870 = P2_STATE_REG & ~n12869;
  assign n12871 = ~n12857 & ~n12870;
  assign n12872 = ~n9616 & ~n12871;
  assign n12873 = n8716 & n12856;
  assign n12874 = n8582 & n10653;
  assign n12875 = ~n12873 & ~n12874;
  assign n12876 = ~n9688 & ~n12875;
  assign n12877 = n8582 & n8722;
  assign n12878 = n8695 & ~n8770;
  assign n12879 = ~n9681 & n12878;
  assign n12880 = n8695 & ~n8844;
  assign n12881 = ~n9560 & n12880;
  assign n12882 = ~n8695 & ~n9616;
  assign n12883 = ~n12879 & ~n12881;
  assign n12884 = ~n12882 & n12883;
  assign n12885 = n12877 & ~n12884;
  assign n12886 = ~n11484 & ~n12885;
  assign n12887 = ~n8634 & n8701;
  assign n12888 = ~n8704 & n12887;
  assign n12889 = n8704 & n8711;
  assign n12890 = ~n12888 & ~n12889;
  assign n12891 = ~n10647 & n12890;
  assign n12892 = ~n9383 & n12891;
  assign n12893 = n9383 & ~n12891;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = ~n9309 & ~n12894;
  assign n12896 = ~n9506 & n12891;
  assign n12897 = n9506 & ~n12891;
  assign n12898 = ~n12896 & ~n12897;
  assign n12899 = n9434 & n12898;
  assign n12900 = ~n9567 & n12891;
  assign n12901 = n9567 & ~n12891;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = n9499 & n12902;
  assign n12904 = ~n12899 & ~n12903;
  assign n12905 = ~n9441 & n12891;
  assign n12906 = n9441 & ~n12891;
  assign n12907 = ~n12905 & ~n12906;
  assign n12908 = n9376 & n12907;
  assign n12909 = n12904 & ~n12908;
  assign n12910 = n12895 & n12909;
  assign n12911 = ~n9499 & ~n12902;
  assign n12912 = ~n9434 & ~n12898;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = ~n9376 & ~n12907;
  assign n12915 = n12904 & n12914;
  assign n12916 = n12913 & ~n12915;
  assign n12917 = ~n12903 & ~n12916;
  assign n12918 = ~n12910 & ~n12917;
  assign n12919 = ~n9630 & n12891;
  assign n12920 = n9630 & ~n12891;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = n9560 & n12921;
  assign n12923 = ~n12918 & ~n12922;
  assign n12924 = ~n9560 & ~n12921;
  assign n12925 = ~n12923 & ~n12924;
  assign n12926 = n9309 & n12894;
  assign n12927 = n12909 & ~n12926;
  assign n12928 = ~n12922 & n12927;
  assign n12929 = ~n9121 & n12891;
  assign n12930 = n9121 & ~n12891;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = ~n9055 & ~n12931;
  assign n12933 = ~n9114 & n12932;
  assign n12934 = ~n9188 & n12891;
  assign n12935 = n9188 & ~n12891;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = n9114 & ~n12932;
  assign n12938 = ~n12936 & ~n12937;
  assign n12939 = ~n9062 & n12891;
  assign n12940 = n9062 & ~n12891;
  assign n12941 = ~n12939 & ~n12940;
  assign n12942 = ~n8989 & ~n12941;
  assign n12943 = n9055 & n12931;
  assign n12944 = n9114 & n12936;
  assign n12945 = ~n12943 & ~n12944;
  assign n12946 = n12942 & n12945;
  assign n12947 = ~n12933 & ~n12938;
  assign n12948 = ~n12946 & n12947;
  assign n12949 = ~n9252 & n12891;
  assign n12950 = n9252 & ~n12891;
  assign n12951 = ~n12949 & ~n12950;
  assign n12952 = n9181 & n12951;
  assign n12953 = ~n12948 & ~n12952;
  assign n12954 = ~n9181 & ~n12951;
  assign n12955 = ~n12953 & ~n12954;
  assign n12956 = n8989 & n12941;
  assign n12957 = n12945 & ~n12956;
  assign n12958 = ~n12952 & n12957;
  assign n12959 = ~n8877 & n12891;
  assign n12960 = n8877 & ~n12891;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = ~n8816 & ~n12961;
  assign n12963 = ~n8870 & n12962;
  assign n12964 = ~n8936 & n12891;
  assign n12965 = n8936 & ~n12891;
  assign n12966 = ~n12964 & ~n12965;
  assign n12967 = n8870 & ~n12962;
  assign n12968 = ~n12966 & ~n12967;
  assign n12969 = ~n12963 & ~n12968;
  assign n12970 = n8816 & n12961;
  assign n12971 = n8870 & n12966;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = ~n8739 & n12891;
  assign n12974 = n8739 & ~n12891;
  assign n12975 = ~n12973 & ~n12974;
  assign n12976 = ~n12891 & ~n12975;
  assign n12977 = ~n8823 & n12891;
  assign n12978 = n8823 & ~n12891;
  assign n12979 = ~n12977 & ~n12978;
  assign n12980 = n8778 & n12979;
  assign n12981 = n12976 & ~n12980;
  assign n12982 = ~n8778 & ~n12979;
  assign n12983 = n12891 & n12975;
  assign n12984 = ~n8762 & ~n12983;
  assign n12985 = ~n12980 & n12984;
  assign n12986 = ~n12981 & ~n12982;
  assign n12987 = ~n12985 & n12986;
  assign n12988 = n12972 & ~n12987;
  assign n12989 = n12969 & ~n12988;
  assign n12990 = ~n8929 & ~n12989;
  assign n12991 = ~n8996 & n12891;
  assign n12992 = n8996 & ~n12891;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = ~n12989 & ~n12993;
  assign n12995 = ~n8929 & ~n12993;
  assign n12996 = ~n12990 & ~n12994;
  assign n12997 = ~n12995 & n12996;
  assign n12998 = n12958 & ~n12997;
  assign n12999 = n12955 & ~n12998;
  assign n13000 = ~n9245 & ~n12999;
  assign n13001 = ~n9316 & n12891;
  assign n13002 = n9316 & ~n12891;
  assign n13003 = ~n13001 & ~n13002;
  assign n13004 = ~n12999 & ~n13003;
  assign n13005 = ~n9245 & ~n13003;
  assign n13006 = ~n13000 & ~n13004;
  assign n13007 = ~n13005 & n13006;
  assign n13008 = n12928 & ~n13007;
  assign n13009 = n12925 & ~n13008;
  assign n13010 = ~n9688 & n12891;
  assign n13011 = n9688 & ~n12891;
  assign n13012 = ~n13010 & ~n13011;
  assign n13013 = n9623 & ~n13012;
  assign n13014 = ~n9623 & n13012;
  assign n13015 = ~n13013 & ~n13014;
  assign n13016 = n13009 & ~n13015;
  assign n13017 = ~n13009 & n13015;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = n8695 & n8719;
  assign n13020 = n8716 & ~n12862;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = n8582 & ~n13021;
  assign n13023 = ~n13018 & n13022;
  assign n13024 = ~n12872 & ~n12876;
  assign n13025 = n12886 & n13024;
  assign n2400 = n13023 | ~n13025;
  assign n13027 = ~n8716 & ~n10663;
  assign n13028 = n12869 & ~n13027;
  assign n13029 = P2_STATE_REG & ~n13028;
  assign n13030 = ~n10246 & n13029;
  assign n13031 = P2_REG3_REG_26_ & ~P2_STATE_REG;
  assign n13032 = ~n10305 & n12878;
  assign n13033 = ~n10195 & n12880;
  assign n13034 = ~n8695 & ~n10246;
  assign n13035 = ~n13032 & ~n13033;
  assign n13036 = ~n13034 & n13035;
  assign n13037 = n12877 & ~n13036;
  assign n13038 = ~n13031 & ~n13037;
  assign n13039 = n8716 & ~n10663;
  assign n13040 = ~n10653 & ~n13039;
  assign n13041 = n8582 & ~n13040;
  assign n13042 = n10307 & n13041;
  assign n13043 = n10255 & n12891;
  assign n13044 = ~n10255 & ~n12891;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = n10195 & n13045;
  assign n13047 = n10307 & n12891;
  assign n13048 = ~n10307 & ~n12891;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = n10253 & ~n13049;
  assign n13051 = ~n10253 & n13049;
  assign n13052 = ~n13050 & ~n13051;
  assign n13053 = n13046 & n13052;
  assign n13054 = ~n10253 & ~n13049;
  assign n13055 = ~n10195 & ~n13045;
  assign n13056 = ~n13054 & n13055;
  assign n13057 = ~n10253 & ~n13046;
  assign n13058 = ~n13046 & ~n13049;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = n13056 & ~n13059;
  assign n13061 = ~n13053 & ~n13060;
  assign n13062 = ~n13054 & ~n13059;
  assign n13063 = n10197 & n12891;
  assign n13064 = ~n10197 & ~n12891;
  assign n13065 = ~n13063 & ~n13064;
  assign n13066 = n10141 & n13065;
  assign n13067 = n10143 & n12891;
  assign n13068 = ~n10143 & ~n12891;
  assign n13069 = ~n13067 & ~n13068;
  assign n13070 = ~n10085 & ~n13069;
  assign n13071 = n10085 & n13069;
  assign n13072 = n10087 & n12891;
  assign n13073 = ~n10087 & ~n12891;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = ~n10031 & ~n13074;
  assign n13076 = n10031 & n13074;
  assign n13077 = n10033 & n12891;
  assign n13078 = ~n10033 & ~n12891;
  assign n13079 = ~n13077 & ~n13078;
  assign n13080 = n9978 & n13079;
  assign n13081 = ~n9978 & ~n13079;
  assign n13082 = n9980 & n12891;
  assign n13083 = ~n9980 & ~n12891;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = ~n9922 & ~n13084;
  assign n13086 = ~n13081 & ~n13085;
  assign n13087 = ~n9926 & n12891;
  assign n13088 = n9926 & ~n12891;
  assign n13089 = ~n13087 & ~n13088;
  assign n13090 = ~n9862 & ~n13089;
  assign n13091 = n9922 & n13084;
  assign n13092 = ~n13080 & ~n13091;
  assign n13093 = n13090 & n13092;
  assign n13094 = n13086 & ~n13093;
  assign n13095 = ~n13080 & ~n13094;
  assign n13096 = n9862 & n13089;
  assign n13097 = n13092 & ~n13096;
  assign n13098 = ~n9869 & n12891;
  assign n13099 = n9869 & ~n12891;
  assign n13100 = ~n13098 & ~n13099;
  assign n13101 = ~n9798 & ~n13100;
  assign n13102 = n9798 & n13100;
  assign n13103 = ~n9744 & n12891;
  assign n13104 = n9744 & ~n12891;
  assign n13105 = ~n13103 & ~n13104;
  assign n13106 = ~n9681 & ~n13105;
  assign n13107 = ~n9737 & n13106;
  assign n13108 = ~n9805 & n12891;
  assign n13109 = n9805 & ~n12891;
  assign n13110 = ~n13108 & ~n13109;
  assign n13111 = n9737 & ~n13106;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = ~n13107 & ~n13112;
  assign n13114 = n9681 & n13105;
  assign n13115 = n9737 & n13110;
  assign n13116 = ~n13114 & ~n13115;
  assign n13117 = n9623 & n13012;
  assign n13118 = ~n12925 & ~n13117;
  assign n13119 = ~n9623 & ~n13012;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = n12928 & ~n13117;
  assign n13122 = ~n13007 & n13121;
  assign n13123 = n13120 & ~n13122;
  assign n13124 = n13116 & ~n13123;
  assign n13125 = n13113 & ~n13124;
  assign n13126 = ~n13102 & ~n13125;
  assign n13127 = ~n13101 & ~n13126;
  assign n13128 = n13097 & ~n13127;
  assign n13129 = ~n13095 & ~n13128;
  assign n13130 = ~n13076 & ~n13129;
  assign n13131 = ~n13075 & ~n13130;
  assign n13132 = ~n13071 & ~n13131;
  assign n13133 = ~n13070 & ~n13132;
  assign n13134 = ~n13066 & ~n13133;
  assign n13135 = n13062 & n13134;
  assign n13136 = ~n10141 & ~n13065;
  assign n13137 = n13062 & n13136;
  assign n13138 = n13052 & ~n13055;
  assign n13139 = ~n13134 & n13138;
  assign n13140 = ~n13136 & n13139;
  assign n13141 = n13061 & ~n13135;
  assign n13142 = ~n13137 & n13141;
  assign n13143 = ~n13140 & n13142;
  assign n13144 = n13022 & n13143;
  assign n13145 = ~n13030 & n13038;
  assign n13146 = ~n13042 & n13145;
  assign n2405 = n13144 | ~n13146;
  assign n13148 = ~n9048 & ~n12871;
  assign n13149 = ~n9121 & ~n12875;
  assign n13150 = ~n9114 & n12878;
  assign n13151 = ~n8989 & n12880;
  assign n13152 = ~n8695 & ~n9048;
  assign n13153 = ~n13150 & ~n13151;
  assign n13154 = ~n13152 & n13153;
  assign n13155 = n12877 & ~n13154;
  assign n13156 = ~n11760 & ~n13155;
  assign n13157 = n9055 & ~n12931;
  assign n13158 = ~n9055 & n12931;
  assign n13159 = ~n13157 & ~n13158;
  assign n13160 = ~n12956 & ~n12997;
  assign n13161 = ~n12942 & ~n13160;
  assign n13162 = ~n13159 & n13161;
  assign n13163 = ~n12932 & ~n12943;
  assign n13164 = ~n13161 & ~n13163;
  assign n13165 = ~n13162 & ~n13164;
  assign n13166 = n13022 & ~n13165;
  assign n13167 = ~n13148 & ~n13149;
  assign n13168 = n13156 & n13167;
  assign n2410 = n13166 | ~n13168;
  assign n13170 = ~n9791 & ~n12871;
  assign n13171 = ~n9869 & ~n12875;
  assign n13172 = ~n9862 & n12878;
  assign n13173 = ~n9737 & n12880;
  assign n13174 = ~n8695 & ~n9791;
  assign n13175 = ~n13172 & ~n13173;
  assign n13176 = ~n13174 & n13175;
  assign n13177 = n12877 & ~n13176;
  assign n13178 = ~n11384 & ~n13177;
  assign n13179 = n9798 & ~n13100;
  assign n13180 = ~n9798 & n13100;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = n13125 & ~n13181;
  assign n13183 = ~n13125 & n13181;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = n13022 & ~n13184;
  assign n13186 = ~n13170 & ~n13171;
  assign n13187 = n13178 & n13186;
  assign n2415 = n13185 | ~n13187;
  assign n13189 = n8816 & ~n12961;
  assign n13190 = ~n8816 & n12961;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = n12987 & ~n13191;
  assign n13193 = ~n12962 & ~n12970;
  assign n13194 = ~n12987 & ~n13193;
  assign n13195 = ~n13192 & ~n13194;
  assign n13196 = n13022 & ~n13195;
  assign n13197 = ~n8877 & ~n12875;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = P2_REG3_REG_2_ & ~n12871;
  assign n13200 = ~n8870 & n12878;
  assign n13201 = ~n8778 & n12880;
  assign n13202 = P2_REG3_REG_2_ & ~n8695;
  assign n13203 = ~n13200 & ~n13201;
  assign n13204 = ~n13202 & n13203;
  assign n13205 = n12877 & ~n13204;
  assign n13206 = ~n11896 & ~n13205;
  assign n13207 = n13198 & ~n13199;
  assign n2420 = ~n13206 | ~n13207;
  assign n13209 = ~n9369 & ~n12871;
  assign n13210 = ~n9441 & ~n12875;
  assign n13211 = ~n9434 & n12878;
  assign n13212 = ~n9309 & n12880;
  assign n13213 = ~n8695 & ~n9369;
  assign n13214 = ~n13211 & ~n13212;
  assign n13215 = ~n13213 & n13214;
  assign n13216 = n12877 & ~n13215;
  assign n13217 = ~n11610 & ~n13216;
  assign n13218 = ~n12926 & ~n13007;
  assign n13219 = ~n12895 & ~n13218;
  assign n13220 = n9376 & ~n12907;
  assign n13221 = ~n9376 & n12907;
  assign n13222 = ~n13220 & ~n13221;
  assign n13223 = n13219 & ~n13222;
  assign n13224 = ~n12908 & ~n12914;
  assign n13225 = ~n13219 & ~n13224;
  assign n13226 = ~n13223 & ~n13225;
  assign n13227 = n13022 & ~n13226;
  assign n13228 = ~n13209 & ~n13210;
  assign n13229 = n13217 & n13228;
  assign n2425 = n13227 | ~n13229;
  assign n13231 = ~n10024 & n13029;
  assign n13232 = P2_REG3_REG_22_ & ~P2_STATE_REG;
  assign n13233 = ~n10085 & n12878;
  assign n13234 = ~n9978 & n12880;
  assign n13235 = ~n8695 & ~n10024;
  assign n13236 = ~n13233 & ~n13234;
  assign n13237 = ~n13235 & n13236;
  assign n13238 = n12877 & ~n13237;
  assign n13239 = ~n13232 & ~n13238;
  assign n13240 = n10087 & n13041;
  assign n13241 = n10031 & ~n13074;
  assign n13242 = ~n10031 & n13074;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = n13129 & ~n13243;
  assign n13245 = ~n13129 & n13243;
  assign n13246 = ~n13244 & ~n13245;
  assign n13247 = n13022 & ~n13246;
  assign n13248 = ~n13231 & n13239;
  assign n13249 = ~n13240 & n13248;
  assign n2430 = n13247 | ~n13249;
  assign n13251 = ~n9492 & ~n12871;
  assign n13252 = ~n9567 & ~n12875;
  assign n13253 = ~n9560 & n12878;
  assign n13254 = ~n9434 & n12880;
  assign n13255 = ~n8695 & ~n9492;
  assign n13256 = ~n13253 & ~n13254;
  assign n13257 = ~n13255 & n13256;
  assign n13258 = n12877 & ~n13257;
  assign n13259 = ~n11544 & ~n13258;
  assign n13260 = n12904 & ~n12911;
  assign n13261 = ~n12908 & ~n13219;
  assign n13262 = ~n12914 & ~n13261;
  assign n13263 = ~n12912 & n13262;
  assign n13264 = n13260 & ~n13263;
  assign n13265 = n9499 & ~n12902;
  assign n13266 = ~n9499 & n12902;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~n12912 & n13267;
  assign n13269 = ~n12899 & ~n13262;
  assign n13270 = n13268 & ~n13269;
  assign n13271 = ~n13264 & ~n13270;
  assign n13272 = n13022 & n13271;
  assign n13273 = ~n13251 & ~n13252;
  assign n13274 = n13259 & n13273;
  assign n2435 = n13272 | ~n13274;
  assign n13276 = ~n9915 & n13029;
  assign n13277 = P2_REG3_REG_20_ & ~P2_STATE_REG;
  assign n13278 = ~n9978 & n12878;
  assign n13279 = ~n9862 & n12880;
  assign n13280 = ~n8695 & ~n9915;
  assign n13281 = ~n13278 & ~n13279;
  assign n13282 = ~n13280 & n13281;
  assign n13283 = n12877 & ~n13282;
  assign n13284 = ~n13277 & ~n13283;
  assign n13285 = n9980 & n13041;
  assign n13286 = n9922 & ~n13084;
  assign n13287 = ~n9922 & n13084;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = ~n13096 & ~n13127;
  assign n13290 = ~n13090 & ~n13289;
  assign n13291 = ~n13288 & n13290;
  assign n13292 = ~n13085 & ~n13091;
  assign n13293 = ~n13290 & ~n13292;
  assign n13294 = ~n13291 & ~n13293;
  assign n13295 = n13022 & ~n13294;
  assign n13296 = ~n13276 & n13284;
  assign n13297 = ~n13285 & n13296;
  assign n2440 = n13295 | ~n13297;
  assign n13299 = ~n8695 & n12877;
  assign n13300 = n12871 & ~n13299;
  assign n13301 = P2_REG3_REG_0_ & ~n13300;
  assign n13302 = ~n12891 & n12975;
  assign n13303 = n12891 & ~n12975;
  assign n13304 = ~n13302 & ~n13303;
  assign n13305 = n8762 & ~n13304;
  assign n13306 = ~n8762 & n13304;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = n13022 & ~n13307;
  assign n13309 = ~n8739 & ~n12875;
  assign n13310 = ~n8778 & n12877;
  assign n13311 = n12878 & n13310;
  assign n13312 = ~n13309 & ~n13311;
  assign n13313 = ~n11956 & ~n13308;
  assign n13314 = n13312 & n13313;
  assign n2445 = n13301 | ~n13314;
  assign n13316 = ~n9238 & ~n12871;
  assign n13317 = ~n9316 & ~n12875;
  assign n13318 = ~n9309 & n12878;
  assign n13319 = ~n9181 & n12880;
  assign n13320 = ~n8695 & ~n9238;
  assign n13321 = ~n13318 & ~n13319;
  assign n13322 = ~n13320 & n13321;
  assign n13323 = n12877 & ~n13322;
  assign n13324 = ~n11670 & ~n13323;
  assign n13325 = n9245 & ~n13003;
  assign n13326 = ~n9245 & n13003;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = n12999 & ~n13327;
  assign n13329 = ~n12999 & n13327;
  assign n13330 = ~n13328 & ~n13329;
  assign n13331 = n13022 & ~n13330;
  assign n13332 = ~n13316 & ~n13317;
  assign n13333 = n13324 & n13332;
  assign n2450 = n13331 | ~n13333;
  assign n13335 = n8929 & ~n12993;
  assign n13336 = ~n8929 & n12993;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = n12989 & ~n13337;
  assign n13339 = ~n12989 & n13337;
  assign n13340 = ~n13338 & ~n13339;
  assign n13341 = n13022 & ~n13340;
  assign n13342 = ~n8996 & ~n12875;
  assign n13343 = ~n13341 & ~n13342;
  assign n13344 = ~n8922 & ~n12871;
  assign n13345 = ~n8989 & n12878;
  assign n13346 = ~n8870 & n12880;
  assign n13347 = ~n8695 & ~n8922;
  assign n13348 = ~n13345 & ~n13346;
  assign n13349 = ~n13347 & n13348;
  assign n13350 = n12877 & ~n13349;
  assign n13351 = ~n11826 & ~n13350;
  assign n13352 = n13343 & ~n13344;
  assign n2455 = ~n13351 | ~n13352;
  assign n13354 = ~n10134 & n13029;
  assign n13355 = P2_REG3_REG_24_ & ~P2_STATE_REG;
  assign n13356 = ~n10195 & n12878;
  assign n13357 = ~n10085 & n12880;
  assign n13358 = ~n8695 & ~n10134;
  assign n13359 = ~n13356 & ~n13357;
  assign n13360 = ~n13358 & n13359;
  assign n13361 = n12877 & ~n13360;
  assign n13362 = ~n13355 & ~n13361;
  assign n13363 = n10197 & n13041;
  assign n13364 = n10141 & ~n13065;
  assign n13365 = ~n10141 & n13065;
  assign n13366 = ~n13364 & ~n13365;
  assign n13367 = n13133 & ~n13366;
  assign n13368 = ~n13066 & ~n13136;
  assign n13369 = ~n13133 & ~n13368;
  assign n13370 = ~n13367 & ~n13369;
  assign n13371 = n13022 & ~n13370;
  assign n13372 = ~n13354 & n13362;
  assign n13373 = ~n13363 & n13372;
  assign n2460 = n13371 | ~n13373;
  assign n13375 = ~n9730 & ~n12871;
  assign n13376 = ~n9805 & ~n12875;
  assign n13377 = ~n9798 & n12878;
  assign n13378 = ~n9681 & n12880;
  assign n13379 = ~n8695 & ~n9730;
  assign n13380 = ~n13377 & ~n13378;
  assign n13381 = ~n13379 & n13380;
  assign n13382 = n12877 & ~n13381;
  assign n13383 = ~n11414 & ~n13382;
  assign n13384 = ~n9737 & ~n13110;
  assign n13385 = n13116 & ~n13384;
  assign n13386 = ~n13106 & n13123;
  assign n13387 = n13385 & ~n13386;
  assign n13388 = n9737 & ~n13110;
  assign n13389 = ~n9737 & n13110;
  assign n13390 = ~n13388 & ~n13389;
  assign n13391 = ~n13106 & n13390;
  assign n13392 = ~n13114 & ~n13123;
  assign n13393 = n13391 & ~n13392;
  assign n13394 = ~n13387 & ~n13393;
  assign n13395 = n13022 & n13394;
  assign n13396 = ~n13375 & ~n13376;
  assign n13397 = n13383 & n13396;
  assign n2465 = n13395 | ~n13397;
  assign n13399 = ~n8982 & ~n12871;
  assign n13400 = ~n9062 & ~n12875;
  assign n13401 = ~n9055 & n12878;
  assign n13402 = ~n8929 & n12880;
  assign n13403 = ~n8695 & ~n8982;
  assign n13404 = ~n13401 & ~n13402;
  assign n13405 = ~n13403 & n13404;
  assign n13406 = n12877 & ~n13405;
  assign n13407 = ~n11797 & ~n13406;
  assign n13408 = n8989 & ~n12941;
  assign n13409 = ~n8989 & n12941;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = n12997 & ~n13410;
  assign n13412 = ~n12997 & n13410;
  assign n13413 = ~n13411 & ~n13412;
  assign n13414 = n13022 & ~n13413;
  assign n13415 = ~n13399 & ~n13400;
  assign n13416 = n13407 & n13415;
  assign n2470 = n13414 | ~n13416;
  assign n13418 = ~n9674 & ~n12871;
  assign n13419 = ~n9744 & ~n12875;
  assign n13420 = ~n9737 & n12878;
  assign n13421 = ~n9623 & n12880;
  assign n13422 = ~n8695 & ~n9674;
  assign n13423 = ~n13420 & ~n13421;
  assign n13424 = ~n13422 & n13423;
  assign n13425 = n12877 & ~n13424;
  assign n13426 = ~n11450 & ~n13425;
  assign n13427 = n9681 & ~n13105;
  assign n13428 = ~n9681 & n13105;
  assign n13429 = ~n13427 & ~n13428;
  assign n13430 = n13123 & ~n13429;
  assign n13431 = ~n13106 & ~n13114;
  assign n13432 = ~n13123 & ~n13431;
  assign n13433 = ~n13430 & ~n13432;
  assign n13434 = n13022 & ~n13433;
  assign n13435 = ~n13418 & ~n13419;
  assign n13436 = n13426 & n13435;
  assign n2475 = n13434 | ~n13436;
  assign n13438 = ~n10188 & n13029;
  assign n13439 = P2_REG3_REG_25_ & ~P2_STATE_REG;
  assign n13440 = ~n10253 & n12878;
  assign n13441 = ~n10141 & n12880;
  assign n13442 = ~n8695 & ~n10188;
  assign n13443 = ~n13440 & ~n13441;
  assign n13444 = ~n13442 & n13443;
  assign n13445 = n12877 & ~n13444;
  assign n13446 = ~n13439 & ~n13445;
  assign n13447 = n10255 & n13041;
  assign n13448 = ~n13134 & ~n13136;
  assign n13449 = n10195 & ~n13045;
  assign n13450 = ~n10195 & n13045;
  assign n13451 = ~n13449 & ~n13450;
  assign n13452 = n13448 & ~n13451;
  assign n13453 = ~n13046 & ~n13055;
  assign n13454 = ~n13448 & ~n13453;
  assign n13455 = ~n13452 & ~n13454;
  assign n13456 = n13022 & ~n13455;
  assign n13457 = ~n13438 & n13446;
  assign n13458 = ~n13447 & n13457;
  assign n2480 = n13456 | ~n13458;
  assign n13460 = ~n9427 & ~n12871;
  assign n13461 = ~n9506 & ~n12875;
  assign n13462 = ~n9499 & n12878;
  assign n13463 = ~n9376 & n12880;
  assign n13464 = ~n8695 & ~n9427;
  assign n13465 = ~n13462 & ~n13463;
  assign n13466 = ~n13464 & n13465;
  assign n13467 = n12877 & ~n13466;
  assign n13468 = ~n11574 & ~n13467;
  assign n13469 = n9434 & ~n12898;
  assign n13470 = ~n9434 & n12898;
  assign n13471 = ~n13469 & ~n13470;
  assign n13472 = n13262 & ~n13471;
  assign n13473 = ~n12899 & ~n12912;
  assign n13474 = ~n13262 & ~n13473;
  assign n13475 = ~n13472 & ~n13474;
  assign n13476 = n13022 & ~n13475;
  assign n13477 = ~n13460 & ~n13461;
  assign n13478 = n13468 & n13477;
  assign n2485 = n13476 | ~n13478;
  assign n13480 = ~n9971 & n13029;
  assign n13481 = P2_REG3_REG_21_ & ~P2_STATE_REG;
  assign n13482 = ~n10031 & n12878;
  assign n13483 = ~n9922 & n12880;
  assign n13484 = ~n8695 & ~n9971;
  assign n13485 = ~n13482 & ~n13483;
  assign n13486 = ~n13484 & n13485;
  assign n13487 = n12877 & ~n13486;
  assign n13488 = ~n13481 & ~n13487;
  assign n13489 = n10033 & n13041;
  assign n13490 = ~n13081 & n13092;
  assign n13491 = ~n13085 & n13290;
  assign n13492 = n13490 & ~n13491;
  assign n13493 = n9978 & ~n13079;
  assign n13494 = ~n9978 & n13079;
  assign n13495 = ~n13493 & ~n13494;
  assign n13496 = ~n13085 & n13495;
  assign n13497 = ~n13091 & ~n13290;
  assign n13498 = n13496 & ~n13497;
  assign n13499 = ~n13492 & ~n13498;
  assign n13500 = n13022 & n13499;
  assign n13501 = ~n13480 & n13488;
  assign n13502 = ~n13489 & n13501;
  assign n2490 = n13500 | ~n13502;
  assign n13504 = ~n12976 & ~n12984;
  assign n13505 = n8778 & ~n12979;
  assign n13506 = ~n8778 & n12979;
  assign n13507 = ~n13505 & ~n13506;
  assign n13508 = n13504 & ~n13507;
  assign n13509 = ~n13504 & n13507;
  assign n13510 = ~n13508 & ~n13509;
  assign n13511 = n13022 & ~n13510;
  assign n13512 = ~n8823 & ~n12875;
  assign n13513 = ~n13511 & ~n13512;
  assign n13514 = P2_REG3_REG_1_ & ~n12871;
  assign n13515 = ~n8816 & n12878;
  assign n13516 = ~n8762 & n12880;
  assign n13517 = P2_REG3_REG_1_ & ~n8695;
  assign n13518 = ~n13515 & ~n13516;
  assign n13519 = ~n13517 & n13518;
  assign n13520 = n12877 & ~n13519;
  assign n13521 = ~n11932 & ~n13520;
  assign n13522 = n13513 & ~n13514;
  assign n2495 = ~n13521 | ~n13522;
  assign n13524 = ~n9174 & ~n12871;
  assign n13525 = ~n9252 & ~n12875;
  assign n13526 = ~n9245 & n12878;
  assign n13527 = ~n9114 & n12880;
  assign n13528 = ~n8695 & ~n9174;
  assign n13529 = ~n13526 & ~n13527;
  assign n13530 = ~n13528 & n13529;
  assign n13531 = n12877 & ~n13530;
  assign n13532 = ~n11679 & ~n13531;
  assign n13533 = n12957 & ~n12997;
  assign n13534 = n12948 & ~n13533;
  assign n13535 = n9181 & ~n12951;
  assign n13536 = ~n9181 & n12951;
  assign n13537 = ~n13535 & ~n13536;
  assign n13538 = n13534 & ~n13537;
  assign n13539 = ~n13534 & n13537;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = n13022 & ~n13540;
  assign n13542 = ~n13524 & ~n13525;
  assign n13543 = n13532 & n13542;
  assign n2500 = n13541 | ~n13543;
  assign n13545 = ~n10352 & n13029;
  assign n13546 = P2_REG3_REG_28_ & ~P2_STATE_REG;
  assign n13547 = ~n10409 & n12878;
  assign n13548 = ~n10305 & n12880;
  assign n13549 = ~n8695 & ~n10352;
  assign n13550 = ~n13547 & ~n13548;
  assign n13551 = ~n13549 & n13550;
  assign n13552 = n12877 & ~n13551;
  assign n13553 = ~n13546 & ~n13552;
  assign n13554 = n10411 & n13041;
  assign n13555 = n10361 & n12891;
  assign n13556 = ~n10361 & ~n12891;
  assign n13557 = ~n13555 & ~n13556;
  assign n13558 = n10305 & n13557;
  assign n13559 = ~n13055 & ~n13136;
  assign n13560 = ~n13054 & n13559;
  assign n13561 = ~n13558 & ~n13560;
  assign n13562 = ~n13054 & ~n13058;
  assign n13563 = ~n13057 & n13562;
  assign n13564 = n13561 & ~n13563;
  assign n13565 = ~n10305 & ~n13557;
  assign n13566 = ~n13564 & ~n13565;
  assign n13567 = n13057 & ~n13066;
  assign n13568 = ~n13046 & ~n13066;
  assign n13569 = ~n13049 & n13568;
  assign n13570 = ~n13567 & ~n13569;
  assign n13571 = ~n13558 & ~n13570;
  assign n13572 = ~n13133 & n13571;
  assign n13573 = ~n10359 & n12891;
  assign n13574 = n10359 & ~n12891;
  assign n13575 = ~n13573 & ~n13574;
  assign n13576 = ~n10411 & ~n13575;
  assign n13577 = n10411 & n13575;
  assign n13578 = ~n13576 & ~n13577;
  assign n13579 = n13566 & ~n13572;
  assign n13580 = ~n13578 & n13579;
  assign n13581 = ~n13560 & ~n13563;
  assign n13582 = ~n13565 & ~n13581;
  assign n13583 = ~n13133 & ~n13570;
  assign n13584 = n13582 & ~n13583;
  assign n13585 = ~n13558 & ~n13584;
  assign n13586 = n13578 & n13585;
  assign n13587 = ~n13580 & ~n13586;
  assign n13588 = n13022 & ~n13587;
  assign n13589 = ~n13545 & n13553;
  assign n13590 = ~n13554 & n13589;
  assign n2505 = n13588 | ~n13590;
  assign n13592 = ~n9855 & ~n12871;
  assign n13593 = ~n9922 & n12878;
  assign n13594 = ~n9798 & n12880;
  assign n13595 = ~n8695 & ~n9855;
  assign n13596 = ~n13593 & ~n13594;
  assign n13597 = ~n13595 & n13596;
  assign n13598 = n12877 & ~n13597;
  assign n13599 = ~n11351 & ~n13598;
  assign n13600 = ~n9926 & ~n12875;
  assign n13601 = n9862 & ~n13089;
  assign n13602 = ~n9862 & n13089;
  assign n13603 = ~n13601 & ~n13602;
  assign n13604 = n13127 & ~n13603;
  assign n13605 = ~n13090 & ~n13096;
  assign n13606 = ~n13127 & ~n13605;
  assign n13607 = ~n13604 & ~n13606;
  assign n13608 = n13022 & ~n13607;
  assign n13609 = ~n13592 & n13599;
  assign n13610 = ~n13600 & n13609;
  assign n2510 = n13608 | ~n13610;
  assign n13612 = ~n8870 & ~n12966;
  assign n13613 = n12972 & ~n13612;
  assign n13614 = ~n12962 & n12987;
  assign n13615 = n13613 & ~n13614;
  assign n13616 = n8870 & ~n12966;
  assign n13617 = ~n8870 & n12966;
  assign n13618 = ~n13616 & ~n13617;
  assign n13619 = ~n12962 & n13618;
  assign n13620 = ~n12970 & ~n12987;
  assign n13621 = n13619 & ~n13620;
  assign n13622 = ~n13615 & ~n13621;
  assign n13623 = n13022 & n13622;
  assign n13624 = ~n8936 & ~n12875;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = ~P2_REG3_REG_3_ & ~n12871;
  assign n13627 = ~n8929 & n12878;
  assign n13628 = ~n8816 & n12880;
  assign n13629 = ~P2_REG3_REG_3_ & ~n8695;
  assign n13630 = ~n13627 & ~n13628;
  assign n13631 = ~n13629 & n13630;
  assign n13632 = n12877 & ~n13631;
  assign n13633 = ~n11856 & ~n13632;
  assign n13634 = n13625 & ~n13626;
  assign n2515 = ~n13633 | ~n13634;
  assign n13636 = ~n9302 & ~n12871;
  assign n13637 = ~n9383 & ~n12875;
  assign n13638 = ~n9376 & n12878;
  assign n13639 = ~n9245 & n12880;
  assign n13640 = ~n8695 & ~n9302;
  assign n13641 = ~n13638 & ~n13639;
  assign n13642 = ~n13640 & n13641;
  assign n13643 = n12877 & ~n13642;
  assign n13644 = ~n11640 & ~n13643;
  assign n13645 = n9309 & ~n12894;
  assign n13646 = ~n9309 & n12894;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = n13007 & ~n13647;
  assign n13649 = ~n13007 & n13647;
  assign n13650 = ~n13648 & ~n13649;
  assign n13651 = n13022 & ~n13650;
  assign n13652 = ~n13636 & ~n13637;
  assign n13653 = n13644 & n13652;
  assign n2520 = n13651 | ~n13653;
  assign n13655 = ~n10078 & n13029;
  assign n13656 = P2_REG3_REG_23_ & ~P2_STATE_REG;
  assign n13657 = ~n10141 & n12878;
  assign n13658 = ~n10031 & n12880;
  assign n13659 = ~n8695 & ~n10078;
  assign n13660 = ~n13657 & ~n13658;
  assign n13661 = ~n13659 & n13660;
  assign n13662 = n12877 & ~n13661;
  assign n13663 = ~n13656 & ~n13662;
  assign n13664 = n10143 & n13041;
  assign n13665 = n10085 & ~n13069;
  assign n13666 = ~n10085 & n13069;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = n13131 & ~n13667;
  assign n13669 = ~n13131 & n13667;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = n13022 & ~n13670;
  assign n13672 = ~n13655 & n13663;
  assign n13673 = ~n13664 & n13672;
  assign n2525 = n13671 | ~n13673;
  assign n13675 = ~n9553 & ~n12871;
  assign n13676 = ~n9630 & ~n12875;
  assign n13677 = ~n9623 & n12878;
  assign n13678 = ~n9499 & n12880;
  assign n13679 = ~n8695 & ~n9553;
  assign n13680 = ~n13677 & ~n13678;
  assign n13681 = ~n13679 & n13680;
  assign n13682 = n12877 & ~n13681;
  assign n13683 = ~n11514 & ~n13682;
  assign n13684 = n12927 & ~n13007;
  assign n13685 = n12918 & ~n13684;
  assign n13686 = n9560 & ~n12921;
  assign n13687 = ~n9560 & n12921;
  assign n13688 = ~n13686 & ~n13687;
  assign n13689 = n13685 & ~n13688;
  assign n13690 = ~n13685 & n13688;
  assign n13691 = ~n13689 & ~n13690;
  assign n13692 = n13022 & ~n13691;
  assign n13693 = ~n13675 & ~n13676;
  assign n13694 = n13683 & n13693;
  assign n2530 = n13692 | ~n13694;
  assign n13696 = ~n10298 & n13029;
  assign n13697 = P2_REG3_REG_27_ & ~P2_STATE_REG;
  assign n13698 = ~n10359 & n12878;
  assign n13699 = ~n10253 & n12880;
  assign n13700 = ~n8695 & ~n10298;
  assign n13701 = ~n13698 & ~n13699;
  assign n13702 = ~n13700 & n13701;
  assign n13703 = n12877 & ~n13702;
  assign n13704 = ~n13697 & ~n13703;
  assign n13705 = n10361 & n13041;
  assign n13706 = ~n13581 & ~n13583;
  assign n13707 = n10305 & ~n13557;
  assign n13708 = ~n10305 & n13557;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = n13706 & ~n13709;
  assign n13711 = ~n13706 & n13709;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = n13022 & ~n13712;
  assign n13714 = ~n13696 & n13704;
  assign n13715 = ~n13705 & n13714;
  assign n2535 = n13713 | ~n13715;
  assign n13717 = ~n9107 & ~n12871;
  assign n13718 = ~n9188 & ~n12875;
  assign n13719 = ~n9181 & n12878;
  assign n13720 = ~n9055 & n12880;
  assign n13721 = ~n8695 & ~n9107;
  assign n13722 = ~n13719 & ~n13720;
  assign n13723 = ~n13721 & n13722;
  assign n13724 = n12877 & ~n13723;
  assign n13725 = ~n11714 & ~n13724;
  assign n13726 = ~n9114 & ~n12936;
  assign n13727 = n12945 & ~n13726;
  assign n13728 = ~n12932 & n13161;
  assign n13729 = n13727 & ~n13728;
  assign n13730 = n9114 & ~n12936;
  assign n13731 = ~n9114 & n12936;
  assign n13732 = ~n13730 & ~n13731;
  assign n13733 = ~n12932 & n13732;
  assign n13734 = ~n12943 & ~n13161;
  assign n13735 = n13733 & ~n13734;
  assign n13736 = ~n13729 & ~n13735;
  assign n13737 = n13022 & n13736;
  assign n13738 = ~n13717 & ~n13718;
  assign n13739 = n13725 & n13738;
  assign n2540 = n13737 | ~n13739;
  assign n13741 = P2_STATE_REG & ~n11002;
  assign n13742 = n8581 & n11003;
  assign n2550 = ~n13741 | n13742;
  assign n1320 = ~P1_STATE_REG;
  assign n2545 = ~P2_STATE_REG;
  always @ (posedge clock) begin
    P1_IR_REG_0_ <= n110;
    P1_IR_REG_1_ <= n115;
    P1_IR_REG_2_ <= n120;
    P1_IR_REG_3_ <= n125;
    P1_IR_REG_4_ <= n130;
    P1_IR_REG_5_ <= n135;
    P1_IR_REG_6_ <= n140;
    P1_IR_REG_7_ <= n145;
    P1_IR_REG_8_ <= n150;
    P1_IR_REG_9_ <= n155;
    P1_IR_REG_10_ <= n160;
    P1_IR_REG_11_ <= n165;
    P1_IR_REG_12_ <= n170;
    P1_IR_REG_13_ <= n175;
    P1_IR_REG_14_ <= n180;
    P1_IR_REG_15_ <= n185;
    P1_IR_REG_16_ <= n190;
    P1_IR_REG_17_ <= n195;
    P1_IR_REG_18_ <= n200;
    P1_IR_REG_19_ <= n205;
    P1_IR_REG_20_ <= n210;
    P1_IR_REG_21_ <= n215;
    P1_IR_REG_22_ <= n220;
    P1_IR_REG_23_ <= n225;
    P1_IR_REG_24_ <= n230;
    P1_IR_REG_25_ <= n235;
    P1_IR_REG_26_ <= n240;
    P1_IR_REG_27_ <= n245;
    P1_IR_REG_28_ <= n250;
    P1_IR_REG_29_ <= n255;
    P1_IR_REG_30_ <= n260;
    P1_IR_REG_31_ <= n265;
    P1_D_REG_0_ <= n270;
    P1_D_REG_1_ <= n275;
    P1_D_REG_2_ <= n280;
    P1_D_REG_3_ <= n285;
    P1_D_REG_4_ <= n290;
    P1_D_REG_5_ <= n295;
    P1_D_REG_6_ <= n300;
    P1_D_REG_7_ <= n305;
    P1_D_REG_8_ <= n310;
    P1_D_REG_9_ <= n315;
    P1_D_REG_10_ <= n320;
    P1_D_REG_11_ <= n325;
    P1_D_REG_12_ <= n330;
    P1_D_REG_13_ <= n335;
    P1_D_REG_14_ <= n340;
    P1_D_REG_15_ <= n345;
    P1_D_REG_16_ <= n350;
    P1_D_REG_17_ <= n355;
    P1_D_REG_18_ <= n360;
    P1_D_REG_19_ <= n365;
    P1_D_REG_20_ <= n370;
    P1_D_REG_21_ <= n375;
    P1_D_REG_22_ <= n380;
    P1_D_REG_23_ <= n385;
    P1_D_REG_24_ <= n390;
    P1_D_REG_25_ <= n395;
    P1_D_REG_26_ <= n400;
    P1_D_REG_27_ <= n405;
    P1_D_REG_28_ <= n410;
    P1_D_REG_29_ <= n415;
    P1_D_REG_30_ <= n420;
    P1_D_REG_31_ <= n425;
    P1_REG0_REG_0_ <= n430;
    P1_REG0_REG_1_ <= n435;
    P1_REG0_REG_2_ <= n440;
    P1_REG0_REG_3_ <= n445;
    P1_REG0_REG_4_ <= n450;
    P1_REG0_REG_5_ <= n455;
    P1_REG0_REG_6_ <= n460;
    P1_REG0_REG_7_ <= n465;
    P1_REG0_REG_8_ <= n470;
    P1_REG0_REG_9_ <= n475;
    P1_REG0_REG_10_ <= n480;
    P1_REG0_REG_11_ <= n485;
    P1_REG0_REG_12_ <= n490;
    P1_REG0_REG_13_ <= n495;
    P1_REG0_REG_14_ <= n500;
    P1_REG0_REG_15_ <= n505;
    P1_REG0_REG_16_ <= n510;
    P1_REG0_REG_17_ <= n515;
    P1_REG0_REG_18_ <= n520;
    P1_REG0_REG_19_ <= n525;
    P1_REG0_REG_20_ <= n530;
    P1_REG0_REG_21_ <= n535;
    P1_REG0_REG_22_ <= n540;
    P1_REG0_REG_23_ <= n545;
    P1_REG0_REG_24_ <= n550;
    P1_REG0_REG_25_ <= n555;
    P1_REG0_REG_26_ <= n560;
    P1_REG0_REG_27_ <= n565;
    P1_REG0_REG_28_ <= n570;
    P1_REG0_REG_29_ <= n575;
    P1_REG0_REG_30_ <= n580;
    P1_REG0_REG_31_ <= n585;
    P1_REG1_REG_0_ <= n590;
    P1_REG1_REG_1_ <= n595;
    P1_REG1_REG_2_ <= n600;
    P1_REG1_REG_3_ <= n605;
    P1_REG1_REG_4_ <= n610;
    P1_REG1_REG_5_ <= n615;
    P1_REG1_REG_6_ <= n620;
    P1_REG1_REG_7_ <= n625;
    P1_REG1_REG_8_ <= n630;
    P1_REG1_REG_9_ <= n635;
    P1_REG1_REG_10_ <= n640;
    P1_REG1_REG_11_ <= n645;
    P1_REG1_REG_12_ <= n650;
    P1_REG1_REG_13_ <= n655;
    P1_REG1_REG_14_ <= n660;
    P1_REG1_REG_15_ <= n665;
    P1_REG1_REG_16_ <= n670;
    P1_REG1_REG_17_ <= n675;
    P1_REG1_REG_18_ <= n680;
    P1_REG1_REG_19_ <= n685;
    P1_REG1_REG_20_ <= n690;
    P1_REG1_REG_21_ <= n695;
    P1_REG1_REG_22_ <= n700;
    P1_REG1_REG_23_ <= n705;
    P1_REG1_REG_24_ <= n710;
    P1_REG1_REG_25_ <= n715;
    P1_REG1_REG_26_ <= n720;
    P1_REG1_REG_27_ <= n725;
    P1_REG1_REG_28_ <= n730;
    P1_REG1_REG_29_ <= n735;
    P1_REG1_REG_30_ <= n740;
    P1_REG1_REG_31_ <= n745;
    P1_REG2_REG_0_ <= n750;
    P1_REG2_REG_1_ <= n755;
    P1_REG2_REG_2_ <= n760;
    P1_REG2_REG_3_ <= n765;
    P1_REG2_REG_4_ <= n770;
    P1_REG2_REG_5_ <= n775;
    P1_REG2_REG_6_ <= n780;
    P1_REG2_REG_7_ <= n785;
    P1_REG2_REG_8_ <= n790;
    P1_REG2_REG_9_ <= n795;
    P1_REG2_REG_10_ <= n800;
    P1_REG2_REG_11_ <= n805;
    P1_REG2_REG_12_ <= n810;
    P1_REG2_REG_13_ <= n815;
    P1_REG2_REG_14_ <= n820;
    P1_REG2_REG_15_ <= n825;
    P1_REG2_REG_16_ <= n830;
    P1_REG2_REG_17_ <= n835;
    P1_REG2_REG_18_ <= n840;
    P1_REG2_REG_19_ <= n845;
    P1_REG2_REG_20_ <= n850;
    P1_REG2_REG_21_ <= n855;
    P1_REG2_REG_22_ <= n860;
    P1_REG2_REG_23_ <= n865;
    P1_REG2_REG_24_ <= n870;
    P1_REG2_REG_25_ <= n875;
    P1_REG2_REG_26_ <= n880;
    P1_REG2_REG_27_ <= n885;
    P1_REG2_REG_28_ <= n890;
    P1_REG2_REG_29_ <= n895;
    P1_REG2_REG_30_ <= n900;
    P1_REG2_REG_31_ <= n905;
    P1_ADDR_REG_19_ <= n910;
    P1_ADDR_REG_18_ <= n915;
    P1_ADDR_REG_17_ <= n920;
    P1_ADDR_REG_16_ <= n925;
    P1_ADDR_REG_15_ <= n930;
    P1_ADDR_REG_14_ <= n935;
    P1_ADDR_REG_13_ <= n940;
    P1_ADDR_REG_12_ <= n945;
    P1_ADDR_REG_11_ <= n950;
    P1_ADDR_REG_10_ <= n955;
    P1_ADDR_REG_9_ <= n960;
    P1_ADDR_REG_8_ <= n965;
    P1_ADDR_REG_7_ <= n970;
    P1_ADDR_REG_6_ <= n975;
    P1_ADDR_REG_5_ <= n980;
    P1_ADDR_REG_4_ <= n985;
    P1_ADDR_REG_3_ <= n990;
    P1_ADDR_REG_2_ <= n995;
    P1_ADDR_REG_1_ <= n1000;
    P1_ADDR_REG_0_ <= n1005;
    P1_DATAO_REG_0_ <= n1010;
    P1_DATAO_REG_1_ <= n1015;
    P1_DATAO_REG_2_ <= n1020;
    P1_DATAO_REG_3_ <= n1025;
    P1_DATAO_REG_4_ <= n1030;
    P1_DATAO_REG_5_ <= n1035;
    P1_DATAO_REG_6_ <= n1040;
    P1_DATAO_REG_7_ <= n1045;
    P1_DATAO_REG_8_ <= n1050;
    P1_DATAO_REG_9_ <= n1055;
    P1_DATAO_REG_10_ <= n1060;
    P1_DATAO_REG_11_ <= n1065;
    P1_DATAO_REG_12_ <= n1070;
    P1_DATAO_REG_13_ <= n1075;
    P1_DATAO_REG_14_ <= n1080;
    P1_DATAO_REG_15_ <= n1085;
    P1_DATAO_REG_16_ <= n1090;
    P1_DATAO_REG_17_ <= n1095;
    P1_DATAO_REG_18_ <= n1100;
    P1_DATAO_REG_19_ <= n1105;
    P1_DATAO_REG_20_ <= n1110;
    P1_DATAO_REG_21_ <= n1115;
    P1_DATAO_REG_22_ <= n1120;
    P1_DATAO_REG_23_ <= n1125;
    P1_DATAO_REG_24_ <= n1130;
    P1_DATAO_REG_25_ <= n1135;
    P1_DATAO_REG_26_ <= n1140;
    P1_DATAO_REG_27_ <= n1145;
    P1_DATAO_REG_28_ <= n1150;
    P1_DATAO_REG_29_ <= n1155;
    P1_DATAO_REG_30_ <= n1160;
    P1_DATAO_REG_31_ <= n1165;
    P1_B_REG <= n1170;
    P1_REG3_REG_15_ <= n1175;
    P1_REG3_REG_26_ <= n1180;
    P1_REG3_REG_6_ <= n1185;
    P1_REG3_REG_18_ <= n1190;
    P1_REG3_REG_2_ <= n1195;
    P1_REG3_REG_11_ <= n1200;
    P1_REG3_REG_22_ <= n1205;
    P1_REG3_REG_13_ <= n1210;
    P1_REG3_REG_20_ <= n1215;
    P1_REG3_REG_0_ <= n1220;
    P1_REG3_REG_9_ <= n1225;
    P1_REG3_REG_4_ <= n1230;
    P1_REG3_REG_24_ <= n1235;
    P1_REG3_REG_17_ <= n1240;
    P1_REG3_REG_5_ <= n1245;
    P1_REG3_REG_16_ <= n1250;
    P1_REG3_REG_25_ <= n1255;
    P1_REG3_REG_12_ <= n1260;
    P1_REG3_REG_21_ <= n1265;
    P1_REG3_REG_1_ <= n1270;
    P1_REG3_REG_8_ <= n1275;
    P1_REG3_REG_28_ <= n1280;
    P1_REG3_REG_19_ <= n1285;
    P1_REG3_REG_3_ <= n1290;
    P1_REG3_REG_10_ <= n1295;
    P1_REG3_REG_23_ <= n1300;
    P1_REG3_REG_14_ <= n1305;
    P1_REG3_REG_27_ <= n1310;
    P1_REG3_REG_7_ <= n1315;
    P1_STATE_REG <= n1320;
    P1_RD_REG <= n1325;
    P1_WR_REG <= n1330;
    P2_IR_REG_0_ <= n1335;
    P2_IR_REG_1_ <= n1340;
    P2_IR_REG_2_ <= n1345;
    P2_IR_REG_3_ <= n1350;
    P2_IR_REG_4_ <= n1355;
    P2_IR_REG_5_ <= n1360;
    P2_IR_REG_6_ <= n1365;
    P2_IR_REG_7_ <= n1370;
    P2_IR_REG_8_ <= n1375;
    P2_IR_REG_9_ <= n1380;
    P2_IR_REG_10_ <= n1385;
    P2_IR_REG_11_ <= n1390;
    P2_IR_REG_12_ <= n1395;
    P2_IR_REG_13_ <= n1400;
    P2_IR_REG_14_ <= n1405;
    P2_IR_REG_15_ <= n1410;
    P2_IR_REG_16_ <= n1415;
    P2_IR_REG_17_ <= n1420;
    P2_IR_REG_18_ <= n1425;
    P2_IR_REG_19_ <= n1430;
    P2_IR_REG_20_ <= n1435;
    P2_IR_REG_21_ <= n1440;
    P2_IR_REG_22_ <= n1445;
    P2_IR_REG_23_ <= n1450;
    P2_IR_REG_24_ <= n1455;
    P2_IR_REG_25_ <= n1460;
    P2_IR_REG_26_ <= n1465;
    P2_IR_REG_27_ <= n1470;
    P2_IR_REG_28_ <= n1475;
    P2_IR_REG_29_ <= n1480;
    P2_IR_REG_30_ <= n1485;
    P2_IR_REG_31_ <= n1490;
    P2_D_REG_0_ <= n1495;
    P2_D_REG_1_ <= n1500;
    P2_D_REG_2_ <= n1505;
    P2_D_REG_3_ <= n1510;
    P2_D_REG_4_ <= n1515;
    P2_D_REG_5_ <= n1520;
    P2_D_REG_6_ <= n1525;
    P2_D_REG_7_ <= n1530;
    P2_D_REG_8_ <= n1535;
    P2_D_REG_9_ <= n1540;
    P2_D_REG_10_ <= n1545;
    P2_D_REG_11_ <= n1550;
    P2_D_REG_12_ <= n1555;
    P2_D_REG_13_ <= n1560;
    P2_D_REG_14_ <= n1565;
    P2_D_REG_15_ <= n1570;
    P2_D_REG_16_ <= n1575;
    P2_D_REG_17_ <= n1580;
    P2_D_REG_18_ <= n1585;
    P2_D_REG_19_ <= n1590;
    P2_D_REG_20_ <= n1595;
    P2_D_REG_21_ <= n1600;
    P2_D_REG_22_ <= n1605;
    P2_D_REG_23_ <= n1610;
    P2_D_REG_24_ <= n1615;
    P2_D_REG_25_ <= n1620;
    P2_D_REG_26_ <= n1625;
    P2_D_REG_27_ <= n1630;
    P2_D_REG_28_ <= n1635;
    P2_D_REG_29_ <= n1640;
    P2_D_REG_30_ <= n1645;
    P2_D_REG_31_ <= n1650;
    P2_REG0_REG_0_ <= n1655;
    P2_REG0_REG_1_ <= n1660;
    P2_REG0_REG_2_ <= n1665;
    P2_REG0_REG_3_ <= n1670;
    P2_REG0_REG_4_ <= n1675;
    P2_REG0_REG_5_ <= n1680;
    P2_REG0_REG_6_ <= n1685;
    P2_REG0_REG_7_ <= n1690;
    P2_REG0_REG_8_ <= n1695;
    P2_REG0_REG_9_ <= n1700;
    P2_REG0_REG_10_ <= n1705;
    P2_REG0_REG_11_ <= n1710;
    P2_REG0_REG_12_ <= n1715;
    P2_REG0_REG_13_ <= n1720;
    P2_REG0_REG_14_ <= n1725;
    P2_REG0_REG_15_ <= n1730;
    P2_REG0_REG_16_ <= n1735;
    P2_REG0_REG_17_ <= n1740;
    P2_REG0_REG_18_ <= n1745;
    P2_REG0_REG_19_ <= n1750;
    P2_REG0_REG_20_ <= n1755;
    P2_REG0_REG_21_ <= n1760;
    P2_REG0_REG_22_ <= n1765;
    P2_REG0_REG_23_ <= n1770;
    P2_REG0_REG_24_ <= n1775;
    P2_REG0_REG_25_ <= n1780;
    P2_REG0_REG_26_ <= n1785;
    P2_REG0_REG_27_ <= n1790;
    P2_REG0_REG_28_ <= n1795;
    P2_REG0_REG_29_ <= n1800;
    P2_REG0_REG_30_ <= n1805;
    P2_REG0_REG_31_ <= n1810;
    P2_REG1_REG_0_ <= n1815;
    P2_REG1_REG_1_ <= n1820;
    P2_REG1_REG_2_ <= n1825;
    P2_REG1_REG_3_ <= n1830;
    P2_REG1_REG_4_ <= n1835;
    P2_REG1_REG_5_ <= n1840;
    P2_REG1_REG_6_ <= n1845;
    P2_REG1_REG_7_ <= n1850;
    P2_REG1_REG_8_ <= n1855;
    P2_REG1_REG_9_ <= n1860;
    P2_REG1_REG_10_ <= n1865;
    P2_REG1_REG_11_ <= n1870;
    P2_REG1_REG_12_ <= n1875;
    P2_REG1_REG_13_ <= n1880;
    P2_REG1_REG_14_ <= n1885;
    P2_REG1_REG_15_ <= n1890;
    P2_REG1_REG_16_ <= n1895;
    P2_REG1_REG_17_ <= n1900;
    P2_REG1_REG_18_ <= n1905;
    P2_REG1_REG_19_ <= n1910;
    P2_REG1_REG_20_ <= n1915;
    P2_REG1_REG_21_ <= n1920;
    P2_REG1_REG_22_ <= n1925;
    P2_REG1_REG_23_ <= n1930;
    P2_REG1_REG_24_ <= n1935;
    P2_REG1_REG_25_ <= n1940;
    P2_REG1_REG_26_ <= n1945;
    P2_REG1_REG_27_ <= n1950;
    P2_REG1_REG_28_ <= n1955;
    P2_REG1_REG_29_ <= n1960;
    P2_REG1_REG_30_ <= n1965;
    P2_REG1_REG_31_ <= n1970;
    P2_REG2_REG_0_ <= n1975;
    P2_REG2_REG_1_ <= n1980;
    P2_REG2_REG_2_ <= n1985;
    P2_REG2_REG_3_ <= n1990;
    P2_REG2_REG_4_ <= n1995;
    P2_REG2_REG_5_ <= n2000;
    P2_REG2_REG_6_ <= n2005;
    P2_REG2_REG_7_ <= n2010;
    P2_REG2_REG_8_ <= n2015;
    P2_REG2_REG_9_ <= n2020;
    P2_REG2_REG_10_ <= n2025;
    P2_REG2_REG_11_ <= n2030;
    P2_REG2_REG_12_ <= n2035;
    P2_REG2_REG_13_ <= n2040;
    P2_REG2_REG_14_ <= n2045;
    P2_REG2_REG_15_ <= n2050;
    P2_REG2_REG_16_ <= n2055;
    P2_REG2_REG_17_ <= n2060;
    P2_REG2_REG_18_ <= n2065;
    P2_REG2_REG_19_ <= n2070;
    P2_REG2_REG_20_ <= n2075;
    P2_REG2_REG_21_ <= n2080;
    P2_REG2_REG_22_ <= n2085;
    P2_REG2_REG_23_ <= n2090;
    P2_REG2_REG_24_ <= n2095;
    P2_REG2_REG_25_ <= n2100;
    P2_REG2_REG_26_ <= n2105;
    P2_REG2_REG_27_ <= n2110;
    P2_REG2_REG_28_ <= n2115;
    P2_REG2_REG_29_ <= n2120;
    P2_REG2_REG_30_ <= n2125;
    P2_REG2_REG_31_ <= n2130;
    P2_ADDR_REG_19_ <= n2135;
    P2_ADDR_REG_18_ <= n2140;
    P2_ADDR_REG_17_ <= n2145;
    P2_ADDR_REG_16_ <= n2150;
    P2_ADDR_REG_15_ <= n2155;
    P2_ADDR_REG_14_ <= n2160;
    P2_ADDR_REG_13_ <= n2165;
    P2_ADDR_REG_12_ <= n2170;
    P2_ADDR_REG_11_ <= n2175;
    P2_ADDR_REG_10_ <= n2180;
    P2_ADDR_REG_9_ <= n2185;
    P2_ADDR_REG_8_ <= n2190;
    P2_ADDR_REG_7_ <= n2195;
    P2_ADDR_REG_6_ <= n2200;
    P2_ADDR_REG_5_ <= n2205;
    P2_ADDR_REG_4_ <= n2210;
    P2_ADDR_REG_3_ <= n2215;
    P2_ADDR_REG_2_ <= n2220;
    P2_ADDR_REG_1_ <= n2225;
    P2_ADDR_REG_0_ <= n2230;
    P2_DATAO_REG_0_ <= n2235;
    P2_DATAO_REG_1_ <= n2240;
    P2_DATAO_REG_2_ <= n2245;
    P2_DATAO_REG_3_ <= n2250;
    P2_DATAO_REG_4_ <= n2255;
    P2_DATAO_REG_5_ <= n2260;
    P2_DATAO_REG_6_ <= n2265;
    P2_DATAO_REG_7_ <= n2270;
    P2_DATAO_REG_8_ <= n2275;
    P2_DATAO_REG_9_ <= n2280;
    P2_DATAO_REG_10_ <= n2285;
    P2_DATAO_REG_11_ <= n2290;
    P2_DATAO_REG_12_ <= n2295;
    P2_DATAO_REG_13_ <= n2300;
    P2_DATAO_REG_14_ <= n2305;
    P2_DATAO_REG_15_ <= n2310;
    P2_DATAO_REG_16_ <= n2315;
    P2_DATAO_REG_17_ <= n2320;
    P2_DATAO_REG_18_ <= n2325;
    P2_DATAO_REG_19_ <= n2330;
    P2_DATAO_REG_20_ <= n2335;
    P2_DATAO_REG_21_ <= n2340;
    P2_DATAO_REG_22_ <= n2345;
    P2_DATAO_REG_23_ <= n2350;
    P2_DATAO_REG_24_ <= n2355;
    P2_DATAO_REG_25_ <= n2360;
    P2_DATAO_REG_26_ <= n2365;
    P2_DATAO_REG_27_ <= n2370;
    P2_DATAO_REG_28_ <= n2375;
    P2_DATAO_REG_29_ <= n2380;
    P2_DATAO_REG_30_ <= n2385;
    P2_DATAO_REG_31_ <= n2390;
    P2_B_REG <= n2395;
    P2_REG3_REG_15_ <= n2400;
    P2_REG3_REG_26_ <= n2405;
    P2_REG3_REG_6_ <= n2410;
    P2_REG3_REG_18_ <= n2415;
    P2_REG3_REG_2_ <= n2420;
    P2_REG3_REG_11_ <= n2425;
    P2_REG3_REG_22_ <= n2430;
    P2_REG3_REG_13_ <= n2435;
    P2_REG3_REG_20_ <= n2440;
    P2_REG3_REG_0_ <= n2445;
    P2_REG3_REG_9_ <= n2450;
    P2_REG3_REG_4_ <= n2455;
    P2_REG3_REG_24_ <= n2460;
    P2_REG3_REG_17_ <= n2465;
    P2_REG3_REG_5_ <= n2470;
    P2_REG3_REG_16_ <= n2475;
    P2_REG3_REG_25_ <= n2480;
    P2_REG3_REG_12_ <= n2485;
    P2_REG3_REG_21_ <= n2490;
    P2_REG3_REG_1_ <= n2495;
    P2_REG3_REG_8_ <= n2500;
    P2_REG3_REG_28_ <= n2505;
    P2_REG3_REG_19_ <= n2510;
    P2_REG3_REG_3_ <= n2515;
    P2_REG3_REG_10_ <= n2520;
    P2_REG3_REG_23_ <= n2525;
    P2_REG3_REG_14_ <= n2530;
    P2_REG3_REG_27_ <= n2535;
    P2_REG3_REG_7_ <= n2540;
    P2_STATE_REG <= n2545;
    P2_RD_REG <= n2550;
    P2_WR_REG <= n2555;
  end
endmodule


