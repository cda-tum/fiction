// Benchmark "top" written by ABC on Mon Nov 27 16:54:28 2023

module top ( 
    \1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \11 , \14 , \15 , \16 , \19 ,
    \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \32 , \33 ,
    \34 , \35 , \36 , \37 , \40 , \43 , \44 , \47 , \48 , \49 , \50 , \51 ,
    \52 , \53 , \54 , \55 , \56 , \57 , \60 , \61 , \62 , \63 , \64 , \65 ,
    \66 , \67 , \68 , \69 , \72 , \73 , \74 , \75 , \76 , \77 , \78 , \79 ,
    \80 , \81 , \82 , \85 , \86 , \87 , \88 , \89 , \90 , \91 , \92 , \93 ,
    \94 , \95 , \96 , \99 , \100 , \101 , \102 , \103 , \104 , \105 ,
    \106 , \107 , \108 , \111 , \112 , \113 , \114 , \115 , \116 , \117 ,
    \118 , \119 , \120 , \123 , \124 , \125 , \126 , \127 , \128 , \129 ,
    \130 , \131 , \132 , \135 , \136 , \137 , \138 , \139 , \140 , \141 ,
    \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 ,
    \152 , \153 , \154 , \155 , \156 , \157 , \158 , \159 , \160 , \161 ,
    \162 , \163 , \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 ,
    \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 ,
    \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 ,
    \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 ,
    \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 ,
    \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \224 , \227 ,
    \230 , \231 , \234 , \237 , \241 , \246 , \253 , \256 , \259 , \262 ,
    \263 , \266 , \269 , \272 , \275 , \278 , \281 , \284 , \287 , \290 ,
    \294 , \297 , \301 , \305 , \309 , \313 , \316 , \319 , \322 , \325 ,
    \328 , \331 , \334 , \337 , \340 , \343 , \346 , \349 , \352 , \355 ,
    \398 , \400 , \401 , \419 , \420 , \456 , \457 , \458 , \487 , \488 ,
    \489 , \490 , \491 , \492 , \493 , \494 , \792 , \799 , \805 , \1026 ,
    \1028 , \1029 , \1269 , \1277 , \1448 , \1726 , \1816 , \1817 , \1818 ,
    \1819 , \1820 , \1821 , \1969 , \1970 , \1971 , \2010 , \2012 , \2014 ,
    \2016 , \2018 , \2020 , \2022 , \2387 , \2388 , \2389 , \2390 , \2496 ,
    \2643 , \2644 , \2891 , \2925 , \2970 , \2971 , \3038 , \3079 , \3546 ,
    \3671 , \3803 , \3804 , \3809 , \3851 , \3875 , \3881 , \3882   );
  input  \1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \11 , \14 , \15 , \16 ,
    \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \32 ,
    \33 , \34 , \35 , \36 , \37 , \40 , \43 , \44 , \47 , \48 , \49 , \50 ,
    \51 , \52 , \53 , \54 , \55 , \56 , \57 , \60 , \61 , \62 , \63 , \64 ,
    \65 , \66 , \67 , \68 , \69 , \72 , \73 , \74 , \75 , \76 , \77 , \78 ,
    \79 , \80 , \81 , \82 , \85 , \86 , \87 , \88 , \89 , \90 , \91 , \92 ,
    \93 , \94 , \95 , \96 , \99 , \100 , \101 , \102 , \103 , \104 , \105 ,
    \106 , \107 , \108 , \111 , \112 , \113 , \114 , \115 , \116 , \117 ,
    \118 , \119 , \120 , \123 , \124 , \125 , \126 , \127 , \128 , \129 ,
    \130 , \131 , \132 , \135 , \136 , \137 , \138 , \139 , \140 , \141 ,
    \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 ,
    \152 , \153 , \154 , \155 , \156 , \157 , \158 , \159 , \160 , \161 ,
    \162 , \163 , \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 ,
    \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 ,
    \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 ,
    \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 ,
    \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 ,
    \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \224 , \227 ,
    \230 , \231 , \234 , \237 , \241 , \246 , \253 , \256 , \259 , \262 ,
    \263 , \266 , \269 , \272 , \275 , \278 , \281 , \284 , \287 , \290 ,
    \294 , \297 , \301 , \305 , \309 , \313 , \316 , \319 , \322 , \325 ,
    \328 , \331 , \334 , \337 , \340 , \343 , \346 , \349 , \352 , \355 ;
  output \398 , \400 , \401 , \419 , \420 , \456 , \457 , \458 , \487 , \488 ,
    \489 , \490 , \491 , \492 , \493 , \494 , \792 , \799 , \805 , \1026 ,
    \1028 , \1029 , \1269 , \1277 , \1448 , \1726 , \1816 , \1817 , \1818 ,
    \1819 , \1820 , \1821 , \1969 , \1970 , \1971 , \2010 , \2012 , \2014 ,
    \2016 , \2018 , \2020 , \2022 , \2387 , \2388 , \2389 , \2390 , \2496 ,
    \2643 , \2644 , \2891 , \2925 , \2970 , \2971 , \3038 , \3079 , \3546 ,
    \3671 , \3803 , \3804 , \3809 , \3851 , \3875 , \3881 , \3882 ;
  wire new_n299, new_n300, new_n302, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n315, new_n316, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n376,
    new_n377, new_n379, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n388, new_n389, new_n390, new_n391, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n417, new_n418,
    new_n420, new_n422, new_n423, new_n424, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814;
  assign new_n299 = \301  & \309 ;
  assign new_n300 = \297  & \305 ;
  assign \792  = ~new_n299 | ~new_n300;
  assign new_n302 = \2  & \15 ;
  assign \799  = ~\237  | ~new_n302;
  assign \1026  = \94  & \219 ;
  assign \1028  = ~\7  | ~\237 ;
  assign \1029  = ~\231  | \1028 ;
  assign \1269  = ~\325  | \1028 ;
  assign new_n308 = \44  & \82 ;
  assign new_n309 = \96  & \132 ;
  assign new_n310 = new_n308 & new_n309;
  assign new_n311 = \57  & \69 ;
  assign new_n312 = \108  & \120 ;
  assign new_n313 = new_n311 & new_n312;
  assign \1277  = new_n310 & new_n313;
  assign new_n315 = \231  & ~new_n313;
  assign new_n316 = \325  & ~new_n310;
  assign \1726  = ~new_n315 & ~new_n316;
  assign new_n318 = \319  & \322 ;
  assign new_n319 = \113  & new_n318;
  assign new_n320 = \319  & ~\322 ;
  assign new_n321 = \101  & new_n320;
  assign new_n322 = ~\319  & ~\322 ;
  assign new_n323 = \137  & new_n322;
  assign new_n324 = ~\319  & \322 ;
  assign new_n325 = \125  & new_n324;
  assign new_n326 = ~new_n319 & ~new_n321;
  assign new_n327 = ~new_n323 & ~new_n325;
  assign \1816  = new_n326 & new_n327;
  assign new_n329 = \124  & new_n324;
  assign new_n330 = \112  & new_n318;
  assign new_n331 = \100  & new_n320;
  assign new_n332 = \136  & new_n322;
  assign new_n333 = ~new_n329 & ~new_n330;
  assign new_n334 = ~new_n331 & ~new_n332;
  assign \1817  = new_n333 & new_n334;
  assign new_n336 = \114  & new_n318;
  assign new_n337 = \102  & new_n320;
  assign new_n338 = \138  & new_n322;
  assign new_n339 = \126  & new_n324;
  assign new_n340 = ~new_n336 & ~new_n337;
  assign new_n341 = ~new_n338 & ~new_n339;
  assign \1818  = new_n340 & new_n341;
  assign new_n343 = \227  & \234 ;
  assign new_n344 = \75  & new_n343;
  assign new_n345 = ~\227  & \234 ;
  assign new_n346 = \62  & new_n345;
  assign new_n347 = \227  & ~\234 ;
  assign new_n348 = \50  & new_n347;
  assign new_n349 = ~\227  & ~\234 ;
  assign new_n350 = \88  & new_n349;
  assign new_n351 = ~new_n344 & ~new_n346;
  assign new_n352 = ~new_n348 & ~new_n350;
  assign \1819  = new_n351 & new_n352;
  assign new_n354 = \76  & new_n343;
  assign new_n355 = \63  & new_n345;
  assign new_n356 = \51  & new_n347;
  assign new_n357 = \89  & new_n349;
  assign new_n358 = ~new_n354 & ~new_n355;
  assign new_n359 = ~new_n356 & ~new_n357;
  assign \1820  = new_n358 & new_n359;
  assign new_n361 = \90  & new_n349;
  assign new_n362 = \77  & new_n343;
  assign new_n363 = \64  & new_n345;
  assign new_n364 = \52  & new_n347;
  assign new_n365 = ~new_n361 & ~new_n362;
  assign new_n366 = ~new_n363 & ~new_n364;
  assign \1821  = new_n365 & new_n366;
  assign new_n368 = \81  & new_n349;
  assign new_n369 = \68  & new_n343;
  assign new_n370 = \43  & new_n347;
  assign new_n371 = \56  & new_n345;
  assign new_n372 = ~new_n368 & ~new_n369;
  assign new_n373 = ~new_n370 & ~new_n371;
  assign new_n374 = new_n372 & new_n373;
  assign \1969  = ~\241  | ~new_n374;
  assign new_n376 = \224  & \237 ;
  assign new_n377 = \1726  & new_n376;
  assign \1970  = ~\36  | ~new_n377;
  assign new_n379 = \1  & \3 ;
  assign \1971  = ~new_n377 | new_n379;
  assign new_n381 = \78  & new_n343;
  assign new_n382 = \65  & new_n345;
  assign new_n383 = \53  & new_n347;
  assign new_n384 = \91  & new_n349;
  assign new_n385 = ~new_n381 & ~new_n382;
  assign new_n386 = ~new_n383 & ~new_n384;
  assign \2010  = ~new_n385 | ~new_n386;
  assign new_n388 = ~\49  & new_n347;
  assign new_n389 = ~\87  & new_n349;
  assign new_n390 = ~\74  & new_n343;
  assign new_n391 = ~new_n388 & ~new_n389;
  assign \2018  = ~new_n390 & new_n391;
  assign new_n393 = \86  & new_n349;
  assign new_n394 = \73  & new_n343;
  assign new_n395 = \48  & new_n347;
  assign new_n396 = \61  & new_n345;
  assign new_n397 = ~new_n393 & ~new_n394;
  assign new_n398 = ~new_n395 & ~new_n396;
  assign \2020  = ~new_n397 | ~new_n398;
  assign new_n400 = \72  & new_n343;
  assign new_n401 = \60  & new_n345;
  assign new_n402 = \47  & new_n347;
  assign new_n403 = \85  & new_n349;
  assign new_n404 = ~new_n400 & ~new_n401;
  assign new_n405 = ~new_n402 & ~new_n403;
  assign \2022  = ~new_n404 | ~new_n405;
  assign new_n407 = \79  & new_n343;
  assign new_n408 = \66  & new_n345;
  assign new_n409 = \54  & new_n347;
  assign new_n410 = \92  & new_n349;
  assign new_n411 = ~new_n407 & ~new_n408;
  assign new_n412 = ~new_n409 & ~new_n410;
  assign new_n413 = new_n411 & new_n412;
  assign new_n414 = ~\246  & ~new_n413;
  assign new_n415 = \246  & ~\1821 ;
  assign \2387  = new_n414 | new_n415;
  assign new_n417 = ~\246  & \2010 ;
  assign new_n418 = \246  & ~\1820 ;
  assign \2389  = new_n417 | new_n418;
  assign new_n420 = \230  & ~\241 ;
  assign \2496  = ~new_n413 | new_n420;
  assign new_n422 = ~\246  & ~new_n374;
  assign new_n423 = ~\230  & new_n413;
  assign new_n424 = \246  & ~new_n423;
  assign \2643  = new_n422 | new_n424;
  assign new_n426 = \123  & new_n324;
  assign new_n427 = \111  & new_n318;
  assign new_n428 = \99  & new_n320;
  assign new_n429 = \135  & new_n322;
  assign new_n430 = ~new_n426 & ~new_n427;
  assign new_n431 = ~new_n428 & ~new_n429;
  assign new_n432 = new_n430 & new_n431;
  assign new_n433 = \313  & ~new_n432;
  assign new_n434 = ~\313  & new_n432;
  assign new_n435 = ~\316  & ~new_n433;
  assign \2891  = new_n434 | ~new_n435;
  assign new_n437 = \259  & ~\337 ;
  assign new_n438 = ~\259  & \337 ;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = ~\340  & ~\343 ;
  assign new_n441 = \340  & \343 ;
  assign new_n442 = ~new_n440 & ~new_n441;
  assign new_n443 = \256  & ~\331 ;
  assign new_n444 = ~\256  & \331 ;
  assign new_n445 = ~new_n443 & ~new_n444;
  assign new_n446 = new_n442 & new_n445;
  assign new_n447 = ~new_n442 & ~new_n445;
  assign new_n448 = ~new_n446 & ~new_n447;
  assign new_n449 = ~\334  & ~\346 ;
  assign new_n450 = \334  & \346 ;
  assign new_n451 = ~new_n449 & ~new_n450;
  assign new_n452 = ~\328  & ~\349 ;
  assign new_n453 = \328  & \349 ;
  assign new_n454 = ~new_n452 & ~new_n453;
  assign new_n455 = new_n451 & ~new_n454;
  assign new_n456 = ~new_n451 & new_n454;
  assign new_n457 = ~new_n455 & ~new_n456;
  assign new_n458 = ~new_n448 & ~new_n457;
  assign new_n459 = new_n448 & new_n457;
  assign new_n460 = ~new_n458 & ~new_n459;
  assign new_n461 = new_n439 & new_n460;
  assign new_n462 = ~new_n439 & ~new_n460;
  assign new_n463 = \14  & ~new_n461;
  assign \2925  = ~new_n462 & new_n463;
  assign new_n465 = ~\301  & ~\309 ;
  assign new_n466 = ~new_n299 & ~new_n465;
  assign new_n467 = ~\316  & ~\355 ;
  assign new_n468 = \316  & \355 ;
  assign new_n469 = ~new_n467 & ~new_n468;
  assign new_n470 = new_n466 & ~new_n469;
  assign new_n471 = ~new_n466 & new_n469;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = ~\294  & ~\297 ;
  assign new_n474 = \294  & \297 ;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = \305  & ~\313 ;
  assign new_n477 = ~\305  & \313 ;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = new_n475 & ~new_n478;
  assign new_n480 = ~new_n475 & new_n478;
  assign new_n481 = ~new_n479 & ~new_n480;
  assign new_n482 = new_n472 & new_n481;
  assign new_n483 = ~new_n472 & ~new_n481;
  assign \2970  = ~new_n482 & ~new_n483;
  assign new_n485 = \275  & ~\278 ;
  assign new_n486 = ~\275  & \278 ;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = ~\281  & ~\284 ;
  assign new_n489 = \281  & \284 ;
  assign new_n490 = ~new_n488 & ~new_n489;
  assign new_n491 = \263  & ~\266 ;
  assign new_n492 = ~\263  & \266 ;
  assign new_n493 = ~new_n491 & ~new_n492;
  assign new_n494 = ~\269  & ~\272 ;
  assign new_n495 = \269  & \272 ;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = ~\287  & ~\352 ;
  assign new_n498 = \287  & \352 ;
  assign new_n499 = ~new_n497 & ~new_n498;
  assign new_n500 = new_n496 & ~new_n499;
  assign new_n501 = ~new_n496 & new_n499;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = new_n493 & new_n502;
  assign new_n504 = ~new_n493 & ~new_n502;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = new_n490 & ~new_n505;
  assign new_n507 = ~new_n490 & new_n505;
  assign new_n508 = ~new_n506 & ~new_n507;
  assign new_n509 = new_n487 & new_n508;
  assign new_n510 = ~new_n487 & ~new_n508;
  assign \2971  = new_n509 | new_n510;
  assign new_n512 = ~\29  & \34 ;
  assign new_n513 = \29  & ~\1816 ;
  assign new_n514 = ~new_n512 & ~new_n513;
  assign new_n515 = \305  & ~new_n514;
  assign new_n516 = ~\29  & \35 ;
  assign new_n517 = \29  & ~\1817 ;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = \309  & ~new_n518;
  assign new_n520 = ~\16  & \21 ;
  assign new_n521 = \16  & ~\1820 ;
  assign new_n522 = ~new_n520 & ~new_n521;
  assign new_n523 = ~\269  & new_n522;
  assign new_n524 = ~\309  & new_n518;
  assign new_n525 = ~\16  & \20 ;
  assign new_n526 = \16  & \2010 ;
  assign new_n527 = ~new_n525 & ~new_n526;
  assign new_n528 = \263  & ~new_n527;
  assign new_n529 = \23  & \275 ;
  assign new_n530 = ~\6  & ~\278 ;
  assign new_n531 = ~\24  & ~\281 ;
  assign new_n532 = \24  & \281 ;
  assign new_n533 = \6  & \278 ;
  assign new_n534 = ~\23  & ~\275 ;
  assign new_n535 = ~new_n529 & ~new_n530;
  assign new_n536 = ~new_n531 & ~new_n532;
  assign new_n537 = ~new_n533 & ~new_n534;
  assign new_n538 = new_n536 & new_n537;
  assign new_n539 = new_n535 & new_n538;
  assign new_n540 = ~\16  & ~new_n539;
  assign new_n541 = ~\16  & \19 ;
  assign new_n542 = \16  & ~new_n374;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign new_n544 = \256  & ~new_n543;
  assign new_n545 = \25  & \284 ;
  assign new_n546 = ~\32  & ~\287 ;
  assign new_n547 = ~\33  & ~\297 ;
  assign new_n548 = \33  & \297 ;
  assign new_n549 = ~\25  & ~\284 ;
  assign new_n550 = \32  & \287 ;
  assign new_n551 = \28  & ~new_n545;
  assign new_n552 = ~new_n546 & ~new_n547;
  assign new_n553 = ~new_n548 & ~new_n549;
  assign new_n554 = ~new_n550 & new_n553;
  assign new_n555 = new_n551 & new_n552;
  assign new_n556 = new_n554 & new_n555;
  assign new_n557 = ~\29  & ~new_n556;
  assign new_n558 = ~\305  & new_n514;
  assign new_n559 = ~\139  & new_n322;
  assign new_n560 = ~\127  & new_n324;
  assign new_n561 = ~\103  & new_n320;
  assign new_n562 = ~\115  & new_n318;
  assign new_n563 = ~new_n559 & ~new_n560;
  assign new_n564 = ~new_n561 & ~new_n562;
  assign new_n565 = new_n563 & new_n564;
  assign new_n566 = \297  & new_n565;
  assign new_n567 = \119  & new_n324;
  assign new_n568 = \107  & new_n318;
  assign new_n569 = \95  & new_n320;
  assign new_n570 = \131  & new_n322;
  assign new_n571 = ~new_n567 & ~new_n568;
  assign new_n572 = ~new_n569 & ~new_n570;
  assign new_n573 = new_n571 & new_n572;
  assign new_n574 = \284  & ~new_n573;
  assign new_n575 = ~\141  & new_n322;
  assign new_n576 = ~\129  & new_n324;
  assign new_n577 = ~\105  & new_n320;
  assign new_n578 = ~\117  & new_n318;
  assign new_n579 = ~new_n575 & ~new_n576;
  assign new_n580 = ~new_n577 & ~new_n578;
  assign new_n581 = new_n579 & new_n580;
  assign new_n582 = ~\287  & ~new_n581;
  assign new_n583 = ~\284  & new_n573;
  assign new_n584 = ~new_n582 & ~new_n583;
  assign new_n585 = \287  & new_n581;
  assign new_n586 = ~\297  & ~new_n565;
  assign new_n587 = ~new_n432 & ~new_n566;
  assign new_n588 = ~new_n574 & ~new_n585;
  assign new_n589 = ~new_n586 & new_n588;
  assign new_n590 = new_n584 & new_n587;
  assign new_n591 = new_n589 & new_n590;
  assign new_n592 = \29  & ~new_n591;
  assign new_n593 = ~\275  & ~\2018 ;
  assign new_n594 = \278  & \2020 ;
  assign new_n595 = \275  & \2018 ;
  assign new_n596 = ~new_n593 & ~new_n594;
  assign new_n597 = ~new_n595 & new_n596;
  assign new_n598 = ~\281  & ~\2022 ;
  assign new_n599 = ~\278  & ~\2020 ;
  assign new_n600 = \281  & \2022 ;
  assign new_n601 = ~new_n598 & ~new_n599;
  assign new_n602 = ~new_n600 & new_n601;
  assign new_n603 = new_n597 & new_n602;
  assign new_n604 = \16  & ~new_n603;
  assign new_n605 = \4  & ~\16 ;
  assign new_n606 = \16  & ~new_n413;
  assign new_n607 = ~new_n605 & ~new_n606;
  assign new_n608 = \259  & ~new_n607;
  assign new_n609 = \5  & ~\16 ;
  assign new_n610 = \16  & ~\1821 ;
  assign new_n611 = ~new_n609 & ~new_n610;
  assign new_n612 = \266  & ~new_n611;
  assign new_n613 = ~\259  & new_n607;
  assign new_n614 = ~\266  & new_n611;
  assign new_n615 = ~\27  & ~\29 ;
  assign new_n616 = \29  & \1818 ;
  assign new_n617 = ~new_n615 & ~new_n616;
  assign new_n618 = ~\301  & ~new_n617;
  assign new_n619 = ~\26  & ~\29 ;
  assign new_n620 = ~\140  & new_n322;
  assign new_n621 = ~\128  & new_n324;
  assign new_n622 = ~\104  & new_n320;
  assign new_n623 = ~\116  & new_n318;
  assign new_n624 = ~new_n620 & ~new_n621;
  assign new_n625 = ~new_n622 & ~new_n623;
  assign new_n626 = new_n624 & new_n625;
  assign new_n627 = \29  & ~new_n626;
  assign new_n628 = ~new_n619 & ~new_n627;
  assign new_n629 = \294  & new_n628;
  assign new_n630 = ~\294  & ~new_n628;
  assign new_n631 = ~\256  & new_n543;
  assign new_n632 = ~\263  & new_n527;
  assign new_n633 = ~\16  & ~\22 ;
  assign new_n634 = \16  & \1819 ;
  assign new_n635 = ~new_n633 & ~new_n634;
  assign new_n636 = \272  & new_n635;
  assign new_n637 = ~\272  & ~new_n635;
  assign new_n638 = \301  & new_n617;
  assign new_n639 = \269  & ~new_n522;
  assign new_n640 = \11  & ~new_n540;
  assign new_n641 = ~new_n557 & new_n640;
  assign new_n642 = ~new_n515 & new_n641;
  assign new_n643 = ~new_n519 & ~new_n523;
  assign new_n644 = ~new_n524 & ~new_n528;
  assign new_n645 = ~new_n544 & ~new_n558;
  assign new_n646 = ~new_n608 & ~new_n612;
  assign new_n647 = ~new_n613 & ~new_n614;
  assign new_n648 = ~new_n618 & ~new_n629;
  assign new_n649 = ~new_n630 & ~new_n631;
  assign new_n650 = ~new_n632 & ~new_n636;
  assign new_n651 = ~new_n637 & ~new_n638;
  assign new_n652 = ~new_n639 & new_n651;
  assign new_n653 = new_n649 & new_n650;
  assign new_n654 = new_n647 & new_n648;
  assign new_n655 = new_n645 & new_n646;
  assign new_n656 = new_n643 & new_n644;
  assign new_n657 = new_n642 & new_n656;
  assign new_n658 = new_n654 & new_n655;
  assign new_n659 = new_n652 & new_n653;
  assign new_n660 = ~new_n592 & ~new_n604;
  assign new_n661 = new_n659 & new_n660;
  assign new_n662 = new_n657 & new_n658;
  assign \3038  = new_n661 & new_n662;
  assign new_n664 = \93  & new_n349;
  assign new_n665 = \80  & new_n343;
  assign new_n666 = \67  & new_n345;
  assign new_n667 = \55  & new_n347;
  assign new_n668 = ~new_n664 & ~new_n665;
  assign new_n669 = ~new_n666 & ~new_n667;
  assign new_n670 = new_n668 & new_n669;
  assign new_n671 = \230  & new_n413;
  assign new_n672 = new_n374 & new_n671;
  assign new_n673 = ~new_n374 & ~new_n671;
  assign new_n674 = ~\241  & ~new_n672;
  assign new_n675 = ~new_n673 & new_n674;
  assign new_n676 = new_n670 & ~new_n675;
  assign new_n677 = ~new_n670 & new_n675;
  assign \3546  = ~new_n676 & ~new_n677;
  assign new_n679 = \130  & new_n324;
  assign new_n680 = \118  & new_n318;
  assign new_n681 = \106  & new_n320;
  assign new_n682 = \142  & new_n322;
  assign new_n683 = ~new_n679 & ~new_n680;
  assign new_n684 = ~new_n681 & ~new_n682;
  assign new_n685 = new_n683 & new_n684;
  assign new_n686 = \1818  & ~new_n685;
  assign new_n687 = ~\1818  & new_n685;
  assign new_n688 = ~new_n686 & ~new_n687;
  assign new_n689 = ~\1816  & ~new_n581;
  assign new_n690 = \1816  & new_n581;
  assign new_n691 = ~new_n689 & ~new_n690;
  assign new_n692 = new_n573 & ~new_n691;
  assign new_n693 = ~new_n573 & new_n691;
  assign new_n694 = ~new_n692 & ~new_n693;
  assign new_n695 = new_n688 & new_n694;
  assign new_n696 = ~new_n688 & ~new_n694;
  assign new_n697 = ~new_n695 & ~new_n696;
  assign new_n698 = \1817  & ~new_n565;
  assign new_n699 = ~\1817  & new_n565;
  assign new_n700 = ~new_n698 & ~new_n699;
  assign new_n701 = new_n432 & ~new_n626;
  assign new_n702 = ~new_n432 & new_n626;
  assign new_n703 = ~new_n701 & ~new_n702;
  assign new_n704 = new_n700 & new_n703;
  assign new_n705 = ~new_n700 & ~new_n703;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = new_n697 & new_n706;
  assign new_n708 = ~new_n697 & ~new_n706;
  assign new_n709 = ~\37  & ~new_n707;
  assign \3671  = ~new_n708 & new_n709;
  assign new_n711 = \1819  & ~new_n670;
  assign new_n712 = ~\1819  & new_n670;
  assign new_n713 = ~new_n711 & ~new_n712;
  assign new_n714 = ~\2020  & ~new_n713;
  assign new_n715 = \2020  & new_n713;
  assign new_n716 = ~new_n714 & ~new_n715;
  assign new_n717 = ~new_n374 & ~\2018 ;
  assign new_n718 = new_n374 & \2018 ;
  assign new_n719 = ~new_n717 & ~new_n718;
  assign new_n720 = \2010  & ~new_n413;
  assign new_n721 = ~\2010  & new_n413;
  assign new_n722 = ~new_n720 & ~new_n721;
  assign new_n723 = ~\2022  & ~new_n722;
  assign new_n724 = \2022  & new_n722;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = new_n719 & ~new_n725;
  assign new_n727 = ~new_n719 & new_n725;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = new_n716 & new_n728;
  assign new_n730 = ~new_n716 & ~new_n728;
  assign new_n731 = ~new_n729 & ~new_n730;
  assign new_n732 = ~new_n423 & new_n731;
  assign new_n733 = new_n423 & ~new_n731;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = \246  & ~new_n734;
  assign new_n736 = ~\246  & ~new_n670;
  assign \3803  = new_n735 | new_n736;
  assign new_n738 = \1820  & new_n731;
  assign new_n739 = ~\1820  & ~new_n731;
  assign new_n740 = ~new_n738 & ~new_n739;
  assign new_n741 = ~\1821  & ~new_n740;
  assign new_n742 = \1821  & new_n740;
  assign new_n743 = ~\37  & ~new_n741;
  assign \3809  = ~new_n742 & new_n743;
  assign new_n745 = ~\262  & ~\1818 ;
  assign new_n746 = \40  & \1816 ;
  assign new_n747 = ~new_n745 & new_n746;
  assign new_n748 = \294  & new_n626;
  assign new_n749 = ~new_n585 & ~new_n748;
  assign new_n750 = ~new_n574 & new_n598;
  assign new_n751 = new_n584 & ~new_n750;
  assign new_n752 = new_n749 & ~new_n751;
  assign new_n753 = ~\294  & ~new_n626;
  assign new_n754 = ~new_n752 & ~new_n753;
  assign new_n755 = new_n747 & ~new_n754;
  assign new_n756 = new_n745 & new_n746;
  assign new_n757 = ~new_n597 & ~new_n756;
  assign new_n758 = \272  & ~new_n756;
  assign new_n759 = \309  & new_n756;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = ~\1819  & ~new_n760;
  assign new_n762 = \1819  & new_n760;
  assign new_n763 = \269  & ~new_n756;
  assign new_n764 = \305  & new_n756;
  assign new_n765 = ~new_n763 & ~new_n764;
  assign new_n766 = ~\1820  & ~new_n765;
  assign new_n767 = ~new_n762 & new_n766;
  assign new_n768 = ~new_n757 & ~new_n761;
  assign new_n769 = ~new_n767 & new_n768;
  assign new_n770 = \8  & ~new_n769;
  assign new_n771 = \263  & ~new_n756;
  assign new_n772 = \297  & new_n756;
  assign new_n773 = ~new_n771 & ~new_n772;
  assign new_n774 = \2010  & ~new_n773;
  assign new_n775 = \266  & ~new_n756;
  assign new_n776 = \301  & new_n756;
  assign new_n777 = ~new_n775 & ~new_n776;
  assign new_n778 = ~\1821  & ~new_n777;
  assign new_n779 = ~\2010  & new_n773;
  assign new_n780 = \287  & new_n756;
  assign new_n781 = \256  & ~new_n756;
  assign new_n782 = new_n374 & ~new_n780;
  assign new_n783 = ~new_n781 & new_n782;
  assign new_n784 = new_n413 & new_n783;
  assign new_n785 = \294  & new_n756;
  assign new_n786 = ~new_n413 & ~new_n783;
  assign new_n787 = \259  & ~new_n756;
  assign new_n788 = ~new_n785 & ~new_n787;
  assign new_n789 = ~new_n786 & new_n788;
  assign new_n790 = ~new_n779 & ~new_n784;
  assign new_n791 = ~new_n789 & new_n790;
  assign new_n792 = ~new_n774 & ~new_n778;
  assign new_n793 = ~new_n791 & new_n792;
  assign new_n794 = \1821  & new_n777;
  assign new_n795 = \1820  & new_n765;
  assign new_n796 = ~new_n762 & ~new_n795;
  assign new_n797 = \8  & ~new_n796;
  assign new_n798 = ~new_n794 & ~new_n797;
  assign new_n799 = ~new_n793 & new_n798;
  assign new_n800 = ~new_n770 & ~new_n799;
  assign new_n801 = ~new_n593 & ~new_n599;
  assign new_n802 = \8  & ~new_n594;
  assign new_n803 = ~new_n756 & new_n802;
  assign new_n804 = ~new_n801 & new_n803;
  assign new_n805 = ~new_n800 & ~new_n804;
  assign new_n806 = ~new_n574 & ~new_n600;
  assign new_n807 = new_n749 & new_n806;
  assign new_n808 = new_n747 & ~new_n807;
  assign new_n809 = ~new_n805 & ~new_n808;
  assign \3851  = new_n755 | new_n809;
  assign new_n811 = \1726  & ~\2970 ;
  assign new_n812 = ~\2925  & new_n811;
  assign new_n813 = ~\2971  & new_n812;
  assign new_n814 = ~\3671  & new_n813;
  assign \3881  = ~\3809  & new_n814;
  assign \3875  = 1'b0;
  assign \487  = ~\44 ;
  assign \488  = ~\132 ;
  assign \489  = ~\82 ;
  assign \490  = ~\96 ;
  assign \491  = ~\69 ;
  assign \492  = ~\120 ;
  assign \493  = ~\57 ;
  assign \494  = ~\108 ;
  assign \1448  = ~\1277 ;
  assign \2012  = ~\1821 ;
  assign \2014  = ~\1820 ;
  assign \2016  = ~\1819 ;
  assign \3079  = ~\3038 ;
  assign \3882  = ~\3881 ;
  assign \398  = \219 ;
  assign \400  = \219 ;
  assign \401  = \219 ;
  assign \419  = \253 ;
  assign \420  = \253 ;
  assign \456  = \290 ;
  assign \457  = \290 ;
  assign \458  = \290 ;
  assign \805  = \219 ;
  assign \2388  = \2387 ;
  assign \2390  = \2389 ;
  assign \2644  = \2643 ;
  assign \3804  = \3803 ;
endmodule


