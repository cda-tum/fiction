// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_, pv88_7_,
    pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_, pv56_15_,
    pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_, pv88_2_,
    pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_, pv88_16_,
    pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_, pv88_13_,
    pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_,
    pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_, pv56_7_,
    pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_, pv56_8_,
    pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_, pv56_1_,
    pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_, pv9_1_,
    pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_, pv24_12_,
    pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_, pv56_29_,
    pv9_0_, pv56_19_, pv56_28_,
    pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_, pv151_18_,
    pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_, pv119_20_,
    pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_, pv119_8_,
    pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_, pv151_28_,
    pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_, pv119_29_,
    pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_, pv151_21_,
    pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_, pv151_22_,
    pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_, pv151_31_,
    pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_, pv151_15_,
    pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_, pv151_10_,
    pv151_8_, pv151_11_  );
  input  pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_,
    pv88_7_, pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_,
    pv56_15_, pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_,
    pv88_2_, pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_,
    pv88_16_, pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_,
    pv88_13_, pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_,
    pv88_23_, pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_,
    pv56_7_, pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_,
    pv56_8_, pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_,
    pv56_1_, pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_,
    pv9_1_, pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_,
    pv24_12_, pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_,
    pv56_29_, pv9_0_, pv56_19_, pv56_28_;
  output pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_,
    pv151_18_, pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_,
    pv119_20_, pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_,
    pv119_8_, pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_,
    pv151_28_, pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_,
    pv119_29_, pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_,
    pv151_21_, pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_,
    pv151_22_, pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_,
    pv151_31_, pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_,
    pv151_15_, pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_,
    pv151_10_, pv151_8_, pv151_11_;
  wire new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n455, new_n456, new_n457, new_n458,
    new_n459, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769;
  assign new_n152 = pv9_8_ & pv9_1_;
  assign new_n153 = ~pv9_10_ & new_n152;
  assign new_n154 = ~pv9_6_ & ~pv9_2_;
  assign new_n155 = ~pv9_5_ & new_n154;
  assign new_n156 = pv9_1_ & new_n155;
  assign new_n157 = ~pv9_10_ & new_n156;
  assign new_n158 = pv9_2_ & pv9_0_;
  assign new_n159 = ~pv9_5_ & new_n158;
  assign new_n160 = ~pv9_1_ & new_n159;
  assign new_n161 = ~pv9_10_ & new_n160;
  assign new_n162 = ~pv9_6_ & new_n161;
  assign new_n163 = pv9_2_ & ~pv9_3_;
  assign new_n164 = pv9_1_ & new_n163;
  assign new_n165 = ~pv9_10_ & new_n164;
  assign new_n166 = pv9_8_ & pv9_2_;
  assign new_n167 = ~pv9_1_ & new_n166;
  assign new_n168 = ~pv9_10_ & new_n167;
  assign new_n169 = ~pv9_1_ & ~pv9_2_;
  assign new_n170 = pv9_10_ & new_n169;
  assign new_n171 = ~pv9_5_ & ~pv9_2_;
  assign new_n172 = ~pv9_1_ & new_n171;
  assign new_n173 = ~pv9_6_ & new_n172;
  assign new_n174 = pv9_7_ & new_n169;
  assign new_n175 = pv9_10_ & pv9_2_;
  assign new_n176 = pv9_1_ & pv9_2_;
  assign new_n177 = pv9_3_ & new_n176;
  assign new_n178 = pv9_10_ & pv9_1_;
  assign new_n179 = ~pv9_5_ & ~pv9_0_;
  assign new_n180 = ~pv9_10_ & new_n179;
  assign new_n181 = pv9_7_ & ~pv9_0_;
  assign new_n182 = ~pv9_10_ & new_n181;
  assign new_n183 = ~new_n153 & ~new_n157;
  assign new_n184 = ~new_n162 & ~new_n165;
  assign new_n185 = new_n183 & new_n184;
  assign new_n186 = ~new_n168 & ~new_n170;
  assign new_n187 = ~new_n173 & new_n186;
  assign new_n188 = new_n185 & new_n187;
  assign new_n189 = ~new_n178 & ~new_n180;
  assign new_n190 = ~new_n182 & new_n189;
  assign new_n191 = ~new_n174 & ~new_n175;
  assign new_n192 = ~new_n177 & new_n191;
  assign new_n193 = new_n190 & new_n192;
  assign new_n194 = new_n188 & new_n193;
  assign new_n195 = ~new_n157 & ~new_n180;
  assign new_n196 = ~new_n173 & ~new_n174;
  assign new_n197 = new_n195 & new_n196;
  assign new_n198 = ~new_n170 & ~new_n182;
  assign new_n199 = ~new_n153 & new_n198;
  assign new_n200 = new_n197 & new_n199;
  assign new_n201 = ~new_n170 & ~new_n174;
  assign new_n202 = ~new_n168 & new_n201;
  assign new_n203 = ~new_n173 & new_n184;
  assign new_n204 = new_n202 & new_n203;
  assign new_n205 = ~new_n194 & new_n200;
  assign new_n206 = new_n204 & new_n205;
  assign new_n207 = pv56_2_ & new_n206;
  assign new_n208 = ~new_n204 & new_n205;
  assign new_n209 = pv88_2_ & new_n208;
  assign new_n210 = ~new_n200 & new_n204;
  assign new_n211 = ~new_n194 & new_n210;
  assign new_n212 = ~new_n194 & ~new_n200;
  assign new_n213 = ~new_n204 & new_n212;
  assign new_n214 = pv24_1_ & new_n213;
  assign new_n215 = ~new_n211 & ~new_n214;
  assign new_n216 = ~new_n194 & ~new_n207;
  assign new_n217 = ~new_n209 & new_n216;
  assign pv119_1_ = ~new_n215 | ~new_n217;
  assign new_n219 = pv56_1_ & new_n206;
  assign new_n220 = pv88_1_ & new_n208;
  assign new_n221 = pv24_0_ & new_n213;
  assign new_n222 = ~new_n211 & ~new_n221;
  assign new_n223 = ~new_n194 & ~new_n219;
  assign new_n224 = ~new_n220 & new_n223;
  assign pv119_0_ = ~new_n222 | ~new_n224;
  assign new_n226 = pv56_4_ & new_n206;
  assign new_n227 = pv88_4_ & new_n208;
  assign new_n228 = pv24_3_ & new_n213;
  assign new_n229 = ~new_n211 & ~new_n228;
  assign new_n230 = ~new_n194 & ~new_n226;
  assign new_n231 = ~new_n227 & new_n230;
  assign pv119_3_ = ~new_n229 | ~new_n231;
  assign new_n233 = pv56_31_ & new_n206;
  assign new_n234 = pv56_20_ & new_n208;
  assign new_n235 = pv56_23_ & new_n211;
  assign new_n236 = pv56_16_ & new_n213;
  assign new_n237 = ~new_n235 & ~new_n236;
  assign new_n238 = ~new_n194 & ~new_n233;
  assign new_n239 = ~new_n234 & new_n238;
  assign pv119_30_ = ~new_n237 | ~new_n239;
  assign new_n241 = pv56_3_ & new_n206;
  assign new_n242 = pv88_3_ & new_n208;
  assign new_n243 = pv24_2_ & new_n213;
  assign new_n244 = ~new_n211 & ~new_n243;
  assign new_n245 = ~new_n194 & ~new_n241;
  assign new_n246 = ~new_n242 & new_n245;
  assign pv119_2_ = ~new_n244 | ~new_n246;
  assign new_n248 = pv88_1_ & new_n206;
  assign new_n249 = ~new_n200 & ~new_n204;
  assign new_n250 = new_n194 & new_n249;
  assign new_n251 = pv56_22_ & new_n208;
  assign new_n252 = new_n204 & new_n212;
  assign new_n253 = pv56_25_ & new_n252;
  assign new_n254 = pv56_18_ & new_n213;
  assign new_n255 = new_n200 & new_n204;
  assign new_n256 = new_n194 & new_n255;
  assign new_n257 = new_n200 & ~new_n204;
  assign new_n258 = new_n194 & new_n257;
  assign new_n259 = new_n194 & new_n210;
  assign new_n260 = ~new_n258 & ~new_n259;
  assign new_n261 = ~new_n254 & ~new_n256;
  assign new_n262 = new_n260 & new_n261;
  assign new_n263 = ~new_n248 & ~new_n250;
  assign new_n264 = ~new_n251 & ~new_n253;
  assign new_n265 = new_n263 & new_n264;
  assign pv151_1_ = ~new_n262 | ~new_n265;
  assign new_n267 = pv88_18_ & new_n206;
  assign new_n268 = pv88_7_ & new_n208;
  assign new_n269 = pv88_10_ & new_n252;
  assign new_n270 = pv88_3_ & new_n213;
  assign new_n271 = ~new_n256 & ~new_n270;
  assign new_n272 = new_n260 & new_n271;
  assign new_n273 = ~new_n250 & ~new_n267;
  assign new_n274 = ~new_n268 & ~new_n269;
  assign new_n275 = new_n273 & new_n274;
  assign pv151_18_ = ~new_n272 | ~new_n275;
  assign new_n277 = pv88_0_ & new_n206;
  assign new_n278 = pv56_21_ & new_n208;
  assign new_n279 = pv56_24_ & new_n252;
  assign new_n280 = pv56_17_ & new_n213;
  assign new_n281 = ~new_n256 & ~new_n280;
  assign new_n282 = new_n260 & new_n281;
  assign new_n283 = ~new_n250 & ~new_n277;
  assign new_n284 = ~new_n278 & ~new_n279;
  assign new_n285 = new_n283 & new_n284;
  assign pv151_0_ = ~new_n282 | ~new_n285;
  assign new_n287 = pv88_19_ & new_n206;
  assign new_n288 = pv88_8_ & new_n208;
  assign new_n289 = pv88_11_ & new_n252;
  assign new_n290 = pv88_4_ & new_n213;
  assign new_n291 = ~new_n256 & ~new_n290;
  assign new_n292 = new_n260 & new_n291;
  assign new_n293 = ~new_n250 & ~new_n287;
  assign new_n294 = ~new_n288 & ~new_n289;
  assign new_n295 = new_n293 & new_n294;
  assign pv151_19_ = ~new_n292 | ~new_n295;
  assign new_n297 = pv56_22_ & new_n206;
  assign new_n298 = pv56_11_ & new_n208;
  assign new_n299 = pv56_14_ & new_n211;
  assign new_n300 = pv56_7_ & new_n213;
  assign new_n301 = ~new_n299 & ~new_n300;
  assign new_n302 = ~new_n194 & ~new_n297;
  assign new_n303 = ~new_n298 & new_n302;
  assign pv119_21_ = ~new_n301 | ~new_n303;
  assign new_n305 = pv88_3_ & new_n206;
  assign new_n306 = pv56_24_ & new_n208;
  assign new_n307 = pv56_27_ & new_n252;
  assign new_n308 = pv56_20_ & new_n213;
  assign new_n309 = ~new_n256 & ~new_n308;
  assign new_n310 = new_n260 & new_n309;
  assign new_n311 = ~new_n250 & ~new_n305;
  assign new_n312 = ~new_n306 & ~new_n307;
  assign new_n313 = new_n311 & new_n312;
  assign pv151_3_ = ~new_n310 | ~new_n313;
  assign new_n315 = pv88_16_ & new_n206;
  assign new_n316 = pv88_5_ & new_n208;
  assign new_n317 = pv88_8_ & new_n252;
  assign new_n318 = pv88_1_ & new_n213;
  assign new_n319 = ~new_n256 & ~new_n318;
  assign new_n320 = new_n260 & new_n319;
  assign new_n321 = ~new_n250 & ~new_n315;
  assign new_n322 = ~new_n316 & ~new_n317;
  assign new_n323 = new_n321 & new_n322;
  assign pv151_16_ = ~new_n320 | ~new_n323;
  assign new_n325 = pv56_21_ & new_n206;
  assign new_n326 = pv56_10_ & new_n208;
  assign new_n327 = pv56_13_ & new_n211;
  assign new_n328 = pv56_6_ & new_n213;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = ~new_n194 & ~new_n325;
  assign new_n331 = ~new_n326 & new_n330;
  assign pv119_20_ = ~new_n329 | ~new_n331;
  assign new_n333 = pv88_2_ & new_n206;
  assign new_n334 = pv56_23_ & new_n208;
  assign new_n335 = pv56_26_ & new_n252;
  assign new_n336 = pv56_19_ & new_n213;
  assign new_n337 = ~new_n256 & ~new_n336;
  assign new_n338 = new_n260 & new_n337;
  assign new_n339 = ~new_n250 & ~new_n333;
  assign new_n340 = ~new_n334 & ~new_n335;
  assign new_n341 = new_n339 & new_n340;
  assign pv151_2_ = ~new_n338 | ~new_n341;
  assign new_n343 = pv88_17_ & new_n206;
  assign new_n344 = pv88_6_ & new_n208;
  assign new_n345 = pv88_9_ & new_n252;
  assign new_n346 = pv88_2_ & new_n213;
  assign new_n347 = ~new_n256 & ~new_n346;
  assign new_n348 = new_n260 & new_n347;
  assign new_n349 = ~new_n250 & ~new_n343;
  assign new_n350 = ~new_n344 & ~new_n345;
  assign new_n351 = new_n349 & new_n350;
  assign pv151_17_ = ~new_n348 | ~new_n351;
  assign new_n353 = pv56_10_ & new_n206;
  assign new_n354 = pv88_10_ & new_n208;
  assign new_n355 = pv56_2_ & new_n211;
  assign new_n356 = pv24_9_ & new_n213;
  assign new_n357 = ~new_n355 & ~new_n356;
  assign new_n358 = ~new_n194 & ~new_n353;
  assign new_n359 = ~new_n354 & new_n358;
  assign pv119_9_ = ~new_n357 | ~new_n359;
  assign new_n361 = pv56_24_ & new_n206;
  assign new_n362 = pv56_13_ & new_n208;
  assign new_n363 = pv56_16_ & new_n211;
  assign new_n364 = pv56_9_ & new_n213;
  assign new_n365 = ~new_n363 & ~new_n364;
  assign new_n366 = ~new_n194 & ~new_n361;
  assign new_n367 = ~new_n362 & new_n366;
  assign pv119_23_ = ~new_n365 | ~new_n367;
  assign new_n369 = pv88_27_ & new_n206;
  assign new_n370 = pv88_16_ & new_n208;
  assign new_n371 = pv88_19_ & new_n252;
  assign new_n372 = pv88_12_ & new_n213;
  assign new_n373 = ~new_n256 & ~new_n372;
  assign new_n374 = new_n260 & new_n373;
  assign new_n375 = ~new_n250 & ~new_n369;
  assign new_n376 = ~new_n370 & ~new_n371;
  assign new_n377 = new_n375 & new_n376;
  assign pv151_27_ = ~new_n374 | ~new_n377;
  assign new_n379 = pv56_9_ & new_n206;
  assign new_n380 = pv88_9_ & new_n208;
  assign new_n381 = pv56_1_ & new_n211;
  assign new_n382 = pv24_8_ & new_n213;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = ~new_n194 & ~new_n379;
  assign new_n385 = ~new_n380 & new_n384;
  assign pv119_8_ = ~new_n383 | ~new_n385;
  assign new_n387 = pv56_23_ & new_n206;
  assign new_n388 = pv56_12_ & new_n208;
  assign new_n389 = pv56_15_ & new_n211;
  assign new_n390 = pv56_8_ & new_n213;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = ~new_n194 & ~new_n387;
  assign new_n393 = ~new_n388 & new_n392;
  assign pv119_22_ = ~new_n391 | ~new_n393;
  assign new_n395 = pv88_26_ & new_n206;
  assign new_n396 = pv88_15_ & new_n208;
  assign new_n397 = pv88_18_ & new_n252;
  assign new_n398 = pv88_11_ & new_n213;
  assign new_n399 = ~new_n256 & ~new_n398;
  assign new_n400 = new_n260 & new_n399;
  assign new_n401 = ~new_n250 & ~new_n395;
  assign new_n402 = ~new_n396 & ~new_n397;
  assign new_n403 = new_n401 & new_n402;
  assign pv151_26_ = ~new_n400 | ~new_n403;
  assign new_n405 = pv56_26_ & new_n206;
  assign new_n406 = pv56_15_ & new_n208;
  assign new_n407 = pv56_18_ & new_n211;
  assign new_n408 = pv56_11_ & new_n213;
  assign new_n409 = ~new_n407 & ~new_n408;
  assign new_n410 = ~new_n194 & ~new_n405;
  assign new_n411 = ~new_n406 & new_n410;
  assign pv119_25_ = ~new_n409 | ~new_n411;
  assign new_n413 = pv88_29_ & new_n206;
  assign new_n414 = pv88_18_ & new_n208;
  assign new_n415 = pv88_21_ & new_n252;
  assign new_n416 = pv88_14_ & new_n213;
  assign new_n417 = ~new_n256 & ~new_n416;
  assign new_n418 = new_n260 & new_n417;
  assign new_n419 = ~new_n250 & ~new_n413;
  assign new_n420 = ~new_n414 & ~new_n415;
  assign new_n421 = new_n419 & new_n420;
  assign pv151_29_ = ~new_n418 | ~new_n421;
  assign new_n423 = pv56_25_ & new_n206;
  assign new_n424 = pv56_14_ & new_n208;
  assign new_n425 = pv56_17_ & new_n211;
  assign new_n426 = pv56_10_ & new_n213;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = ~new_n194 & ~new_n423;
  assign new_n429 = ~new_n424 & new_n428;
  assign pv119_24_ = ~new_n427 | ~new_n429;
  assign new_n431 = pv88_28_ & new_n206;
  assign new_n432 = pv88_17_ & new_n208;
  assign new_n433 = pv88_20_ & new_n252;
  assign new_n434 = pv88_13_ & new_n213;
  assign new_n435 = ~new_n256 & ~new_n434;
  assign new_n436 = new_n260 & new_n435;
  assign new_n437 = ~new_n250 & ~new_n431;
  assign new_n438 = ~new_n432 & ~new_n433;
  assign new_n439 = new_n437 & new_n438;
  assign pv151_28_ = ~new_n436 | ~new_n439;
  assign new_n441 = pv56_6_ & new_n206;
  assign new_n442 = pv24_5_ & new_n213;
  assign new_n443 = ~new_n211 & ~new_n442;
  assign new_n444 = ~new_n194 & ~new_n441;
  assign new_n445 = ~new_n344 & new_n444;
  assign pv119_5_ = ~new_n443 | ~new_n445;
  assign new_n447 = pv56_28_ & new_n206;
  assign new_n448 = pv56_17_ & new_n208;
  assign new_n449 = pv56_20_ & new_n211;
  assign new_n450 = pv56_13_ & new_n213;
  assign new_n451 = ~new_n449 & ~new_n450;
  assign new_n452 = ~new_n194 & ~new_n447;
  assign new_n453 = ~new_n448 & new_n452;
  assign pv119_27_ = ~new_n451 | ~new_n453;
  assign new_n455 = pv56_5_ & new_n206;
  assign new_n456 = pv24_4_ & new_n213;
  assign new_n457 = ~new_n211 & ~new_n456;
  assign new_n458 = ~new_n194 & ~new_n455;
  assign new_n459 = ~new_n316 & new_n458;
  assign pv119_4_ = ~new_n457 | ~new_n459;
  assign new_n461 = pv56_27_ & new_n206;
  assign new_n462 = pv56_16_ & new_n208;
  assign new_n463 = pv56_19_ & new_n211;
  assign new_n464 = pv56_12_ & new_n213;
  assign new_n465 = ~new_n463 & ~new_n464;
  assign new_n466 = ~new_n194 & ~new_n461;
  assign new_n467 = ~new_n462 & new_n466;
  assign pv119_26_ = ~new_n465 | ~new_n467;
  assign new_n469 = pv56_8_ & new_n206;
  assign new_n470 = pv56_0_ & new_n211;
  assign new_n471 = pv24_7_ & new_n213;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = ~new_n194 & ~new_n469;
  assign new_n474 = ~new_n288 & new_n473;
  assign pv119_7_ = ~new_n472 | ~new_n474;
  assign new_n476 = pv56_30_ & new_n206;
  assign new_n477 = pv56_19_ & new_n208;
  assign new_n478 = pv56_22_ & new_n211;
  assign new_n479 = pv56_15_ & new_n213;
  assign new_n480 = ~new_n478 & ~new_n479;
  assign new_n481 = ~new_n194 & ~new_n476;
  assign new_n482 = ~new_n477 & new_n481;
  assign pv119_29_ = ~new_n480 | ~new_n482;
  assign new_n484 = pv56_7_ & new_n206;
  assign new_n485 = pv24_6_ & new_n213;
  assign new_n486 = ~new_n211 & ~new_n485;
  assign new_n487 = ~new_n194 & ~new_n484;
  assign new_n488 = ~new_n268 & new_n487;
  assign pv119_6_ = ~new_n486 | ~new_n488;
  assign new_n490 = pv56_29_ & new_n206;
  assign new_n491 = pv56_18_ & new_n208;
  assign new_n492 = pv56_21_ & new_n211;
  assign new_n493 = pv56_14_ & new_n213;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = ~new_n194 & ~new_n490;
  assign new_n496 = ~new_n491 & new_n495;
  assign pv119_28_ = ~new_n494 | ~new_n496;
  assign new_n498 = pv56_19_ & new_n206;
  assign new_n499 = pv56_8_ & new_n208;
  assign new_n500 = pv56_11_ & new_n211;
  assign new_n501 = pv56_4_ & new_n213;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = ~new_n194 & ~new_n498;
  assign new_n504 = ~new_n499 & new_n503;
  assign pv119_18_ = ~new_n502 | ~new_n504;
  assign new_n506 = pv56_20_ & new_n206;
  assign new_n507 = pv56_9_ & new_n208;
  assign new_n508 = pv56_12_ & new_n211;
  assign new_n509 = pv56_5_ & new_n213;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = ~new_n194 & ~new_n506;
  assign new_n512 = ~new_n507 & new_n511;
  assign pv119_19_ = ~new_n510 | ~new_n512;
  assign new_n514 = pv56_17_ & new_n206;
  assign new_n515 = pv56_6_ & new_n208;
  assign new_n516 = pv56_9_ & new_n211;
  assign new_n517 = pv56_2_ & new_n213;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = ~new_n194 & ~new_n514;
  assign new_n520 = ~new_n515 & new_n519;
  assign pv119_16_ = ~new_n518 | ~new_n520;
  assign new_n522 = pv88_21_ & new_n206;
  assign new_n523 = pv88_13_ & new_n252;
  assign new_n524 = pv88_6_ & new_n213;
  assign new_n525 = ~new_n256 & ~new_n524;
  assign new_n526 = new_n260 & new_n525;
  assign new_n527 = ~new_n250 & ~new_n522;
  assign new_n528 = ~new_n354 & ~new_n523;
  assign new_n529 = new_n527 & new_n528;
  assign pv151_21_ = ~new_n526 | ~new_n529;
  assign new_n531 = pv56_18_ & new_n206;
  assign new_n532 = pv56_7_ & new_n208;
  assign new_n533 = pv56_10_ & new_n211;
  assign new_n534 = pv56_3_ & new_n213;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign new_n536 = ~new_n194 & ~new_n531;
  assign new_n537 = ~new_n532 & new_n536;
  assign pv119_17_ = ~new_n535 | ~new_n537;
  assign new_n539 = pv88_20_ & new_n206;
  assign new_n540 = pv88_12_ & new_n252;
  assign new_n541 = pv88_5_ & new_n213;
  assign new_n542 = ~new_n256 & ~new_n541;
  assign new_n543 = new_n260 & new_n542;
  assign new_n544 = ~new_n250 & ~new_n539;
  assign new_n545 = ~new_n380 & ~new_n540;
  assign new_n546 = new_n544 & new_n545;
  assign pv151_20_ = ~new_n543 | ~new_n546;
  assign new_n548 = pv56_15_ & new_n206;
  assign new_n549 = pv56_4_ & new_n208;
  assign new_n550 = pv56_7_ & new_n211;
  assign new_n551 = pv24_14_ & new_n213;
  assign new_n552 = ~new_n550 & ~new_n551;
  assign new_n553 = ~new_n194 & ~new_n548;
  assign new_n554 = ~new_n549 & new_n553;
  assign pv119_14_ = ~new_n552 | ~new_n554;
  assign new_n556 = pv88_23_ & new_n206;
  assign new_n557 = pv88_12_ & new_n208;
  assign new_n558 = pv88_15_ & new_n252;
  assign new_n559 = pv88_8_ & new_n213;
  assign new_n560 = ~new_n256 & ~new_n559;
  assign new_n561 = new_n260 & new_n560;
  assign new_n562 = ~new_n250 & ~new_n556;
  assign new_n563 = ~new_n557 & ~new_n558;
  assign new_n564 = new_n562 & new_n563;
  assign pv151_23_ = ~new_n561 | ~new_n564;
  assign new_n566 = pv56_16_ & new_n206;
  assign new_n567 = pv56_5_ & new_n208;
  assign new_n568 = pv56_8_ & new_n211;
  assign new_n569 = pv56_1_ & new_n213;
  assign new_n570 = ~new_n568 & ~new_n569;
  assign new_n571 = ~new_n194 & ~new_n566;
  assign new_n572 = ~new_n567 & new_n571;
  assign pv119_15_ = ~new_n570 | ~new_n572;
  assign new_n574 = pv88_22_ & new_n206;
  assign new_n575 = pv88_11_ & new_n208;
  assign new_n576 = pv88_14_ & new_n252;
  assign new_n577 = pv88_7_ & new_n213;
  assign new_n578 = ~new_n256 & ~new_n577;
  assign new_n579 = new_n260 & new_n578;
  assign new_n580 = ~new_n250 & ~new_n574;
  assign new_n581 = ~new_n575 & ~new_n576;
  assign new_n582 = new_n580 & new_n581;
  assign pv151_22_ = ~new_n579 | ~new_n582;
  assign new_n584 = pv56_13_ & new_n206;
  assign new_n585 = pv56_2_ & new_n208;
  assign new_n586 = pv56_5_ & new_n211;
  assign new_n587 = pv24_12_ & new_n213;
  assign new_n588 = ~new_n586 & ~new_n587;
  assign new_n589 = ~new_n194 & ~new_n584;
  assign new_n590 = ~new_n585 & new_n589;
  assign pv119_12_ = ~new_n588 | ~new_n590;
  assign new_n592 = pv88_25_ & new_n206;
  assign new_n593 = pv88_14_ & new_n208;
  assign new_n594 = pv88_17_ & new_n252;
  assign new_n595 = pv88_10_ & new_n213;
  assign new_n596 = ~new_n256 & ~new_n595;
  assign new_n597 = new_n260 & new_n596;
  assign new_n598 = ~new_n250 & ~new_n592;
  assign new_n599 = ~new_n593 & ~new_n594;
  assign new_n600 = new_n598 & new_n599;
  assign pv151_25_ = ~new_n597 | ~new_n600;
  assign new_n602 = pv88_30_ & new_n206;
  assign new_n603 = pv88_19_ & new_n208;
  assign new_n604 = pv88_22_ & new_n252;
  assign new_n605 = pv88_15_ & new_n213;
  assign new_n606 = ~new_n256 & ~new_n605;
  assign new_n607 = new_n260 & new_n606;
  assign new_n608 = ~new_n250 & ~new_n602;
  assign new_n609 = ~new_n603 & ~new_n604;
  assign new_n610 = new_n608 & new_n609;
  assign pv151_30_ = ~new_n607 | ~new_n610;
  assign new_n612 = pv56_14_ & new_n206;
  assign new_n613 = pv56_3_ & new_n208;
  assign new_n614 = pv56_6_ & new_n211;
  assign new_n615 = pv24_13_ & new_n213;
  assign new_n616 = ~new_n614 & ~new_n615;
  assign new_n617 = ~new_n194 & ~new_n612;
  assign new_n618 = ~new_n613 & new_n617;
  assign pv119_13_ = ~new_n616 | ~new_n618;
  assign new_n620 = pv88_24_ & new_n206;
  assign new_n621 = pv88_13_ & new_n208;
  assign new_n622 = pv88_16_ & new_n252;
  assign new_n623 = pv88_9_ & new_n213;
  assign new_n624 = ~new_n256 & ~new_n623;
  assign new_n625 = new_n260 & new_n624;
  assign new_n626 = ~new_n250 & ~new_n620;
  assign new_n627 = ~new_n621 & ~new_n622;
  assign new_n628 = new_n626 & new_n627;
  assign pv151_24_ = ~new_n625 | ~new_n628;
  assign new_n630 = pv88_31_ & new_n206;
  assign new_n631 = pv88_20_ & new_n208;
  assign new_n632 = pv88_23_ & new_n252;
  assign new_n633 = pv88_16_ & new_n213;
  assign new_n634 = ~new_n256 & ~new_n633;
  assign new_n635 = new_n260 & new_n634;
  assign new_n636 = ~new_n250 & ~new_n630;
  assign new_n637 = ~new_n631 & ~new_n632;
  assign new_n638 = new_n636 & new_n637;
  assign pv151_31_ = ~new_n635 | ~new_n638;
  assign new_n640 = pv56_11_ & new_n206;
  assign new_n641 = pv56_3_ & new_n211;
  assign new_n642 = pv24_10_ & new_n213;
  assign new_n643 = ~new_n641 & ~new_n642;
  assign new_n644 = ~new_n194 & ~new_n640;
  assign new_n645 = ~new_n575 & new_n644;
  assign pv119_10_ = ~new_n643 | ~new_n645;
  assign new_n647 = pv88_5_ & new_n206;
  assign new_n648 = pv56_26_ & new_n208;
  assign new_n649 = pv56_29_ & new_n252;
  assign new_n650 = pv56_22_ & new_n213;
  assign new_n651 = ~new_n256 & ~new_n650;
  assign new_n652 = new_n260 & new_n651;
  assign new_n653 = ~new_n250 & ~new_n647;
  assign new_n654 = ~new_n648 & ~new_n649;
  assign new_n655 = new_n653 & new_n654;
  assign pv151_5_ = ~new_n652 | ~new_n655;
  assign new_n657 = pv88_14_ & new_n206;
  assign new_n658 = pv88_6_ & new_n252;
  assign new_n659 = pv56_31_ & new_n213;
  assign new_n660 = ~new_n256 & ~new_n659;
  assign new_n661 = new_n260 & new_n660;
  assign new_n662 = ~new_n250 & ~new_n657;
  assign new_n663 = ~new_n242 & ~new_n658;
  assign new_n664 = new_n662 & new_n663;
  assign pv151_14_ = ~new_n661 | ~new_n664;
  assign new_n666 = pv56_12_ & new_n206;
  assign new_n667 = pv56_1_ & new_n208;
  assign new_n668 = pv56_4_ & new_n211;
  assign new_n669 = pv24_11_ & new_n213;
  assign new_n670 = ~new_n668 & ~new_n669;
  assign new_n671 = ~new_n194 & ~new_n666;
  assign new_n672 = ~new_n667 & new_n671;
  assign pv119_11_ = ~new_n670 | ~new_n672;
  assign new_n674 = pv88_4_ & new_n206;
  assign new_n675 = pv56_25_ & new_n208;
  assign new_n676 = pv56_28_ & new_n252;
  assign new_n677 = pv56_21_ & new_n213;
  assign new_n678 = ~new_n256 & ~new_n677;
  assign new_n679 = new_n260 & new_n678;
  assign new_n680 = ~new_n250 & ~new_n674;
  assign new_n681 = ~new_n675 & ~new_n676;
  assign new_n682 = new_n680 & new_n681;
  assign pv151_4_ = ~new_n679 | ~new_n682;
  assign new_n684 = pv88_15_ & new_n206;
  assign new_n685 = pv88_7_ & new_n252;
  assign new_n686 = pv88_0_ & new_n213;
  assign new_n687 = ~new_n256 & ~new_n686;
  assign new_n688 = new_n260 & new_n687;
  assign new_n689 = ~new_n250 & ~new_n684;
  assign new_n690 = ~new_n227 & ~new_n685;
  assign new_n691 = new_n689 & new_n690;
  assign pv151_15_ = ~new_n688 | ~new_n691;
  assign new_n693 = pv88_7_ & new_n206;
  assign new_n694 = pv56_28_ & new_n208;
  assign new_n695 = pv56_31_ & new_n252;
  assign new_n696 = pv56_24_ & new_n213;
  assign new_n697 = ~new_n256 & ~new_n696;
  assign new_n698 = new_n260 & new_n697;
  assign new_n699 = ~new_n250 & ~new_n693;
  assign new_n700 = ~new_n694 & ~new_n695;
  assign new_n701 = new_n699 & new_n700;
  assign pv151_7_ = ~new_n698 | ~new_n701;
  assign new_n703 = pv88_12_ & new_n206;
  assign new_n704 = pv88_4_ & new_n252;
  assign new_n705 = pv56_29_ & new_n213;
  assign new_n706 = ~new_n256 & ~new_n705;
  assign new_n707 = new_n260 & new_n706;
  assign new_n708 = ~new_n250 & ~new_n703;
  assign new_n709 = ~new_n220 & ~new_n704;
  assign new_n710 = new_n708 & new_n709;
  assign pv151_12_ = ~new_n707 | ~new_n710;
  assign new_n712 = pv88_6_ & new_n206;
  assign new_n713 = pv56_27_ & new_n208;
  assign new_n714 = pv56_30_ & new_n252;
  assign new_n715 = pv56_23_ & new_n213;
  assign new_n716 = ~new_n256 & ~new_n715;
  assign new_n717 = new_n260 & new_n716;
  assign new_n718 = ~new_n250 & ~new_n712;
  assign new_n719 = ~new_n713 & ~new_n714;
  assign new_n720 = new_n718 & new_n719;
  assign pv151_6_ = ~new_n717 | ~new_n720;
  assign new_n722 = pv88_13_ & new_n206;
  assign new_n723 = pv88_5_ & new_n252;
  assign new_n724 = pv56_30_ & new_n213;
  assign new_n725 = ~new_n256 & ~new_n724;
  assign new_n726 = new_n260 & new_n725;
  assign new_n727 = ~new_n250 & ~new_n722;
  assign new_n728 = ~new_n209 & ~new_n723;
  assign new_n729 = new_n727 & new_n728;
  assign pv151_13_ = ~new_n726 | ~new_n729;
  assign new_n731 = pv88_9_ & new_n206;
  assign new_n732 = pv56_30_ & new_n208;
  assign new_n733 = pv88_1_ & new_n252;
  assign new_n734 = pv56_26_ & new_n213;
  assign new_n735 = ~new_n256 & ~new_n734;
  assign new_n736 = new_n260 & new_n735;
  assign new_n737 = ~new_n250 & ~new_n731;
  assign new_n738 = ~new_n732 & ~new_n733;
  assign new_n739 = new_n737 & new_n738;
  assign pv151_9_ = ~new_n736 | ~new_n739;
  assign new_n741 = pv88_10_ & new_n206;
  assign new_n742 = pv56_31_ & new_n208;
  assign new_n743 = pv88_2_ & new_n252;
  assign new_n744 = pv56_27_ & new_n213;
  assign new_n745 = ~new_n256 & ~new_n744;
  assign new_n746 = new_n260 & new_n745;
  assign new_n747 = ~new_n250 & ~new_n741;
  assign new_n748 = ~new_n742 & ~new_n743;
  assign new_n749 = new_n747 & new_n748;
  assign pv151_10_ = ~new_n746 | ~new_n749;
  assign new_n751 = pv88_8_ & new_n206;
  assign new_n752 = pv56_29_ & new_n208;
  assign new_n753 = pv88_0_ & new_n252;
  assign new_n754 = pv56_25_ & new_n213;
  assign new_n755 = ~new_n256 & ~new_n754;
  assign new_n756 = new_n260 & new_n755;
  assign new_n757 = ~new_n250 & ~new_n751;
  assign new_n758 = ~new_n752 & ~new_n753;
  assign new_n759 = new_n757 & new_n758;
  assign pv151_8_ = ~new_n756 | ~new_n759;
  assign new_n761 = pv88_11_ & new_n206;
  assign new_n762 = pv88_0_ & new_n208;
  assign new_n763 = pv88_3_ & new_n252;
  assign new_n764 = pv56_28_ & new_n213;
  assign new_n765 = ~new_n256 & ~new_n764;
  assign new_n766 = new_n260 & new_n765;
  assign new_n767 = ~new_n250 & ~new_n761;
  assign new_n768 = ~new_n762 & ~new_n763;
  assign new_n769 = new_n767 & new_n768;
  assign pv151_11_ = ~new_n766 | ~new_n769;
endmodule


