// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    p0, q1, r2, s3, a, p1, q0, r3, s2, b, p2, q3, r0, s1, c, p3, q2, r1,
    s0, d, t0, u1, v2, w3, e, t1, u0, v3, w2, f, t2, u3, v0, w1, g, t3, u2,
    v1, w0, h, x0, y1, z2, i, x1, y0, z3, j, x2, y3, z0, k, x3, y2, z1, l,
    m, n, o, a1, b2, c3, d4, p, a0, b3, c2, e4, q, a3, b0, c1, r, a2, b1,
    c0, s, d0, e1, f2, g3, t, a4, d1, e0, f3, g2, u, b4, d2, e3, f0, g1, v,
    c4, d3, e2, f1, g0, w, h0, i1, j2, k3, x, h1, i0, j3, k2, y, h2, i3,
    j0, k1, z, h3, i2, j1, k0, l0, m1, n2, o3, l1, m0, n3, o2, l2, m3, n0,
    o1, l3, m2, n1, o0,
    t4, u5, v6, w7, t5, u4, v7, w6, t6, u7, v4, w5, t7, u6, v5, w4, p4, q5,
    r6, s7, p5, q4, r7, s6, p6, q7, r4, s5, p7, q6, r5, s4, x4, y5, z6, x5,
    y4, z7, x6, y7, z4, x7, y6, z5, e5, f6, g7, h8, d5, f7, g6, d6, e7, f4,
    g5, d7, e6, f5, g4, a5, b6, c7, b7, c6, a7, c5, a6, b5, l4, m5, n6, o7,
    a8, l5, m4, n7, o6, b8, l6, m7, n4, o5, c8, l7, m6, n5, o4, d8, h4, i5,
    j6, k7, e8, h5, i4, j7, k6, f8, h6, i7, j4, k5, g8, h7, i6, j5, k4  );
  input  p0, q1, r2, s3, a, p1, q0, r3, s2, b, p2, q3, r0, s1, c, p3, q2,
    r1, s0, d, t0, u1, v2, w3, e, t1, u0, v3, w2, f, t2, u3, v0, w1, g, t3,
    u2, v1, w0, h, x0, y1, z2, i, x1, y0, z3, j, x2, y3, z0, k, x3, y2, z1,
    l, m, n, o, a1, b2, c3, d4, p, a0, b3, c2, e4, q, a3, b0, c1, r, a2,
    b1, c0, s, d0, e1, f2, g3, t, a4, d1, e0, f3, g2, u, b4, d2, e3, f0,
    g1, v, c4, d3, e2, f1, g0, w, h0, i1, j2, k3, x, h1, i0, j3, k2, y, h2,
    i3, j0, k1, z, h3, i2, j1, k0, l0, m1, n2, o3, l1, m0, n3, o2, l2, m3,
    n0, o1, l3, m2, n1, o0;
  output t4, u5, v6, w7, t5, u4, v7, w6, t6, u7, v4, w5, t7, u6, v5, w4, p4,
    q5, r6, s7, p5, q4, r7, s6, p6, q7, r4, s5, p7, q6, r5, s4, x4, y5, z6,
    x5, y4, z7, x6, y7, z4, x7, y6, z5, e5, f6, g7, h8, d5, f7, g6, d6, e7,
    f4, g5, d7, e6, f5, g4, a5, b6, c7, b7, c6, a7, c5, a6, b5, l4, m5, n6,
    o7, a8, l5, m4, n7, o6, b8, l6, m7, n4, o5, c8, l7, m6, n5, o4, d8, h4,
    i5, j6, k7, e8, h5, i4, j7, k6, f8, h6, i7, j4, k5, g8, h7, i6, j5, k4;
  wire new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n342, new_n343, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378, new_n379, new_n380, new_n381, new_n382, new_n383, new_n384,
    new_n385, new_n386, new_n387, new_n388, new_n389, new_n390, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414, new_n415, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1076, new_n1077, new_n1079, new_n1080,
    new_n1081, new_n1083, new_n1085, new_n1086, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1122, new_n1123, new_n1125, new_n1126, new_n1127, new_n1129,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1202,
    new_n1204, new_n1205, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1237, new_n1238, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1260, new_n1261, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1327,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1346;
  assign new_n243 = d & f;
  assign new_n244 = e & new_n243;
  assign new_n245 = a & new_n244;
  assign new_n246 = a & ~s1;
  assign new_n247 = a & ~n;
  assign new_n248 = a & r1;
  assign new_n249 = ~new_n245 & ~new_n246;
  assign new_n250 = ~new_n247 & ~new_n248;
  assign new_n251 = new_n249 & new_n250;
  assign new_n252 = o2 & ~new_n251;
  assign new_n253 = n2 & ~new_n251;
  assign new_n254 = ~new_n252 & ~new_n253;
  assign new_n255 = z1 & o2;
  assign new_n256 = r1 & new_n255;
  assign new_n257 = ~s1 & new_n256;
  assign new_n258 = ~p1 & new_n257;
  assign new_n259 = h2 & new_n258;
  assign new_n260 = ~g2 & ~h2;
  assign new_n261 = f2 & new_n260;
  assign new_n262 = ~g2 & h2;
  assign new_n263 = ~f2 & new_n262;
  assign new_n264 = ~new_n261 & ~new_n263;
  assign new_n265 = o2 & l2;
  assign new_n266 = ~r1 & new_n265;
  assign new_n267 = s1 & new_n266;
  assign new_n268 = ~p1 & new_n267;
  assign new_n269 = ~new_n264 & new_n268;
  assign new_n270 = f2 & new_n269;
  assign new_n271 = f2 & new_n258;
  assign new_n272 = ~r1 & new_n255;
  assign new_n273 = s1 & new_n272;
  assign new_n274 = ~p1 & new_n273;
  assign new_n275 = h2 & new_n274;
  assign new_n276 = f2 & new_n274;
  assign new_n277 = r1 & new_n265;
  assign new_n278 = ~s1 & new_n277;
  assign new_n279 = ~p1 & new_n278;
  assign new_n280 = ~new_n264 & new_n279;
  assign new_n281 = h2 & new_n280;
  assign new_n282 = f2 & new_n280;
  assign new_n283 = h2 & new_n269;
  assign new_n284 = ~new_n259 & ~new_n270;
  assign new_n285 = ~new_n271 & ~new_n275;
  assign new_n286 = new_n284 & new_n285;
  assign new_n287 = ~new_n282 & ~new_n283;
  assign new_n288 = ~new_n276 & ~new_n281;
  assign new_n289 = new_n287 & new_n288;
  assign new_n290 = new_n286 & new_n289;
  assign new_n291 = s0 & u2;
  assign new_n292 = u & new_n291;
  assign new_n293 = ~s0 & u2;
  assign new_n294 = h0 & new_n293;
  assign new_n295 = y1 & x1;
  assign new_n296 = m2 & new_n295;
  assign new_n297 = x2 & ~new_n296;
  assign new_n298 = u3 & ~i;
  assign new_n299 = u3 & new_n291;
  assign new_n300 = ~u & new_n299;
  assign new_n301 = ~h & new_n300;
  assign new_n302 = ~j & d0;
  assign new_n303 = ~l & ~d0;
  assign new_n304 = x2 & ~h0;
  assign new_n305 = ~d0 & new_n304;
  assign new_n306 = ~w2 & new_n305;
  assign new_n307 = ~m & new_n306;
  assign new_n308 = u2 & new_n307;
  assign new_n309 = ~s0 & new_n308;
  assign new_n310 = x2 & ~u;
  assign new_n311 = ~d0 & new_n310;
  assign new_n312 = ~w2 & new_n311;
  assign new_n313 = ~m & new_n312;
  assign new_n314 = u2 & new_n313;
  assign new_n315 = s0 & new_n314;
  assign new_n316 = d0 & new_n304;
  assign new_n317 = ~w2 & new_n316;
  assign new_n318 = ~k & new_n317;
  assign new_n319 = u2 & new_n318;
  assign new_n320 = ~s0 & new_n319;
  assign new_n321 = u3 & new_n293;
  assign new_n322 = ~h0 & new_n321;
  assign new_n323 = ~h & new_n322;
  assign new_n324 = d0 & new_n310;
  assign new_n325 = ~w2 & new_n324;
  assign new_n326 = ~k & new_n325;
  assign new_n327 = u2 & new_n326;
  assign new_n328 = s0 & new_n327;
  assign new_n329 = g & ~new_n303;
  assign new_n330 = ~new_n298 & ~new_n301;
  assign new_n331 = ~new_n302 & new_n330;
  assign new_n332 = new_n329 & new_n331;
  assign new_n333 = ~new_n323 & ~new_n328;
  assign new_n334 = ~new_n309 & ~new_n315;
  assign new_n335 = ~new_n320 & new_n334;
  assign new_n336 = new_n333 & new_n335;
  assign new_n337 = new_n332 & new_n336;
  assign new_n338 = w2 & new_n337;
  assign new_n339 = w2 & ~x2;
  assign new_n340 = ~new_n297 & ~new_n338;
  assign d8 = new_n339 | ~new_n340;
  assign new_n342 = c2 & d8;
  assign new_n343 = ~new_n292 & ~new_n294;
  assign j4 = new_n342 | ~new_n343;
  assign new_n345 = ~new_n290 & ~j4;
  assign new_n346 = a & f0;
  assign new_n347 = ~new_n345 & ~new_n346;
  assign new_n348 = r2 & new_n347;
  assign new_n349 = s0 & ~b2;
  assign new_n350 = s0 & d8;
  assign new_n351 = s1 & s0;
  assign new_n352 = ~new_n349 & ~new_n350;
  assign new_n353 = ~new_n351 & new_n352;
  assign new_n354 = ~z3 & ~new_n353;
  assign new_n355 = ~d8 & new_n354;
  assign new_n356 = u2 & new_n355;
  assign new_n357 = n1 & d8;
  assign new_n358 = ~s1 & n1;
  assign new_n359 = ~b2 & n1;
  assign new_n360 = r1 & n1;
  assign new_n361 = ~new_n357 & ~new_n358;
  assign new_n362 = ~new_n359 & ~new_n360;
  assign new_n363 = new_n361 & new_n362;
  assign new_n364 = ~z3 & ~new_n363;
  assign new_n365 = ~d8 & new_n364;
  assign new_n366 = v2 & new_n365;
  assign new_n367 = new_n296 & new_n337;
  assign new_n368 = w2 & new_n367;
  assign new_n369 = ~z3 & ~y3;
  assign new_n370 = ~d8 & new_n369;
  assign new_n371 = v2 & new_n370;
  assign new_n372 = ~s & ~l3;
  assign new_n373 = ~d8 & new_n372;
  assign new_n374 = ~z3 & new_n373;
  assign new_n375 = u2 & new_n374;
  assign new_n376 = b2 & ~d8;
  assign new_n377 = v1 & new_n376;
  assign new_n378 = i3 & ~new_n377;
  assign new_n379 = m3 & new_n378;
  assign new_n380 = ~h3 & new_n379;
  assign new_n381 = f3 & ~new_n377;
  assign new_n382 = ~new_n380 & ~new_n381;
  assign new_n383 = ~i3 & ~new_n377;
  assign new_n384 = m3 & new_n383;
  assign new_n385 = h3 & new_n384;
  assign new_n386 = e3 & ~new_n377;
  assign new_n387 = ~new_n385 & ~new_n386;
  assign new_n388 = new_n382 & new_n387;
  assign new_n389 = r1 & ~new_n290;
  assign new_n390 = ~new_n377 & ~new_n388;
  assign new_n391 = ~new_n389 & new_n390;
  assign new_n392 = g3 & new_n391;
  assign new_n393 = ~new_n388 & new_n392;
  assign new_n394 = ~d8 & new_n393;
  assign new_n395 = ~new_n389 & new_n394;
  assign new_n396 = y2 & new_n395;
  assign new_n397 = ~z3 & new_n396;
  assign new_n398 = ~new_n356 & ~new_n366;
  assign new_n399 = ~new_n368 & ~new_n371;
  assign new_n400 = new_n398 & new_n399;
  assign new_n401 = ~new_n339 & ~new_n375;
  assign new_n402 = ~new_n397 & new_n401;
  assign new_n403 = new_n400 & new_n402;
  assign new_n404 = ~new_n348 & ~new_n403;
  assign new_n405 = ~n2 & ~new_n254;
  assign new_n406 = ~new_n404 & new_n405;
  assign new_n407 = n2 & new_n254;
  assign new_n408 = ~new_n404 & new_n407;
  assign new_n409 = s0 & u;
  assign new_n410 = u2 & new_n409;
  assign new_n411 = ~t & new_n410;
  assign new_n412 = ~s0 & h0;
  assign new_n413 = u2 & new_n412;
  assign new_n414 = ~g0 & new_n413;
  assign new_n415 = ~new_n411 & ~new_n414;
  assign i4 = d8 | ~new_n415;
  assign h4 = v2 | d8;
  assign new_n418 = i4 & ~h4;
  assign new_n419 = new_n404 & new_n418;
  assign new_n420 = y2 & ~new_n388;
  assign new_n421 = new_n404 & new_n420;
  assign new_n422 = ~i4 & h4;
  assign new_n423 = new_n404 & new_n422;
  assign new_n424 = s0 & v;
  assign new_n425 = ~i4 & new_n424;
  assign new_n426 = new_n404 & new_n425;
  assign new_n427 = ~s0 & i0;
  assign new_n428 = ~i4 & new_n427;
  assign new_n429 = new_n404 & new_n428;
  assign new_n430 = ~new_n406 & ~new_n408;
  assign new_n431 = ~new_n419 & ~new_n421;
  assign new_n432 = new_n430 & new_n431;
  assign new_n433 = ~new_n423 & ~new_n426;
  assign new_n434 = ~new_n429 & new_n433;
  assign t4 = ~new_n432 | ~new_n434;
  assign new_n436 = l2 & ~new_n264;
  assign new_n437 = u2 & ~new_n348;
  assign new_n438 = l0 & new_n437;
  assign new_n439 = ~s0 & l0;
  assign new_n440 = ~t3 & ~o3;
  assign new_n441 = ~n3 & new_n440;
  assign new_n442 = a2 & ~new_n441;
  assign new_n443 = l0 & ~new_n442;
  assign new_n444 = ~z1 & ~new_n443;
  assign new_n445 = ~new_n436 & ~new_n438;
  assign new_n446 = ~new_n439 & new_n445;
  assign u5 = ~new_n444 | ~new_n446;
  assign v6 = ~y0 & ~z0;
  assign new_n449 = ~z2 & ~a3;
  assign new_n450 = k0 & ~new_n449;
  assign new_n451 = k0 & ~new_n442;
  assign new_n452 = h0 & k0;
  assign new_n453 = ~new_n450 & ~new_n451;
  assign new_n454 = ~l2 & ~new_n452;
  assign t5 = ~new_n453 | ~new_n454;
  assign new_n456 = o2 & new_n254;
  assign new_n457 = ~new_n404 & new_n456;
  assign new_n458 = y2 & ~new_n382;
  assign new_n459 = ~new_n387 & new_n458;
  assign new_n460 = new_n404 & new_n459;
  assign new_n461 = n2 & o2;
  assign new_n462 = ~new_n404 & new_n461;
  assign new_n463 = ~o2 & new_n405;
  assign new_n464 = ~new_n404 & new_n463;
  assign new_n465 = ~new_n457 & ~new_n460;
  assign new_n466 = ~new_n419 & new_n465;
  assign new_n467 = ~new_n423 & ~new_n462;
  assign new_n468 = ~new_n464 & new_n467;
  assign u4 = ~new_n466 | ~new_n468;
  assign new_n470 = ~p & ~q;
  assign new_n471 = o & new_n470;
  assign new_n472 = l2 & new_n471;
  assign new_n473 = ~k2 & new_n472;
  assign new_n474 = ~x0 & ~z0;
  assign new_n475 = y0 & new_n474;
  assign new_n476 = ~w0 & new_n475;
  assign new_n477 = x0 & ~z0;
  assign new_n478 = ~y0 & new_n477;
  assign new_n479 = ~w0 & new_n478;
  assign new_n480 = w0 & z0;
  assign new_n481 = ~new_n476 & ~new_n479;
  assign new_n482 = ~new_n480 & new_n481;
  assign new_n483 = u1 & ~z0;
  assign new_n484 = ~x0 & new_n483;
  assign new_n485 = ~y0 & new_n484;
  assign new_n486 = ~w0 & new_n485;
  assign new_n487 = u1 & z0;
  assign new_n488 = x0 & new_n487;
  assign new_n489 = ~y0 & new_n488;
  assign new_n490 = ~w0 & new_n489;
  assign new_n491 = y0 & new_n484;
  assign new_n492 = w0 & new_n491;
  assign new_n493 = y0 & new_n488;
  assign new_n494 = w0 & new_n493;
  assign new_n495 = ~new_n486 & ~new_n490;
  assign new_n496 = ~new_n492 & ~new_n494;
  assign new_n497 = new_n495 & new_n496;
  assign new_n498 = new_n482 & new_n497;
  assign new_n499 = j2 & new_n498;
  assign t6 = new_n473 | new_n499;
  assign new_n501 = n2 & new_n347;
  assign new_n502 = ~new_n403 & new_n501;
  assign new_n503 = o2 & new_n347;
  assign new_n504 = r2 & new_n503;
  assign new_n505 = new_n347 & ~new_n403;
  assign new_n506 = new_n251 & new_n505;
  assign new_n507 = r2 & new_n501;
  assign new_n508 = new_n251 & new_n347;
  assign new_n509 = r2 & new_n508;
  assign new_n510 = ~new_n403 & new_n503;
  assign new_n511 = ~new_n502 & ~new_n504;
  assign new_n512 = ~new_n506 & new_n511;
  assign new_n513 = ~new_n507 & ~new_n509;
  assign new_n514 = ~new_n510 & new_n513;
  assign v4 = ~new_n512 | ~new_n514;
  assign new_n516 = j2 & ~new_n497;
  assign new_n517 = j2 & ~new_n482;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = l0 & new_n518;
  assign new_n520 = m0 & new_n519;
  assign new_n521 = k0 & new_n520;
  assign new_n522 = t0 & n3;
  assign new_n523 = ~h0 & new_n522;
  assign new_n524 = new_n521 & ~new_n523;
  assign new_n525 = new_n442 & new_n524;
  assign new_n526 = j0 & new_n521;
  assign new_n527 = ~new_n525 & ~new_n526;
  assign w5 = n3 & ~new_n527;
  assign new_n529 = t0 & new_n497;
  assign u6 = g0 & new_n529;
  assign new_n531 = h0 & ~l3;
  assign new_n532 = t0 & new_n531;
  assign new_n533 = ~g0 & new_n532;
  assign new_n534 = ~q & l2;
  assign new_n535 = ~o & new_n534;
  assign new_n536 = p & new_n535;
  assign new_n537 = ~new_n533 & new_n536;
  assign new_n538 = h3 & new_n537;
  assign new_n539 = ~i3 & new_n537;
  assign new_n540 = ~y1 & m2;
  assign new_n541 = ~w1 & new_n540;
  assign new_n542 = x1 & new_n541;
  assign new_n543 = ~new_n533 & new_n542;
  assign new_n544 = p2 & l2;
  assign new_n545 = p & new_n544;
  assign new_n546 = ~q & new_n545;
  assign new_n547 = ~new_n533 & new_n546;
  assign new_n548 = m0 & ~new_n533;
  assign new_n549 = ~new_n547 & ~new_n548;
  assign new_n550 = ~new_n538 & ~new_n539;
  assign new_n551 = ~new_n543 & new_n550;
  assign v5 = ~new_n549 | ~new_n551;
  assign new_n553 = ~b & ~new_n251;
  assign new_n554 = ~new_n404 & new_n553;
  assign new_n555 = b & new_n251;
  assign new_n556 = ~new_n404 & new_n555;
  assign new_n557 = d2 & new_n404;
  assign new_n558 = ~new_n554 & ~new_n556;
  assign w4 = new_n557 | ~new_n558;
  assign new_n560 = z1 & ~f2;
  assign new_n561 = ~t2 & new_n560;
  assign new_n562 = new_n348 & new_n561;
  assign new_n563 = ~a & new_n562;
  assign new_n564 = z1 & ~g2;
  assign new_n565 = t1 & new_n564;
  assign new_n566 = ~new_n403 & new_n565;
  assign new_n567 = ~a & new_n566;
  assign new_n568 = ~new_n403 & new_n561;
  assign new_n569 = ~a & new_n568;
  assign new_n570 = t1 & new_n560;
  assign new_n571 = new_n348 & new_n570;
  assign new_n572 = ~a & new_n571;
  assign new_n573 = ~new_n403 & new_n570;
  assign new_n574 = ~a & new_n573;
  assign new_n575 = ~t2 & new_n260;
  assign new_n576 = new_n348 & new_n575;
  assign new_n577 = ~a & new_n576;
  assign new_n578 = l2 & new_n577;
  assign new_n579 = z1 & ~l2;
  assign new_n580 = t1 & new_n579;
  assign new_n581 = ~new_n403 & new_n580;
  assign new_n582 = ~a & new_n581;
  assign new_n583 = t1 & new_n260;
  assign new_n584 = new_n348 & new_n583;
  assign new_n585 = ~a & new_n584;
  assign new_n586 = l2 & new_n585;
  assign new_n587 = ~t2 & new_n579;
  assign new_n588 = ~new_n403 & new_n587;
  assign new_n589 = ~a & new_n588;
  assign new_n590 = new_n348 & new_n580;
  assign new_n591 = ~a & new_n590;
  assign new_n592 = new_n348 & new_n587;
  assign new_n593 = ~a & new_n592;
  assign new_n594 = ~f2 & ~g2;
  assign new_n595 = ~t2 & new_n594;
  assign new_n596 = new_n348 & new_n595;
  assign new_n597 = ~a & new_n596;
  assign new_n598 = l2 & new_n597;
  assign new_n599 = ~f2 & ~h2;
  assign new_n600 = t1 & new_n599;
  assign new_n601 = ~new_n403 & new_n600;
  assign new_n602 = ~a & new_n601;
  assign new_n603 = t1 & new_n594;
  assign new_n604 = new_n348 & new_n603;
  assign new_n605 = ~a & new_n604;
  assign new_n606 = l2 & new_n605;
  assign new_n607 = ~t2 & new_n599;
  assign new_n608 = ~new_n403 & new_n607;
  assign new_n609 = ~a & new_n608;
  assign new_n610 = ~new_n403 & new_n575;
  assign new_n611 = ~a & new_n610;
  assign new_n612 = l2 & new_n611;
  assign new_n613 = new_n348 & new_n600;
  assign new_n614 = ~a & new_n613;
  assign new_n615 = ~new_n403 & new_n583;
  assign new_n616 = ~a & new_n615;
  assign new_n617 = l2 & new_n616;
  assign new_n618 = new_n348 & new_n607;
  assign new_n619 = ~a & new_n618;
  assign new_n620 = ~new_n403 & new_n595;
  assign new_n621 = ~a & new_n620;
  assign new_n622 = l2 & new_n621;
  assign new_n623 = z1 & ~h2;
  assign new_n624 = t1 & new_n623;
  assign new_n625 = new_n348 & new_n624;
  assign new_n626 = ~a & new_n625;
  assign new_n627 = ~new_n403 & new_n603;
  assign new_n628 = ~a & new_n627;
  assign new_n629 = l2 & new_n628;
  assign new_n630 = ~t2 & new_n623;
  assign new_n631 = new_n348 & new_n630;
  assign new_n632 = ~a & new_n631;
  assign new_n633 = ~new_n403 & new_n630;
  assign new_n634 = ~a & new_n633;
  assign new_n635 = ~t2 & new_n564;
  assign new_n636 = new_n348 & new_n635;
  assign new_n637 = ~a & new_n636;
  assign new_n638 = ~new_n403 & new_n624;
  assign new_n639 = ~a & new_n638;
  assign new_n640 = ~new_n403 & new_n635;
  assign new_n641 = ~a & new_n640;
  assign new_n642 = new_n348 & new_n565;
  assign new_n643 = ~a & new_n642;
  assign new_n644 = ~new_n639 & ~new_n641;
  assign new_n645 = ~new_n643 & new_n644;
  assign new_n646 = ~new_n629 & ~new_n632;
  assign new_n647 = ~new_n634 & ~new_n637;
  assign new_n648 = new_n646 & new_n647;
  assign new_n649 = new_n645 & new_n648;
  assign new_n650 = ~new_n619 & ~new_n622;
  assign new_n651 = ~new_n626 & new_n650;
  assign new_n652 = ~new_n614 & ~new_n617;
  assign new_n653 = ~new_n609 & ~new_n612;
  assign new_n654 = new_n652 & new_n653;
  assign new_n655 = new_n651 & new_n654;
  assign new_n656 = new_n649 & new_n655;
  assign new_n657 = ~new_n598 & ~new_n602;
  assign new_n658 = ~new_n606 & new_n657;
  assign new_n659 = ~new_n586 & ~new_n589;
  assign new_n660 = ~new_n591 & ~new_n593;
  assign new_n661 = new_n659 & new_n660;
  assign new_n662 = new_n658 & new_n661;
  assign new_n663 = ~new_n563 & ~new_n567;
  assign new_n664 = ~new_n569 & ~new_n572;
  assign new_n665 = new_n663 & new_n664;
  assign new_n666 = ~new_n574 & ~new_n578;
  assign new_n667 = ~new_n582 & new_n666;
  assign new_n668 = new_n665 & new_n667;
  assign new_n669 = new_n662 & new_n668;
  assign p4 = ~new_n656 | ~new_n669;
  assign new_n671 = new_n442 & ~new_n521;
  assign new_n672 = j0 & new_n523;
  assign new_n673 = ~i3 & h3;
  assign new_n674 = i3 & ~h3;
  assign new_n675 = ~new_n673 & ~new_n674;
  assign new_n676 = l2 & o0;
  assign new_n677 = d3 & new_n676;
  assign new_n678 = new_n449 & new_n677;
  assign new_n679 = z2 & new_n678;
  assign new_n680 = ~a3 & new_n678;
  assign new_n681 = ~d3 & new_n449;
  assign new_n682 = ~b3 & new_n681;
  assign new_n683 = ~c3 & new_n682;
  assign new_n684 = ~a3 & new_n683;
  assign new_n685 = ~new_n389 & new_n449;
  assign new_n686 = ~c3 & new_n685;
  assign new_n687 = ~d3 & new_n686;
  assign new_n688 = ~b3 & new_n687;
  assign new_n689 = z2 & new_n683;
  assign new_n690 = o0 & new_n449;
  assign new_n691 = b3 & new_n690;
  assign new_n692 = ~c3 & new_n691;
  assign new_n693 = ~a3 & new_n692;
  assign new_n694 = l2 & new_n693;
  assign new_n695 = ~c3 & new_n690;
  assign new_n696 = ~new_n389 & new_n695;
  assign new_n697 = b3 & new_n696;
  assign new_n698 = l2 & new_n697;
  assign new_n699 = ~new_n389 & new_n676;
  assign new_n700 = new_n449 & new_n699;
  assign new_n701 = d3 & new_n700;
  assign new_n702 = z2 & new_n692;
  assign new_n703 = l2 & new_n702;
  assign new_n704 = ~new_n688 & ~new_n689;
  assign new_n705 = ~new_n679 & ~new_n680;
  assign new_n706 = ~new_n684 & new_n705;
  assign new_n707 = new_n704 & new_n706;
  assign new_n708 = ~new_n701 & ~new_n703;
  assign new_n709 = ~new_n694 & ~new_n698;
  assign new_n710 = new_n708 & new_n709;
  assign new_n711 = new_n707 & new_n710;
  assign new_n712 = new_n685 & new_n711;
  assign new_n713 = m3 & new_n712;
  assign new_n714 = i3 & new_n449;
  assign new_n715 = new_n711 & new_n714;
  assign new_n716 = h3 & new_n715;
  assign new_n717 = ~new_n713 & ~new_n716;
  assign new_n718 = ~new_n675 & new_n717;
  assign new_n719 = t0 & ~new_n497;
  assign new_n720 = ~l2 & new_n719;
  assign new_n721 = g0 & new_n720;
  assign new_n722 = new_n442 & new_n721;
  assign new_n723 = ~new_n471 & ~new_n518;
  assign new_n724 = new_n482 & ~new_n518;
  assign new_n725 = ~l2 & ~new_n518;
  assign new_n726 = new_n348 & new_n442;
  assign new_n727 = t0 & new_n726;
  assign new_n728 = ~l3 & new_n727;
  assign new_n729 = t0 & new_n449;
  assign new_n730 = ~l3 & new_n729;
  assign new_n731 = new_n442 & new_n730;
  assign new_n732 = ~h0 & new_n731;
  assign new_n733 = ~u2 & new_n442;
  assign new_n734 = t0 & new_n733;
  assign new_n735 = ~l3 & new_n734;
  assign new_n736 = ~s0 & d8;
  assign new_n737 = ~h0 & new_n736;
  assign new_n738 = ~s0 & z3;
  assign new_n739 = ~h0 & new_n738;
  assign new_n740 = ~u & new_n350;
  assign new_n741 = s0 & z3;
  assign new_n742 = ~u & new_n741;
  assign new_n743 = ~new_n739 & ~new_n740;
  assign new_n744 = ~new_n742 & new_n743;
  assign new_n745 = ~new_n732 & ~new_n735;
  assign new_n746 = ~new_n737 & new_n745;
  assign new_n747 = new_n744 & new_n746;
  assign new_n748 = ~new_n718 & ~new_n722;
  assign new_n749 = ~new_n723 & new_n748;
  assign new_n750 = ~new_n724 & ~new_n725;
  assign new_n751 = ~new_n728 & new_n750;
  assign new_n752 = new_n749 & new_n751;
  assign new_n753 = new_n747 & new_n752;
  assign new_n754 = new_n442 & ~new_n753;
  assign new_n755 = j0 & ~new_n521;
  assign new_n756 = j0 & ~new_n753;
  assign new_n757 = new_n442 & new_n523;
  assign new_n758 = ~new_n671 & ~new_n672;
  assign new_n759 = ~new_n754 & new_n758;
  assign new_n760 = ~new_n755 & ~new_n756;
  assign new_n761 = ~new_n757 & new_n760;
  assign q5 = ~new_n759 | ~new_n761;
  assign new_n763 = c3 & o0;
  assign new_n764 = b3 & o0;
  assign new_n765 = ~new_n763 & ~new_n764;
  assign new_n766 = c3 & new_n711;
  assign new_n767 = new_n765 & new_n766;
  assign new_n768 = b3 & new_n767;
  assign new_n769 = ~new_n389 & new_n765;
  assign new_n770 = new_n711 & new_n769;
  assign new_n771 = c3 & new_n770;
  assign new_n772 = a3 & ~new_n711;
  assign new_n773 = ~new_n768 & ~new_n771;
  assign r6 = new_n772 | ~new_n773;
  assign new_n775 = g2 & ~h2;
  assign new_n776 = g2 & l2;
  assign new_n777 = f2 & ~h2;
  assign new_n778 = f2 & l2;
  assign new_n779 = ~h2 & ~l2;
  assign new_n780 = ~new_n778 & ~new_n779;
  assign new_n781 = ~new_n775 & ~new_n776;
  assign new_n782 = ~new_n777 & new_n781;
  assign p5 = ~new_n780 | ~new_n782;
  assign new_n784 = ~a & new_n599;
  assign new_n785 = ~t1 & new_n784;
  assign new_n786 = t2 & new_n785;
  assign new_n787 = t2 & a1;
  assign q4 = new_n786 | new_n787;
  assign new_n789 = new_n296 & ~new_n337;
  assign new_n790 = s1 & new_n789;
  assign new_n791 = ~r1 & new_n790;
  assign new_n792 = s1 & d4;
  assign new_n793 = ~r1 & new_n792;
  assign new_n794 = s1 & d8;
  assign new_n795 = ~r1 & new_n794;
  assign new_n796 = ~new_n791 & ~new_n793;
  assign r7 = new_n795 | ~new_n796;
  assign new_n798 = ~o0 & new_n711;
  assign new_n799 = d3 & new_n798;
  assign new_n800 = c3 & ~new_n765;
  assign s6 = new_n799 | new_n800;
  assign new_n802 = i3 & ~new_n449;
  assign new_n803 = h3 & new_n802;
  assign new_n804 = ~new_n389 & ~new_n711;
  assign new_n805 = ~new_n675 & new_n804;
  assign new_n806 = m3 & new_n805;
  assign new_n807 = new_n711 & new_n729;
  assign new_n808 = ~h0 & new_n807;
  assign new_n809 = ~new_n449 & new_n808;
  assign new_n810 = i3 & ~new_n711;
  assign new_n811 = h3 & new_n810;
  assign new_n812 = ~new_n711 & new_n808;
  assign new_n813 = ~new_n389 & ~new_n449;
  assign new_n814 = ~new_n675 & new_n813;
  assign new_n815 = m3 & new_n814;
  assign new_n816 = ~new_n803 & ~new_n806;
  assign new_n817 = ~new_n809 & new_n816;
  assign new_n818 = ~new_n811 & ~new_n812;
  assign new_n819 = ~new_n815 & new_n818;
  assign new_n820 = new_n817 & new_n819;
  assign new_n821 = a3 & new_n711;
  assign new_n822 = new_n820 & new_n821;
  assign new_n823 = z2 & new_n822;
  assign new_n824 = new_n711 & new_n820;
  assign new_n825 = ~new_n389 & new_n824;
  assign new_n826 = a3 & new_n825;
  assign new_n827 = new_n424 & ~new_n820;
  assign new_n828 = ~u & new_n827;
  assign new_n829 = new_n427 & ~new_n820;
  assign new_n830 = ~h0 & new_n829;
  assign new_n831 = ~new_n675 & ~new_n820;
  assign new_n832 = ~s0 & new_n711;
  assign new_n833 = a3 & new_n832;
  assign new_n834 = ~new_n389 & new_n833;
  assign new_n835 = h0 & new_n834;
  assign new_n836 = s0 & new_n711;
  assign new_n837 = a3 & new_n836;
  assign new_n838 = ~new_n389 & new_n837;
  assign new_n839 = u & new_n838;
  assign new_n840 = z2 & new_n832;
  assign new_n841 = a3 & new_n840;
  assign new_n842 = h0 & new_n841;
  assign new_n843 = z2 & new_n836;
  assign new_n844 = a3 & new_n843;
  assign new_n845 = u & new_n844;
  assign new_n846 = ~s0 & ~new_n820;
  assign new_n847 = z2 & new_n846;
  assign new_n848 = a3 & new_n847;
  assign new_n849 = h0 & new_n848;
  assign new_n850 = ~s0 & ~new_n389;
  assign new_n851 = a3 & new_n850;
  assign new_n852 = ~new_n820 & new_n851;
  assign new_n853 = h0 & new_n852;
  assign new_n854 = s0 & ~new_n820;
  assign new_n855 = z2 & new_n854;
  assign new_n856 = a3 & new_n855;
  assign new_n857 = u & new_n856;
  assign new_n858 = s0 & ~new_n389;
  assign new_n859 = a3 & new_n858;
  assign new_n860 = ~new_n820 & new_n859;
  assign new_n861 = u & new_n860;
  assign new_n862 = ~new_n823 & ~new_n826;
  assign new_n863 = ~new_n828 & ~new_n830;
  assign new_n864 = new_n862 & new_n863;
  assign new_n865 = ~new_n831 & ~new_n835;
  assign new_n866 = ~new_n839 & new_n865;
  assign new_n867 = new_n864 & new_n866;
  assign new_n868 = ~new_n853 & ~new_n857;
  assign new_n869 = ~new_n861 & new_n868;
  assign new_n870 = ~new_n842 & ~new_n845;
  assign new_n871 = ~new_n849 & new_n870;
  assign new_n872 = new_n869 & new_n871;
  assign p6 = ~new_n867 | ~new_n872;
  assign new_n874 = ~s1 & new_n789;
  assign new_n875 = ~s1 & d4;
  assign new_n876 = ~s1 & d8;
  assign new_n877 = ~new_n874 & ~new_n875;
  assign q7 = new_n876 | ~new_n877;
  assign new_n879 = ~g1 & ~h1;
  assign new_n880 = o0 & new_n879;
  assign new_n881 = ~f1 & new_n880;
  assign new_n882 = a & new_n881;
  assign new_n883 = g2 & new_n882;
  assign new_n884 = new_n264 & new_n881;
  assign new_n885 = g2 & new_n884;
  assign new_n886 = h2 & new_n470;
  assign new_n887 = ~o & new_n886;
  assign new_n888 = ~l2 & new_n887;
  assign new_n889 = ~q1 & ~r1;
  assign new_n890 = ~l2 & new_n889;
  assign new_n891 = ~h2 & new_n890;
  assign new_n892 = a & new_n891;
  assign new_n893 = ~s1 & new_n892;
  assign new_n894 = ~l2 & o0;
  assign new_n895 = ~s1 & ~r1;
  assign new_n896 = h2 & new_n895;
  assign new_n897 = ~q1 & new_n896;
  assign new_n898 = new_n264 & new_n897;
  assign new_n899 = ~p & new_n898;
  assign new_n900 = ~q & new_n899;
  assign new_n901 = ~g2 & new_n900;
  assign new_n902 = ~o & new_n901;
  assign new_n903 = h2 & new_n879;
  assign new_n904 = ~f1 & new_n903;
  assign new_n905 = new_n264 & new_n904;
  assign new_n906 = ~p & new_n905;
  assign new_n907 = ~q & new_n906;
  assign new_n908 = g2 & new_n907;
  assign new_n909 = ~o & new_n908;
  assign new_n910 = a & new_n897;
  assign new_n911 = ~p & new_n910;
  assign new_n912 = ~q & new_n911;
  assign new_n913 = ~g2 & new_n912;
  assign new_n914 = ~o & new_n913;
  assign new_n915 = a & new_n904;
  assign new_n916 = ~p & new_n915;
  assign new_n917 = ~q & new_n916;
  assign new_n918 = g2 & new_n917;
  assign new_n919 = ~o & new_n918;
  assign new_n920 = ~h2 & new_n895;
  assign new_n921 = ~q1 & new_n920;
  assign new_n922 = a & new_n921;
  assign new_n923 = ~g2 & new_n922;
  assign new_n924 = ~h2 & new_n879;
  assign new_n925 = ~f1 & new_n924;
  assign new_n926 = a & new_n925;
  assign new_n927 = ~s1 & new_n926;
  assign new_n928 = g2 & new_n927;
  assign new_n929 = ~q1 & new_n928;
  assign new_n930 = ~r1 & new_n929;
  assign new_n931 = o0 & new_n895;
  assign new_n932 = ~q1 & new_n931;
  assign new_n933 = a & new_n932;
  assign new_n934 = ~g2 & new_n933;
  assign new_n935 = new_n264 & new_n932;
  assign new_n936 = ~g2 & new_n935;
  assign new_n937 = ~new_n883 & ~new_n885;
  assign new_n938 = ~new_n888 & ~new_n893;
  assign new_n939 = new_n937 & new_n938;
  assign new_n940 = ~new_n894 & ~new_n902;
  assign new_n941 = ~new_n909 & new_n940;
  assign new_n942 = new_n939 & new_n941;
  assign new_n943 = ~new_n930 & ~new_n934;
  assign new_n944 = ~new_n936 & new_n943;
  assign new_n945 = ~new_n914 & ~new_n919;
  assign new_n946 = ~new_n923 & new_n945;
  assign new_n947 = new_n944 & new_n946;
  assign r4 = ~new_n942 | ~new_n947;
  assign new_n949 = ~o3 & new_n442;
  assign s5 = new_n499 | new_n949;
  assign new_n951 = a4 & ~d8;
  assign new_n952 = ~new_n348 & new_n951;
  assign new_n953 = ~new_n363 & new_n952;
  assign new_n954 = a4 & new_n392;
  assign new_n955 = ~new_n348 & new_n954;
  assign new_n956 = ~d8 & new_n955;
  assign new_n957 = ~new_n527 & new_n952;
  assign new_n958 = e4 & i1;
  assign new_n959 = new_n952 & new_n958;
  assign new_n960 = ~v2 & new_n951;
  assign new_n961 = ~new_n363 & new_n960;
  assign new_n962 = ~v2 & new_n353;
  assign new_n963 = ~d8 & new_n962;
  assign new_n964 = ~new_n392 & new_n963;
  assign new_n965 = new_n958 & new_n964;
  assign new_n966 = a4 & new_n965;
  assign new_n967 = s & new_n966;
  assign new_n968 = ~new_n527 & new_n964;
  assign new_n969 = a4 & new_n968;
  assign new_n970 = l3 & new_n969;
  assign new_n971 = l3 & new_n966;
  assign new_n972 = y3 & ~new_n392;
  assign new_n973 = new_n363 & new_n972;
  assign new_n974 = ~d8 & new_n973;
  assign new_n975 = ~new_n527 & new_n974;
  assign new_n976 = s & new_n975;
  assign new_n977 = new_n353 & new_n976;
  assign new_n978 = a4 & new_n977;
  assign new_n979 = y3 & new_n388;
  assign new_n980 = ~d8 & new_n979;
  assign new_n981 = new_n392 & new_n980;
  assign new_n982 = new_n363 & new_n981;
  assign new_n983 = a4 & new_n982;
  assign new_n984 = new_n958 & new_n974;
  assign new_n985 = l3 & new_n984;
  assign new_n986 = new_n353 & new_n985;
  assign new_n987 = a4 & new_n986;
  assign new_n988 = ~u2 & ~new_n392;
  assign new_n989 = new_n363 & new_n988;
  assign new_n990 = ~d8 & new_n989;
  assign new_n991 = ~new_n527 & new_n990;
  assign new_n992 = y3 & new_n991;
  assign new_n993 = a4 & new_n992;
  assign new_n994 = new_n958 & new_n990;
  assign new_n995 = y3 & new_n994;
  assign new_n996 = a4 & new_n995;
  assign new_n997 = s & new_n969;
  assign new_n998 = l3 & new_n975;
  assign new_n999 = new_n353 & new_n998;
  assign new_n1000 = a4 & new_n999;
  assign new_n1001 = y3 & ~y2;
  assign new_n1002 = ~d8 & new_n1001;
  assign new_n1003 = new_n392 & new_n1002;
  assign new_n1004 = new_n363 & new_n1003;
  assign new_n1005 = a4 & new_n1004;
  assign new_n1006 = s & new_n984;
  assign new_n1007 = new_n353 & new_n1006;
  assign new_n1008 = a4 & new_n1007;
  assign new_n1009 = y3 & new_n389;
  assign new_n1010 = ~d8 & new_n1009;
  assign new_n1011 = new_n392 & new_n1010;
  assign new_n1012 = new_n363 & new_n1011;
  assign new_n1013 = a4 & new_n1012;
  assign new_n1014 = ~v2 & ~u2;
  assign new_n1015 = ~d8 & new_n1014;
  assign new_n1016 = ~new_n392 & new_n1015;
  assign new_n1017 = new_n958 & new_n1016;
  assign new_n1018 = a4 & new_n1017;
  assign new_n1019 = a4 & new_n388;
  assign new_n1020 = new_n392 & new_n1019;
  assign new_n1021 = ~v2 & new_n1020;
  assign new_n1022 = ~d8 & new_n1021;
  assign new_n1023 = ~new_n527 & new_n1016;
  assign new_n1024 = a4 & new_n1023;
  assign new_n1025 = ~y2 & a4;
  assign new_n1026 = new_n392 & new_n1025;
  assign new_n1027 = ~v2 & new_n1026;
  assign new_n1028 = ~d8 & new_n1027;
  assign new_n1029 = a4 & new_n389;
  assign new_n1030 = new_n392 & new_n1029;
  assign new_n1031 = ~v2 & new_n1030;
  assign new_n1032 = ~d8 & new_n1031;
  assign new_n1033 = ~new_n1028 & ~new_n1032;
  assign new_n1034 = ~new_n1018 & ~new_n1022;
  assign new_n1035 = ~new_n1024 & new_n1034;
  assign new_n1036 = new_n1033 & new_n1035;
  assign new_n1037 = ~new_n1005 & ~new_n1008;
  assign new_n1038 = ~new_n1013 & new_n1037;
  assign new_n1039 = ~new_n996 & ~new_n997;
  assign new_n1040 = ~new_n1000 & new_n1039;
  assign new_n1041 = new_n1038 & new_n1040;
  assign new_n1042 = new_n1036 & new_n1041;
  assign new_n1043 = ~new_n983 & ~new_n987;
  assign new_n1044 = ~new_n993 & new_n1043;
  assign new_n1045 = ~new_n970 & ~new_n971;
  assign new_n1046 = ~new_n978 & new_n1045;
  assign new_n1047 = new_n1044 & new_n1046;
  assign new_n1048 = ~new_n953 & ~new_n956;
  assign new_n1049 = ~new_n957 & new_n1048;
  assign new_n1050 = ~new_n959 & ~new_n961;
  assign new_n1051 = ~new_n967 & new_n1050;
  assign new_n1052 = new_n1049 & new_n1051;
  assign new_n1053 = new_n1047 & new_n1052;
  assign p7 = ~new_n1042 | ~new_n1053;
  assign new_n1055 = new_n711 & new_n765;
  assign new_n1056 = b3 & new_n1055;
  assign new_n1057 = z2 & ~new_n711;
  assign q6 = new_n1056 | new_n1057;
  assign new_n1059 = ~new_n527 & new_n753;
  assign r5 = ~new_n533 & new_n1059;
  assign new_n1061 = ~new_n290 & j4;
  assign new_n1062 = ~a & new_n1061;
  assign new_n1063 = ~a & f0;
  assign s4 = new_n1062 | new_n1063;
  assign new_n1065 = b & ~new_n251;
  assign new_n1066 = ~c & new_n1065;
  assign new_n1067 = ~new_n404 & new_n1066;
  assign new_n1068 = ~b & c;
  assign new_n1069 = ~new_n404 & new_n1068;
  assign new_n1070 = c & new_n251;
  assign new_n1071 = ~new_n404 & new_n1070;
  assign new_n1072 = e2 & new_n404;
  assign new_n1073 = ~new_n1067 & ~new_n1069;
  assign new_n1074 = ~new_n1071 & ~new_n1072;
  assign x4 = ~new_n1073 | ~new_n1074;
  assign new_n1076 = t0 & l3;
  assign new_n1077 = g0 & new_n1076;
  assign y5 = ~new_n518 | new_n1077;
  assign new_n1079 = k2 & ~l2;
  assign new_n1080 = k2 & ~new_n471;
  assign new_n1081 = ~new_n1079 & ~new_n1080;
  assign x5 = new_n721 | ~new_n1081;
  assign new_n1083 = v0 & ~x3;
  assign y4 = a | new_n1083;
  assign new_n1085 = k & ~d0;
  assign new_n1086 = m & d0;
  assign z7 = new_n1085 | new_n1086;
  assign x6 = ~w0 & ~x0;
  assign y7 = p3 & j3;
  assign z4 = v0 & b4;
  assign new_n1091 = r & k3;
  assign new_n1092 = ~p3 & r;
  assign new_n1093 = s2 & u0;
  assign new_n1094 = ~new_n1091 & ~new_n1092;
  assign x7 = new_n1093 | ~new_n1094;
  assign new_n1096 = ~k2 & ~new_n523;
  assign new_n1097 = ~i2 & ~d8;
  assign z5 = ~new_n1096 | ~new_n1097;
  assign new_n1099 = ~e1 & l2;
  assign new_n1100 = ~d1 & new_n1099;
  assign new_n1101 = ~p & q;
  assign new_n1102 = n & new_n1101;
  assign new_n1103 = l2 & ~new_n1102;
  assign e5 = new_n1100 | new_n1103;
  assign new_n1105 = p2 & m2;
  assign new_n1106 = q2 & m2;
  assign new_n1107 = r0 & m2;
  assign new_n1108 = ~new_n1105 & ~new_n1106;
  assign f6 = new_n1107 | ~new_n1108;
  assign new_n1110 = y1 & m2;
  assign new_n1111 = ~x1 & new_n1110;
  assign new_n1112 = ~q2 & new_n1111;
  assign new_n1113 = q2 & ~m2;
  assign new_n1114 = p2 & new_n1113;
  assign new_n1115 = q & new_n1114;
  assign new_n1116 = ~p2 & new_n1111;
  assign new_n1117 = ~new_n1112 & ~new_n1115;
  assign new_n1118 = ~new_n1116 & new_n1117;
  assign new_n1119 = ~k1 & ~new_n1118;
  assign new_n1120 = q3 & new_n1118;
  assign g7 = new_n1119 | new_n1120;
  assign new_n1122 = ~w2 & d8;
  assign new_n1123 = ~w2 & ~x2;
  assign h8 = new_n1122 | new_n1123;
  assign new_n1125 = ~d1 & l2;
  assign new_n1126 = ~e1 & new_n1125;
  assign new_n1127 = ~c1 & new_n1126;
  assign d5 = new_n1103 | new_n1127;
  assign new_n1129 = m1 & m2;
  assign f7 = ~new_n1108 | new_n1129;
  assign new_n1131 = p & new_n1114;
  assign new_n1132 = ~q2 & m2;
  assign new_n1133 = x1 & new_n1132;
  assign new_n1134 = ~y1 & new_n1133;
  assign new_n1135 = r0 & new_n1134;
  assign new_n1136 = ~p2 & m2;
  assign new_n1137 = x1 & new_n1136;
  assign new_n1138 = ~y1 & new_n1137;
  assign new_n1139 = r0 & new_n1138;
  assign new_n1140 = ~new_n1135 & ~new_n1139;
  assign new_n1141 = ~new_n1131 & new_n1140;
  assign new_n1142 = ~p0 & ~new_n1141;
  assign new_n1143 = v3 & new_n1141;
  assign g6 = new_n1142 | new_n1143;
  assign new_n1145 = y3 & l3;
  assign new_n1146 = z3 & new_n1145;
  assign new_n1147 = new_n958 & new_n1146;
  assign new_n1148 = y3 & s;
  assign new_n1149 = z3 & new_n1148;
  assign new_n1150 = new_n958 & new_n1149;
  assign e7 = new_n1147 | new_n1150;
  assign new_n1152 = e0 & y;
  assign new_n1153 = x & ~y;
  assign new_n1154 = j1 & new_n1153;
  assign new_n1155 = e0 & ~x;
  assign new_n1156 = ~new_n1152 & ~new_n1154;
  assign f4 = new_n1155 | ~new_n1156;
  assign g5 = new_n1099 | new_n1103;
  assign new_n1159 = q2 & l2;
  assign new_n1160 = p2 & new_n1159;
  assign new_n1161 = q & new_n1160;
  assign new_n1162 = q2 & ~new_n1161;
  assign new_n1163 = i1 & new_n1162;
  assign new_n1164 = ~s1 & m1;
  assign new_n1165 = ~new_n1161 & new_n1164;
  assign new_n1166 = i1 & new_n1165;
  assign new_n1167 = ~l2 & ~new_n1161;
  assign new_n1168 = i1 & new_n1167;
  assign new_n1169 = p2 & ~new_n1161;
  assign new_n1170 = i1 & new_n1169;
  assign new_n1171 = i1 & ~new_n1161;
  assign new_n1172 = ~q & new_n1171;
  assign new_n1173 = ~y3 & o1;
  assign new_n1174 = ~new_n1161 & new_n1173;
  assign new_n1175 = ~s1 & new_n1174;
  assign new_n1176 = m1 & new_n1175;
  assign new_n1177 = new_n290 & new_n1174;
  assign new_n1178 = m1 & new_n1177;
  assign new_n1179 = ~y3 & ~new_n1161;
  assign new_n1180 = o1 & new_n1179;
  assign new_n1181 = q2 & new_n1180;
  assign new_n1182 = ~l2 & new_n1180;
  assign new_n1183 = p2 & new_n1180;
  assign new_n1184 = m1 & new_n290;
  assign new_n1185 = ~new_n1161 & new_n1184;
  assign new_n1186 = i1 & new_n1185;
  assign new_n1187 = ~q & new_n1180;
  assign new_n1188 = ~new_n1183 & ~new_n1186;
  assign new_n1189 = ~new_n1187 & new_n1188;
  assign new_n1190 = ~new_n1178 & ~new_n1181;
  assign new_n1191 = ~new_n1182 & new_n1190;
  assign new_n1192 = new_n1189 & new_n1191;
  assign new_n1193 = ~new_n1163 & ~new_n1166;
  assign new_n1194 = ~new_n1168 & new_n1193;
  assign new_n1195 = ~new_n1170 & ~new_n1172;
  assign new_n1196 = ~new_n1176 & new_n1195;
  assign new_n1197 = new_n1194 & new_n1196;
  assign d7 = ~new_n1192 | ~new_n1197;
  assign new_n1199 = p2 & ~q2;
  assign new_n1200 = ~p2 & q2;
  assign e6 = new_n1199 | new_n1200;
  assign new_n1202 = ~c1 & new_n1099;
  assign f5 = new_n1103 | new_n1202;
  assign new_n1204 = p0 & ~y1;
  assign new_n1205 = y1 & k1;
  assign g4 = new_n1204 | new_n1205;
  assign new_n1207 = ~new_n1106 & ~new_n1129;
  assign b6 = new_n1107 | ~new_n1207;
  assign new_n1209 = ~y3 & new_n290;
  assign new_n1210 = o1 & new_n1209;
  assign new_n1211 = ~new_n1161 & new_n1210;
  assign new_n1212 = new_n290 & ~new_n1161;
  assign new_n1213 = m1 & new_n1212;
  assign new_n1214 = ~s1 & ~y3;
  assign new_n1215 = o1 & new_n1214;
  assign new_n1216 = ~new_n1161 & new_n1215;
  assign new_n1217 = ~s1 & ~new_n1161;
  assign new_n1218 = m1 & new_n1217;
  assign new_n1219 = ~new_n1211 & ~new_n1213;
  assign new_n1220 = ~new_n1216 & ~new_n1218;
  assign c7 = ~new_n1219 | ~new_n1220;
  assign new_n1222 = x1 & m2;
  assign new_n1223 = ~y1 & new_n1222;
  assign c6 = w1 & new_n1223;
  assign new_n1225 = e1 & ~d1;
  assign new_n1226 = ~e1 & d1;
  assign new_n1227 = c1 & new_n1226;
  assign new_n1228 = ~c1 & e1;
  assign new_n1229 = ~new_n1225 & ~new_n1227;
  assign c5 = new_n1228 | ~new_n1229;
  assign new_n1231 = ~y & n0;
  assign new_n1232 = ~x & y;
  assign new_n1233 = e0 & new_n1232;
  assign new_n1234 = x & n0;
  assign new_n1235 = ~new_n1231 & ~new_n1233;
  assign a6 = new_n1234 | ~new_n1235;
  assign new_n1237 = c1 & ~d1;
  assign new_n1238 = ~c1 & d1;
  assign b5 = new_n1237 | new_n1238;
  assign new_n1240 = s1 & ~r1;
  assign new_n1241 = ~d & new_n1240;
  assign new_n1242 = ~e & new_n1240;
  assign new_n1243 = ~e & b1;
  assign new_n1244 = ~f & b1;
  assign new_n1245 = ~d & b1;
  assign new_n1246 = ~f & new_n1240;
  assign new_n1247 = ~new_n1241 & ~new_n1242;
  assign new_n1248 = ~new_n1243 & new_n1247;
  assign new_n1249 = ~new_n1244 & ~new_n1245;
  assign new_n1250 = ~new_n1246 & new_n1249;
  assign m5 = ~new_n1248 | ~new_n1250;
  assign new_n1252 = i3 & ~new_n717;
  assign new_n1253 = ~i3 & new_n717;
  assign new_n1254 = h3 & new_n1253;
  assign new_n1255 = ~new_n1252 & ~new_n1254;
  assign n6 = new_n808 | ~new_n1255;
  assign new_n1257 = ~new_n392 & new_n441;
  assign o7 = ~new_n363 | new_n1257;
  assign a8 = c4 | new_n789;
  assign new_n1260 = c1 & e1;
  assign new_n1261 = d1 & new_n1260;
  assign l5 = n & new_n1261;
  assign n7 = new_n363 & new_n392;
  assign new_n1264 = z2 & new_n824;
  assign new_n1265 = new_n675 & new_n711;
  assign new_n1266 = z2 & new_n1265;
  assign new_n1267 = ~u & new_n854;
  assign new_n1268 = ~h0 & new_n846;
  assign new_n1269 = new_n675 & ~new_n820;
  assign new_n1270 = z2 & new_n1269;
  assign new_n1271 = ~new_n1268 & ~new_n1270;
  assign new_n1272 = ~new_n1264 & ~new_n1266;
  assign new_n1273 = ~new_n1267 & new_n1272;
  assign o6 = ~new_n1271 | ~new_n1273;
  assign new_n1275 = x2 & new_n337;
  assign new_n1276 = new_n296 & new_n1275;
  assign b8 = ~w2 & new_n1276;
  assign new_n1278 = ~i3 & m2;
  assign new_n1279 = ~k2 & new_n1278;
  assign new_n1280 = p2 & ~k2;
  assign new_n1281 = h3 & m2;
  assign new_n1282 = ~k2 & new_n1281;
  assign k6 = ~k2 & ~m0;
  assign new_n1284 = ~new_n1279 & ~new_n1280;
  assign new_n1285 = ~new_n1282 & ~k6;
  assign l6 = ~new_n1284 | ~new_n1285;
  assign new_n1287 = new_n363 & ~new_n392;
  assign m7 = ~new_n441 & new_n1287;
  assign new_n1289 = d1 & new_n1111;
  assign new_n1290 = e1 & new_n1289;
  assign new_n1291 = c1 & new_n1290;
  assign new_n1292 = ~n & new_n1111;
  assign new_n1293 = ~w1 & new_n296;
  assign new_n1294 = ~new_n1291 & ~new_n1292;
  assign new_n1295 = new_n1140 & ~new_n1293;
  assign n4 = ~new_n1294 | ~new_n1295;
  assign new_n1297 = f2 & ~l2;
  assign new_n1298 = h2 & new_n1297;
  assign new_n1299 = h2 & ~l2;
  assign new_n1300 = ~g2 & new_n1299;
  assign o5 = new_n1298 | new_n1300;
  assign new_n1302 = w2 & ~new_n296;
  assign c8 = ~a4 | new_n1302;
  assign new_n1304 = s & ~l3;
  assign new_n1305 = u2 & new_n404;
  assign new_n1306 = ~new_n1304 & ~new_n1305;
  assign l7 = new_n392 | ~new_n1306;
  assign new_n1308 = h3 & ~new_n717;
  assign new_n1309 = ~new_n808 & ~new_n1308;
  assign m6 = new_n533 | ~new_n1309;
  assign new_n1311 = g2 & ~l2;
  assign new_n1312 = h2 & new_n1311;
  assign new_n1313 = ~f2 & new_n1312;
  assign n5 = a | new_n1313;
  assign o4 = w1 & new_n296;
  assign i5 = new_n1103 | new_n1125;
  assign new_n1317 = ~q2 & ~new_n389;
  assign new_n1318 = r0 & new_n1317;
  assign new_n1319 = ~l2 & ~new_n389;
  assign new_n1320 = r0 & new_n1319;
  assign new_n1321 = ~p2 & ~new_n389;
  assign new_n1322 = r0 & new_n1321;
  assign new_n1323 = ~new_n1318 & ~new_n1320;
  assign new_n1324 = ~new_n533 & ~new_n1322;
  assign j6 = ~new_n1323 | ~new_n1324;
  assign k7 = i1 | new_n1111;
  assign new_n1327 = ~c1 & new_n1125;
  assign h5 = new_n1103 | new_n1327;
  assign j7 = ~m1 & ~d8;
  assign new_n1330 = ~p0 & q0;
  assign new_n1331 = ~new_n1141 & new_n1330;
  assign new_n1332 = p0 & ~q0;
  assign new_n1333 = ~new_n1141 & new_n1332;
  assign new_n1334 = w3 & new_n1141;
  assign new_n1335 = ~new_n1331 & ~new_n1333;
  assign h6 = new_n1334 | ~new_n1335;
  assign i7 = y3 & new_n958;
  assign new_n1338 = ~k1 & l1;
  assign new_n1339 = ~new_n1118 & new_n1338;
  assign new_n1340 = k1 & ~l1;
  assign new_n1341 = ~new_n1118 & new_n1340;
  assign new_n1342 = r3 & new_n1118;
  assign new_n1343 = ~new_n1339 & ~new_n1341;
  assign h7 = new_n1342 | ~new_n1343;
  assign i6 = l3 & ~new_n527;
  assign new_n1346 = ~c1 & l2;
  assign j5 = new_n1103 | new_n1346;
  assign d6 = ~p2;
  assign l4 = ~o3;
  assign w7 = c0;
  assign v7 = b0;
  assign w6 = y0;
  assign u7 = a0;
  assign t7 = z;
  assign s7 = w;
  assign z6 = v6;
  assign y6 = w0;
  assign a5 = m2;
  assign b7 = z0;
  assign a7 = y0;
  assign m4 = t3;
  assign e8 = x6;
  assign f8 = w0;
  assign k5 = l2;
  assign g8 = x0;
  assign k4 = s3;
endmodule


