// Benchmark "top" written by ABC on Mon Feb 19 11:52:45 2024

module top ( 
    pp, pq, pr, ps, pt, pu, pv, pw, px, py, pa, pb, pc, pe, pf, pg, ph, pi,
    pj, pk, pl, pm, pn, po,
    pa0, pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pz, pk0, pl0, pm0,
    pn0, po0, pp0, pq0, pr0, ps0, pt0  );
  input  pp, pq, pr, ps, pt, pu, pv, pw, px, py, pa, pb, pc, pe, pf, pg,
    ph, pi, pj, pk, pl, pm, pn, po;
  output pa0, pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pz, pk0, pl0, pm0,
    pn0, po0, pp0, pq0, pr0, ps0, pt0;
  wire new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52,
    new_n53, new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60,
    new_n61, new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68,
    new_n69, new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76,
    new_n77, new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84,
    new_n85, new_n86, new_n87, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n102, new_n103, new_n104, new_n105, new_n106, new_n107, new_n108,
    new_n109, new_n110, new_n111, new_n112, new_n113, new_n114, new_n115,
    new_n116, new_n117, new_n118, new_n119, new_n120, new_n121, new_n122,
    new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n129,
    new_n130, new_n131, new_n132, new_n133, new_n134, new_n135, new_n136,
    new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n374, new_n375, new_n376, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n396, new_n397, new_n398, new_n399,
    new_n400, new_n401, new_n402, new_n403, new_n404, new_n405, new_n406,
    new_n407, new_n408, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n418, new_n419, new_n420,
    new_n421, new_n422, new_n423, new_n424, new_n425, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553;
  assign new_n46 = pq & pw;
  assign new_n47 = pq & ~pv;
  assign new_n48 = ~new_n46 & ~new_n47;
  assign new_n49 = ~pv & ~py;
  assign new_n50 = pw & new_n48;
  assign new_n51 = ~new_n49 & new_n50;
  assign new_n52 = ps & ~pv;
  assign new_n53 = ps & ~pf;
  assign new_n54 = pt & ~pf;
  assign new_n55 = ~pt & ~pu;
  assign new_n56 = pt & new_n55;
  assign new_n57 = pt & ~pv;
  assign new_n58 = ~pv & py;
  assign new_n59 = pu & new_n58;
  assign new_n60 = ~pu & pv;
  assign new_n61 = ~new_n59 & ~new_n60;
  assign new_n62 = ~pf & new_n61;
  assign new_n63 = new_n55 & new_n61;
  assign new_n64 = ps & new_n55;
  assign new_n65 = ~pv & new_n61;
  assign new_n66 = ~new_n64 & ~new_n65;
  assign new_n67 = ~new_n62 & ~new_n63;
  assign new_n68 = new_n66 & new_n67;
  assign new_n69 = ~new_n56 & ~new_n57;
  assign new_n70 = ~new_n52 & ~new_n53;
  assign new_n71 = ~new_n54 & new_n70;
  assign new_n72 = new_n69 & new_n71;
  assign new_n73 = new_n68 & new_n72;
  assign new_n74 = new_n48 & new_n73;
  assign new_n75 = ~pu & new_n74;
  assign new_n76 = pt & new_n50;
  assign new_n77 = ~ps & new_n50;
  assign new_n78 = ~pu & new_n50;
  assign new_n79 = ~new_n49 & new_n74;
  assign new_n80 = pt & new_n74;
  assign new_n81 = ~ps & new_n74;
  assign new_n82 = ~new_n51 & ~new_n75;
  assign new_n83 = ~new_n76 & ~new_n77;
  assign new_n84 = new_n82 & new_n83;
  assign new_n85 = ~new_n80 & ~new_n81;
  assign new_n86 = ~new_n78 & ~new_n79;
  assign new_n87 = new_n85 & new_n86;
  assign pa0 = ~new_n84 | ~new_n87;
  assign new_n89 = ~pt & py;
  assign new_n90 = ~pv & new_n89;
  assign new_n91 = ~ps & new_n90;
  assign new_n92 = pv & ~pg;
  assign new_n93 = ~pu & ~pv;
  assign new_n94 = ~new_n91 & ~new_n92;
  assign new_n95 = ~new_n55 & ~new_n93;
  assign new_n96 = new_n94 & new_n95;
  assign new_n97 = ~pt & ~py;
  assign new_n98 = new_n52 & new_n97;
  assign new_n99 = new_n96 & new_n98;
  assign new_n100 = ~pw & new_n96;
  assign pb0 = new_n99 | new_n100;
  assign new_n102 = ~ps & new_n58;
  assign new_n103 = pq & new_n102;
  assign new_n104 = ~pt & new_n103;
  assign new_n105 = ~pw & new_n93;
  assign new_n106 = ~new_n104 & ~new_n105;
  assign new_n107 = pw & new_n106;
  assign new_n108 = new_n98 & new_n107;
  assign new_n109 = ~ps & new_n108;
  assign new_n110 = pt & new_n108;
  assign new_n111 = pt & new_n106;
  assign new_n112 = pw & new_n111;
  assign new_n113 = ~pq & new_n112;
  assign new_n114 = pu & new_n106;
  assign new_n115 = pw & new_n114;
  assign new_n116 = ~pq & new_n115;
  assign new_n117 = ~ps & new_n106;
  assign new_n118 = pw & new_n117;
  assign new_n119 = ~pq & new_n118;
  assign new_n120 = pt & pv;
  assign new_n121 = pu & pv;
  assign new_n122 = pt & ~pu;
  assign new_n123 = ~new_n120 & ~new_n121;
  assign new_n124 = ~new_n122 & new_n123;
  assign new_n125 = new_n98 & new_n106;
  assign new_n126 = new_n124 & new_n125;
  assign new_n127 = pt & new_n126;
  assign new_n128 = ph & new_n125;
  assign new_n129 = pu & new_n128;
  assign new_n130 = ~ps & new_n126;
  assign new_n131 = ~pq & pw;
  assign new_n132 = new_n106 & new_n131;
  assign new_n133 = ph & new_n132;
  assign new_n134 = ~pq & new_n133;
  assign new_n135 = new_n124 & new_n132;
  assign new_n136 = ~pq & new_n135;
  assign new_n137 = ~pw & new_n133;
  assign new_n138 = pu & new_n126;
  assign new_n139 = new_n98 & new_n133;
  assign new_n140 = ~pw & new_n106;
  assign new_n141 = new_n124 & new_n140;
  assign new_n142 = ~ps & new_n141;
  assign new_n143 = ph & new_n140;
  assign new_n144 = pt & new_n143;
  assign new_n145 = new_n114 & new_n124;
  assign new_n146 = ~pq & new_n145;
  assign new_n147 = pu & new_n143;
  assign new_n148 = pu & new_n141;
  assign new_n149 = ~ps & new_n128;
  assign new_n150 = pt & new_n141;
  assign new_n151 = pt & new_n128;
  assign new_n152 = ~pw & new_n135;
  assign new_n153 = new_n98 & new_n135;
  assign new_n154 = new_n111 & new_n124;
  assign new_n155 = ~pq & new_n154;
  assign new_n156 = ph & new_n114;
  assign new_n157 = ~pq & new_n156;
  assign new_n158 = new_n117 & new_n124;
  assign new_n159 = ~pq & new_n158;
  assign new_n160 = ~ps & new_n143;
  assign new_n161 = ph & new_n111;
  assign new_n162 = ~pq & new_n161;
  assign new_n163 = new_n125 & new_n131;
  assign new_n164 = pw & new_n163;
  assign new_n165 = ph & new_n117;
  assign new_n166 = ~pq & new_n165;
  assign new_n167 = pu & new_n108;
  assign new_n168 = new_n107 & new_n131;
  assign new_n169 = ~pq & new_n168;
  assign new_n170 = ~new_n144 & ~new_n146;
  assign new_n171 = ~new_n139 & ~new_n142;
  assign new_n172 = new_n170 & new_n171;
  assign new_n173 = ~new_n137 & ~new_n138;
  assign new_n174 = ~new_n134 & ~new_n136;
  assign new_n175 = new_n173 & new_n174;
  assign new_n176 = new_n172 & new_n175;
  assign new_n177 = ~new_n109 & ~new_n110;
  assign new_n178 = ~new_n113 & ~new_n116;
  assign new_n179 = new_n177 & new_n178;
  assign new_n180 = ~new_n129 & ~new_n130;
  assign new_n181 = ~new_n119 & ~new_n127;
  assign new_n182 = new_n180 & new_n181;
  assign new_n183 = new_n179 & new_n182;
  assign new_n184 = new_n176 & new_n183;
  assign new_n185 = ~new_n167 & ~new_n169;
  assign new_n186 = ~new_n164 & ~new_n166;
  assign new_n187 = new_n185 & new_n186;
  assign new_n188 = ~new_n160 & ~new_n162;
  assign new_n189 = ~new_n157 & ~new_n159;
  assign new_n190 = new_n188 & new_n189;
  assign new_n191 = new_n187 & new_n190;
  assign new_n192 = ~new_n153 & ~new_n155;
  assign new_n193 = ~new_n151 & ~new_n152;
  assign new_n194 = new_n192 & new_n193;
  assign new_n195 = ~new_n147 & ~new_n148;
  assign new_n196 = ~new_n149 & ~new_n150;
  assign new_n197 = new_n195 & new_n196;
  assign new_n198 = new_n194 & new_n197;
  assign new_n199 = new_n191 & new_n198;
  assign pc0 = ~new_n184 | ~new_n199;
  assign new_n201 = pu & ~pv;
  assign new_n202 = pv & ~pi;
  assign new_n203 = ~ps & ~pv;
  assign new_n204 = ~new_n201 & ~new_n202;
  assign new_n205 = ~new_n55 & ~new_n203;
  assign new_n206 = new_n204 & new_n205;
  assign pd0 = ~pw & new_n206;
  assign new_n208 = ~pt & pv;
  assign new_n209 = ~pu & new_n208;
  assign new_n210 = ~ps & new_n209;
  assign new_n211 = ~pj & new_n120;
  assign new_n212 = ps & new_n57;
  assign new_n213 = pu & ~pj;
  assign new_n214 = ~new_n210 & ~new_n211;
  assign new_n215 = ~new_n212 & ~new_n213;
  assign new_n216 = new_n214 & new_n215;
  assign new_n217 = ~pw & new_n216;
  assign new_n218 = ~pu & new_n217;
  assign new_n219 = pv & new_n217;
  assign pe0 = new_n218 | new_n219;
  assign pf0 = ~pa & ~pk;
  assign new_n222 = pk & pm;
  assign new_n223 = ~pl & new_n222;
  assign new_n224 = ~pa & new_n223;
  assign new_n225 = pk & ~pn;
  assign new_n226 = ~pl & new_n225;
  assign new_n227 = ~pa & new_n226;
  assign new_n228 = ~pk & pl;
  assign new_n229 = ~pa & new_n228;
  assign new_n230 = ~new_n224 & ~new_n227;
  assign pg0 = new_n229 | ~new_n230;
  assign new_n232 = ~pl & pm;
  assign new_n233 = ~pa & new_n232;
  assign new_n234 = pk & ~pm;
  assign new_n235 = pl & new_n234;
  assign new_n236 = ~pa & new_n235;
  assign new_n237 = ~pk & pm;
  assign new_n238 = ~pa & new_n237;
  assign new_n239 = ~new_n233 & ~new_n236;
  assign ph0 = new_n238 | ~new_n239;
  assign new_n241 = ~pl & ~pm;
  assign new_n242 = pk & new_n241;
  assign new_n243 = pl & pn;
  assign new_n244 = pm & new_n243;
  assign new_n245 = pk & new_n244;
  assign new_n246 = ~new_n242 & ~new_n245;
  assign new_n247 = ~pa & new_n246;
  assign new_n248 = pk & pl;
  assign new_n249 = pm & new_n248;
  assign new_n250 = new_n247 & new_n249;
  assign new_n251 = pn & new_n247;
  assign pi0 = new_n250 | new_n251;
  assign new_n253 = ~pa & po;
  assign new_n254 = ~px & new_n253;
  assign new_n255 = ~pk & new_n254;
  assign new_n256 = pl & new_n254;
  assign new_n257 = ~pa & ~po;
  assign new_n258 = px & new_n257;
  assign new_n259 = pl & new_n258;
  assign new_n260 = pm & new_n258;
  assign new_n261 = ~pk & new_n258;
  assign new_n262 = ~pl & pn;
  assign new_n263 = new_n234 & new_n262;
  assign new_n264 = ~px & ~pa;
  assign new_n265 = new_n263 & new_n264;
  assign new_n266 = pl & new_n265;
  assign new_n267 = pm & new_n265;
  assign new_n268 = pn & po;
  assign new_n269 = ~pa & ~new_n268;
  assign new_n270 = new_n263 & new_n269;
  assign new_n271 = ~po & new_n270;
  assign new_n272 = ~px & new_n270;
  assign new_n273 = new_n257 & new_n263;
  assign new_n274 = pm & new_n273;
  assign new_n275 = ~pk & new_n265;
  assign new_n276 = pl & new_n273;
  assign new_n277 = new_n264 & ~new_n268;
  assign new_n278 = po & new_n277;
  assign new_n279 = ~pk & new_n273;
  assign new_n280 = pm & new_n254;
  assign new_n281 = px & ~pa;
  assign new_n282 = ~new_n268 & new_n281;
  assign new_n283 = ~po & new_n282;
  assign new_n284 = ~new_n280 & ~new_n283;
  assign new_n285 = ~new_n278 & ~new_n279;
  assign new_n286 = new_n284 & new_n285;
  assign new_n287 = ~new_n275 & ~new_n276;
  assign new_n288 = ~new_n272 & ~new_n274;
  assign new_n289 = new_n287 & new_n288;
  assign new_n290 = new_n286 & new_n289;
  assign new_n291 = ~new_n255 & ~new_n256;
  assign new_n292 = ~new_n259 & ~new_n260;
  assign new_n293 = new_n291 & new_n292;
  assign new_n294 = ~new_n267 & ~new_n271;
  assign new_n295 = ~new_n261 & ~new_n266;
  assign new_n296 = new_n294 & new_n295;
  assign new_n297 = new_n293 & new_n296;
  assign pj0 = ~new_n290 | ~new_n297;
  assign new_n299 = ~pe & new_n120;
  assign new_n300 = ~ps & pv;
  assign new_n301 = ~pe & new_n300;
  assign new_n302 = pu & ~pe;
  assign new_n303 = ~new_n301 & ~new_n302;
  assign new_n304 = ~new_n210 & ~new_n299;
  assign new_n305 = ~new_n201 & new_n304;
  assign new_n306 = new_n303 & new_n305;
  assign pz = ~pw & new_n306;
  assign new_n308 = ~pq & pr;
  assign new_n309 = px & new_n308;
  assign new_n310 = po & new_n309;
  assign new_n311 = ~pp & ~po;
  assign new_n312 = pp & px;
  assign new_n313 = po & new_n312;
  assign new_n314 = ~new_n310 & ~new_n311;
  assign new_n315 = ~pa & ~new_n313;
  assign new_n316 = new_n314 & new_n315;
  assign new_n317 = ~pp & ~new_n308;
  assign new_n318 = px & new_n316;
  assign new_n319 = new_n317 & new_n318;
  assign new_n320 = pp & new_n316;
  assign new_n321 = pl & new_n320;
  assign new_n322 = ~pk & new_n318;
  assign new_n323 = ~pm & pn;
  assign new_n324 = po & new_n323;
  assign new_n325 = new_n318 & ~new_n324;
  assign new_n326 = pl & new_n318;
  assign new_n327 = new_n263 & new_n316;
  assign new_n328 = ~new_n324 & new_n327;
  assign new_n329 = new_n317 & new_n327;
  assign new_n330 = ~pk & new_n327;
  assign new_n331 = new_n317 & new_n320;
  assign new_n332 = pl & new_n327;
  assign new_n333 = ~pk & new_n320;
  assign new_n334 = new_n320 & ~new_n324;
  assign new_n335 = ~new_n332 & ~new_n333;
  assign new_n336 = ~new_n334 & new_n335;
  assign new_n337 = ~new_n329 & ~new_n330;
  assign new_n338 = ~new_n331 & new_n337;
  assign new_n339 = new_n336 & new_n338;
  assign new_n340 = ~new_n319 & ~new_n321;
  assign new_n341 = ~new_n322 & new_n340;
  assign new_n342 = ~new_n325 & ~new_n326;
  assign new_n343 = ~new_n328 & new_n342;
  assign new_n344 = new_n341 & new_n343;
  assign pk0 = ~new_n339 | ~new_n344;
  assign new_n346 = ~pq & ~po;
  assign new_n347 = ~pp & ~pq;
  assign new_n348 = ~new_n346 & ~new_n347;
  assign new_n349 = ~pa & new_n348;
  assign new_n350 = px & new_n349;
  assign new_n351 = ~pp & new_n350;
  assign new_n352 = ~pq & new_n350;
  assign new_n353 = pq & new_n349;
  assign new_n354 = ~pp & new_n353;
  assign new_n355 = ~po & new_n350;
  assign new_n356 = ~po & new_n353;
  assign new_n357 = ~pm & new_n262;
  assign new_n358 = pk & new_n357;
  assign new_n359 = ~px & ~new_n358;
  assign new_n360 = new_n349 & new_n359;
  assign new_n361 = new_n263 & new_n360;
  assign new_n362 = px & new_n360;
  assign new_n363 = new_n263 & new_n349;
  assign new_n364 = ~pq & new_n363;
  assign new_n365 = pq & new_n360;
  assign new_n366 = ~po & new_n363;
  assign new_n367 = ~pp & new_n363;
  assign new_n368 = ~new_n351 & ~new_n352;
  assign new_n369 = ~new_n354 & new_n368;
  assign new_n370 = ~new_n355 & ~new_n356;
  assign new_n371 = ~new_n361 & new_n370;
  assign new_n372 = new_n369 & new_n371;
  assign new_n373 = ~new_n366 & ~new_n367;
  assign new_n374 = ~new_n362 & ~new_n364;
  assign new_n375 = ~new_n365 & new_n374;
  assign new_n376 = new_n373 & new_n375;
  assign pl0 = ~new_n372 | ~new_n376;
  assign new_n378 = ~pq & ~pr;
  assign new_n379 = ~pr & ~po;
  assign new_n380 = ~pp & ~pr;
  assign new_n381 = ~new_n378 & ~new_n379;
  assign new_n382 = ~pa & ~new_n380;
  assign new_n383 = new_n381 & new_n382;
  assign new_n384 = ~po & new_n383;
  assign new_n385 = px & new_n384;
  assign new_n386 = ~pk & new_n385;
  assign new_n387 = pl & new_n385;
  assign new_n388 = pq & pr;
  assign new_n389 = pp & new_n388;
  assign new_n390 = ~new_n347 & ~new_n389;
  assign new_n391 = new_n383 & new_n390;
  assign new_n392 = new_n263 & new_n391;
  assign new_n393 = pr & new_n391;
  assign new_n394 = px & new_n391;
  assign new_n395 = ~new_n324 & new_n383;
  assign new_n396 = pr & new_n395;
  assign new_n397 = ~po & new_n396;
  assign new_n398 = ~px & new_n396;
  assign new_n399 = pr & new_n384;
  assign new_n400 = ~pk & new_n399;
  assign new_n401 = pl & new_n399;
  assign new_n402 = ~px & new_n383;
  assign new_n403 = pr & new_n402;
  assign new_n404 = ~pk & new_n403;
  assign new_n405 = pl & new_n403;
  assign new_n406 = new_n263 & new_n383;
  assign new_n407 = ~new_n324 & new_n406;
  assign new_n408 = ~po & new_n407;
  assign new_n409 = ~px & new_n407;
  assign new_n410 = px & new_n383;
  assign new_n411 = ~new_n324 & new_n410;
  assign new_n412 = ~po & new_n411;
  assign new_n413 = new_n263 & new_n402;
  assign new_n414 = ~pk & new_n413;
  assign new_n415 = pl & new_n413;
  assign new_n416 = new_n263 & new_n384;
  assign new_n417 = ~pk & new_n416;
  assign new_n418 = pl & new_n416;
  assign new_n419 = ~new_n417 & ~new_n418;
  assign new_n420 = ~new_n414 & ~new_n415;
  assign new_n421 = new_n419 & new_n420;
  assign new_n422 = ~new_n409 & ~new_n412;
  assign new_n423 = ~new_n404 & ~new_n405;
  assign new_n424 = ~new_n408 & new_n423;
  assign new_n425 = new_n422 & new_n424;
  assign new_n426 = new_n421 & new_n425;
  assign new_n427 = ~new_n400 & ~new_n401;
  assign new_n428 = ~new_n397 & ~new_n398;
  assign new_n429 = new_n427 & new_n428;
  assign new_n430 = ~new_n393 & ~new_n394;
  assign new_n431 = ~new_n386 & ~new_n387;
  assign new_n432 = ~new_n392 & new_n431;
  assign new_n433 = new_n430 & new_n432;
  assign new_n434 = new_n429 & new_n433;
  assign pm0 = ~new_n426 | ~new_n434;
  assign new_n436 = ps & ~pa;
  assign new_n437 = new_n359 & new_n436;
  assign new_n438 = po & ~new_n359;
  assign new_n439 = ~pp & new_n308;
  assign new_n440 = new_n438 & new_n439;
  assign new_n441 = ~pa & new_n440;
  assign new_n442 = pp & new_n441;
  assign new_n443 = ~po & new_n436;
  assign new_n444 = ps & new_n308;
  assign new_n445 = new_n436 & ~new_n444;
  assign new_n446 = pp & new_n436;
  assign new_n447 = new_n359 & new_n441;
  assign new_n448 = ~po & new_n441;
  assign new_n449 = new_n441 & ~new_n444;
  assign new_n450 = ~new_n437 & ~new_n442;
  assign new_n451 = ~new_n443 & ~new_n445;
  assign new_n452 = new_n450 & new_n451;
  assign new_n453 = ~new_n448 & ~new_n449;
  assign new_n454 = ~new_n446 & ~new_n447;
  assign new_n455 = new_n453 & new_n454;
  assign pn0 = ~new_n452 | ~new_n455;
  assign new_n457 = ~pl & new_n234;
  assign new_n458 = pn & new_n457;
  assign new_n459 = ~px & ~new_n458;
  assign new_n460 = ~new_n60 & ~new_n459;
  assign new_n461 = ~pp & po;
  assign new_n462 = ~pq & ps;
  assign new_n463 = pr & ~pt;
  assign new_n464 = new_n462 & new_n463;
  assign new_n465 = new_n460 & new_n461;
  assign new_n466 = new_n464 & new_n465;
  assign new_n467 = ~pa & new_n466;
  assign new_n468 = pr & po;
  assign new_n469 = new_n462 & new_n468;
  assign new_n470 = ~pp & new_n469;
  assign new_n471 = new_n263 & new_n470;
  assign new_n472 = px & new_n470;
  assign new_n473 = ~new_n471 & ~new_n472;
  assign new_n474 = pt & new_n473;
  assign new_n475 = ~pa & new_n474;
  assign po0 = new_n467 | new_n475;
  assign new_n477 = ~px & ~pn;
  assign new_n478 = ~px & pl;
  assign new_n479 = ~px & pm;
  assign new_n480 = ~px & ~pk;
  assign new_n481 = ~new_n477 & ~new_n478;
  assign new_n482 = ~new_n479 & ~new_n480;
  assign new_n483 = new_n481 & new_n482;
  assign new_n484 = ~pq & new_n461;
  assign new_n485 = pr & pt;
  assign new_n486 = ps & ~pu;
  assign new_n487 = new_n485 & new_n486;
  assign new_n488 = new_n483 & new_n484;
  assign new_n489 = new_n487 & new_n488;
  assign new_n490 = ~pa & new_n489;
  assign new_n491 = ps & po;
  assign new_n492 = new_n485 & new_n491;
  assign new_n493 = ~pp & new_n492;
  assign new_n494 = ~pq & new_n493;
  assign new_n495 = new_n263 & new_n494;
  assign new_n496 = px & new_n494;
  assign new_n497 = ~new_n495 & ~new_n496;
  assign new_n498 = pu & new_n497;
  assign new_n499 = ~pa & new_n498;
  assign pp0 = new_n490 | new_n499;
  assign new_n501 = ps & pu;
  assign new_n502 = new_n57 & new_n501;
  assign new_n503 = ~pq & po;
  assign new_n504 = ~pp & pr;
  assign new_n505 = new_n503 & new_n504;
  assign new_n506 = new_n483 & new_n502;
  assign new_n507 = new_n505 & new_n506;
  assign new_n508 = ~pa & new_n507;
  assign new_n509 = pr & ~pu;
  assign new_n510 = ps & new_n509;
  assign new_n511 = ~pt & new_n510;
  assign new_n512 = pr & pu;
  assign new_n513 = ps & new_n512;
  assign new_n514 = pt & new_n513;
  assign new_n515 = ~new_n511 & ~new_n514;
  assign new_n516 = po & ~new_n515;
  assign new_n517 = ~pp & new_n516;
  assign new_n518 = ~pq & new_n517;
  assign new_n519 = new_n263 & new_n518;
  assign new_n520 = px & new_n518;
  assign new_n521 = ~new_n519 & ~new_n520;
  assign new_n522 = pv & new_n521;
  assign new_n523 = ~pa & new_n522;
  assign pq0 = new_n508 | new_n523;
  assign new_n525 = pw & ~pa;
  assign new_n526 = ~new_n49 & new_n525;
  assign new_n527 = ~pt & new_n58;
  assign new_n528 = ~ps & pu;
  assign new_n529 = new_n527 & new_n528;
  assign new_n530 = ~pa & new_n529;
  assign new_n531 = ~pu & new_n530;
  assign new_n532 = pt & new_n525;
  assign new_n533 = ~ps & new_n525;
  assign new_n534 = ~pu & new_n525;
  assign new_n535 = ~new_n49 & new_n530;
  assign new_n536 = pt & new_n530;
  assign new_n537 = ~ps & new_n530;
  assign new_n538 = ~new_n526 & ~new_n531;
  assign new_n539 = ~new_n532 & ~new_n533;
  assign new_n540 = new_n538 & new_n539;
  assign new_n541 = ~new_n536 & ~new_n537;
  assign new_n542 = ~new_n534 & ~new_n535;
  assign new_n543 = new_n541 & new_n542;
  assign pr0 = ~new_n540 | ~new_n543;
  assign new_n545 = ~px & pb;
  assign new_n546 = ~pa & new_n545;
  assign new_n547 = px & ~pb;
  assign new_n548 = ~pa & new_n547;
  assign ps0 = new_n546 | new_n548;
  assign new_n550 = ~py & pc;
  assign new_n551 = ~pa & new_n550;
  assign new_n552 = py & ~pc;
  assign new_n553 = ~pa & new_n552;
  assign pt0 = new_n551 | new_n553;
endmodule


