// Benchmark "top" written by ABC on Mon Feb 19 11:52:45 2024

module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0,
    pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pb, pr0, pc,
    ps0, pd, pt0, pe, pu0, pf, pv0, pg, pw0, ph, px0, pi, py0, pj, pz0, pk,
    pl, pm, pn, po,
    pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, ph1, ph2, pk1, pi2, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1,
    pu1, pt1, pw1, pv1, py1, px1, pz1  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, ph0, pi0, py, pj0, pz, pk0, pl0, pm0, pn0, po0, pp0, pa, pq0, pb,
    pr0, pc, ps0, pd, pt0, pe, pu0, pf, pv0, pg, pw0, ph, px0, pi, py0, pj,
    pz0, pk, pl, pm, pn, po;
  output pa1, pb2, pc2, pc1, pa2, pb1, pe1, pf2, pd1, pg2, pd2, pg1, pe2, pf1,
    pi1, ph1, ph2, pk1, pi2, pj1, pm1, pl1, po1, pn1, pq1, pp1, ps1, pr1,
    pu1, pt1, pw1, pv1, py1, px1, pz1;
  wire new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n102, new_n103, new_n104, new_n105, new_n106, new_n107, new_n108,
    new_n109, new_n110, new_n111, new_n112, new_n113, new_n114, new_n115,
    new_n116, new_n117, new_n118, new_n119, new_n120, new_n121, new_n122,
    new_n123, new_n124, new_n125, new_n126, new_n127, new_n128, new_n130,
    new_n131, new_n132, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n158, new_n159, new_n160, new_n161,
    new_n162, new_n163, new_n164, new_n165, new_n166, new_n167, new_n168,
    new_n169, new_n170, new_n171, new_n172, new_n173, new_n174, new_n175,
    new_n176, new_n177, new_n178, new_n179, new_n180, new_n181, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n195, new_n196, new_n197,
    new_n198, new_n199, new_n200, new_n201, new_n202, new_n203, new_n204,
    new_n205, new_n206, new_n207, new_n208, new_n209, new_n210, new_n211,
    new_n212, new_n213, new_n214, new_n215, new_n216, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n226, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n450, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1409, new_n1410, new_n1411, new_n1412, new_n1413, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1435, new_n1436, new_n1437, new_n1438, new_n1439,
    new_n1440, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1446, new_n1447, new_n1448, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495, new_n1496, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1501, new_n1502, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507, new_n1508, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1640, new_n1641, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655;
  assign new_n87 = pa0 & ~pb;
  assign new_n88 = pf0 & ~pb;
  assign new_n89 = pa0 & pm;
  assign new_n90 = pa0 & ~pl;
  assign new_n91 = pa0 & pn;
  assign new_n92 = ~pb & pr0;
  assign new_n93 = pa0 & ~pr;
  assign new_n94 = ~pv & new_n93;
  assign new_n95 = ~pj & new_n94;
  assign new_n96 = ~new_n87 & ~new_n88;
  assign new_n97 = ~new_n89 & ~new_n90;
  assign new_n98 = new_n96 & new_n97;
  assign new_n99 = ~new_n91 & ~new_n92;
  assign new_n100 = ~new_n95 & new_n99;
  assign pa1 = ~new_n98 | ~new_n100;
  assign new_n102 = ~pm & po;
  assign new_n103 = ~pe & new_n102;
  assign new_n104 = ~pg & new_n103;
  assign new_n105 = ~pa & new_n104;
  assign new_n106 = pp0 & new_n105;
  assign new_n107 = ~pv & new_n106;
  assign new_n108 = ~pw & new_n107;
  assign new_n109 = pp & new_n108;
  assign new_n110 = ~pu & new_n109;
  assign new_n111 = ~pp & po;
  assign new_n112 = ~pe & new_n111;
  assign new_n113 = ~pm & new_n112;
  assign new_n114 = ~pa & new_n113;
  assign new_n115 = ~pw & new_n114;
  assign new_n116 = pp0 & new_n115;
  assign new_n117 = ~pu & new_n116;
  assign new_n118 = ~pv & new_n117;
  assign new_n119 = pe0 & new_n105;
  assign new_n120 = ~pv & new_n119;
  assign new_n121 = ~pw & new_n120;
  assign new_n122 = pp & new_n121;
  assign new_n123 = ~pu & new_n122;
  assign new_n124 = pe0 & new_n115;
  assign new_n125 = ~pu & new_n124;
  assign new_n126 = ~pv & new_n125;
  assign new_n127 = ~new_n110 & ~new_n118;
  assign new_n128 = ~new_n123 & ~new_n126;
  assign pb2 = ~new_n127 | ~new_n128;
  assign new_n130 = pb0 & ~pm;
  assign new_n131 = ~pv & new_n130;
  assign new_n132 = pb0 & pv;
  assign pc1 = new_n131 | new_n132;
  assign pa2 = pf0 | pr0;
  assign new_n135 = ~pm & ~pn;
  assign new_n136 = pb & new_n135;
  assign new_n137 = pj & new_n136;
  assign new_n138 = ~pa & new_n137;
  assign new_n139 = pa0 & new_n138;
  assign new_n140 = ~pk & new_n139;
  assign new_n141 = pl & new_n140;
  assign new_n142 = ~pj & new_n136;
  assign new_n143 = ~pa & new_n142;
  assign new_n144 = pl & new_n143;
  assign new_n145 = pa0 & new_n144;
  assign new_n146 = pv & new_n145;
  assign new_n147 = ~pk & new_n146;
  assign new_n148 = pg0 & pc;
  assign new_n149 = ~pw & new_n148;
  assign new_n150 = pj & new_n149;
  assign new_n151 = pv & new_n143;
  assign new_n152 = pk0 & new_n151;
  assign new_n153 = po0 & pt0;
  assign new_n154 = ~new_n152 & ~new_n153;
  assign new_n155 = ~new_n141 & ~new_n147;
  assign new_n156 = ~new_n150 & new_n155;
  assign pb1 = ~new_n154 | ~new_n156;
  assign new_n158 = pd0 & ~po;
  assign new_n159 = pg & new_n158;
  assign new_n160 = ~pm & new_n159;
  assign new_n161 = pd & new_n160;
  assign new_n162 = pe & new_n161;
  assign new_n163 = pd0 & ~pu;
  assign new_n164 = ~pm & new_n163;
  assign new_n165 = ~po & new_n164;
  assign new_n166 = pd & new_n165;
  assign new_n167 = ~pe & new_n166;
  assign new_n168 = ~pw & new_n167;
  assign new_n169 = pe0 & ~ph;
  assign new_n170 = ~po & new_n169;
  assign new_n171 = ~pa & new_n170;
  assign new_n172 = ~pm & new_n171;
  assign new_n173 = pu & ~po;
  assign new_n174 = pg & new_n173;
  assign new_n175 = ~pm & new_n174;
  assign new_n176 = pd & new_n175;
  assign new_n177 = pd0 & new_n176;
  assign new_n178 = po0 & pu0;
  assign new_n179 = ~new_n177 & ~new_n178;
  assign new_n180 = ~new_n162 & ~new_n168;
  assign new_n181 = ~new_n172 & new_n180;
  assign pe1 = ~new_n179 | ~new_n181;
  assign new_n183 = ~pi0 & ~pm0;
  assign new_n184 = ~pa0 & new_n183;
  assign new_n185 = ~pf0 & new_n184;
  assign new_n186 = po & new_n185;
  assign new_n187 = pd & new_n186;
  assign new_n188 = ~ps0 & new_n187;
  assign new_n189 = ~px0 & new_n188;
  assign new_n190 = ~pp0 & new_n189;
  assign new_n191 = ~pr0 & new_n190;
  assign new_n192 = ~pd0 & new_n183;
  assign new_n193 = ~pf0 & new_n192;
  assign new_n194 = ~pa0 & new_n193;
  assign new_n195 = ~pe0 & new_n194;
  assign new_n196 = ~ps0 & new_n195;
  assign new_n197 = ~px0 & new_n196;
  assign new_n198 = ~pp0 & new_n197;
  assign new_n199 = ~pr0 & new_n198;
  assign new_n200 = ~ph & ~px0;
  assign new_n201 = ~pm0 & new_n200;
  assign new_n202 = ~pr0 & new_n201;
  assign new_n203 = ~pf0 & new_n202;
  assign new_n204 = pz0 & new_n203;
  assign new_n205 = pb & new_n204;
  assign new_n206 = pl & new_n205;
  assign new_n207 = ~pf0 & ~pi0;
  assign new_n208 = ~pa0 & new_n207;
  assign new_n209 = ~pd0 & new_n208;
  assign new_n210 = po & new_n209;
  assign new_n211 = ~px0 & new_n210;
  assign new_n212 = ~pr0 & new_n211;
  assign new_n213 = ~ps0 & new_n212;
  assign new_n214 = ~pm0 & new_n213;
  assign new_n215 = ~pp0 & new_n214;
  assign new_n216 = ~pr0 & ~px0;
  assign new_n217 = ~pf0 & new_n216;
  assign new_n218 = ~pm0 & new_n217;
  assign new_n219 = ~pa0 & new_n218;
  assign new_n220 = ~ph & new_n219;
  assign new_n221 = ~pp0 & ~pr0;
  assign new_n222 = ~pf0 & new_n221;
  assign new_n223 = ~pm0 & new_n222;
  assign new_n224 = po & new_n223;
  assign new_n225 = pl & new_n224;
  assign new_n226 = pz0 & new_n225;
  assign new_n227 = pb & new_n226;
  assign new_n228 = pd & new_n227;
  assign new_n229 = ~pt & new_n228;
  assign new_n230 = ~ps0 & new_n229;
  assign new_n231 = ~px0 & new_n230;
  assign new_n232 = ~pr0 & ~ps0;
  assign new_n233 = ~pm0 & new_n232;
  assign new_n234 = ~pp0 & new_n233;
  assign new_n235 = ~pf0 & new_n234;
  assign new_n236 = ~pm & new_n235;
  assign new_n237 = pr & new_n236;
  assign new_n238 = ~pj & new_n237;
  assign new_n239 = pl & new_n238;
  assign new_n240 = pb & new_n239;
  assign new_n241 = ~pe0 & new_n240;
  assign new_n242 = ~pt & new_n241;
  assign new_n243 = ~px0 & new_n242;
  assign new_n244 = pd & new_n243;
  assign new_n245 = ~pd0 & new_n223;
  assign new_n246 = pl & new_n245;
  assign new_n247 = pz0 & new_n246;
  assign new_n248 = pb & new_n247;
  assign new_n249 = ~pe0 & new_n248;
  assign new_n250 = ~pt & new_n249;
  assign new_n251 = ~ps0 & new_n250;
  assign new_n252 = ~px0 & new_n251;
  assign new_n253 = pl & new_n235;
  assign new_n254 = pz0 & new_n253;
  assign new_n255 = pb & new_n254;
  assign new_n256 = ~pe0 & new_n255;
  assign new_n257 = ~pt & new_n256;
  assign new_n258 = ~px0 & new_n257;
  assign new_n259 = pd & new_n258;
  assign new_n260 = po & new_n193;
  assign new_n261 = ~pm & new_n260;
  assign new_n262 = pr & new_n261;
  assign new_n263 = ~pj & new_n262;
  assign new_n264 = pl & new_n263;
  assign new_n265 = pb & new_n264;
  assign new_n266 = ~ps0 & new_n265;
  assign new_n267 = ~px0 & new_n266;
  assign new_n268 = ~pp0 & new_n267;
  assign new_n269 = ~pr0 & new_n268;
  assign new_n270 = ~pm0 & ~pp0;
  assign new_n271 = ~pd0 & new_n270;
  assign new_n272 = ~pf0 & new_n271;
  assign new_n273 = po & new_n272;
  assign new_n274 = ~pm & new_n273;
  assign new_n275 = pr & new_n274;
  assign new_n276 = ~pj & new_n275;
  assign new_n277 = pl & new_n276;
  assign new_n278 = pb & new_n277;
  assign new_n279 = ~px0 & new_n278;
  assign new_n280 = ~pt & new_n279;
  assign new_n281 = ~pr0 & new_n280;
  assign new_n282 = ~ps0 & new_n281;
  assign new_n283 = ~pf0 & new_n270;
  assign new_n284 = ~pi0 & new_n283;
  assign new_n285 = po & new_n284;
  assign new_n286 = pl & new_n285;
  assign new_n287 = pz0 & new_n286;
  assign new_n288 = pb & new_n287;
  assign new_n289 = ~px0 & new_n288;
  assign new_n290 = pd & new_n289;
  assign new_n291 = ~pr0 & new_n290;
  assign new_n292 = ~ps0 & new_n291;
  assign new_n293 = ~pi0 & new_n221;
  assign new_n294 = ~pm0 & new_n293;
  assign new_n295 = ~pf0 & new_n294;
  assign new_n296 = ~pm & new_n295;
  assign new_n297 = pr & new_n296;
  assign new_n298 = ~pj & new_n297;
  assign new_n299 = pl & new_n298;
  assign new_n300 = pb & new_n299;
  assign new_n301 = pd & new_n300;
  assign new_n302 = ~pe0 & new_n301;
  assign new_n303 = ~ps0 & new_n302;
  assign new_n304 = ~px0 & new_n303;
  assign new_n305 = ~pd0 & new_n284;
  assign new_n306 = pl & new_n305;
  assign new_n307 = pz0 & new_n306;
  assign new_n308 = pb & new_n307;
  assign new_n309 = ~px0 & new_n308;
  assign new_n310 = ~pe0 & new_n309;
  assign new_n311 = ~pr0 & new_n310;
  assign new_n312 = ~ps0 & new_n311;
  assign new_n313 = ~pm & new_n245;
  assign new_n314 = pr & new_n313;
  assign new_n315 = ~pj & new_n314;
  assign new_n316 = pl & new_n315;
  assign new_n317 = pb & new_n316;
  assign new_n318 = ~pe0 & new_n317;
  assign new_n319 = ~pt & new_n318;
  assign new_n320 = ~ps0 & new_n319;
  assign new_n321 = ~px0 & new_n320;
  assign new_n322 = pl & new_n295;
  assign new_n323 = pz0 & new_n322;
  assign new_n324 = pb & new_n323;
  assign new_n325 = pd & new_n324;
  assign new_n326 = ~pe0 & new_n325;
  assign new_n327 = ~ps0 & new_n326;
  assign new_n328 = ~px0 & new_n327;
  assign new_n329 = ~pm & new_n224;
  assign new_n330 = pr & new_n329;
  assign new_n331 = ~pj & new_n330;
  assign new_n332 = pl & new_n331;
  assign new_n333 = pb & new_n332;
  assign new_n334 = pd & new_n333;
  assign new_n335 = ~pt & new_n334;
  assign new_n336 = ~ps0 & new_n335;
  assign new_n337 = ~px0 & new_n336;
  assign new_n338 = pl & new_n273;
  assign new_n339 = pz0 & new_n338;
  assign new_n340 = pb & new_n339;
  assign new_n341 = ~px0 & new_n340;
  assign new_n342 = ~pt & new_n341;
  assign new_n343 = ~pr0 & new_n342;
  assign new_n344 = ~ps0 & new_n343;
  assign new_n345 = ~pm & new_n305;
  assign new_n346 = pr & new_n345;
  assign new_n347 = ~pj & new_n346;
  assign new_n348 = pl & new_n347;
  assign new_n349 = pb & new_n348;
  assign new_n350 = ~px0 & new_n349;
  assign new_n351 = ~pe0 & new_n350;
  assign new_n352 = ~pr0 & new_n351;
  assign new_n353 = ~ps0 & new_n352;
  assign new_n354 = pr & new_n203;
  assign new_n355 = pl & new_n354;
  assign new_n356 = ~pm & new_n355;
  assign new_n357 = pb & new_n356;
  assign new_n358 = ~pj & new_n357;
  assign new_n359 = ~pm & new_n285;
  assign new_n360 = pr & new_n359;
  assign new_n361 = ~pj & new_n360;
  assign new_n362 = pl & new_n361;
  assign new_n363 = pb & new_n362;
  assign new_n364 = ~px0 & new_n363;
  assign new_n365 = pd & new_n364;
  assign new_n366 = ~pr0 & new_n365;
  assign new_n367 = ~ps0 & new_n366;
  assign new_n368 = pl & new_n260;
  assign new_n369 = pz0 & new_n368;
  assign new_n370 = pb & new_n369;
  assign new_n371 = ~ps0 & new_n370;
  assign new_n372 = ~px0 & new_n371;
  assign new_n373 = ~pp0 & new_n372;
  assign new_n374 = ~pr0 & new_n373;
  assign new_n375 = ~pa0 & new_n223;
  assign new_n376 = ~pt & new_n375;
  assign new_n377 = pd & new_n376;
  assign new_n378 = ~pe0 & new_n377;
  assign new_n379 = ~ps0 & new_n378;
  assign new_n380 = ~px0 & new_n379;
  assign new_n381 = ~pa0 & new_n270;
  assign new_n382 = ~pf0 & new_n381;
  assign new_n383 = po & new_n382;
  assign new_n384 = ~pt & new_n383;
  assign new_n385 = ~px0 & new_n384;
  assign new_n386 = pd & new_n385;
  assign new_n387 = ~pr0 & new_n386;
  assign new_n388 = ~ps0 & new_n387;
  assign new_n389 = ~pa0 & new_n272;
  assign new_n390 = ~pt & new_n389;
  assign new_n391 = ~px0 & new_n390;
  assign new_n392 = ~pe0 & new_n391;
  assign new_n393 = ~pr0 & new_n392;
  assign new_n394 = ~ps0 & new_n393;
  assign new_n395 = ~pa0 & new_n284;
  assign new_n396 = ~pe0 & new_n395;
  assign new_n397 = ~px0 & new_n396;
  assign new_n398 = pd & new_n397;
  assign new_n399 = ~pr0 & new_n398;
  assign new_n400 = ~ps0 & new_n399;
  assign new_n401 = ~pf0 & ~pm0;
  assign new_n402 = ~pa0 & new_n401;
  assign new_n403 = ~pd0 & new_n402;
  assign new_n404 = po & new_n403;
  assign new_n405 = ~pt & new_n404;
  assign new_n406 = ~ps0 & new_n405;
  assign new_n407 = ~px0 & new_n406;
  assign new_n408 = ~pp0 & new_n407;
  assign new_n409 = ~pr0 & new_n408;
  assign new_n410 = ~new_n191 & ~new_n199;
  assign new_n411 = ~new_n206 & ~new_n215;
  assign new_n412 = new_n410 & new_n411;
  assign new_n413 = ~new_n220 & ~new_n231;
  assign new_n414 = ~new_n244 & new_n413;
  assign new_n415 = new_n412 & new_n414;
  assign new_n416 = ~new_n292 & ~new_n304;
  assign new_n417 = ~new_n312 & new_n416;
  assign new_n418 = ~new_n269 & ~new_n282;
  assign new_n419 = ~new_n252 & ~new_n259;
  assign new_n420 = new_n418 & new_n419;
  assign new_n421 = new_n417 & new_n420;
  assign new_n422 = new_n415 & new_n421;
  assign new_n423 = ~new_n394 & ~new_n400;
  assign new_n424 = ~new_n409 & new_n423;
  assign new_n425 = ~new_n374 & ~new_n380;
  assign new_n426 = ~new_n388 & new_n425;
  assign new_n427 = new_n424 & new_n426;
  assign new_n428 = ~new_n353 & ~new_n358;
  assign new_n429 = ~new_n367 & new_n428;
  assign new_n430 = ~new_n337 & ~new_n344;
  assign new_n431 = ~new_n321 & ~new_n328;
  assign new_n432 = new_n430 & new_n431;
  assign new_n433 = new_n429 & new_n432;
  assign new_n434 = new_n427 & new_n433;
  assign pf2 = ~new_n422 | ~new_n434;
  assign new_n436 = ~pd & ~ph;
  assign new_n437 = ~pm & new_n436;
  assign new_n438 = ~pa & new_n437;
  assign new_n439 = ~pv & new_n438;
  assign new_n440 = pd0 & new_n439;
  assign new_n441 = ~po & new_n440;
  assign new_n442 = pc0 & ~pm;
  assign new_n443 = ~pv & new_n442;
  assign new_n444 = ~pp & new_n439;
  assign new_n445 = pd0 & new_n444;
  assign new_n446 = pc0 & pv;
  assign new_n447 = ~new_n441 & ~new_n443;
  assign new_n448 = ~new_n445 & ~new_n446;
  assign pd1 = ~new_n447 | ~new_n448;
  assign new_n450 = ~pz0 & new_n89;
  assign new_n451 = pb & new_n450;
  assign new_n452 = pa0 & pj;
  assign new_n453 = ~pz0 & new_n452;
  assign new_n454 = pb & new_n453;
  assign new_n455 = pd0 & ~pd;
  assign new_n456 = ph & new_n455;
  assign new_n457 = pa0 & ~pz0;
  assign new_n458 = ~pr & new_n457;
  assign new_n459 = pb & new_n458;
  assign new_n460 = pe0 & ~po;
  assign new_n461 = ph & new_n460;
  assign new_n462 = pb & new_n90;
  assign new_n463 = pt & pi0;
  assign ps1 = ph & new_n463;
  assign new_n465 = pp0 & ph;
  assign new_n466 = ps0 & ph;
  assign new_n467 = ~pm0 & ~new_n87;
  assign new_n468 = new_n216 & new_n467;
  assign new_n469 = ~pf0 & ~new_n451;
  assign new_n470 = ~new_n454 & new_n469;
  assign new_n471 = new_n468 & new_n470;
  assign new_n472 = ~ps1 & ~new_n465;
  assign new_n473 = ~new_n466 & new_n472;
  assign new_n474 = ~new_n461 & ~new_n462;
  assign new_n475 = ~new_n456 & ~new_n459;
  assign new_n476 = new_n474 & new_n475;
  assign new_n477 = new_n473 & new_n476;
  assign pg2 = ~new_n471 | ~new_n477;
  assign new_n479 = pp0 & pi;
  assign new_n480 = pv & new_n479;
  assign new_n481 = ~pa & new_n480;
  assign new_n482 = ~pv & pq0;
  assign new_n483 = pg & new_n482;
  assign new_n484 = pi & new_n483;
  assign new_n485 = ~pa & new_n484;
  assign new_n486 = ~po & new_n485;
  assign new_n487 = ~pp & new_n485;
  assign new_n488 = pp0 & ~po;
  assign new_n489 = pg & new_n488;
  assign new_n490 = pi & new_n489;
  assign new_n491 = ~pa & new_n490;
  assign new_n492 = ~pq & ~pv;
  assign new_n493 = pg & new_n492;
  assign new_n494 = pi & new_n493;
  assign new_n495 = ~pa & new_n494;
  assign new_n496 = pq0 & new_n495;
  assign new_n497 = ~pq & pp0;
  assign new_n498 = pg & new_n497;
  assign new_n499 = pi & new_n498;
  assign new_n500 = ~pa & new_n499;
  assign new_n501 = ~pp & pp0;
  assign new_n502 = pg & new_n501;
  assign new_n503 = pi & new_n502;
  assign new_n504 = ~pa & new_n503;
  assign new_n505 = ~new_n500 & ~new_n504;
  assign new_n506 = ~new_n487 & ~new_n491;
  assign new_n507 = ~new_n496 & new_n506;
  assign new_n508 = new_n505 & new_n507;
  assign new_n509 = ~pi0 & ~pz;
  assign new_n510 = ~new_n486 & new_n509;
  assign new_n511 = ~py & ~new_n481;
  assign new_n512 = ~ph0 & new_n511;
  assign new_n513 = new_n510 & new_n512;
  assign pd2 = ~new_n508 | ~new_n513;
  assign new_n515 = pp & ~pv;
  assign new_n516 = ~pm & new_n515;
  assign new_n517 = po & new_n516;
  assign new_n518 = pe & new_n517;
  assign new_n519 = pd0 & new_n518;
  assign new_n520 = pg & new_n519;
  assign new_n521 = pu & ~pv;
  assign new_n522 = po & new_n521;
  assign new_n523 = pp & new_n522;
  assign new_n524 = ~pm & new_n523;
  assign new_n525 = pd0 & new_n524;
  assign new_n526 = pg & new_n525;
  assign new_n527 = po0 & pv0;
  assign new_n528 = pp & ~pu;
  assign new_n529 = ~pm & new_n528;
  assign new_n530 = po & new_n529;
  assign new_n531 = ~pe & new_n530;
  assign new_n532 = ~pv & new_n531;
  assign new_n533 = pd0 & new_n532;
  assign new_n534 = pd0 & pv;
  assign new_n535 = ~pa & ~pg;
  assign new_n536 = ~pp & new_n535;
  assign new_n537 = ~pv & new_n536;
  assign new_n538 = ~pm & new_n537;
  assign new_n539 = ~pd & new_n538;
  assign new_n540 = ~ps & new_n539;
  assign new_n541 = ~ph & new_n540;
  assign new_n542 = pp0 & new_n541;
  assign new_n543 = ~ph & new_n498;
  assign new_n544 = ~pa & new_n543;
  assign new_n545 = ~pi & new_n544;
  assign new_n546 = ~ps & new_n545;
  assign new_n547 = ~po & new_n535;
  assign new_n548 = ~pv & new_n547;
  assign new_n549 = ~pm & new_n548;
  assign new_n550 = ~pd & new_n549;
  assign new_n551 = ~ps & new_n550;
  assign new_n552 = ~ph & new_n551;
  assign new_n553 = pp0 & new_n552;
  assign new_n554 = ~pa & ~pc;
  assign new_n555 = ~po & new_n554;
  assign new_n556 = ~pv & new_n555;
  assign new_n557 = ~pm & new_n556;
  assign new_n558 = ~pr & new_n557;
  assign new_n559 = pp0 & new_n558;
  assign new_n560 = ~pg & new_n559;
  assign new_n561 = ~ph & new_n560;
  assign new_n562 = ~pp & new_n554;
  assign new_n563 = ~pv & new_n562;
  assign new_n564 = ~pm & new_n563;
  assign new_n565 = ~pr & new_n564;
  assign new_n566 = pp0 & new_n565;
  assign new_n567 = ~pg & new_n566;
  assign new_n568 = ~ph & new_n567;
  assign new_n569 = ~pg & ~ph;
  assign new_n570 = ~pv & new_n569;
  assign new_n571 = ~pa & new_n570;
  assign new_n572 = ~pm & new_n571;
  assign new_n573 = ~pd & new_n572;
  assign new_n574 = ~ps & new_n573;
  assign new_n575 = ~pq & new_n574;
  assign new_n576 = pp0 & new_n575;
  assign new_n577 = ~pc & ~pg;
  assign new_n578 = ~pv & new_n577;
  assign new_n579 = ~pa & new_n578;
  assign new_n580 = ~pm & new_n579;
  assign new_n581 = ~pr & new_n580;
  assign new_n582 = pp0 & new_n581;
  assign new_n583 = ~ph & new_n582;
  assign new_n584 = ~pq & new_n583;
  assign new_n585 = pp0 & new_n557;
  assign new_n586 = ~ps & new_n585;
  assign new_n587 = ~pg & new_n586;
  assign new_n588 = ~ph & new_n587;
  assign new_n589 = pp0 & ~ph;
  assign new_n590 = pv & new_n589;
  assign new_n591 = ~pa & new_n590;
  assign new_n592 = ~pp & new_n591;
  assign new_n593 = ~pi & new_n592;
  assign new_n594 = ~ps & new_n593;
  assign new_n595 = pp0 & new_n572;
  assign new_n596 = ~pd & new_n595;
  assign new_n597 = ~pq & new_n596;
  assign new_n598 = ~pr & new_n597;
  assign new_n599 = ~pa & new_n589;
  assign new_n600 = pg & new_n599;
  assign new_n601 = ~po & new_n600;
  assign new_n602 = ~pi & new_n601;
  assign new_n603 = ~ps & new_n602;
  assign new_n604 = pp0 & new_n580;
  assign new_n605 = ~ps & new_n604;
  assign new_n606 = ~ph & new_n605;
  assign new_n607 = ~pq & new_n606;
  assign new_n608 = ~pp & new_n600;
  assign new_n609 = ~pi & new_n608;
  assign new_n610 = ~ps & new_n609;
  assign new_n611 = pp0 & new_n564;
  assign new_n612 = ~ps & new_n611;
  assign new_n613 = ~pg & new_n612;
  assign new_n614 = ~ph & new_n613;
  assign new_n615 = ~pa & new_n497;
  assign new_n616 = ~ph & new_n615;
  assign new_n617 = pv & new_n616;
  assign new_n618 = ~pi & new_n617;
  assign new_n619 = ~ps & new_n618;
  assign new_n620 = pp0 & new_n538;
  assign new_n621 = ~pd & new_n620;
  assign new_n622 = ~ph & new_n621;
  assign new_n623 = ~pr & new_n622;
  assign new_n624 = ~pq & ~pr;
  assign new_n625 = pg & new_n624;
  assign new_n626 = ~ph & new_n625;
  assign new_n627 = ~pa & new_n626;
  assign new_n628 = pp0 & new_n627;
  assign new_n629 = ~pi & new_n628;
  assign new_n630 = pp0 & new_n549;
  assign new_n631 = ~pd & new_n630;
  assign new_n632 = ~ph & new_n631;
  assign new_n633 = ~pr & new_n632;
  assign new_n634 = ~po & new_n591;
  assign new_n635 = ~pi & new_n634;
  assign new_n636 = ~ps & new_n635;
  assign new_n637 = ~pa & new_n624;
  assign new_n638 = ~ph & new_n637;
  assign new_n639 = pv & new_n638;
  assign new_n640 = pp0 & new_n639;
  assign new_n641 = ~pi & new_n640;
  assign new_n642 = ~pr & ~ph;
  assign new_n643 = ~pa & new_n642;
  assign new_n644 = pg & new_n643;
  assign new_n645 = ~po & new_n644;
  assign new_n646 = pp0 & new_n645;
  assign new_n647 = ~pi & new_n646;
  assign new_n648 = ~pp & new_n644;
  assign new_n649 = pp0 & new_n648;
  assign new_n650 = ~pi & new_n649;
  assign new_n651 = pv & new_n642;
  assign new_n652 = ~pa & new_n651;
  assign new_n653 = ~po & new_n652;
  assign new_n654 = pp0 & new_n653;
  assign new_n655 = ~pi & new_n654;
  assign new_n656 = ~pp & new_n652;
  assign new_n657 = pp0 & new_n656;
  assign new_n658 = ~pi & new_n657;
  assign new_n659 = ~new_n650 & ~new_n655;
  assign new_n660 = ~new_n658 & new_n659;
  assign new_n661 = ~new_n641 & ~new_n647;
  assign new_n662 = ~new_n633 & ~new_n636;
  assign new_n663 = new_n661 & new_n662;
  assign new_n664 = new_n660 & new_n663;
  assign new_n665 = ~new_n619 & ~new_n623;
  assign new_n666 = ~new_n629 & new_n665;
  assign new_n667 = ~new_n610 & ~new_n614;
  assign new_n668 = ~new_n603 & ~new_n607;
  assign new_n669 = new_n667 & new_n668;
  assign new_n670 = new_n666 & new_n669;
  assign new_n671 = new_n664 & new_n670;
  assign new_n672 = ~new_n520 & ~new_n526;
  assign new_n673 = ~new_n527 & ~new_n533;
  assign new_n674 = new_n672 & new_n673;
  assign new_n675 = ~new_n546 & ~new_n553;
  assign new_n676 = ~new_n534 & ~new_n542;
  assign new_n677 = new_n675 & new_n676;
  assign new_n678 = new_n674 & new_n677;
  assign new_n679 = ~new_n588 & ~new_n594;
  assign new_n680 = ~new_n598 & new_n679;
  assign new_n681 = ~new_n576 & ~new_n584;
  assign new_n682 = ~new_n561 & ~new_n568;
  assign new_n683 = new_n681 & new_n682;
  assign new_n684 = new_n680 & new_n683;
  assign new_n685 = new_n678 & new_n684;
  assign pg1 = ~new_n671 | ~new_n685;
  assign new_n687 = ~pi0 & ~pg;
  assign new_n688 = ~pz & new_n687;
  assign new_n689 = ~ph0 & new_n688;
  assign new_n690 = ~py & new_n689;
  assign new_n691 = ~pp0 & new_n690;
  assign new_n692 = pv & ~pi0;
  assign new_n693 = ~pz & new_n692;
  assign new_n694 = ~ph0 & new_n693;
  assign new_n695 = ~py & new_n694;
  assign new_n696 = ~pp0 & new_n695;
  assign new_n697 = ~pi0 & ~pi;
  assign new_n698 = ~pz & new_n697;
  assign new_n699 = ~ph0 & new_n698;
  assign new_n700 = ~py & new_n699;
  assign new_n701 = ~pv & new_n690;
  assign new_n702 = ~ph0 & ~pi0;
  assign new_n703 = ~py & new_n702;
  assign new_n704 = ~pz & new_n703;
  assign new_n705 = pa & new_n704;
  assign new_n706 = ~pi0 & ~pp0;
  assign new_n707 = ~pz & new_n706;
  assign new_n708 = ~ph0 & new_n707;
  assign new_n709 = ~py & new_n708;
  assign new_n710 = pq & new_n709;
  assign new_n711 = po & new_n710;
  assign new_n712 = pp & new_n711;
  assign new_n713 = ~pq0 & new_n709;
  assign new_n714 = ~pv & ~pi0;
  assign new_n715 = ~pz & new_n714;
  assign new_n716 = ~ph0 & new_n715;
  assign new_n717 = ~py & new_n716;
  assign new_n718 = pq & new_n717;
  assign new_n719 = po & new_n718;
  assign new_n720 = pp & new_n719;
  assign new_n721 = ~new_n691 & ~new_n696;
  assign new_n722 = ~new_n700 & ~new_n701;
  assign new_n723 = new_n721 & new_n722;
  assign new_n724 = ~new_n713 & ~new_n720;
  assign new_n725 = ~new_n705 & ~new_n712;
  assign new_n726 = new_n724 & new_n725;
  assign pe2 = ~new_n723 | ~new_n726;
  assign new_n728 = ~pq & ~pi;
  assign new_n729 = pq0 & new_n728;
  assign new_n730 = pp & ~pm;
  assign new_n731 = ~pa & new_n730;
  assign new_n732 = ~ph & new_n731;
  assign new_n733 = po & new_n732;
  assign new_n734 = pe0 & new_n733;
  assign new_n735 = ~pq & pq0;
  assign new_n736 = ~pg & new_n735;
  assign new_n737 = pq0 & ~pi;
  assign new_n738 = ~po & new_n737;
  assign new_n739 = pq0 & ~po;
  assign new_n740 = ~pg & new_n739;
  assign new_n741 = ~new_n738 & ~new_n740;
  assign new_n742 = ~new_n729 & ~new_n734;
  assign new_n743 = ~new_n736 & new_n742;
  assign pf1 = ~new_n741 | ~new_n743;
  assign new_n745 = ~pu & ~pw;
  assign new_n746 = ~pe & new_n745;
  assign new_n747 = ph & new_n746;
  assign new_n748 = ~pa & new_n747;
  assign new_n749 = ~po & new_n748;
  assign new_n750 = pe0 & new_n749;
  assign new_n751 = pp0 & new_n748;
  assign new_n752 = ~pd & new_n748;
  assign new_n753 = pd0 & new_n752;
  assign new_n754 = ps0 & new_n748;
  assign new_n755 = ~new_n750 & ~new_n751;
  assign new_n756 = ~new_n753 & ~new_n754;
  assign ph1 = ~new_n755 | ~new_n756;
  assign new_n758 = ~pb0 & ~pc0;
  assign new_n759 = ~py & new_n758;
  assign new_n760 = ~pz & new_n759;
  assign new_n761 = ~pi & new_n760;
  assign new_n762 = ~pc & new_n761;
  assign new_n763 = ~pd0 & new_n762;
  assign new_n764 = ~ph0 & new_n763;
  assign new_n765 = ~pb & new_n764;
  assign new_n766 = ~pb0 & ~pz;
  assign new_n767 = ~pl & new_n766;
  assign new_n768 = ~py & new_n767;
  assign new_n769 = ~pj & new_n768;
  assign new_n770 = ~pd0 & new_n769;
  assign new_n771 = ~pi0 & new_n770;
  assign new_n772 = ~pc0 & new_n771;
  assign new_n773 = ~ph0 & new_n772;
  assign new_n774 = ~pj & new_n766;
  assign new_n775 = ~py & new_n774;
  assign new_n776 = ~pi & new_n775;
  assign new_n777 = ~pb & new_n776;
  assign new_n778 = ~pd0 & new_n777;
  assign new_n779 = ~pc0 & new_n778;
  assign new_n780 = ~ph0 & new_n779;
  assign new_n781 = ~pi & new_n768;
  assign new_n782 = ~pc & new_n781;
  assign new_n783 = ~pd0 & new_n782;
  assign new_n784 = ~pc0 & new_n783;
  assign new_n785 = ~ph0 & new_n784;
  assign new_n786 = ~py & ~pz;
  assign new_n787 = ~pj & new_n786;
  assign new_n788 = ~pl & new_n787;
  assign new_n789 = ~pi & new_n788;
  assign new_n790 = ~ph0 & new_n789;
  assign new_n791 = ~pd0 & new_n790;
  assign new_n792 = ~pb0 & new_n791;
  assign new_n793 = ~pc0 & new_n792;
  assign new_n794 = ph & new_n786;
  assign new_n795 = ~pj & new_n794;
  assign new_n796 = ~pd & new_n795;
  assign new_n797 = ~pv & new_n796;
  assign new_n798 = ~ph0 & new_n797;
  assign new_n799 = ~pi0 & new_n798;
  assign new_n800 = ~pb0 & new_n799;
  assign new_n801 = ~pc0 & new_n800;
  assign new_n802 = ~pl & new_n794;
  assign new_n803 = ~pd & new_n802;
  assign new_n804 = ~pi0 & new_n803;
  assign new_n805 = ~ph0 & new_n804;
  assign new_n806 = ~pc & new_n805;
  assign new_n807 = ~pb0 & new_n806;
  assign new_n808 = ~pc0 & new_n807;
  assign new_n809 = ~pd0 & new_n761;
  assign new_n810 = pn & new_n809;
  assign new_n811 = ~ph0 & new_n810;
  assign new_n812 = ~pc & new_n811;
  assign new_n813 = ~pj & new_n760;
  assign new_n814 = ~pi0 & new_n813;
  assign new_n815 = pa & new_n814;
  assign new_n816 = ~ph0 & new_n815;
  assign new_n817 = ~pd0 & new_n816;
  assign new_n818 = ~py & ~pj;
  assign new_n819 = ph & new_n818;
  assign new_n820 = ~pi & new_n819;
  assign new_n821 = ~pd & new_n820;
  assign new_n822 = ~pv & new_n821;
  assign new_n823 = ~pc0 & new_n822;
  assign new_n824 = ~ph0 & new_n823;
  assign new_n825 = ~pz & new_n824;
  assign new_n826 = ~pb0 & new_n825;
  assign new_n827 = ph & new_n766;
  assign new_n828 = ~py & new_n827;
  assign new_n829 = ~pd & new_n828;
  assign new_n830 = ~pi0 & new_n829;
  assign new_n831 = ~pb & new_n830;
  assign new_n832 = ~pc & new_n831;
  assign new_n833 = ~pc0 & new_n832;
  assign new_n834 = ~ph0 & new_n833;
  assign new_n835 = ~pd0 & new_n776;
  assign new_n836 = pn & new_n835;
  assign new_n837 = ~pc0 & new_n836;
  assign new_n838 = ~ph0 & new_n837;
  assign new_n839 = ~pc0 & ~ph0;
  assign new_n840 = ~pz & new_n839;
  assign new_n841 = ~pb0 & new_n840;
  assign new_n842 = ~py & new_n841;
  assign new_n843 = ~pi0 & new_n842;
  assign new_n844 = pa & new_n843;
  assign new_n845 = ~pc & new_n844;
  assign new_n846 = ~pd0 & new_n845;
  assign new_n847 = ~pi & new_n794;
  assign new_n848 = ~pd & new_n847;
  assign new_n849 = ~pk0 & new_n848;
  assign new_n850 = ~pg0 & new_n849;
  assign new_n851 = ~ph0 & new_n850;
  assign new_n852 = ~pa0 & new_n851;
  assign new_n853 = ~pb0 & new_n852;
  assign new_n854 = ~pc0 & new_n853;
  assign new_n855 = pj & new_n760;
  assign new_n856 = ~pg0 & new_n855;
  assign new_n857 = ~pi0 & new_n856;
  assign new_n858 = ~pa0 & new_n857;
  assign new_n859 = ~ph0 & new_n858;
  assign new_n860 = ~pd0 & new_n859;
  assign new_n861 = ~py & ~pl;
  assign new_n862 = ph & new_n861;
  assign new_n863 = ~pj & new_n862;
  assign new_n864 = ~pd & new_n863;
  assign new_n865 = ~pi0 & new_n864;
  assign new_n866 = ~pc0 & new_n865;
  assign new_n867 = ~ph0 & new_n866;
  assign new_n868 = ~pz & new_n867;
  assign new_n869 = ~pb0 & new_n868;
  assign new_n870 = pn & new_n843;
  assign new_n871 = ~pc & new_n870;
  assign new_n872 = ~pd0 & new_n871;
  assign new_n873 = ~pg0 & new_n761;
  assign new_n874 = pa & new_n873;
  assign new_n875 = ~ph0 & new_n874;
  assign new_n876 = ~pd0 & new_n875;
  assign new_n877 = ~pk0 & new_n829;
  assign new_n878 = ~pg0 & new_n877;
  assign new_n879 = ~pi0 & new_n878;
  assign new_n880 = ~pa0 & new_n879;
  assign new_n881 = ~pc0 & new_n880;
  assign new_n882 = ~ph0 & new_n881;
  assign new_n883 = pj & new_n766;
  assign new_n884 = ~py & new_n883;
  assign new_n885 = ~pi & new_n884;
  assign new_n886 = ~pg0 & new_n885;
  assign new_n887 = ~pd0 & new_n886;
  assign new_n888 = ~pa0 & new_n887;
  assign new_n889 = ~pc0 & new_n888;
  assign new_n890 = ~ph0 & new_n889;
  assign new_n891 = ~pi0 & new_n796;
  assign new_n892 = ~ph0 & new_n891;
  assign new_n893 = ~pb & new_n892;
  assign new_n894 = ~pb0 & new_n893;
  assign new_n895 = ~pc0 & new_n894;
  assign new_n896 = pn & new_n814;
  assign new_n897 = ~ph0 & new_n896;
  assign new_n898 = ~pd0 & new_n897;
  assign new_n899 = ~pg0 & new_n842;
  assign new_n900 = pa & new_n899;
  assign new_n901 = ~pd0 & new_n900;
  assign new_n902 = ~pi0 & new_n901;
  assign new_n903 = pj & new_n794;
  assign new_n904 = ~pd & new_n903;
  assign new_n905 = ~pg0 & new_n904;
  assign new_n906 = ~pa0 & new_n905;
  assign new_n907 = ~ph0 & new_n906;
  assign new_n908 = ~pi0 & new_n907;
  assign new_n909 = ~pb0 & new_n908;
  assign new_n910 = ~pc0 & new_n909;
  assign new_n911 = pn & new_n848;
  assign new_n912 = ~ph0 & new_n911;
  assign new_n913 = ~pg0 & new_n912;
  assign new_n914 = ~pb0 & new_n913;
  assign new_n915 = ~pc0 & new_n914;
  assign new_n916 = ~pg0 & new_n829;
  assign new_n917 = ~pb & new_n916;
  assign new_n918 = ~pi0 & new_n917;
  assign new_n919 = ~pc0 & new_n918;
  assign new_n920 = ~ph0 & new_n919;
  assign new_n921 = ~pi & new_n862;
  assign new_n922 = ~pd & new_n921;
  assign new_n923 = ~pc & new_n922;
  assign new_n924 = ~pc0 & new_n923;
  assign new_n925 = ~ph0 & new_n924;
  assign new_n926 = ~pz & new_n925;
  assign new_n927 = ~pb0 & new_n926;
  assign new_n928 = pm & new_n843;
  assign new_n929 = ~pc & new_n928;
  assign new_n930 = ~pd0 & new_n929;
  assign new_n931 = ~pv & new_n835;
  assign new_n932 = ~pc0 & new_n931;
  assign new_n933 = ~ph0 & new_n932;
  assign new_n934 = ~py & pj;
  assign new_n935 = ph & new_n934;
  assign new_n936 = ~pi & new_n935;
  assign new_n937 = ~pd & new_n936;
  assign new_n938 = ~pg0 & new_n937;
  assign new_n939 = ~pa0 & new_n938;
  assign new_n940 = ~pc0 & new_n939;
  assign new_n941 = ~ph0 & new_n940;
  assign new_n942 = ~pz & new_n941;
  assign new_n943 = ~pb0 & new_n942;
  assign new_n944 = pn & new_n829;
  assign new_n945 = ~pi0 & new_n944;
  assign new_n946 = ~pg0 & new_n945;
  assign new_n947 = ~pc0 & new_n946;
  assign new_n948 = ~ph0 & new_n947;
  assign new_n949 = ~pg0 & new_n803;
  assign new_n950 = ~ph0 & new_n949;
  assign new_n951 = ~pi0 & new_n950;
  assign new_n952 = ~pb0 & new_n951;
  assign new_n953 = ~pc0 & new_n952;
  assign new_n954 = ~pc & new_n848;
  assign new_n955 = ~ph0 & new_n954;
  assign new_n956 = ~pb & new_n955;
  assign new_n957 = ~pb0 & new_n956;
  assign new_n958 = ~pc0 & new_n957;
  assign new_n959 = pm & new_n814;
  assign new_n960 = ~ph0 & new_n959;
  assign new_n961 = ~pd0 & new_n960;
  assign new_n962 = ~pv & new_n814;
  assign new_n963 = ~ph0 & new_n962;
  assign new_n964 = ~pd0 & new_n963;
  assign new_n965 = pm & new_n848;
  assign new_n966 = ~ph0 & new_n965;
  assign new_n967 = ~pc & new_n966;
  assign new_n968 = ~pb0 & new_n967;
  assign new_n969 = ~pc0 & new_n968;
  assign new_n970 = ~pv & new_n761;
  assign new_n971 = ~pd0 & new_n970;
  assign new_n972 = ~pa0 & new_n971;
  assign new_n973 = ~ph0 & new_n972;
  assign new_n974 = ~pc & new_n973;
  assign new_n975 = ~pg0 & new_n848;
  assign new_n976 = ~ph0 & new_n975;
  assign new_n977 = ~pb & new_n976;
  assign new_n978 = ~pb0 & new_n977;
  assign new_n979 = ~pc0 & new_n978;
  assign new_n980 = ~pj & ~pl;
  assign new_n981 = ph & new_n980;
  assign new_n982 = ~pi & new_n981;
  assign new_n983 = ~pd & new_n982;
  assign new_n984 = ~ph0 & new_n983;
  assign new_n985 = ~pb0 & new_n984;
  assign new_n986 = ~pc0 & new_n985;
  assign new_n987 = ~py & new_n986;
  assign new_n988 = ~pz & new_n987;
  assign new_n989 = pm & new_n899;
  assign new_n990 = ~pd0 & new_n989;
  assign new_n991 = ~pi0 & new_n990;
  assign new_n992 = pa & new_n835;
  assign new_n993 = ~pc0 & new_n992;
  assign new_n994 = ~ph0 & new_n993;
  assign new_n995 = pm & new_n821;
  assign new_n996 = ~pc0 & new_n995;
  assign new_n997 = ~ph0 & new_n996;
  assign new_n998 = ~pz & new_n997;
  assign new_n999 = ~pb0 & new_n998;
  assign new_n1000 = ~pv & new_n842;
  assign new_n1001 = ~pi0 & new_n1000;
  assign new_n1002 = ~pa0 & new_n1001;
  assign new_n1003 = ~pc & new_n1002;
  assign new_n1004 = ~pd0 & new_n1003;
  assign new_n1005 = ~pg0 & new_n922;
  assign new_n1006 = ~pc0 & new_n1005;
  assign new_n1007 = ~ph0 & new_n1006;
  assign new_n1008 = ~pz & new_n1007;
  assign new_n1009 = ~pb0 & new_n1008;
  assign new_n1010 = ~pb & new_n821;
  assign new_n1011 = ~pc0 & new_n1010;
  assign new_n1012 = ~ph0 & new_n1011;
  assign new_n1013 = ~pz & new_n1012;
  assign new_n1014 = ~pb0 & new_n1013;
  assign new_n1015 = pm & new_n873;
  assign new_n1016 = ~ph0 & new_n1015;
  assign new_n1017 = ~pd0 & new_n1016;
  assign new_n1018 = pa & new_n809;
  assign new_n1019 = ~ph0 & new_n1018;
  assign new_n1020 = ~pc & new_n1019;
  assign new_n1021 = ~pv & new_n829;
  assign new_n1022 = ~pg0 & new_n1021;
  assign new_n1023 = ~pi0 & new_n1022;
  assign new_n1024 = ~pa0 & new_n1023;
  assign new_n1025 = ~pc0 & new_n1024;
  assign new_n1026 = ~ph0 & new_n1025;
  assign new_n1027 = ~pk0 & new_n813;
  assign new_n1028 = ~pi0 & new_n1027;
  assign new_n1029 = ~pa0 & new_n1028;
  assign new_n1030 = ~ph0 & new_n1029;
  assign new_n1031 = ~pd0 & new_n1030;
  assign new_n1032 = pm & new_n829;
  assign new_n1033 = ~pc & new_n1032;
  assign new_n1034 = ~pi0 & new_n1033;
  assign new_n1035 = ~pc0 & new_n1034;
  assign new_n1036 = ~ph0 & new_n1035;
  assign new_n1037 = ~pa0 & new_n970;
  assign new_n1038 = ~pg0 & new_n1037;
  assign new_n1039 = ~ph0 & new_n1038;
  assign new_n1040 = ~pd0 & new_n1039;
  assign new_n1041 = ~pa0 & new_n855;
  assign new_n1042 = ~pd0 & new_n1041;
  assign new_n1043 = ~pi0 & new_n1042;
  assign new_n1044 = ~ph0 & new_n1043;
  assign new_n1045 = ~pc & new_n1044;
  assign new_n1046 = pn & new_n873;
  assign new_n1047 = ~ph0 & new_n1046;
  assign new_n1048 = ~pd0 & new_n1047;
  assign new_n1049 = ~pv & new_n848;
  assign new_n1050 = ~pg0 & new_n1049;
  assign new_n1051 = ~ph0 & new_n1050;
  assign new_n1052 = ~pa0 & new_n1051;
  assign new_n1053 = ~pb0 & new_n1052;
  assign new_n1054 = ~pc0 & new_n1053;
  assign new_n1055 = ~pk0 & new_n842;
  assign new_n1056 = ~pi0 & new_n1055;
  assign new_n1057 = ~pa0 & new_n1056;
  assign new_n1058 = ~pc & new_n1057;
  assign new_n1059 = ~pd0 & new_n1058;
  assign new_n1060 = pm & new_n796;
  assign new_n1061 = ~ph0 & new_n1060;
  assign new_n1062 = ~pi0 & new_n1061;
  assign new_n1063 = ~pb0 & new_n1062;
  assign new_n1064 = ~pc0 & new_n1063;
  assign new_n1065 = ~pa0 & new_n1000;
  assign new_n1066 = ~pg0 & new_n1065;
  assign new_n1067 = ~pd0 & new_n1066;
  assign new_n1068 = ~pi0 & new_n1067;
  assign new_n1069 = ~pa0 & new_n885;
  assign new_n1070 = ~pc & new_n1069;
  assign new_n1071 = ~pd0 & new_n1070;
  assign new_n1072 = ~pc0 & new_n1071;
  assign new_n1073 = ~ph0 & new_n1072;
  assign new_n1074 = pn & new_n899;
  assign new_n1075 = ~pd0 & new_n1074;
  assign new_n1076 = ~pi0 & new_n1075;
  assign new_n1077 = ~pa0 & new_n1021;
  assign new_n1078 = ~pc & new_n1077;
  assign new_n1079 = ~pi0 & new_n1078;
  assign new_n1080 = ~pc0 & new_n1079;
  assign new_n1081 = ~ph0 & new_n1080;
  assign new_n1082 = ~pk0 & new_n776;
  assign new_n1083 = ~pd0 & new_n1082;
  assign new_n1084 = ~pa0 & new_n1083;
  assign new_n1085 = ~pc0 & new_n1084;
  assign new_n1086 = ~ph0 & new_n1085;
  assign new_n1087 = ~pi0 & new_n1032;
  assign new_n1088 = ~pg0 & new_n1087;
  assign new_n1089 = ~pc0 & new_n1088;
  assign new_n1090 = ~ph0 & new_n1089;
  assign new_n1091 = pa & new_n821;
  assign new_n1092 = ~pc0 & new_n1091;
  assign new_n1093 = ~ph0 & new_n1092;
  assign new_n1094 = ~pz & new_n1093;
  assign new_n1095 = ~pb0 & new_n1094;
  assign new_n1096 = pm & new_n809;
  assign new_n1097 = ~ph0 & new_n1096;
  assign new_n1098 = ~pc & new_n1097;
  assign new_n1099 = ~pl & new_n760;
  assign new_n1100 = ~pi0 & new_n1099;
  assign new_n1101 = ~pg0 & new_n1100;
  assign new_n1102 = ~ph0 & new_n1101;
  assign new_n1103 = ~pd0 & new_n1102;
  assign new_n1104 = ~pa0 & new_n1049;
  assign new_n1105 = ~ph0 & new_n1104;
  assign new_n1106 = ~pc & new_n1105;
  assign new_n1107 = ~pb0 & new_n1106;
  assign new_n1108 = ~pc0 & new_n1107;
  assign new_n1109 = ~pk0 & new_n761;
  assign new_n1110 = ~pd0 & new_n1109;
  assign new_n1111 = ~pa0 & new_n1110;
  assign new_n1112 = ~ph0 & new_n1111;
  assign new_n1113 = ~pc & new_n1112;
  assign new_n1114 = ~pg0 & new_n966;
  assign new_n1115 = ~pb0 & new_n1114;
  assign new_n1116 = ~pc0 & new_n1115;
  assign new_n1117 = pa & new_n848;
  assign new_n1118 = ~ph0 & new_n1117;
  assign new_n1119 = ~pc & new_n1118;
  assign new_n1120 = ~pb0 & new_n1119;
  assign new_n1121 = ~pc0 & new_n1120;
  assign new_n1122 = pm & new_n835;
  assign new_n1123 = ~pc0 & new_n1122;
  assign new_n1124 = ~ph0 & new_n1123;
  assign new_n1125 = ~pg0 & new_n843;
  assign new_n1126 = ~pb & new_n1125;
  assign new_n1127 = ~pd0 & new_n1126;
  assign new_n1128 = ~pa0 & new_n877;
  assign new_n1129 = ~pc & new_n1128;
  assign new_n1130 = ~pi0 & new_n1129;
  assign new_n1131 = ~pc0 & new_n1130;
  assign new_n1132 = ~ph0 & new_n1131;
  assign new_n1133 = ~pa0 & new_n937;
  assign new_n1134 = ~pc & new_n1133;
  assign new_n1135 = ~pc0 & new_n1134;
  assign new_n1136 = ~ph0 & new_n1135;
  assign new_n1137 = ~pz & new_n1136;
  assign new_n1138 = ~pb0 & new_n1137;
  assign new_n1139 = ~pc & new_n912;
  assign new_n1140 = ~pb0 & new_n1139;
  assign new_n1141 = ~pc0 & new_n1140;
  assign new_n1142 = pa & new_n796;
  assign new_n1143 = ~ph0 & new_n1142;
  assign new_n1144 = ~pi0 & new_n1143;
  assign new_n1145 = ~pb0 & new_n1144;
  assign new_n1146 = ~pc0 & new_n1145;
  assign new_n1147 = ~pk0 & new_n796;
  assign new_n1148 = ~pa0 & new_n1147;
  assign new_n1149 = ~ph0 & new_n1148;
  assign new_n1150 = ~pi0 & new_n1149;
  assign new_n1151 = ~pb0 & new_n1150;
  assign new_n1152 = ~pc0 & new_n1151;
  assign new_n1153 = ~pa0 & new_n904;
  assign new_n1154 = ~pi0 & new_n1153;
  assign new_n1155 = ~ph0 & new_n1154;
  assign new_n1156 = ~pc & new_n1155;
  assign new_n1157 = ~pb0 & new_n1156;
  assign new_n1158 = ~pc0 & new_n1157;
  assign new_n1159 = pn & new_n821;
  assign new_n1160 = ~pc0 & new_n1159;
  assign new_n1161 = ~ph0 & new_n1160;
  assign new_n1162 = ~pz & new_n1161;
  assign new_n1163 = ~pb0 & new_n1162;
  assign new_n1164 = pa & new_n829;
  assign new_n1165 = ~pc & new_n1164;
  assign new_n1166 = ~pi0 & new_n1165;
  assign new_n1167 = ~pc0 & new_n1166;
  assign new_n1168 = ~ph0 & new_n1167;
  assign new_n1169 = ~pa0 & new_n849;
  assign new_n1170 = ~ph0 & new_n1169;
  assign new_n1171 = ~pc & new_n1170;
  assign new_n1172 = ~pb0 & new_n1171;
  assign new_n1173 = ~pc0 & new_n1172;
  assign new_n1174 = ~pa0 & new_n1109;
  assign new_n1175 = ~pg0 & new_n1174;
  assign new_n1176 = ~ph0 & new_n1175;
  assign new_n1177 = ~pd0 & new_n1176;
  assign new_n1178 = ~pc & new_n944;
  assign new_n1179 = ~pi0 & new_n1178;
  assign new_n1180 = ~pc0 & new_n1179;
  assign new_n1181 = ~ph0 & new_n1180;
  assign new_n1182 = ~pg0 & new_n1118;
  assign new_n1183 = ~pb0 & new_n1182;
  assign new_n1184 = ~pc0 & new_n1183;
  assign new_n1185 = ~pk0 & new_n821;
  assign new_n1186 = ~pa0 & new_n1185;
  assign new_n1187 = ~pc0 & new_n1186;
  assign new_n1188 = ~ph0 & new_n1187;
  assign new_n1189 = ~pz & new_n1188;
  assign new_n1190 = ~pb0 & new_n1189;
  assign new_n1191 = ~pa0 & new_n1055;
  assign new_n1192 = ~pg0 & new_n1191;
  assign new_n1193 = ~pd0 & new_n1192;
  assign new_n1194 = ~pi0 & new_n1193;
  assign new_n1195 = pn & new_n796;
  assign new_n1196 = ~ph0 & new_n1195;
  assign new_n1197 = ~pi0 & new_n1196;
  assign new_n1198 = ~pb0 & new_n1197;
  assign new_n1199 = ~pc0 & new_n1198;
  assign new_n1200 = ~pi0 & new_n1164;
  assign new_n1201 = ~pg0 & new_n1200;
  assign new_n1202 = ~pc0 & new_n1201;
  assign new_n1203 = ~ph0 & new_n1202;
  assign new_n1204 = ~pg0 & new_n809;
  assign new_n1205 = ~ph0 & new_n1204;
  assign new_n1206 = ~pb & new_n1205;
  assign new_n1207 = ~pd0 & new_n842;
  assign new_n1208 = ~pi0 & new_n1207;
  assign new_n1209 = ~pb & new_n1208;
  assign new_n1210 = ~pc & new_n1209;
  assign new_n1211 = ~pd0 & new_n781;
  assign new_n1212 = ~pg0 & new_n1211;
  assign new_n1213 = ~pc0 & new_n1212;
  assign new_n1214 = ~ph0 & new_n1213;
  assign new_n1215 = ~pd0 & new_n813;
  assign new_n1216 = ~pi0 & new_n1215;
  assign new_n1217 = ~ph0 & new_n1216;
  assign new_n1218 = ~pb & new_n1217;
  assign new_n1219 = ~pd0 & new_n1099;
  assign new_n1220 = ~pi0 & new_n1219;
  assign new_n1221 = ~ph0 & new_n1220;
  assign new_n1222 = ~pc & new_n1221;
  assign new_n1223 = ~new_n1218 & ~new_n1222;
  assign new_n1224 = ~new_n1206 & ~new_n1210;
  assign new_n1225 = ~new_n1214 & new_n1224;
  assign new_n1226 = new_n1223 & new_n1225;
  assign new_n1227 = ~new_n1194 & ~new_n1199;
  assign new_n1228 = ~new_n1203 & new_n1227;
  assign new_n1229 = ~new_n1181 & ~new_n1184;
  assign new_n1230 = ~new_n1190 & new_n1229;
  assign new_n1231 = new_n1228 & new_n1230;
  assign new_n1232 = new_n1226 & new_n1231;
  assign new_n1233 = ~new_n1168 & ~new_n1173;
  assign new_n1234 = ~new_n1177 & new_n1233;
  assign new_n1235 = ~new_n1152 & ~new_n1158;
  assign new_n1236 = ~new_n1163 & new_n1235;
  assign new_n1237 = new_n1234 & new_n1236;
  assign new_n1238 = ~new_n1138 & ~new_n1141;
  assign new_n1239 = ~new_n1146 & new_n1238;
  assign new_n1240 = ~new_n1124 & ~new_n1127;
  assign new_n1241 = ~new_n1132 & new_n1240;
  assign new_n1242 = new_n1239 & new_n1241;
  assign new_n1243 = new_n1237 & new_n1242;
  assign new_n1244 = new_n1232 & new_n1243;
  assign new_n1245 = ~new_n1116 & ~new_n1121;
  assign new_n1246 = ~new_n1103 & ~new_n1108;
  assign new_n1247 = ~new_n1113 & new_n1246;
  assign new_n1248 = new_n1245 & new_n1247;
  assign new_n1249 = ~new_n1090 & ~new_n1095;
  assign new_n1250 = ~new_n1098 & new_n1249;
  assign new_n1251 = ~new_n1076 & ~new_n1081;
  assign new_n1252 = ~new_n1086 & new_n1251;
  assign new_n1253 = new_n1250 & new_n1252;
  assign new_n1254 = new_n1248 & new_n1253;
  assign new_n1255 = ~new_n1064 & ~new_n1068;
  assign new_n1256 = ~new_n1073 & new_n1255;
  assign new_n1257 = ~new_n1048 & ~new_n1054;
  assign new_n1258 = ~new_n1059 & new_n1257;
  assign new_n1259 = new_n1256 & new_n1258;
  assign new_n1260 = ~new_n1036 & ~new_n1040;
  assign new_n1261 = ~new_n1045 & new_n1260;
  assign new_n1262 = ~new_n1020 & ~new_n1026;
  assign new_n1263 = ~new_n1031 & new_n1262;
  assign new_n1264 = new_n1261 & new_n1263;
  assign new_n1265 = new_n1259 & new_n1264;
  assign new_n1266 = new_n1254 & new_n1265;
  assign new_n1267 = new_n1244 & new_n1266;
  assign new_n1268 = ~new_n1014 & ~new_n1017;
  assign new_n1269 = ~new_n999 & ~new_n1004;
  assign new_n1270 = ~new_n1009 & new_n1269;
  assign new_n1271 = new_n1268 & new_n1270;
  assign new_n1272 = ~new_n988 & ~new_n991;
  assign new_n1273 = ~new_n994 & new_n1272;
  assign new_n1274 = ~new_n969 & ~new_n974;
  assign new_n1275 = ~new_n979 & new_n1274;
  assign new_n1276 = new_n1273 & new_n1275;
  assign new_n1277 = new_n1271 & new_n1276;
  assign new_n1278 = ~new_n958 & ~new_n961;
  assign new_n1279 = ~new_n964 & new_n1278;
  assign new_n1280 = ~new_n943 & ~new_n948;
  assign new_n1281 = ~new_n953 & new_n1280;
  assign new_n1282 = new_n1279 & new_n1281;
  assign new_n1283 = ~new_n927 & ~new_n930;
  assign new_n1284 = ~new_n933 & new_n1283;
  assign new_n1285 = ~new_n910 & ~new_n915;
  assign new_n1286 = ~new_n920 & new_n1285;
  assign new_n1287 = new_n1284 & new_n1286;
  assign new_n1288 = new_n1282 & new_n1287;
  assign new_n1289 = new_n1277 & new_n1288;
  assign new_n1290 = ~new_n898 & ~new_n902;
  assign new_n1291 = ~new_n882 & ~new_n890;
  assign new_n1292 = ~new_n895 & new_n1291;
  assign new_n1293 = new_n1290 & new_n1292;
  assign new_n1294 = ~new_n846 & ~new_n854;
  assign new_n1295 = ~new_n860 & new_n1294;
  assign new_n1296 = ~new_n869 & ~new_n872;
  assign new_n1297 = ~new_n876 & new_n1296;
  assign new_n1298 = new_n1295 & new_n1297;
  assign new_n1299 = new_n1293 & new_n1298;
  assign new_n1300 = ~new_n785 & ~new_n793;
  assign new_n1301 = ~new_n801 & new_n1300;
  assign new_n1302 = ~new_n765 & ~new_n773;
  assign new_n1303 = ~new_n780 & new_n1302;
  assign new_n1304 = new_n1301 & new_n1303;
  assign new_n1305 = ~new_n808 & ~new_n812;
  assign new_n1306 = ~new_n817 & new_n1305;
  assign new_n1307 = ~new_n826 & ~new_n834;
  assign new_n1308 = ~new_n838 & new_n1307;
  assign new_n1309 = new_n1306 & new_n1308;
  assign new_n1310 = new_n1304 & new_n1309;
  assign new_n1311 = new_n1299 & new_n1310;
  assign new_n1312 = new_n1289 & new_n1311;
  assign ph2 = ~new_n1267 | ~new_n1312;
  assign new_n1314 = pb & pr0;
  assign new_n1315 = pk0 & pm;
  assign new_n1316 = pg0 & pm;
  assign new_n1317 = ph0 & pm;
  assign new_n1318 = pe0 & pm;
  assign new_n1319 = pd0 & ~pv;
  assign new_n1320 = pm & new_n1319;
  assign new_n1321 = ~pv & pp0;
  assign new_n1322 = pm & new_n1321;
  assign new_n1323 = pc0 & ~pv;
  assign new_n1324 = pm & new_n1323;
  assign new_n1325 = pb0 & ~pv;
  assign new_n1326 = pm & new_n1325;
  assign new_n1327 = pa & ~pj;
  assign new_n1328 = pg0 & new_n1327;
  assign new_n1329 = pa & pq0;
  assign new_n1330 = pa & new_n463;
  assign new_n1331 = pa & ps0;
  assign new_n1332 = pa0 & pa;
  assign new_n1333 = pw & new_n1319;
  assign new_n1334 = pd & new_n1333;
  assign new_n1335 = pj0 & pa;
  assign new_n1336 = ps & pl0;
  assign new_n1337 = pr & new_n1336;
  assign new_n1338 = pp0 & pa;
  assign new_n1339 = pr & ps;
  assign new_n1340 = pp0 & new_n1339;
  assign new_n1341 = pk0 & pa;
  assign new_n1342 = pd0 & pa;
  assign new_n1343 = pe0 & pa;
  assign new_n1344 = ph0 & pa;
  assign new_n1345 = pq0 & pm;
  assign new_n1346 = ps0 & pm;
  assign new_n1347 = ~new_n1341 & ~new_n1342;
  assign new_n1348 = ~new_n1343 & new_n1347;
  assign new_n1349 = ~new_n1344 & ~new_n1345;
  assign new_n1350 = ~new_n1346 & new_n1349;
  assign new_n1351 = new_n1348 & new_n1350;
  assign new_n1352 = ~new_n1337 & ~new_n1338;
  assign new_n1353 = ~new_n1340 & new_n1352;
  assign new_n1354 = ~new_n1332 & ~new_n1334;
  assign new_n1355 = ~new_n1335 & new_n1354;
  assign new_n1356 = new_n1353 & new_n1355;
  assign new_n1357 = new_n1351 & new_n1356;
  assign new_n1358 = ~new_n1329 & ~new_n1330;
  assign new_n1359 = ~new_n1331 & new_n1358;
  assign new_n1360 = ~new_n1324 & ~new_n1326;
  assign new_n1361 = ~new_n1328 & new_n1360;
  assign new_n1362 = new_n1359 & new_n1361;
  assign new_n1363 = ~new_n1314 & ~new_n1315;
  assign new_n1364 = ~new_n1316 & ~new_n1317;
  assign new_n1365 = new_n1363 & new_n1364;
  assign new_n1366 = ~new_n1318 & ~new_n1320;
  assign new_n1367 = ~new_n1322 & new_n1366;
  assign new_n1368 = new_n1365 & new_n1367;
  assign new_n1369 = new_n1362 & new_n1368;
  assign pk1 = ~new_n1357 | ~new_n1369;
  assign new_n1371 = pb & pl;
  assign new_n1372 = pg0 & new_n1371;
  assign new_n1373 = ~pa & new_n1372;
  assign new_n1374 = pc & new_n1373;
  assign new_n1375 = pv & new_n1374;
  assign new_n1376 = pk0 & new_n1375;
  assign new_n1377 = ~pm & new_n1376;
  assign new_n1378 = ~pn & new_n1377;
  assign new_n1379 = pl & new_n136;
  assign new_n1380 = ~pa & new_n1379;
  assign new_n1381 = pv & new_n1380;
  assign new_n1382 = pa0 & new_n1381;
  assign new_n1383 = pl & ~pm;
  assign new_n1384 = ~pa & new_n1383;
  assign new_n1385 = pb & new_n1384;
  assign new_n1386 = ~pj & new_n1385;
  assign new_n1387 = pk0 & new_n1386;
  assign new_n1388 = ~pn & new_n1387;
  assign new_n1389 = pv & new_n1388;
  assign new_n1390 = pj & new_n1385;
  assign new_n1391 = ~pn & new_n1390;
  assign new_n1392 = pa0 & new_n1391;
  assign new_n1393 = pd0 & pd;
  assign new_n1394 = pg0 & pj;
  assign new_n1395 = pc & new_n1394;
  assign new_n1396 = pi0 & pi;
  assign new_n1397 = pd0 & ~ph;
  assign new_n1398 = ~new_n1395 & ~new_n1396;
  assign new_n1399 = ~new_n1397 & new_n1398;
  assign new_n1400 = ~new_n1389 & ~new_n1392;
  assign new_n1401 = ~new_n1393 & new_n1400;
  assign new_n1402 = new_n1399 & new_n1401;
  assign new_n1403 = ~pb0 & ~py;
  assign new_n1404 = new_n839 & new_n1403;
  assign new_n1405 = ~pz & ~new_n1378;
  assign new_n1406 = ~new_n1382 & new_n1405;
  assign new_n1407 = new_n1404 & new_n1406;
  assign pi2 = ~new_n1402 | ~new_n1407;
  assign new_n1409 = pd & new_n102;
  assign new_n1410 = ~pe & new_n1409;
  assign new_n1411 = ~pa & new_n1410;
  assign new_n1412 = pd0 & new_n1411;
  assign new_n1413 = ~pv & new_n1412;
  assign new_n1414 = ~pw & new_n1413;
  assign new_n1415 = ~pp & new_n1414;
  assign new_n1416 = ~pu & new_n1415;
  assign new_n1417 = ph0 & pj;
  assign pm1 = new_n1416 | new_n1417;
  assign new_n1419 = pf0 & pb;
  assign new_n1420 = pd0 & pu;
  assign new_n1421 = ph & new_n1420;
  assign new_n1422 = ph0 & pe;
  assign new_n1423 = pw & ph0;
  assign new_n1424 = pu & ph0;
  assign new_n1425 = pe & new_n111;
  assign new_n1426 = ~pa & new_n1425;
  assign new_n1427 = ~ph & new_n1426;
  assign new_n1428 = ~pv & new_n1427;
  assign new_n1429 = pe0 & new_n1428;
  assign new_n1430 = ~pa & pd;
  assign new_n1431 = pu & new_n1430;
  assign new_n1432 = pd0 & new_n1431;
  assign new_n1433 = ~ph & new_n1432;
  assign new_n1434 = ~pv & new_n1433;
  assign new_n1435 = po & new_n1434;
  assign new_n1436 = ~pp & new_n1435;
  assign new_n1437 = pd0 & new_n1430;
  assign new_n1438 = pe & new_n1437;
  assign new_n1439 = ~ph & new_n1438;
  assign new_n1440 = ~pv & new_n1439;
  assign new_n1441 = po & new_n1440;
  assign new_n1442 = ~pp & new_n1441;
  assign new_n1443 = ~pa & ~pd;
  assign new_n1444 = pu & new_n1443;
  assign new_n1445 = pd0 & new_n1444;
  assign new_n1446 = ~ph & new_n1445;
  assign new_n1447 = pp & new_n1446;
  assign new_n1448 = ~pv & new_n1447;
  assign new_n1449 = ~pg & new_n1448;
  assign new_n1450 = po & new_n1449;
  assign new_n1451 = ~pv & ~pg;
  assign new_n1452 = pe & new_n1451;
  assign new_n1453 = ~pa & new_n1452;
  assign new_n1454 = ~ph & new_n1453;
  assign new_n1455 = pe0 & new_n1454;
  assign new_n1456 = ~pg & new_n1433;
  assign new_n1457 = ~pv & new_n1456;
  assign new_n1458 = ~pg & new_n1439;
  assign new_n1459 = ~pv & new_n1458;
  assign new_n1460 = pu & new_n111;
  assign new_n1461 = ~pa & new_n1460;
  assign new_n1462 = ~ph & new_n1461;
  assign new_n1463 = ~pv & new_n1462;
  assign new_n1464 = pe0 & new_n1463;
  assign new_n1465 = pp & pq0;
  assign new_n1466 = pq & new_n1465;
  assign new_n1467 = po & new_n1466;
  assign new_n1468 = pd0 & new_n1443;
  assign new_n1469 = pe & new_n1468;
  assign new_n1470 = ~ph & new_n1469;
  assign new_n1471 = pp & new_n1470;
  assign new_n1472 = ~pv & new_n1471;
  assign new_n1473 = ~pg & new_n1472;
  assign new_n1474 = po & new_n1473;
  assign new_n1475 = pu & new_n1451;
  assign new_n1476 = ~pa & new_n1475;
  assign new_n1477 = ~ph & new_n1476;
  assign new_n1478 = pe0 & new_n1477;
  assign new_n1479 = pp & pp0;
  assign new_n1480 = pq & new_n1479;
  assign new_n1481 = po & new_n1480;
  assign new_n1482 = pe0 & pe;
  assign new_n1483 = ph & new_n1482;
  assign new_n1484 = pa0 & pk;
  assign new_n1485 = pb & new_n1484;
  assign new_n1486 = pd0 & pe;
  assign new_n1487 = ph & new_n1486;
  assign new_n1488 = pe0 & pu;
  assign new_n1489 = ph & new_n1488;
  assign new_n1490 = ~new_n1487 & ~new_n1489;
  assign new_n1491 = ~new_n1481 & ~new_n1483;
  assign new_n1492 = ~new_n1485 & new_n1491;
  assign new_n1493 = new_n1490 & new_n1492;
  assign new_n1494 = ~new_n1474 & ~new_n1478;
  assign new_n1495 = ~new_n1459 & ~new_n1464;
  assign new_n1496 = ~new_n1467 & new_n1495;
  assign new_n1497 = new_n1494 & new_n1496;
  assign new_n1498 = new_n1493 & new_n1497;
  assign new_n1499 = ~new_n1455 & ~new_n1457;
  assign new_n1500 = ~new_n1436 & ~new_n1442;
  assign new_n1501 = ~new_n1450 & new_n1500;
  assign new_n1502 = new_n1499 & new_n1501;
  assign new_n1503 = ~new_n1423 & ~new_n1424;
  assign new_n1504 = ~new_n1429 & new_n1503;
  assign new_n1505 = ~new_n1419 & ~new_n1421;
  assign new_n1506 = ~new_n1422 & new_n1505;
  assign new_n1507 = new_n1504 & new_n1506;
  assign new_n1508 = new_n1502 & new_n1507;
  assign pl1 = ~new_n1498 | ~new_n1508;
  assign new_n1510 = ~pq & pg;
  assign new_n1511 = pi & new_n1510;
  assign new_n1512 = ~pv & new_n1511;
  assign new_n1513 = ~pa & new_n1512;
  assign new_n1514 = pq0 & new_n1513;
  assign new_n1515 = pp0 & pg;
  assign new_n1516 = pi & new_n1515;
  assign new_n1517 = ~pv & new_n1516;
  assign new_n1518 = ~pa & new_n1517;
  assign new_n1519 = ~pp & new_n1518;
  assign new_n1520 = ~pq & new_n1518;
  assign new_n1521 = pi0 & ~ph;
  assign new_n1522 = pi & new_n1521;
  assign new_n1523 = ~pa & new_n1522;
  assign new_n1524 = pq0 & pg;
  assign new_n1525 = pi & new_n1524;
  assign new_n1526 = ~pv & new_n1525;
  assign new_n1527 = ~pa & new_n1526;
  assign new_n1528 = ~po & new_n1527;
  assign new_n1529 = ~pp & new_n1527;
  assign new_n1530 = ~po & new_n1518;
  assign new_n1531 = ~new_n1514 & ~new_n1519;
  assign new_n1532 = ~new_n481 & ~new_n1520;
  assign new_n1533 = new_n1531 & new_n1532;
  assign new_n1534 = ~new_n1529 & ~new_n1530;
  assign new_n1535 = ~new_n1523 & ~new_n1528;
  assign new_n1536 = new_n1534 & new_n1535;
  assign po1 = ~new_n1533 | ~new_n1536;
  assign new_n1538 = ~pu & ~pe;
  assign new_n1539 = ~ph & new_n1538;
  assign new_n1540 = ~pm & new_n1539;
  assign new_n1541 = ~pa & new_n1540;
  assign new_n1542 = ~pw & new_n1541;
  assign new_n1543 = ps0 & new_n1542;
  assign new_n1544 = ~pm & new_n745;
  assign new_n1545 = ~pe & new_n1544;
  assign new_n1546 = ~pa & new_n1545;
  assign new_n1547 = po0 & new_n1546;
  assign new_n1548 = pw0 & new_n1547;
  assign new_n1549 = ~pc & ~ph;
  assign new_n1550 = pj & new_n1549;
  assign new_n1551 = pg0 & new_n1550;
  assign new_n1552 = ~pa & new_n1551;
  assign new_n1553 = ~pm & new_n1552;
  assign new_n1554 = ~pj & new_n1538;
  assign new_n1555 = ~pm & new_n1554;
  assign new_n1556 = ~pa & new_n1555;
  assign new_n1557 = ~pw & new_n1556;
  assign new_n1558 = ph0 & new_n1557;
  assign new_n1559 = pv & pg0;
  assign new_n1560 = pf & new_n1559;
  assign new_n1561 = ~pj & new_n1560;
  assign new_n1562 = ~pa & new_n1561;
  assign new_n1563 = ~pe & ~pm;
  assign new_n1564 = ~pv & new_n1563;
  assign new_n1565 = pc & new_n1564;
  assign new_n1566 = ~pa & new_n1565;
  assign new_n1567 = pp0 & new_n1566;
  assign new_n1568 = ~pg & new_n1567;
  assign new_n1569 = pd & new_n1568;
  assign new_n1570 = ~pu & new_n1569;
  assign new_n1571 = ~pw & new_n1570;
  assign new_n1572 = ~pm & new_n111;
  assign new_n1573 = ~pe & new_n1572;
  assign new_n1574 = ~pa & new_n1573;
  assign new_n1575 = pe0 & new_n1574;
  assign new_n1576 = ~pu & new_n1575;
  assign new_n1577 = ~pw & new_n1576;
  assign new_n1578 = pp & po;
  assign new_n1579 = ~pm & new_n1578;
  assign new_n1580 = ~pe & new_n1579;
  assign new_n1581 = ~pa & new_n1580;
  assign new_n1582 = pq0 & new_n1581;
  assign new_n1583 = ~pg & new_n1582;
  assign new_n1584 = ~pq & new_n1583;
  assign new_n1585 = ~pu & new_n1584;
  assign new_n1586 = ~pw & new_n1585;
  assign new_n1587 = ~new_n1543 & ~new_n1548;
  assign new_n1588 = ~new_n1553 & ~new_n1558;
  assign new_n1589 = new_n1587 & new_n1588;
  assign new_n1590 = ~new_n1577 & ~new_n1586;
  assign new_n1591 = ~new_n1562 & ~new_n1571;
  assign new_n1592 = new_n1590 & new_n1591;
  assign pn1 = ~new_n1589 | ~new_n1592;
  assign new_n1594 = pr & ~pm;
  assign new_n1595 = pb & new_n1594;
  assign new_n1596 = ~pj & new_n1595;
  assign new_n1597 = ~pa & new_n1596;
  assign new_n1598 = pk0 & new_n1597;
  assign new_n1599 = ~ps & new_n1598;
  assign new_n1600 = ~pv & new_n1599;
  assign new_n1601 = pa0 & new_n1597;
  assign new_n1602 = ~pk & new_n1601;
  assign new_n1603 = pl & new_n1602;
  assign new_n1604 = ~ps & new_n1603;
  assign new_n1605 = ~pv & new_n1604;
  assign new_n1606 = ~pi & new_n1521;
  assign new_n1607 = ~pa & new_n1606;
  assign new_n1608 = ~pt & pi0;
  assign new_n1609 = ~ph & new_n1608;
  assign new_n1610 = ~pi & new_n1609;
  assign new_n1611 = pa & new_n1610;
  assign new_n1612 = pj0 & ~pa;
  assign new_n1613 = ~new_n1611 & ~new_n1612;
  assign new_n1614 = ~new_n1600 & ~new_n1605;
  assign new_n1615 = ~new_n1607 & new_n1614;
  assign pr1 = ~new_n1613 | ~new_n1615;
  assign new_n1617 = ps & pk0;
  assign new_n1618 = pr & new_n1617;
  assign new_n1619 = pa0 & ps;
  assign new_n1620 = pr & new_n1619;
  assign pw1 = new_n1618 | new_n1620;
  assign new_n1622 = ~pj & new_n1559;
  assign new_n1623 = ~pm & new_n1622;
  assign new_n1624 = ~pa & new_n1623;
  assign new_n1625 = ~pf & new_n1624;
  assign new_n1626 = pv & pn;
  assign new_n1627 = ~pj & new_n1626;
  assign new_n1628 = ~pm & new_n1627;
  assign new_n1629 = ~pa & new_n1628;
  assign new_n1630 = pk0 & new_n1629;
  assign new_n1631 = ~pv & pk0;
  assign new_n1632 = ~pj & new_n1631;
  assign new_n1633 = ~pm & new_n1632;
  assign new_n1634 = ~pa & new_n1633;
  assign new_n1635 = ~pr & new_n1634;
  assign new_n1636 = ~pv & pg0;
  assign new_n1637 = ~pj & new_n1636;
  assign new_n1638 = ~pm & new_n1637;
  assign new_n1639 = ~pa & new_n1638;
  assign new_n1640 = ~new_n1625 & ~new_n1630;
  assign new_n1641 = ~new_n1635 & ~new_n1639;
  assign pv1 = ~new_n1640 | ~new_n1641;
  assign new_n1643 = ~pg0 & ~pr0;
  assign new_n1644 = ~ph0 & new_n1643;
  assign new_n1645 = ~pf0 & new_n1644;
  assign new_n1646 = ~pz & new_n1645;
  assign new_n1647 = ~ph0 & ~pz;
  assign new_n1648 = pj & new_n1647;
  assign py1 = new_n1646 | new_n1648;
  assign new_n1650 = pf0 & ~pj;
  assign new_n1651 = pr0 & ~pj;
  assign new_n1652 = pg0 & ~pj;
  assign new_n1653 = ~pz & ~new_n1652;
  assign new_n1654 = ~new_n1650 & ~new_n1651;
  assign new_n1655 = ~ph0 & new_n1654;
  assign px1 = ~new_n1653 | ~new_n1655;
  assign pz1 = pc0 | pd0;
  assign pc2 = ph0;
  assign pi1 = pm0;
  assign pj1 = pn0;
  assign pq1 = pz;
  assign pp1 = py;
  assign pu1 = py0;
  assign pt1 = px0;
endmodule


