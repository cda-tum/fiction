// Benchmark "top" written by ABC on Mon Nov 27 16:57:47 2023

module top ( 
    a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15,
    a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29,
    a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43,
    a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57,
    a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71,
    a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85,
    a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99,
    a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111,
    a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123,
    a124, a125, a126, a127, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10,
    b11, b12, b13, b14, b15, b16, b17, b18, b19, b20, b21, b22, b23, b24,
    b25, b26, b27, b28, b29, b30, b31, b32, b33, b34, b35, b36, b37, b38,
    b39, b40, b41, b42, b43, b44, b45, b46, b47, b48, b49, b50, b51, b52,
    b53, b54, b55, b56, b57, b58, b59, b60, b61, b62, b63, b64, b65, b66,
    b67, b68, b69, b70, b71, b72, b73, b74, b75, b76, b77, b78, b79, b80,
    b81, b82, b83, b84, b85, b86, b87, b88, b89, b90, b91, b92, b93, b94,
    b95, b96, b97, b98, b99, b100, b101, b102, b103, b104, b105, b106,
    b107, b108, b109, b110, b111, b112, b113, b114, b115, b116, b117, b118,
    b119, b120, b121, b122, b123, b124, b125, b126, b127,
    f0, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26, f27, f28, f29,
    f30, f31, f32, f33, f34, f35, f36, f37, f38, f39, f40, f41, f42, f43,
    f44, f45, f46, f47, f48, f49, f50, f51, f52, f53, f54, f55, f56, f57,
    f58, f59, f60, f61, f62, f63, f64, f65, f66, f67, f68, f69, f70, f71,
    f72, f73, f74, f75, f76, f77, f78, f79, f80, f81, f82, f83, f84, f85,
    f86, f87, f88, f89, f90, f91, f92, f93, f94, f95, f96, f97, f98, f99,
    f100, f101, f102, f103, f104, f105, f106, f107, f108, f109, f110, f111,
    f112, f113, f114, f115, f116, f117, f118, f119, f120, f121, f122, f123,
    f124, f125, f126, f127, cOut  );
  input  a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14,
    a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28,
    a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42,
    a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56,
    a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70,
    a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84,
    a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98,
    a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110,
    a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122,
    a123, a124, a125, a126, a127, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9,
    b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b20, b21, b22, b23,
    b24, b25, b26, b27, b28, b29, b30, b31, b32, b33, b34, b35, b36, b37,
    b38, b39, b40, b41, b42, b43, b44, b45, b46, b47, b48, b49, b50, b51,
    b52, b53, b54, b55, b56, b57, b58, b59, b60, b61, b62, b63, b64, b65,
    b66, b67, b68, b69, b70, b71, b72, b73, b74, b75, b76, b77, b78, b79,
    b80, b81, b82, b83, b84, b85, b86, b87, b88, b89, b90, b91, b92, b93,
    b94, b95, b96, b97, b98, b99, b100, b101, b102, b103, b104, b105, b106,
    b107, b108, b109, b110, b111, b112, b113, b114, b115, b116, b117, b118,
    b119, b120, b121, b122, b123, b124, b125, b126, b127;
  output f0, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15,
    f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26, f27, f28, f29,
    f30, f31, f32, f33, f34, f35, f36, f37, f38, f39, f40, f41, f42, f43,
    f44, f45, f46, f47, f48, f49, f50, f51, f52, f53, f54, f55, f56, f57,
    f58, f59, f60, f61, f62, f63, f64, f65, f66, f67, f68, f69, f70, f71,
    f72, f73, f74, f75, f76, f77, f78, f79, f80, f81, f82, f83, f84, f85,
    f86, f87, f88, f89, f90, f91, f92, f93, f94, f95, f96, f97, f98, f99,
    f100, f101, f102, f103, f104, f105, f106, f107, f108, f109, f110, f111,
    f112, f113, f114, f115, f116, f117, f118, f119, f120, f121, f122, f123,
    f124, f125, f126, f127, cOut;
  wire new_n386, new_n387, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n430, new_n431, new_n432, new_n433, new_n434,
    new_n435, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275;
  assign new_n386 = a0 & b0;
  assign new_n387 = ~a0 & ~b0;
  assign f0 = ~new_n386 & ~new_n387;
  assign new_n389 = a1 & b1;
  assign new_n390 = ~a1 & ~b1;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = new_n386 & ~new_n391;
  assign new_n393 = ~new_n386 & new_n391;
  assign f1 = new_n392 | new_n393;
  assign new_n395 = ~new_n390 & ~new_n393;
  assign new_n396 = a2 & b2;
  assign new_n397 = ~a2 & ~b2;
  assign new_n398 = ~new_n396 & ~new_n397;
  assign new_n399 = new_n395 & new_n398;
  assign new_n400 = ~new_n395 & ~new_n398;
  assign f2 = ~new_n399 & ~new_n400;
  assign new_n402 = ~new_n396 & ~new_n399;
  assign new_n403 = a3 & b3;
  assign new_n404 = ~a3 & ~b3;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = ~new_n402 & new_n405;
  assign new_n407 = new_n402 & ~new_n405;
  assign f3 = ~new_n406 & ~new_n407;
  assign new_n409 = ~new_n403 & ~new_n406;
  assign new_n410 = a4 & b4;
  assign new_n411 = ~a4 & ~b4;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign new_n413 = new_n409 & new_n412;
  assign new_n414 = ~new_n409 & ~new_n412;
  assign f4 = new_n413 | new_n414;
  assign new_n416 = ~new_n411 & ~new_n413;
  assign new_n417 = a5 & b5;
  assign new_n418 = ~a5 & ~b5;
  assign new_n419 = ~new_n417 & ~new_n418;
  assign new_n420 = ~new_n416 & new_n419;
  assign new_n421 = new_n416 & ~new_n419;
  assign f5 = new_n420 | new_n421;
  assign new_n423 = ~new_n418 & ~new_n420;
  assign new_n424 = a6 & b6;
  assign new_n425 = ~a6 & ~b6;
  assign new_n426 = ~new_n424 & ~new_n425;
  assign new_n427 = ~new_n423 & new_n426;
  assign new_n428 = new_n423 & ~new_n426;
  assign f6 = new_n427 | new_n428;
  assign new_n430 = ~new_n425 & ~new_n427;
  assign new_n431 = a7 & b7;
  assign new_n432 = ~a7 & ~b7;
  assign new_n433 = ~new_n431 & ~new_n432;
  assign new_n434 = ~new_n430 & new_n433;
  assign new_n435 = new_n430 & ~new_n433;
  assign f7 = new_n434 | new_n435;
  assign new_n437 = ~new_n432 & ~new_n434;
  assign new_n438 = a8 & b8;
  assign new_n439 = ~a8 & ~b8;
  assign new_n440 = ~new_n438 & ~new_n439;
  assign new_n441 = ~new_n437 & new_n440;
  assign new_n442 = new_n437 & ~new_n440;
  assign f8 = new_n441 | new_n442;
  assign new_n444 = ~new_n439 & ~new_n441;
  assign new_n445 = a9 & b9;
  assign new_n446 = ~a9 & ~b9;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign new_n448 = ~new_n444 & new_n447;
  assign new_n449 = new_n444 & ~new_n447;
  assign f9 = new_n448 | new_n449;
  assign new_n451 = ~new_n446 & ~new_n448;
  assign new_n452 = a10 & b10;
  assign new_n453 = ~a10 & ~b10;
  assign new_n454 = ~new_n452 & ~new_n453;
  assign new_n455 = ~new_n451 & new_n454;
  assign new_n456 = new_n451 & ~new_n454;
  assign f10 = new_n455 | new_n456;
  assign new_n458 = ~new_n453 & ~new_n455;
  assign new_n459 = a11 & b11;
  assign new_n460 = ~a11 & ~b11;
  assign new_n461 = ~new_n459 & ~new_n460;
  assign new_n462 = ~new_n458 & new_n461;
  assign new_n463 = new_n458 & ~new_n461;
  assign f11 = new_n462 | new_n463;
  assign new_n465 = ~new_n460 & ~new_n462;
  assign new_n466 = a12 & b12;
  assign new_n467 = ~a12 & ~b12;
  assign new_n468 = ~new_n466 & ~new_n467;
  assign new_n469 = ~new_n465 & new_n468;
  assign new_n470 = new_n465 & ~new_n468;
  assign f12 = new_n469 | new_n470;
  assign new_n472 = ~new_n467 & ~new_n469;
  assign new_n473 = a13 & b13;
  assign new_n474 = ~a13 & ~b13;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = ~new_n472 & new_n475;
  assign new_n477 = new_n472 & ~new_n475;
  assign f13 = new_n476 | new_n477;
  assign new_n479 = ~new_n474 & ~new_n476;
  assign new_n480 = a14 & b14;
  assign new_n481 = ~a14 & ~b14;
  assign new_n482 = ~new_n480 & ~new_n481;
  assign new_n483 = ~new_n479 & new_n482;
  assign new_n484 = new_n479 & ~new_n482;
  assign f14 = new_n483 | new_n484;
  assign new_n486 = ~new_n481 & ~new_n483;
  assign new_n487 = a15 & b15;
  assign new_n488 = ~a15 & ~b15;
  assign new_n489 = ~new_n487 & ~new_n488;
  assign new_n490 = ~new_n486 & new_n489;
  assign new_n491 = new_n486 & ~new_n489;
  assign f15 = new_n490 | new_n491;
  assign new_n493 = ~new_n488 & ~new_n490;
  assign new_n494 = a16 & b16;
  assign new_n495 = ~a16 & ~b16;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = ~new_n493 & new_n496;
  assign new_n498 = new_n493 & ~new_n496;
  assign f16 = new_n497 | new_n498;
  assign new_n500 = ~new_n495 & ~new_n497;
  assign new_n501 = a17 & b17;
  assign new_n502 = ~a17 & ~b17;
  assign new_n503 = ~new_n501 & ~new_n502;
  assign new_n504 = ~new_n500 & new_n503;
  assign new_n505 = new_n500 & ~new_n503;
  assign f17 = new_n504 | new_n505;
  assign new_n507 = ~new_n502 & ~new_n504;
  assign new_n508 = a18 & b18;
  assign new_n509 = ~a18 & ~b18;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = ~new_n507 & new_n510;
  assign new_n512 = new_n507 & ~new_n510;
  assign f18 = new_n511 | new_n512;
  assign new_n514 = ~new_n509 & ~new_n511;
  assign new_n515 = a19 & b19;
  assign new_n516 = ~a19 & ~b19;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = ~new_n514 & new_n517;
  assign new_n519 = new_n514 & ~new_n517;
  assign f19 = new_n518 | new_n519;
  assign new_n521 = ~new_n516 & ~new_n518;
  assign new_n522 = a20 & b20;
  assign new_n523 = ~a20 & ~b20;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = ~new_n521 & new_n524;
  assign new_n526 = new_n521 & ~new_n524;
  assign f20 = new_n525 | new_n526;
  assign new_n528 = ~new_n523 & ~new_n525;
  assign new_n529 = a21 & b21;
  assign new_n530 = ~a21 & ~b21;
  assign new_n531 = ~new_n529 & ~new_n530;
  assign new_n532 = ~new_n528 & new_n531;
  assign new_n533 = new_n528 & ~new_n531;
  assign f21 = new_n532 | new_n533;
  assign new_n535 = ~new_n530 & ~new_n532;
  assign new_n536 = a22 & b22;
  assign new_n537 = ~a22 & ~b22;
  assign new_n538 = ~new_n536 & ~new_n537;
  assign new_n539 = ~new_n535 & new_n538;
  assign new_n540 = new_n535 & ~new_n538;
  assign f22 = new_n539 | new_n540;
  assign new_n542 = ~new_n537 & ~new_n539;
  assign new_n543 = a23 & b23;
  assign new_n544 = ~a23 & ~b23;
  assign new_n545 = ~new_n543 & ~new_n544;
  assign new_n546 = ~new_n542 & new_n545;
  assign new_n547 = new_n542 & ~new_n545;
  assign f23 = new_n546 | new_n547;
  assign new_n549 = ~new_n544 & ~new_n546;
  assign new_n550 = a24 & b24;
  assign new_n551 = ~a24 & ~b24;
  assign new_n552 = ~new_n550 & ~new_n551;
  assign new_n553 = ~new_n549 & new_n552;
  assign new_n554 = new_n549 & ~new_n552;
  assign f24 = new_n553 | new_n554;
  assign new_n556 = ~new_n551 & ~new_n553;
  assign new_n557 = a25 & b25;
  assign new_n558 = ~a25 & ~b25;
  assign new_n559 = ~new_n557 & ~new_n558;
  assign new_n560 = ~new_n556 & new_n559;
  assign new_n561 = new_n556 & ~new_n559;
  assign f25 = new_n560 | new_n561;
  assign new_n563 = ~new_n558 & ~new_n560;
  assign new_n564 = a26 & b26;
  assign new_n565 = ~a26 & ~b26;
  assign new_n566 = ~new_n564 & ~new_n565;
  assign new_n567 = ~new_n563 & new_n566;
  assign new_n568 = new_n563 & ~new_n566;
  assign f26 = new_n567 | new_n568;
  assign new_n570 = ~new_n565 & ~new_n567;
  assign new_n571 = a27 & b27;
  assign new_n572 = ~a27 & ~b27;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = ~new_n570 & new_n573;
  assign new_n575 = new_n570 & ~new_n573;
  assign f27 = new_n574 | new_n575;
  assign new_n577 = ~new_n572 & ~new_n574;
  assign new_n578 = a28 & b28;
  assign new_n579 = ~a28 & ~b28;
  assign new_n580 = ~new_n578 & ~new_n579;
  assign new_n581 = ~new_n577 & new_n580;
  assign new_n582 = new_n577 & ~new_n580;
  assign f28 = new_n581 | new_n582;
  assign new_n584 = ~new_n579 & ~new_n581;
  assign new_n585 = a29 & b29;
  assign new_n586 = ~a29 & ~b29;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = ~new_n584 & new_n587;
  assign new_n589 = new_n584 & ~new_n587;
  assign f29 = new_n588 | new_n589;
  assign new_n591 = ~new_n586 & ~new_n588;
  assign new_n592 = a30 & b30;
  assign new_n593 = ~a30 & ~b30;
  assign new_n594 = ~new_n592 & ~new_n593;
  assign new_n595 = ~new_n591 & new_n594;
  assign new_n596 = new_n591 & ~new_n594;
  assign f30 = new_n595 | new_n596;
  assign new_n598 = ~new_n593 & ~new_n595;
  assign new_n599 = a31 & b31;
  assign new_n600 = ~a31 & ~b31;
  assign new_n601 = ~new_n599 & ~new_n600;
  assign new_n602 = ~new_n598 & new_n601;
  assign new_n603 = new_n598 & ~new_n601;
  assign f31 = new_n602 | new_n603;
  assign new_n605 = ~new_n600 & ~new_n602;
  assign new_n606 = a32 & b32;
  assign new_n607 = ~a32 & ~b32;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = ~new_n605 & new_n608;
  assign new_n610 = new_n605 & ~new_n608;
  assign f32 = new_n609 | new_n610;
  assign new_n612 = ~new_n607 & ~new_n609;
  assign new_n613 = a33 & b33;
  assign new_n614 = ~a33 & ~b33;
  assign new_n615 = ~new_n613 & ~new_n614;
  assign new_n616 = ~new_n612 & new_n615;
  assign new_n617 = new_n612 & ~new_n615;
  assign f33 = new_n616 | new_n617;
  assign new_n619 = ~new_n614 & ~new_n616;
  assign new_n620 = a34 & b34;
  assign new_n621 = ~a34 & ~b34;
  assign new_n622 = ~new_n620 & ~new_n621;
  assign new_n623 = ~new_n619 & new_n622;
  assign new_n624 = new_n619 & ~new_n622;
  assign f34 = new_n623 | new_n624;
  assign new_n626 = ~new_n621 & ~new_n623;
  assign new_n627 = a35 & b35;
  assign new_n628 = ~a35 & ~b35;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = ~new_n626 & new_n629;
  assign new_n631 = new_n626 & ~new_n629;
  assign f35 = new_n630 | new_n631;
  assign new_n633 = ~new_n628 & ~new_n630;
  assign new_n634 = a36 & b36;
  assign new_n635 = ~a36 & ~b36;
  assign new_n636 = ~new_n634 & ~new_n635;
  assign new_n637 = ~new_n633 & new_n636;
  assign new_n638 = new_n633 & ~new_n636;
  assign f36 = new_n637 | new_n638;
  assign new_n640 = ~new_n635 & ~new_n637;
  assign new_n641 = a37 & b37;
  assign new_n642 = ~a37 & ~b37;
  assign new_n643 = ~new_n641 & ~new_n642;
  assign new_n644 = ~new_n640 & new_n643;
  assign new_n645 = new_n640 & ~new_n643;
  assign f37 = new_n644 | new_n645;
  assign new_n647 = ~new_n642 & ~new_n644;
  assign new_n648 = a38 & b38;
  assign new_n649 = ~a38 & ~b38;
  assign new_n650 = ~new_n648 & ~new_n649;
  assign new_n651 = ~new_n647 & new_n650;
  assign new_n652 = new_n647 & ~new_n650;
  assign f38 = new_n651 | new_n652;
  assign new_n654 = ~new_n649 & ~new_n651;
  assign new_n655 = a39 & b39;
  assign new_n656 = ~a39 & ~b39;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign new_n658 = ~new_n654 & new_n657;
  assign new_n659 = new_n654 & ~new_n657;
  assign f39 = new_n658 | new_n659;
  assign new_n661 = ~new_n656 & ~new_n658;
  assign new_n662 = a40 & b40;
  assign new_n663 = ~a40 & ~b40;
  assign new_n664 = ~new_n662 & ~new_n663;
  assign new_n665 = ~new_n661 & new_n664;
  assign new_n666 = new_n661 & ~new_n664;
  assign f40 = new_n665 | new_n666;
  assign new_n668 = ~new_n663 & ~new_n665;
  assign new_n669 = a41 & b41;
  assign new_n670 = ~a41 & ~b41;
  assign new_n671 = ~new_n669 & ~new_n670;
  assign new_n672 = ~new_n668 & new_n671;
  assign new_n673 = new_n668 & ~new_n671;
  assign f41 = new_n672 | new_n673;
  assign new_n675 = ~new_n670 & ~new_n672;
  assign new_n676 = a42 & b42;
  assign new_n677 = ~a42 & ~b42;
  assign new_n678 = ~new_n676 & ~new_n677;
  assign new_n679 = ~new_n675 & new_n678;
  assign new_n680 = new_n675 & ~new_n678;
  assign f42 = new_n679 | new_n680;
  assign new_n682 = ~new_n677 & ~new_n679;
  assign new_n683 = a43 & b43;
  assign new_n684 = ~a43 & ~b43;
  assign new_n685 = ~new_n683 & ~new_n684;
  assign new_n686 = ~new_n682 & new_n685;
  assign new_n687 = new_n682 & ~new_n685;
  assign f43 = new_n686 | new_n687;
  assign new_n689 = ~new_n684 & ~new_n686;
  assign new_n690 = a44 & b44;
  assign new_n691 = ~a44 & ~b44;
  assign new_n692 = ~new_n690 & ~new_n691;
  assign new_n693 = ~new_n689 & new_n692;
  assign new_n694 = new_n689 & ~new_n692;
  assign f44 = new_n693 | new_n694;
  assign new_n696 = ~new_n691 & ~new_n693;
  assign new_n697 = a45 & b45;
  assign new_n698 = ~a45 & ~b45;
  assign new_n699 = ~new_n697 & ~new_n698;
  assign new_n700 = ~new_n696 & new_n699;
  assign new_n701 = new_n696 & ~new_n699;
  assign f45 = new_n700 | new_n701;
  assign new_n703 = ~new_n698 & ~new_n700;
  assign new_n704 = a46 & b46;
  assign new_n705 = ~a46 & ~b46;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = ~new_n703 & new_n706;
  assign new_n708 = new_n703 & ~new_n706;
  assign f46 = new_n707 | new_n708;
  assign new_n710 = ~new_n705 & ~new_n707;
  assign new_n711 = a47 & b47;
  assign new_n712 = ~a47 & ~b47;
  assign new_n713 = ~new_n711 & ~new_n712;
  assign new_n714 = ~new_n710 & new_n713;
  assign new_n715 = new_n710 & ~new_n713;
  assign f47 = new_n714 | new_n715;
  assign new_n717 = ~new_n712 & ~new_n714;
  assign new_n718 = a48 & b48;
  assign new_n719 = ~a48 & ~b48;
  assign new_n720 = ~new_n718 & ~new_n719;
  assign new_n721 = ~new_n717 & new_n720;
  assign new_n722 = new_n717 & ~new_n720;
  assign f48 = new_n721 | new_n722;
  assign new_n724 = ~new_n719 & ~new_n721;
  assign new_n725 = a49 & b49;
  assign new_n726 = ~a49 & ~b49;
  assign new_n727 = ~new_n725 & ~new_n726;
  assign new_n728 = ~new_n724 & new_n727;
  assign new_n729 = new_n724 & ~new_n727;
  assign f49 = new_n728 | new_n729;
  assign new_n731 = ~new_n726 & ~new_n728;
  assign new_n732 = a50 & b50;
  assign new_n733 = ~a50 & ~b50;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = ~new_n731 & new_n734;
  assign new_n736 = new_n731 & ~new_n734;
  assign f50 = new_n735 | new_n736;
  assign new_n738 = ~new_n733 & ~new_n735;
  assign new_n739 = a51 & b51;
  assign new_n740 = ~a51 & ~b51;
  assign new_n741 = ~new_n739 & ~new_n740;
  assign new_n742 = ~new_n738 & new_n741;
  assign new_n743 = new_n738 & ~new_n741;
  assign f51 = new_n742 | new_n743;
  assign new_n745 = ~new_n740 & ~new_n742;
  assign new_n746 = a52 & b52;
  assign new_n747 = ~a52 & ~b52;
  assign new_n748 = ~new_n746 & ~new_n747;
  assign new_n749 = ~new_n745 & new_n748;
  assign new_n750 = new_n745 & ~new_n748;
  assign f52 = new_n749 | new_n750;
  assign new_n752 = ~new_n747 & ~new_n749;
  assign new_n753 = a53 & b53;
  assign new_n754 = ~a53 & ~b53;
  assign new_n755 = ~new_n753 & ~new_n754;
  assign new_n756 = ~new_n752 & new_n755;
  assign new_n757 = new_n752 & ~new_n755;
  assign f53 = new_n756 | new_n757;
  assign new_n759 = ~new_n754 & ~new_n756;
  assign new_n760 = a54 & b54;
  assign new_n761 = ~a54 & ~b54;
  assign new_n762 = ~new_n760 & ~new_n761;
  assign new_n763 = ~new_n759 & new_n762;
  assign new_n764 = new_n759 & ~new_n762;
  assign f54 = new_n763 | new_n764;
  assign new_n766 = ~new_n761 & ~new_n763;
  assign new_n767 = a55 & b55;
  assign new_n768 = ~a55 & ~b55;
  assign new_n769 = ~new_n767 & ~new_n768;
  assign new_n770 = ~new_n766 & new_n769;
  assign new_n771 = new_n766 & ~new_n769;
  assign f55 = new_n770 | new_n771;
  assign new_n773 = ~new_n768 & ~new_n770;
  assign new_n774 = a56 & b56;
  assign new_n775 = ~a56 & ~b56;
  assign new_n776 = ~new_n774 & ~new_n775;
  assign new_n777 = ~new_n773 & new_n776;
  assign new_n778 = new_n773 & ~new_n776;
  assign f56 = new_n777 | new_n778;
  assign new_n780 = ~new_n775 & ~new_n777;
  assign new_n781 = a57 & b57;
  assign new_n782 = ~a57 & ~b57;
  assign new_n783 = ~new_n781 & ~new_n782;
  assign new_n784 = ~new_n780 & new_n783;
  assign new_n785 = new_n780 & ~new_n783;
  assign f57 = new_n784 | new_n785;
  assign new_n787 = ~new_n782 & ~new_n784;
  assign new_n788 = a58 & b58;
  assign new_n789 = ~a58 & ~b58;
  assign new_n790 = ~new_n788 & ~new_n789;
  assign new_n791 = ~new_n787 & new_n790;
  assign new_n792 = new_n787 & ~new_n790;
  assign f58 = new_n791 | new_n792;
  assign new_n794 = ~new_n789 & ~new_n791;
  assign new_n795 = a59 & b59;
  assign new_n796 = ~a59 & ~b59;
  assign new_n797 = ~new_n795 & ~new_n796;
  assign new_n798 = ~new_n794 & new_n797;
  assign new_n799 = new_n794 & ~new_n797;
  assign f59 = new_n798 | new_n799;
  assign new_n801 = ~new_n796 & ~new_n798;
  assign new_n802 = a60 & b60;
  assign new_n803 = ~a60 & ~b60;
  assign new_n804 = ~new_n802 & ~new_n803;
  assign new_n805 = ~new_n801 & new_n804;
  assign new_n806 = new_n801 & ~new_n804;
  assign f60 = new_n805 | new_n806;
  assign new_n808 = ~new_n803 & ~new_n805;
  assign new_n809 = a61 & b61;
  assign new_n810 = ~a61 & ~b61;
  assign new_n811 = ~new_n809 & ~new_n810;
  assign new_n812 = ~new_n808 & new_n811;
  assign new_n813 = new_n808 & ~new_n811;
  assign f61 = new_n812 | new_n813;
  assign new_n815 = ~new_n810 & ~new_n812;
  assign new_n816 = a62 & b62;
  assign new_n817 = ~a62 & ~b62;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = ~new_n815 & new_n818;
  assign new_n820 = new_n815 & ~new_n818;
  assign f62 = new_n819 | new_n820;
  assign new_n822 = ~new_n817 & ~new_n819;
  assign new_n823 = a63 & b63;
  assign new_n824 = ~a63 & ~b63;
  assign new_n825 = ~new_n823 & ~new_n824;
  assign new_n826 = ~new_n822 & new_n825;
  assign new_n827 = new_n822 & ~new_n825;
  assign f63 = new_n826 | new_n827;
  assign new_n829 = ~new_n824 & ~new_n826;
  assign new_n830 = a64 & b64;
  assign new_n831 = ~a64 & ~b64;
  assign new_n832 = ~new_n830 & ~new_n831;
  assign new_n833 = ~new_n829 & new_n832;
  assign new_n834 = new_n829 & ~new_n832;
  assign f64 = new_n833 | new_n834;
  assign new_n836 = ~new_n831 & ~new_n833;
  assign new_n837 = a65 & b65;
  assign new_n838 = ~a65 & ~b65;
  assign new_n839 = ~new_n837 & ~new_n838;
  assign new_n840 = ~new_n836 & new_n839;
  assign new_n841 = new_n836 & ~new_n839;
  assign f65 = new_n840 | new_n841;
  assign new_n843 = ~new_n838 & ~new_n840;
  assign new_n844 = a66 & b66;
  assign new_n845 = ~a66 & ~b66;
  assign new_n846 = ~new_n844 & ~new_n845;
  assign new_n847 = ~new_n843 & new_n846;
  assign new_n848 = new_n843 & ~new_n846;
  assign f66 = new_n847 | new_n848;
  assign new_n850 = ~new_n845 & ~new_n847;
  assign new_n851 = a67 & b67;
  assign new_n852 = ~a67 & ~b67;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = ~new_n850 & new_n853;
  assign new_n855 = new_n850 & ~new_n853;
  assign f67 = new_n854 | new_n855;
  assign new_n857 = ~new_n852 & ~new_n854;
  assign new_n858 = a68 & b68;
  assign new_n859 = ~a68 & ~b68;
  assign new_n860 = ~new_n858 & ~new_n859;
  assign new_n861 = ~new_n857 & new_n860;
  assign new_n862 = new_n857 & ~new_n860;
  assign f68 = new_n861 | new_n862;
  assign new_n864 = ~new_n859 & ~new_n861;
  assign new_n865 = a69 & b69;
  assign new_n866 = ~a69 & ~b69;
  assign new_n867 = ~new_n865 & ~new_n866;
  assign new_n868 = ~new_n864 & new_n867;
  assign new_n869 = new_n864 & ~new_n867;
  assign f69 = new_n868 | new_n869;
  assign new_n871 = ~new_n866 & ~new_n868;
  assign new_n872 = a70 & b70;
  assign new_n873 = ~a70 & ~b70;
  assign new_n874 = ~new_n872 & ~new_n873;
  assign new_n875 = ~new_n871 & new_n874;
  assign new_n876 = new_n871 & ~new_n874;
  assign f70 = new_n875 | new_n876;
  assign new_n878 = ~new_n873 & ~new_n875;
  assign new_n879 = a71 & b71;
  assign new_n880 = ~a71 & ~b71;
  assign new_n881 = ~new_n879 & ~new_n880;
  assign new_n882 = ~new_n878 & new_n881;
  assign new_n883 = new_n878 & ~new_n881;
  assign f71 = new_n882 | new_n883;
  assign new_n885 = ~new_n880 & ~new_n882;
  assign new_n886 = a72 & b72;
  assign new_n887 = ~a72 & ~b72;
  assign new_n888 = ~new_n886 & ~new_n887;
  assign new_n889 = ~new_n885 & new_n888;
  assign new_n890 = new_n885 & ~new_n888;
  assign f72 = new_n889 | new_n890;
  assign new_n892 = ~new_n887 & ~new_n889;
  assign new_n893 = a73 & b73;
  assign new_n894 = ~a73 & ~b73;
  assign new_n895 = ~new_n893 & ~new_n894;
  assign new_n896 = ~new_n892 & new_n895;
  assign new_n897 = new_n892 & ~new_n895;
  assign f73 = new_n896 | new_n897;
  assign new_n899 = ~new_n894 & ~new_n896;
  assign new_n900 = a74 & b74;
  assign new_n901 = ~a74 & ~b74;
  assign new_n902 = ~new_n900 & ~new_n901;
  assign new_n903 = ~new_n899 & new_n902;
  assign new_n904 = new_n899 & ~new_n902;
  assign f74 = new_n903 | new_n904;
  assign new_n906 = ~new_n901 & ~new_n903;
  assign new_n907 = a75 & b75;
  assign new_n908 = ~a75 & ~b75;
  assign new_n909 = ~new_n907 & ~new_n908;
  assign new_n910 = ~new_n906 & new_n909;
  assign new_n911 = new_n906 & ~new_n909;
  assign f75 = new_n910 | new_n911;
  assign new_n913 = ~new_n908 & ~new_n910;
  assign new_n914 = a76 & b76;
  assign new_n915 = ~a76 & ~b76;
  assign new_n916 = ~new_n914 & ~new_n915;
  assign new_n917 = ~new_n913 & new_n916;
  assign new_n918 = new_n913 & ~new_n916;
  assign f76 = new_n917 | new_n918;
  assign new_n920 = ~new_n915 & ~new_n917;
  assign new_n921 = a77 & b77;
  assign new_n922 = ~a77 & ~b77;
  assign new_n923 = ~new_n921 & ~new_n922;
  assign new_n924 = ~new_n920 & new_n923;
  assign new_n925 = new_n920 & ~new_n923;
  assign f77 = new_n924 | new_n925;
  assign new_n927 = ~new_n922 & ~new_n924;
  assign new_n928 = a78 & b78;
  assign new_n929 = ~a78 & ~b78;
  assign new_n930 = ~new_n928 & ~new_n929;
  assign new_n931 = ~new_n927 & new_n930;
  assign new_n932 = new_n927 & ~new_n930;
  assign f78 = new_n931 | new_n932;
  assign new_n934 = ~new_n929 & ~new_n931;
  assign new_n935 = a79 & b79;
  assign new_n936 = ~a79 & ~b79;
  assign new_n937 = ~new_n935 & ~new_n936;
  assign new_n938 = ~new_n934 & new_n937;
  assign new_n939 = new_n934 & ~new_n937;
  assign f79 = new_n938 | new_n939;
  assign new_n941 = ~new_n936 & ~new_n938;
  assign new_n942 = a80 & b80;
  assign new_n943 = ~a80 & ~b80;
  assign new_n944 = ~new_n942 & ~new_n943;
  assign new_n945 = ~new_n941 & new_n944;
  assign new_n946 = new_n941 & ~new_n944;
  assign f80 = new_n945 | new_n946;
  assign new_n948 = ~new_n943 & ~new_n945;
  assign new_n949 = a81 & b81;
  assign new_n950 = ~a81 & ~b81;
  assign new_n951 = ~new_n949 & ~new_n950;
  assign new_n952 = ~new_n948 & new_n951;
  assign new_n953 = new_n948 & ~new_n951;
  assign f81 = new_n952 | new_n953;
  assign new_n955 = ~new_n950 & ~new_n952;
  assign new_n956 = a82 & b82;
  assign new_n957 = ~a82 & ~b82;
  assign new_n958 = ~new_n956 & ~new_n957;
  assign new_n959 = ~new_n955 & new_n958;
  assign new_n960 = new_n955 & ~new_n958;
  assign f82 = new_n959 | new_n960;
  assign new_n962 = ~new_n957 & ~new_n959;
  assign new_n963 = a83 & b83;
  assign new_n964 = ~a83 & ~b83;
  assign new_n965 = ~new_n963 & ~new_n964;
  assign new_n966 = ~new_n962 & new_n965;
  assign new_n967 = new_n962 & ~new_n965;
  assign f83 = new_n966 | new_n967;
  assign new_n969 = ~new_n964 & ~new_n966;
  assign new_n970 = a84 & b84;
  assign new_n971 = ~a84 & ~b84;
  assign new_n972 = ~new_n970 & ~new_n971;
  assign new_n973 = ~new_n969 & new_n972;
  assign new_n974 = new_n969 & ~new_n972;
  assign f84 = new_n973 | new_n974;
  assign new_n976 = ~new_n971 & ~new_n973;
  assign new_n977 = a85 & b85;
  assign new_n978 = ~a85 & ~b85;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980 = ~new_n976 & new_n979;
  assign new_n981 = new_n976 & ~new_n979;
  assign f85 = new_n980 | new_n981;
  assign new_n983 = ~new_n978 & ~new_n980;
  assign new_n984 = a86 & b86;
  assign new_n985 = ~a86 & ~b86;
  assign new_n986 = ~new_n984 & ~new_n985;
  assign new_n987 = ~new_n983 & new_n986;
  assign new_n988 = new_n983 & ~new_n986;
  assign f86 = new_n987 | new_n988;
  assign new_n990 = ~new_n985 & ~new_n987;
  assign new_n991 = a87 & b87;
  assign new_n992 = ~a87 & ~b87;
  assign new_n993 = ~new_n991 & ~new_n992;
  assign new_n994 = ~new_n990 & new_n993;
  assign new_n995 = new_n990 & ~new_n993;
  assign f87 = new_n994 | new_n995;
  assign new_n997 = ~new_n992 & ~new_n994;
  assign new_n998 = a88 & b88;
  assign new_n999 = ~a88 & ~b88;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = ~new_n997 & new_n1000;
  assign new_n1002 = new_n997 & ~new_n1000;
  assign f88 = new_n1001 | new_n1002;
  assign new_n1004 = ~new_n999 & ~new_n1001;
  assign new_n1005 = a89 & b89;
  assign new_n1006 = ~a89 & ~b89;
  assign new_n1007 = ~new_n1005 & ~new_n1006;
  assign new_n1008 = ~new_n1004 & new_n1007;
  assign new_n1009 = new_n1004 & ~new_n1007;
  assign f89 = new_n1008 | new_n1009;
  assign new_n1011 = ~new_n1006 & ~new_n1008;
  assign new_n1012 = a90 & b90;
  assign new_n1013 = ~a90 & ~b90;
  assign new_n1014 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = ~new_n1011 & new_n1014;
  assign new_n1016 = new_n1011 & ~new_n1014;
  assign f90 = new_n1015 | new_n1016;
  assign new_n1018 = ~new_n1013 & ~new_n1015;
  assign new_n1019 = a91 & b91;
  assign new_n1020 = ~a91 & ~b91;
  assign new_n1021 = ~new_n1019 & ~new_n1020;
  assign new_n1022 = ~new_n1018 & new_n1021;
  assign new_n1023 = new_n1018 & ~new_n1021;
  assign f91 = new_n1022 | new_n1023;
  assign new_n1025 = ~new_n1020 & ~new_n1022;
  assign new_n1026 = a92 & b92;
  assign new_n1027 = ~a92 & ~b92;
  assign new_n1028 = ~new_n1026 & ~new_n1027;
  assign new_n1029 = ~new_n1025 & new_n1028;
  assign new_n1030 = new_n1025 & ~new_n1028;
  assign f92 = new_n1029 | new_n1030;
  assign new_n1032 = ~new_n1027 & ~new_n1029;
  assign new_n1033 = a93 & b93;
  assign new_n1034 = ~a93 & ~b93;
  assign new_n1035 = ~new_n1033 & ~new_n1034;
  assign new_n1036 = ~new_n1032 & new_n1035;
  assign new_n1037 = new_n1032 & ~new_n1035;
  assign f93 = new_n1036 | new_n1037;
  assign new_n1039 = ~new_n1034 & ~new_n1036;
  assign new_n1040 = a94 & b94;
  assign new_n1041 = ~a94 & ~b94;
  assign new_n1042 = ~new_n1040 & ~new_n1041;
  assign new_n1043 = ~new_n1039 & new_n1042;
  assign new_n1044 = new_n1039 & ~new_n1042;
  assign f94 = new_n1043 | new_n1044;
  assign new_n1046 = ~new_n1041 & ~new_n1043;
  assign new_n1047 = a95 & b95;
  assign new_n1048 = ~a95 & ~b95;
  assign new_n1049 = ~new_n1047 & ~new_n1048;
  assign new_n1050 = ~new_n1046 & new_n1049;
  assign new_n1051 = new_n1046 & ~new_n1049;
  assign f95 = new_n1050 | new_n1051;
  assign new_n1053 = ~new_n1048 & ~new_n1050;
  assign new_n1054 = a96 & b96;
  assign new_n1055 = ~a96 & ~b96;
  assign new_n1056 = ~new_n1054 & ~new_n1055;
  assign new_n1057 = ~new_n1053 & new_n1056;
  assign new_n1058 = new_n1053 & ~new_n1056;
  assign f96 = new_n1057 | new_n1058;
  assign new_n1060 = ~new_n1055 & ~new_n1057;
  assign new_n1061 = a97 & b97;
  assign new_n1062 = ~a97 & ~b97;
  assign new_n1063 = ~new_n1061 & ~new_n1062;
  assign new_n1064 = ~new_n1060 & new_n1063;
  assign new_n1065 = new_n1060 & ~new_n1063;
  assign f97 = new_n1064 | new_n1065;
  assign new_n1067 = ~new_n1062 & ~new_n1064;
  assign new_n1068 = a98 & b98;
  assign new_n1069 = ~a98 & ~b98;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = ~new_n1067 & new_n1070;
  assign new_n1072 = new_n1067 & ~new_n1070;
  assign f98 = new_n1071 | new_n1072;
  assign new_n1074 = ~new_n1069 & ~new_n1071;
  assign new_n1075 = a99 & b99;
  assign new_n1076 = ~a99 & ~b99;
  assign new_n1077 = ~new_n1075 & ~new_n1076;
  assign new_n1078 = ~new_n1074 & new_n1077;
  assign new_n1079 = new_n1074 & ~new_n1077;
  assign f99 = new_n1078 | new_n1079;
  assign new_n1081 = ~new_n1076 & ~new_n1078;
  assign new_n1082 = a100 & b100;
  assign new_n1083 = ~a100 & ~b100;
  assign new_n1084 = ~new_n1082 & ~new_n1083;
  assign new_n1085 = ~new_n1081 & new_n1084;
  assign new_n1086 = new_n1081 & ~new_n1084;
  assign f100 = new_n1085 | new_n1086;
  assign new_n1088 = ~new_n1083 & ~new_n1085;
  assign new_n1089 = a101 & b101;
  assign new_n1090 = ~a101 & ~b101;
  assign new_n1091 = ~new_n1089 & ~new_n1090;
  assign new_n1092 = ~new_n1088 & new_n1091;
  assign new_n1093 = new_n1088 & ~new_n1091;
  assign f101 = new_n1092 | new_n1093;
  assign new_n1095 = ~new_n1090 & ~new_n1092;
  assign new_n1096 = a102 & b102;
  assign new_n1097 = ~a102 & ~b102;
  assign new_n1098 = ~new_n1096 & ~new_n1097;
  assign new_n1099 = ~new_n1095 & new_n1098;
  assign new_n1100 = new_n1095 & ~new_n1098;
  assign f102 = new_n1099 | new_n1100;
  assign new_n1102 = ~new_n1097 & ~new_n1099;
  assign new_n1103 = a103 & b103;
  assign new_n1104 = ~a103 & ~b103;
  assign new_n1105 = ~new_n1103 & ~new_n1104;
  assign new_n1106 = ~new_n1102 & new_n1105;
  assign new_n1107 = new_n1102 & ~new_n1105;
  assign f103 = new_n1106 | new_n1107;
  assign new_n1109 = ~new_n1104 & ~new_n1106;
  assign new_n1110 = a104 & b104;
  assign new_n1111 = ~a104 & ~b104;
  assign new_n1112 = ~new_n1110 & ~new_n1111;
  assign new_n1113 = ~new_n1109 & new_n1112;
  assign new_n1114 = new_n1109 & ~new_n1112;
  assign f104 = new_n1113 | new_n1114;
  assign new_n1116 = ~new_n1111 & ~new_n1113;
  assign new_n1117 = a105 & b105;
  assign new_n1118 = ~a105 & ~b105;
  assign new_n1119 = ~new_n1117 & ~new_n1118;
  assign new_n1120 = ~new_n1116 & new_n1119;
  assign new_n1121 = new_n1116 & ~new_n1119;
  assign f105 = new_n1120 | new_n1121;
  assign new_n1123 = ~new_n1118 & ~new_n1120;
  assign new_n1124 = a106 & b106;
  assign new_n1125 = ~a106 & ~b106;
  assign new_n1126 = ~new_n1124 & ~new_n1125;
  assign new_n1127 = ~new_n1123 & new_n1126;
  assign new_n1128 = new_n1123 & ~new_n1126;
  assign f106 = new_n1127 | new_n1128;
  assign new_n1130 = ~new_n1125 & ~new_n1127;
  assign new_n1131 = a107 & b107;
  assign new_n1132 = ~a107 & ~b107;
  assign new_n1133 = ~new_n1131 & ~new_n1132;
  assign new_n1134 = ~new_n1130 & new_n1133;
  assign new_n1135 = new_n1130 & ~new_n1133;
  assign f107 = new_n1134 | new_n1135;
  assign new_n1137 = ~new_n1132 & ~new_n1134;
  assign new_n1138 = a108 & b108;
  assign new_n1139 = ~a108 & ~b108;
  assign new_n1140 = ~new_n1138 & ~new_n1139;
  assign new_n1141 = ~new_n1137 & new_n1140;
  assign new_n1142 = new_n1137 & ~new_n1140;
  assign f108 = new_n1141 | new_n1142;
  assign new_n1144 = ~new_n1139 & ~new_n1141;
  assign new_n1145 = a109 & b109;
  assign new_n1146 = ~a109 & ~b109;
  assign new_n1147 = ~new_n1145 & ~new_n1146;
  assign new_n1148 = ~new_n1144 & new_n1147;
  assign new_n1149 = new_n1144 & ~new_n1147;
  assign f109 = new_n1148 | new_n1149;
  assign new_n1151 = ~new_n1146 & ~new_n1148;
  assign new_n1152 = a110 & b110;
  assign new_n1153 = ~a110 & ~b110;
  assign new_n1154 = ~new_n1152 & ~new_n1153;
  assign new_n1155 = ~new_n1151 & new_n1154;
  assign new_n1156 = new_n1151 & ~new_n1154;
  assign f110 = new_n1155 | new_n1156;
  assign new_n1158 = ~new_n1153 & ~new_n1155;
  assign new_n1159 = a111 & b111;
  assign new_n1160 = ~a111 & ~b111;
  assign new_n1161 = ~new_n1159 & ~new_n1160;
  assign new_n1162 = ~new_n1158 & new_n1161;
  assign new_n1163 = new_n1158 & ~new_n1161;
  assign f111 = new_n1162 | new_n1163;
  assign new_n1165 = ~new_n1160 & ~new_n1162;
  assign new_n1166 = a112 & b112;
  assign new_n1167 = ~a112 & ~b112;
  assign new_n1168 = ~new_n1166 & ~new_n1167;
  assign new_n1169 = ~new_n1165 & new_n1168;
  assign new_n1170 = new_n1165 & ~new_n1168;
  assign f112 = new_n1169 | new_n1170;
  assign new_n1172 = ~new_n1167 & ~new_n1169;
  assign new_n1173 = a113 & b113;
  assign new_n1174 = ~a113 & ~b113;
  assign new_n1175 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = ~new_n1172 & new_n1175;
  assign new_n1177 = new_n1172 & ~new_n1175;
  assign f113 = new_n1176 | new_n1177;
  assign new_n1179 = ~new_n1174 & ~new_n1176;
  assign new_n1180 = a114 & b114;
  assign new_n1181 = ~a114 & ~b114;
  assign new_n1182 = ~new_n1180 & ~new_n1181;
  assign new_n1183 = ~new_n1179 & new_n1182;
  assign new_n1184 = new_n1179 & ~new_n1182;
  assign f114 = new_n1183 | new_n1184;
  assign new_n1186 = ~new_n1181 & ~new_n1183;
  assign new_n1187 = a115 & b115;
  assign new_n1188 = ~a115 & ~b115;
  assign new_n1189 = ~new_n1187 & ~new_n1188;
  assign new_n1190 = ~new_n1186 & new_n1189;
  assign new_n1191 = new_n1186 & ~new_n1189;
  assign f115 = new_n1190 | new_n1191;
  assign new_n1193 = ~new_n1188 & ~new_n1190;
  assign new_n1194 = a116 & b116;
  assign new_n1195 = ~a116 & ~b116;
  assign new_n1196 = ~new_n1194 & ~new_n1195;
  assign new_n1197 = ~new_n1193 & new_n1196;
  assign new_n1198 = new_n1193 & ~new_n1196;
  assign f116 = new_n1197 | new_n1198;
  assign new_n1200 = ~new_n1195 & ~new_n1197;
  assign new_n1201 = a117 & b117;
  assign new_n1202 = ~a117 & ~b117;
  assign new_n1203 = ~new_n1201 & ~new_n1202;
  assign new_n1204 = ~new_n1200 & new_n1203;
  assign new_n1205 = new_n1200 & ~new_n1203;
  assign f117 = new_n1204 | new_n1205;
  assign new_n1207 = ~new_n1202 & ~new_n1204;
  assign new_n1208 = a118 & b118;
  assign new_n1209 = ~a118 & ~b118;
  assign new_n1210 = ~new_n1208 & ~new_n1209;
  assign new_n1211 = ~new_n1207 & new_n1210;
  assign new_n1212 = new_n1207 & ~new_n1210;
  assign f118 = new_n1211 | new_n1212;
  assign new_n1214 = ~new_n1209 & ~new_n1211;
  assign new_n1215 = a119 & b119;
  assign new_n1216 = ~a119 & ~b119;
  assign new_n1217 = ~new_n1215 & ~new_n1216;
  assign new_n1218 = ~new_n1214 & new_n1217;
  assign new_n1219 = new_n1214 & ~new_n1217;
  assign f119 = new_n1218 | new_n1219;
  assign new_n1221 = ~new_n1216 & ~new_n1218;
  assign new_n1222 = a120 & b120;
  assign new_n1223 = ~a120 & ~b120;
  assign new_n1224 = ~new_n1222 & ~new_n1223;
  assign new_n1225 = ~new_n1221 & new_n1224;
  assign new_n1226 = new_n1221 & ~new_n1224;
  assign f120 = new_n1225 | new_n1226;
  assign new_n1228 = ~new_n1223 & ~new_n1225;
  assign new_n1229 = a121 & b121;
  assign new_n1230 = ~a121 & ~b121;
  assign new_n1231 = ~new_n1229 & ~new_n1230;
  assign new_n1232 = ~new_n1228 & new_n1231;
  assign new_n1233 = new_n1228 & ~new_n1231;
  assign f121 = new_n1232 | new_n1233;
  assign new_n1235 = ~new_n1230 & ~new_n1232;
  assign new_n1236 = a122 & b122;
  assign new_n1237 = ~a122 & ~b122;
  assign new_n1238 = ~new_n1236 & ~new_n1237;
  assign new_n1239 = ~new_n1235 & new_n1238;
  assign new_n1240 = new_n1235 & ~new_n1238;
  assign f122 = new_n1239 | new_n1240;
  assign new_n1242 = ~new_n1237 & ~new_n1239;
  assign new_n1243 = a123 & b123;
  assign new_n1244 = ~a123 & ~b123;
  assign new_n1245 = ~new_n1243 & ~new_n1244;
  assign new_n1246 = ~new_n1242 & new_n1245;
  assign new_n1247 = new_n1242 & ~new_n1245;
  assign f123 = new_n1246 | new_n1247;
  assign new_n1249 = ~new_n1244 & ~new_n1246;
  assign new_n1250 = a124 & b124;
  assign new_n1251 = ~a124 & ~b124;
  assign new_n1252 = ~new_n1250 & ~new_n1251;
  assign new_n1253 = ~new_n1249 & new_n1252;
  assign new_n1254 = new_n1249 & ~new_n1252;
  assign f124 = new_n1253 | new_n1254;
  assign new_n1256 = ~new_n1251 & ~new_n1253;
  assign new_n1257 = a125 & b125;
  assign new_n1258 = ~a125 & ~b125;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = ~new_n1256 & new_n1259;
  assign new_n1261 = new_n1256 & ~new_n1259;
  assign f125 = new_n1260 | new_n1261;
  assign new_n1263 = ~new_n1258 & ~new_n1260;
  assign new_n1264 = a126 & b126;
  assign new_n1265 = ~a126 & ~b126;
  assign new_n1266 = ~new_n1264 & ~new_n1265;
  assign new_n1267 = ~new_n1263 & new_n1266;
  assign new_n1268 = new_n1263 & ~new_n1266;
  assign f126 = new_n1267 | new_n1268;
  assign new_n1270 = ~new_n1265 & ~new_n1267;
  assign new_n1271 = a127 & b127;
  assign new_n1272 = ~a127 & ~b127;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = ~new_n1270 & new_n1273;
  assign new_n1275 = new_n1270 & ~new_n1273;
  assign f127 = new_n1274 | new_n1275;
  assign cOut = ~new_n1272 & ~new_n1274;
endmodule


