// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_, i_10_,
    i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_,
    i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_, i_24_,
    i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_, i_32_,
    i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_, i_19_,
    i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_,
    i_29_, i_51_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_  );
  input  i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_,
    i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_,
    i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_,
    i_24_, i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_,
    i_32_, i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_,
    i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_,
    i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_;
  wire new_n131, new_n132, new_n133, new_n134, new_n135, new_n136, new_n137,
    new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n424, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n473, new_n474, new_n475,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898;
  assign new_n131 = ~i_59_ & ~i_60_;
  assign new_n132 = ~i_58_ & new_n131;
  assign new_n133 = ~i_61_ & ~i_62_;
  assign new_n134 = ~i_56_ & ~i_55_;
  assign new_n135 = ~i_54_ & new_n134;
  assign new_n136 = new_n132 & new_n133;
  assign new_n137 = new_n135 & new_n136;
  assign new_n138 = ~i_46_ & ~i_47_;
  assign new_n139 = ~i_43_ & new_n138;
  assign new_n140 = ~i_53_ & ~i_51_;
  assign new_n141 = ~i_50_ & new_n140;
  assign new_n142 = ~i_41_ & ~i_42_;
  assign new_n143 = ~i_40_ & new_n142;
  assign new_n144 = new_n139 & new_n141;
  assign new_n145 = new_n143 & new_n144;
  assign new_n146 = new_n137 & new_n145;
  assign new_n147 = ~i_18_ & ~i_22_;
  assign new_n148 = ~i_17_ & new_n147;
  assign new_n149 = ~i_25_ & ~i_26_;
  assign new_n150 = ~i_24_ & new_n149;
  assign new_n151 = ~i_14_ & ~i_15_;
  assign new_n152 = ~i_11_ & new_n151;
  assign new_n153 = new_n148 & new_n150;
  assign new_n154 = new_n152 & new_n153;
  assign new_n155 = ~i_34_ & ~i_33_;
  assign new_n156 = ~i_31_ & new_n155;
  assign new_n157 = ~i_39_ & ~i_37_;
  assign new_n158 = ~i_35_ & new_n157;
  assign new_n159 = ~i_30_ & i_29_;
  assign new_n160 = ~i_28_ & new_n159;
  assign new_n161 = new_n156 & new_n158;
  assign new_n162 = new_n160 & new_n161;
  assign new_n163 = ~i_7_ & ~i_6_;
  assign new_n164 = i_5_ & new_n163;
  assign new_n165 = ~i_9_ & ~i_10_;
  assign new_n166 = ~i_8_ & new_n165;
  assign new_n167 = ~i_3_ & ~i_4_;
  assign new_n168 = ~i_0_ & new_n167;
  assign new_n169 = new_n164 & new_n166;
  assign new_n170 = new_n168 & new_n169;
  assign new_n171 = new_n154 & new_n162;
  assign new_n172 = new_n170 & new_n171;
  assign o_1_ = new_n146 & new_n172;
  assign new_n174 = ~i_54_ & ~i_53_;
  assign new_n175 = ~i_51_ & new_n174;
  assign new_n176 = ~i_57_ & ~i_56_;
  assign new_n177 = ~i_55_ & new_n176;
  assign new_n178 = ~i_50_ & ~i_49_;
  assign new_n179 = ~i_48_ & new_n178;
  assign new_n180 = new_n175 & new_n177;
  assign new_n181 = new_n179 & new_n180;
  assign new_n182 = i_64_ & ~i_62_;
  assign new_n183 = ~i_61_ & new_n182;
  assign new_n184 = new_n132 & new_n183;
  assign new_n185 = ~i_42_ & ~i_43_;
  assign new_n186 = ~i_41_ & new_n185;
  assign new_n187 = ~i_45_ & new_n138;
  assign new_n188 = ~i_40_ & ~i_39_;
  assign new_n189 = ~i_37_ & new_n188;
  assign new_n190 = new_n186 & new_n187;
  assign new_n191 = new_n189 & new_n190;
  assign new_n192 = new_n181 & new_n184;
  assign new_n193 = new_n191 & new_n192;
  assign new_n194 = ~i_17_ & ~i_15_;
  assign new_n195 = ~i_14_ & new_n194;
  assign new_n196 = ~i_24_ & ~i_22_;
  assign new_n197 = ~i_18_ & new_n196;
  assign new_n198 = ~i_10_ & ~i_11_;
  assign new_n199 = ~i_9_ & new_n198;
  assign new_n200 = new_n195 & new_n197;
  assign new_n201 = new_n199 & new_n200;
  assign new_n202 = ~i_30_ & ~i_31_;
  assign new_n203 = i_29_ & new_n202;
  assign new_n204 = ~i_34_ & ~i_35_;
  assign new_n205 = ~i_33_ & new_n204;
  assign new_n206 = ~i_28_ & ~i_26_;
  assign new_n207 = ~i_25_ & new_n206;
  assign new_n208 = new_n203 & new_n205;
  assign new_n209 = new_n207 & new_n208;
  assign new_n210 = ~i_5_ & ~i_4_;
  assign new_n211 = ~i_3_ & new_n210;
  assign new_n212 = ~i_7_ & ~i_8_;
  assign new_n213 = ~i_6_ & new_n212;
  assign new_n214 = ~i_1_ & ~i_2_;
  assign new_n215 = ~i_0_ & new_n214;
  assign new_n216 = new_n211 & new_n213;
  assign new_n217 = new_n215 & new_n216;
  assign new_n218 = new_n201 & new_n209;
  assign new_n219 = new_n217 & new_n218;
  assign o_19_ = new_n193 & new_n219;
  assign new_n221 = ~i_40_ & ~i_41_;
  assign new_n222 = ~i_39_ & new_n221;
  assign new_n223 = ~i_43_ & ~i_44_;
  assign new_n224 = ~i_42_ & new_n223;
  assign new_n225 = ~i_38_ & ~i_37_;
  assign new_n226 = ~i_36_ & new_n225;
  assign new_n227 = new_n222 & new_n224;
  assign new_n228 = new_n226 & new_n227;
  assign new_n229 = ~i_53_ & ~i_52_;
  assign new_n230 = ~i_51_ & new_n229;
  assign new_n231 = new_n179 & new_n230;
  assign new_n232 = new_n187 & new_n231;
  assign new_n233 = ~i_32_ & ~i_31_;
  assign new_n234 = ~i_30_ & new_n233;
  assign new_n235 = ~i_28_ & i_29_;
  assign new_n236 = i_27_ & new_n235;
  assign new_n237 = new_n205 & new_n234;
  assign new_n238 = new_n236 & new_n237;
  assign new_n239 = new_n228 & new_n232;
  assign new_n240 = new_n238 & new_n239;
  assign new_n241 = ~i_63_ & ~i_64_;
  assign new_n242 = ~i_59_ & ~i_58_;
  assign new_n243 = ~i_57_ & new_n242;
  assign new_n244 = ~i_60_ & new_n133;
  assign new_n245 = new_n243 & new_n244;
  assign new_n246 = new_n135 & new_n245;
  assign new_n247 = new_n241 & new_n246;
  assign new_n248 = ~i_14_ & ~i_13_;
  assign new_n249 = ~i_12_ & new_n248;
  assign new_n250 = ~i_17_ & ~i_16_;
  assign new_n251 = ~i_15_ & new_n250;
  assign new_n252 = new_n249 & new_n251;
  assign new_n253 = new_n199 & new_n252;
  assign new_n254 = ~i_23_ & ~i_22_;
  assign new_n255 = ~i_21_ & new_n254;
  assign new_n256 = ~i_20_ & ~i_19_;
  assign new_n257 = ~i_18_ & new_n256;
  assign new_n258 = new_n150 & new_n255;
  assign new_n259 = new_n257 & new_n258;
  assign new_n260 = new_n253 & new_n259;
  assign new_n261 = new_n217 & new_n260;
  assign new_n262 = new_n240 & new_n247;
  assign o_2_ = new_n261 & new_n262;
  assign new_n264 = ~i_56_ & new_n242;
  assign new_n265 = ~i_55_ & ~i_54_;
  assign new_n266 = ~i_53_ & new_n265;
  assign new_n267 = new_n244 & new_n264;
  assign new_n268 = new_n266 & new_n267;
  assign new_n269 = i_45_ & ~i_46_;
  assign new_n270 = ~i_43_ & new_n269;
  assign new_n271 = ~i_50_ & ~i_51_;
  assign new_n272 = ~i_47_ & new_n271;
  assign new_n273 = new_n270 & new_n272;
  assign new_n274 = new_n143 & new_n273;
  assign new_n275 = new_n268 & new_n274;
  assign new_n276 = ~i_5_ & new_n163;
  assign new_n277 = new_n166 & new_n276;
  assign new_n278 = new_n168 & new_n277;
  assign new_n279 = new_n171 & new_n278;
  assign o_0_ = new_n275 & new_n279;
  assign new_n281 = ~i_50_ & ~i_58_;
  assign new_n282 = ~i_46_ & new_n281;
  assign new_n283 = i_60_ & new_n282;
  assign new_n284 = i_29_ & ~i_37_;
  assign new_n285 = ~i_28_ & new_n284;
  assign new_n286 = ~i_40_ & ~i_43_;
  assign new_n287 = ~i_39_ & new_n286;
  assign new_n288 = ~i_10_ & new_n151;
  assign new_n289 = new_n285 & new_n287;
  assign new_n290 = new_n288 & new_n289;
  assign o_29_ = new_n283 & new_n290;
  assign new_n292 = ~i_50_ & ~i_47_;
  assign new_n293 = ~i_46_ & new_n292;
  assign new_n294 = ~i_30_ & ~i_37_;
  assign new_n295 = i_29_ & new_n294;
  assign new_n296 = new_n287 & new_n293;
  assign new_n297 = new_n295 & new_n296;
  assign new_n298 = ~i_58_ & ~i_60_;
  assign new_n299 = ~i_56_ & new_n298;
  assign new_n300 = ~i_28_ & ~i_25_;
  assign new_n301 = ~i_24_ & new_n300;
  assign new_n302 = ~i_10_ & ~i_8_;
  assign new_n303 = i_7_ & new_n302;
  assign new_n304 = new_n152 & new_n301;
  assign new_n305 = new_n303 & new_n304;
  assign new_n306 = new_n297 & new_n299;
  assign o_60_ = new_n305 & new_n306;
  assign new_n308 = ~i_55_ & ~i_51_;
  assign new_n309 = ~i_50_ & new_n308;
  assign new_n310 = new_n133 & new_n299;
  assign new_n311 = new_n309 & new_n310;
  assign new_n312 = ~i_15_ & new_n147;
  assign new_n313 = new_n150 & new_n160;
  assign new_n314 = new_n312 & new_n313;
  assign new_n315 = ~i_41_ & i_42_;
  assign new_n316 = ~i_40_ & new_n315;
  assign new_n317 = new_n139 & new_n316;
  assign new_n318 = new_n158 & new_n317;
  assign new_n319 = ~i_14_ & ~i_11_;
  assign new_n320 = ~i_10_ & new_n319;
  assign new_n321 = new_n213 & new_n320;
  assign new_n322 = new_n168 & new_n321;
  assign new_n323 = new_n314 & new_n318;
  assign new_n324 = new_n322 & new_n323;
  assign o_39_ = new_n311 & new_n324;
  assign new_n326 = i_59_ & ~i_58_;
  assign new_n327 = ~i_56_ & new_n326;
  assign new_n328 = new_n244 & new_n327;
  assign new_n329 = new_n309 & new_n328;
  assign new_n330 = new_n139 & new_n143;
  assign new_n331 = new_n158 & new_n330;
  assign new_n332 = new_n314 & new_n331;
  assign new_n333 = new_n322 & new_n332;
  assign o_38_ = new_n329 & new_n333;
  assign new_n335 = ~i_50_ & new_n298;
  assign new_n336 = ~i_46_ & ~i_43_;
  assign new_n337 = ~i_40_ & new_n336;
  assign new_n338 = new_n335 & new_n337;
  assign new_n339 = i_24_ & new_n300;
  assign new_n340 = i_29_ & new_n157;
  assign new_n341 = new_n339 & new_n340;
  assign new_n342 = new_n288 & new_n341;
  assign o_25_ = new_n338 & new_n342;
  assign new_n344 = new_n222 & new_n295;
  assign new_n345 = new_n207 & new_n344;
  assign new_n346 = ~i_58_ & ~i_56_;
  assign new_n347 = ~i_50_ & new_n346;
  assign new_n348 = ~i_62_ & ~i_60_;
  assign new_n349 = new_n347 & new_n348;
  assign new_n350 = new_n139 & new_n349;
  assign new_n351 = ~i_8_ & new_n198;
  assign new_n352 = ~i_24_ & ~i_15_;
  assign new_n353 = ~i_14_ & new_n352;
  assign new_n354 = ~i_7_ & i_6_;
  assign new_n355 = ~i_3_ & new_n354;
  assign new_n356 = new_n351 & new_n353;
  assign new_n357 = new_n355 & new_n356;
  assign new_n358 = new_n345 & new_n350;
  assign o_12_ = new_n357 & new_n358;
  assign new_n360 = ~i_45_ & ~i_43_;
  assign new_n361 = ~i_42_ & new_n360;
  assign new_n362 = ~i_47_ & ~i_48_;
  assign new_n363 = ~i_46_ & new_n362;
  assign new_n364 = new_n361 & new_n363;
  assign new_n365 = new_n222 & new_n364;
  assign new_n366 = ~i_52_ & new_n174;
  assign new_n367 = ~i_49_ & new_n271;
  assign new_n368 = new_n177 & new_n366;
  assign new_n369 = new_n367 & new_n368;
  assign new_n370 = ~i_32_ & new_n155;
  assign new_n371 = ~i_36_ & ~i_37_;
  assign new_n372 = ~i_35_ & new_n371;
  assign new_n373 = new_n370 & new_n372;
  assign new_n374 = new_n203 & new_n373;
  assign new_n375 = new_n365 & new_n369;
  assign new_n376 = new_n374 & new_n375;
  assign new_n377 = ~i_63_ & ~i_62_;
  assign new_n378 = ~i_61_ & new_n377;
  assign new_n379 = ~i_64_ & new_n378;
  assign new_n380 = new_n132 & new_n379;
  assign new_n381 = ~i_21_ & new_n196;
  assign new_n382 = ~i_20_ & i_19_;
  assign new_n383 = ~i_18_ & new_n382;
  assign new_n384 = new_n207 & new_n381;
  assign new_n385 = new_n383 & new_n384;
  assign new_n386 = new_n253 & new_n385;
  assign new_n387 = new_n217 & new_n386;
  assign new_n388 = new_n376 & new_n380;
  assign o_37_ = new_n387 & new_n388;
  assign new_n390 = ~i_45_ & ~i_46_;
  assign new_n391 = ~i_43_ & new_n390;
  assign new_n392 = ~i_49_ & ~i_48_;
  assign new_n393 = ~i_47_ & new_n392;
  assign new_n394 = new_n391 & new_n393;
  assign new_n395 = new_n143 & new_n394;
  assign new_n396 = ~i_58_ & ~i_57_;
  assign new_n397 = ~i_56_ & new_n396;
  assign new_n398 = ~i_52_ & ~i_51_;
  assign new_n399 = ~i_50_ & new_n398;
  assign new_n400 = new_n266 & new_n397;
  assign new_n401 = new_n399 & new_n400;
  assign new_n402 = ~i_36_ & new_n157;
  assign new_n403 = i_32_ & ~i_31_;
  assign new_n404 = ~i_30_ & new_n403;
  assign new_n405 = new_n205 & new_n402;
  assign new_n406 = new_n404 & new_n405;
  assign new_n407 = new_n395 & new_n401;
  assign new_n408 = new_n406 & new_n407;
  assign new_n409 = ~i_62_ & new_n241;
  assign new_n410 = ~i_61_ & ~i_60_;
  assign new_n411 = ~i_59_ & new_n410;
  assign new_n412 = new_n409 & new_n411;
  assign new_n413 = ~i_25_ & ~i_24_;
  assign new_n414 = ~i_22_ & new_n413;
  assign new_n415 = ~i_26_ & new_n235;
  assign new_n416 = ~i_20_ & ~i_21_;
  assign new_n417 = ~i_18_ & new_n416;
  assign new_n418 = new_n414 & new_n415;
  assign new_n419 = new_n417 & new_n418;
  assign new_n420 = new_n253 & new_n419;
  assign new_n421 = new_n217 & new_n420;
  assign new_n422 = new_n408 & new_n412;
  assign o_26_ = new_n421 & new_n422;
  assign new_n424 = i_29_ & i_37_;
  assign o_11_ = ~i_15_ & new_n424;
  assign new_n426 = i_57_ & ~i_56_;
  assign new_n427 = ~i_55_ & new_n426;
  assign new_n428 = new_n175 & new_n427;
  assign new_n429 = new_n179 & new_n428;
  assign new_n430 = new_n136 & new_n429;
  assign new_n431 = new_n191 & new_n430;
  assign o_50_ = new_n219 & new_n431;
  assign new_n433 = i_61_ & ~i_62_;
  assign new_n434 = ~i_60_ & new_n433;
  assign new_n435 = ~i_55_ & new_n346;
  assign new_n436 = new_n434 & new_n435;
  assign new_n437 = ~i_30_ & ~i_35_;
  assign new_n438 = i_29_ & new_n437;
  assign new_n439 = new_n207 & new_n438;
  assign new_n440 = new_n197 & new_n439;
  assign new_n441 = ~i_41_ & new_n336;
  assign new_n442 = new_n272 & new_n441;
  assign new_n443 = new_n189 & new_n442;
  assign new_n444 = ~i_7_ & new_n302;
  assign new_n445 = ~i_6_ & ~i_3_;
  assign new_n446 = ~i_0_ & new_n445;
  assign new_n447 = new_n152 & new_n444;
  assign new_n448 = new_n446 & new_n447;
  assign new_n449 = new_n440 & new_n443;
  assign new_n450 = new_n448 & new_n449;
  assign o_36_ = new_n436 & new_n450;
  assign new_n452 = new_n179 & new_n187;
  assign new_n453 = new_n186 & new_n452;
  assign new_n454 = new_n135 & new_n243;
  assign new_n455 = new_n230 & new_n454;
  assign new_n456 = ~i_36_ & ~i_35_;
  assign new_n457 = ~i_34_ & new_n456;
  assign new_n458 = ~i_31_ & ~i_33_;
  assign new_n459 = ~i_30_ & new_n458;
  assign new_n460 = new_n189 & new_n457;
  assign new_n461 = new_n459 & new_n460;
  assign new_n462 = new_n453 & new_n455;
  assign new_n463 = new_n461 & new_n462;
  assign new_n464 = new_n241 & new_n244;
  assign new_n465 = ~i_14_ & i_13_;
  assign new_n466 = ~i_12_ & new_n465;
  assign new_n467 = new_n251 & new_n466;
  assign new_n468 = new_n199 & new_n467;
  assign new_n469 = new_n419 & new_n468;
  assign new_n470 = new_n217 & new_n469;
  assign new_n471 = new_n463 & new_n464;
  assign o_27_ = new_n470 & new_n471;
  assign new_n473 = i_50_ & ~i_58_;
  assign new_n474 = ~i_43_ & new_n473;
  assign new_n475 = new_n285 & new_n474;
  assign o_14_ = new_n288 & new_n475;
  assign new_n477 = ~i_58_ & new_n410;
  assign new_n478 = ~i_51_ & new_n134;
  assign new_n479 = ~i_62_ & new_n477;
  assign new_n480 = new_n478 & new_n479;
  assign new_n481 = ~i_41_ & ~i_43_;
  assign new_n482 = ~i_40_ & new_n481;
  assign new_n483 = new_n293 & new_n482;
  assign new_n484 = new_n158 & new_n483;
  assign new_n485 = ~i_3_ & i_4_;
  assign new_n486 = ~i_0_ & new_n485;
  assign new_n487 = new_n321 & new_n486;
  assign new_n488 = new_n314 & new_n484;
  assign new_n489 = new_n487 & new_n488;
  assign o_35_ = new_n480 & new_n489;
  assign new_n491 = ~i_50_ & ~i_46_;
  assign new_n492 = ~i_43_ & new_n491;
  assign new_n493 = new_n298 & new_n492;
  assign new_n494 = i_25_ & new_n235;
  assign new_n495 = new_n189 & new_n494;
  assign new_n496 = new_n288 & new_n495;
  assign o_28_ = new_n493 & new_n496;
  assign new_n498 = ~i_30_ & new_n157;
  assign new_n499 = i_41_ & ~i_43_;
  assign new_n500 = ~i_40_ & new_n499;
  assign new_n501 = new_n498 & new_n500;
  assign new_n502 = new_n415 & new_n501;
  assign new_n503 = ~i_62_ & new_n299;
  assign new_n504 = new_n293 & new_n503;
  assign new_n505 = ~i_15_ & new_n413;
  assign new_n506 = ~i_3_ & new_n212;
  assign new_n507 = new_n320 & new_n505;
  assign new_n508 = new_n506 & new_n507;
  assign new_n509 = new_n502 & new_n504;
  assign o_13_ = new_n508 & new_n509;
  assign new_n511 = ~i_43_ & ~i_37_;
  assign new_n512 = i_29_ & new_n511;
  assign new_n513 = ~i_28_ & ~i_15_;
  assign new_n514 = ~i_14_ & new_n513;
  assign new_n515 = i_58_ & new_n512;
  assign o_34_ = new_n514 & new_n515;
  assign new_n517 = new_n207 & new_n295;
  assign new_n518 = new_n197 & new_n517;
  assign new_n519 = new_n139 & new_n347;
  assign new_n520 = new_n222 & new_n519;
  assign new_n521 = i_0_ & new_n445;
  assign new_n522 = new_n447 & new_n521;
  assign new_n523 = new_n518 & new_n520;
  assign new_n524 = new_n522 & new_n523;
  assign o_21_ = new_n348 & new_n524;
  assign new_n526 = i_26_ & new_n235;
  assign new_n527 = new_n337 & new_n498;
  assign new_n528 = new_n526 & new_n527;
  assign new_n529 = ~i_58_ & new_n348;
  assign new_n530 = ~i_50_ & ~i_56_;
  assign new_n531 = ~i_47_ & new_n530;
  assign new_n532 = new_n529 & new_n531;
  assign new_n533 = new_n528 & new_n532;
  assign o_16_ = new_n508 & new_n533;
  assign new_n535 = i_54_ & new_n134;
  assign new_n536 = ~i_42_ & new_n336;
  assign new_n537 = new_n272 & new_n535;
  assign new_n538 = new_n536 & new_n537;
  assign new_n539 = new_n136 & new_n538;
  assign new_n540 = new_n197 & new_n207;
  assign new_n541 = new_n195 & new_n540;
  assign new_n542 = ~i_35_ & ~i_37_;
  assign new_n543 = ~i_34_ & new_n542;
  assign new_n544 = ~i_30_ & ~i_33_;
  assign new_n545 = i_29_ & new_n544;
  assign new_n546 = new_n222 & new_n543;
  assign new_n547 = new_n545 & new_n546;
  assign new_n548 = new_n199 & new_n213;
  assign new_n549 = new_n168 & new_n548;
  assign new_n550 = new_n541 & new_n547;
  assign new_n551 = new_n549 & new_n550;
  assign o_40_ = new_n539 & new_n551;
  assign new_n553 = i_39_ & new_n286;
  assign new_n554 = new_n285 & new_n553;
  assign new_n555 = new_n288 & new_n554;
  assign o_33_ = new_n281 & new_n555;
  assign new_n557 = new_n266 & new_n367;
  assign new_n558 = new_n363 & new_n557;
  assign new_n559 = new_n397 & new_n412;
  assign new_n560 = i_36_ & ~i_37_;
  assign new_n561 = ~i_35_ & new_n560;
  assign new_n562 = new_n222 & new_n361;
  assign new_n563 = new_n561 & new_n562;
  assign new_n564 = new_n558 & new_n559;
  assign new_n565 = new_n563 & new_n564;
  assign new_n566 = ~i_12_ & new_n151;
  assign new_n567 = new_n148 & new_n566;
  assign new_n568 = new_n199 & new_n567;
  assign new_n569 = new_n156 & new_n160;
  assign new_n570 = new_n150 & new_n569;
  assign new_n571 = new_n568 & new_n570;
  assign new_n572 = new_n217 & new_n571;
  assign o_22_ = new_n565 & new_n572;
  assign new_n574 = ~i_58_ & ~i_43_;
  assign new_n575 = i_10_ & new_n151;
  assign new_n576 = new_n285 & new_n574;
  assign o_15_ = new_n575 & new_n576;
  assign new_n578 = i_46_ & new_n281;
  assign o_32_ = new_n290 & new_n578;
  assign new_n580 = new_n393 & new_n399;
  assign new_n581 = new_n391 & new_n580;
  assign new_n582 = new_n397 & new_n411;
  assign new_n583 = new_n266 & new_n582;
  assign new_n584 = new_n143 & new_n402;
  assign new_n585 = new_n205 & new_n584;
  assign new_n586 = new_n581 & new_n583;
  assign new_n587 = new_n585 & new_n586;
  assign new_n588 = ~i_18_ & ~i_17_;
  assign new_n589 = i_16_ & new_n588;
  assign new_n590 = new_n566 & new_n589;
  assign new_n591 = new_n199 & new_n590;
  assign new_n592 = new_n203 & new_n207;
  assign new_n593 = new_n381 & new_n592;
  assign new_n594 = new_n591 & new_n593;
  assign new_n595 = new_n217 & new_n594;
  assign new_n596 = new_n409 & new_n587;
  assign o_23_ = new_n595 & new_n596;
  assign new_n598 = i_62_ & new_n299;
  assign new_n599 = new_n304 & new_n444;
  assign new_n600 = new_n297 & new_n598;
  assign o_18_ = new_n599 & new_n600;
  assign new_n602 = new_n175 & new_n179;
  assign new_n603 = new_n187 & new_n602;
  assign new_n604 = new_n132 & new_n378;
  assign new_n605 = new_n177 & new_n604;
  assign new_n606 = new_n186 & new_n189;
  assign new_n607 = new_n457 & new_n606;
  assign new_n608 = new_n603 & new_n605;
  assign new_n609 = new_n607 & new_n608;
  assign new_n610 = ~i_18_ & i_21_;
  assign new_n611 = ~i_17_ & new_n610;
  assign new_n612 = new_n566 & new_n611;
  assign new_n613 = new_n199 & new_n612;
  assign new_n614 = new_n415 & new_n459;
  assign new_n615 = new_n414 & new_n614;
  assign new_n616 = new_n613 & new_n615;
  assign new_n617 = new_n217 & new_n616;
  assign new_n618 = ~i_64_ & new_n609;
  assign o_31_ = new_n617 & new_n618;
  assign new_n620 = ~i_60_ & new_n282;
  assign new_n621 = new_n287 & new_n620;
  assign new_n622 = ~i_14_ & i_11_;
  assign new_n623 = ~i_10_ & new_n622;
  assign new_n624 = new_n285 & new_n505;
  assign new_n625 = new_n623 & new_n624;
  assign o_24_ = new_n621 & new_n625;
  assign new_n627 = new_n139 & new_n189;
  assign new_n628 = new_n160 & new_n627;
  assign new_n629 = i_3_ & new_n212;
  assign new_n630 = new_n507 & new_n629;
  assign new_n631 = new_n349 & new_n628;
  assign o_17_ = new_n630 & new_n631;
  assign new_n633 = new_n363 & new_n367;
  assign new_n634 = new_n361 & new_n633;
  assign new_n635 = new_n132 & new_n177;
  assign new_n636 = new_n366 & new_n635;
  assign new_n637 = new_n222 & new_n372;
  assign new_n638 = new_n156 & new_n637;
  assign new_n639 = new_n634 & new_n636;
  assign new_n640 = new_n638 & new_n639;
  assign new_n641 = ~i_16_ & new_n588;
  assign new_n642 = new_n566 & new_n641;
  assign new_n643 = new_n199 & new_n642;
  assign new_n644 = ~i_21_ & ~i_22_;
  assign new_n645 = i_20_ & new_n644;
  assign new_n646 = new_n313 & new_n645;
  assign new_n647 = new_n643 & new_n646;
  assign new_n648 = new_n217 & new_n647;
  assign new_n649 = new_n379 & new_n640;
  assign o_56_ = new_n648 & new_n649;
  assign new_n651 = new_n132 & new_n135;
  assign new_n652 = new_n141 & new_n651;
  assign new_n653 = new_n133 & new_n652;
  assign new_n654 = new_n191 & new_n653;
  assign new_n655 = i_1_ & ~i_2_;
  assign new_n656 = ~i_0_ & new_n655;
  assign new_n657 = new_n216 & new_n656;
  assign new_n658 = new_n218 & new_n657;
  assign o_43_ = new_n654 & new_n658;
  assign new_n660 = ~i_53_ & i_52_;
  assign new_n661 = ~i_51_ & new_n660;
  assign new_n662 = new_n179 & new_n661;
  assign new_n663 = new_n187 & new_n662;
  assign new_n664 = new_n246 & new_n663;
  assign new_n665 = new_n607 & new_n664;
  assign new_n666 = ~i_18_ & ~i_21_;
  assign new_n667 = ~i_17_ & new_n666;
  assign new_n668 = new_n566 & new_n667;
  assign new_n669 = new_n199 & new_n668;
  assign new_n670 = new_n615 & new_n669;
  assign new_n671 = new_n217 & new_n670;
  assign new_n672 = new_n241 & new_n665;
  assign o_30_ = new_n671 & new_n672;
  assign new_n674 = ~i_30_ & i_35_;
  assign new_n675 = i_29_ & new_n674;
  assign new_n676 = new_n207 & new_n675;
  assign new_n677 = new_n197 & new_n676;
  assign new_n678 = new_n443 & new_n677;
  assign new_n679 = new_n448 & new_n678;
  assign o_55_ = new_n503 & new_n679;
  assign new_n681 = new_n411 & new_n435;
  assign new_n682 = new_n175 & new_n681;
  assign new_n683 = new_n293 & new_n361;
  assign new_n684 = new_n222 & new_n683;
  assign new_n685 = ~i_62_ & new_n682;
  assign new_n686 = new_n684 & new_n685;
  assign new_n687 = ~i_15_ & new_n588;
  assign new_n688 = new_n414 & new_n687;
  assign new_n689 = new_n320 & new_n688;
  assign new_n690 = new_n459 & new_n543;
  assign new_n691 = new_n415 & new_n690;
  assign new_n692 = ~i_5_ & ~i_6_;
  assign new_n693 = ~i_4_ & new_n692;
  assign new_n694 = ~i_9_ & ~i_8_;
  assign new_n695 = ~i_7_ & new_n694;
  assign new_n696 = ~i_3_ & i_2_;
  assign new_n697 = ~i_0_ & new_n696;
  assign new_n698 = new_n693 & new_n695;
  assign new_n699 = new_n697 & new_n698;
  assign new_n700 = new_n689 & new_n691;
  assign new_n701 = new_n699 & new_n700;
  assign o_44_ = new_n686 & new_n701;
  assign new_n703 = new_n160 & new_n189;
  assign new_n704 = new_n150 & new_n703;
  assign new_n705 = new_n441 & new_n532;
  assign new_n706 = i_22_ & ~i_15_;
  assign new_n707 = ~i_14_ & new_n706;
  assign new_n708 = ~i_3_ & new_n163;
  assign new_n709 = new_n351 & new_n707;
  assign new_n710 = new_n708 & new_n709;
  assign new_n711 = new_n704 & new_n705;
  assign o_58_ = new_n710 & new_n711;
  assign new_n713 = ~i_62_ & new_n411;
  assign new_n714 = new_n272 & new_n435;
  assign new_n715 = new_n536 & new_n714;
  assign new_n716 = new_n713 & new_n715;
  assign new_n717 = ~i_30_ & i_33_;
  assign new_n718 = i_29_ & new_n717;
  assign new_n719 = new_n546 & new_n718;
  assign new_n720 = new_n541 & new_n719;
  assign new_n721 = new_n549 & new_n720;
  assign o_41_ = new_n716 & new_n721;
  assign new_n723 = new_n415 & new_n498;
  assign new_n724 = new_n414 & new_n723;
  assign new_n725 = new_n293 & new_n299;
  assign new_n726 = new_n482 & new_n725;
  assign new_n727 = i_18_ & ~i_15_;
  assign new_n728 = ~i_14_ & new_n727;
  assign new_n729 = new_n351 & new_n728;
  assign new_n730 = new_n708 & new_n729;
  assign new_n731 = new_n724 & new_n726;
  assign new_n732 = new_n730 & new_n731;
  assign o_57_ = ~i_62_ & new_n732;
  assign new_n734 = i_49_ & new_n271;
  assign new_n735 = new_n264 & new_n266;
  assign new_n736 = new_n734 & new_n735;
  assign new_n737 = new_n244 & new_n736;
  assign new_n738 = new_n191 & new_n737;
  assign o_42_ = new_n219 & new_n738;
  assign new_n740 = ~i_56_ & i_51_;
  assign new_n741 = ~i_50_ & new_n740;
  assign new_n742 = new_n139 & new_n741;
  assign new_n743 = new_n222 & new_n742;
  assign new_n744 = new_n518 & new_n743;
  assign new_n745 = new_n448 & new_n744;
  assign o_20_ = new_n529 & new_n745;
  assign new_n747 = new_n135 & new_n141;
  assign new_n748 = new_n393 & new_n747;
  assign new_n749 = new_n243 & new_n464;
  assign new_n750 = new_n143 & new_n391;
  assign new_n751 = new_n158 & new_n750;
  assign new_n752 = new_n748 & new_n749;
  assign new_n753 = new_n751 & new_n752;
  assign new_n754 = i_12_ & new_n151;
  assign new_n755 = new_n148 & new_n754;
  assign new_n756 = new_n199 & new_n755;
  assign new_n757 = new_n570 & new_n756;
  assign new_n758 = new_n217 & new_n757;
  assign o_52_ = new_n753 & new_n758;
  assign new_n760 = new_n272 & new_n681;
  assign new_n761 = ~i_62_ & new_n760;
  assign new_n762 = ~i_18_ & i_17_;
  assign new_n763 = ~i_15_ & new_n762;
  assign new_n764 = new_n418 & new_n763;
  assign new_n765 = ~i_30_ & new_n542;
  assign new_n766 = new_n222 & new_n536;
  assign new_n767 = new_n765 & new_n766;
  assign new_n768 = new_n764 & new_n767;
  assign new_n769 = new_n322 & new_n768;
  assign o_47_ = new_n761 & new_n769;
  assign new_n771 = i_48_ & new_n178;
  assign new_n772 = new_n175 & new_n435;
  assign new_n773 = new_n771 & new_n772;
  assign new_n774 = new_n713 & new_n773;
  assign new_n775 = new_n191 & new_n774;
  assign o_51_ = new_n219 & new_n775;
  assign new_n777 = new_n435 & new_n713;
  assign new_n778 = new_n175 & new_n293;
  assign new_n779 = new_n186 & new_n778;
  assign new_n780 = new_n777 & new_n779;
  assign new_n781 = ~i_30_ & i_31_;
  assign new_n782 = i_29_ & new_n781;
  assign new_n783 = new_n189 & new_n205;
  assign new_n784 = new_n782 & new_n783;
  assign new_n785 = new_n541 & new_n784;
  assign new_n786 = new_n549 & new_n785;
  assign o_48_ = new_n780 & new_n786;
  assign new_n788 = i_55_ & new_n346;
  assign new_n789 = new_n348 & new_n788;
  assign o_54_ = new_n450 & new_n789;
  assign new_n791 = new_n264 & new_n309;
  assign new_n792 = new_n139 & new_n791;
  assign new_n793 = new_n244 & new_n792;
  assign new_n794 = ~i_30_ & i_34_;
  assign new_n795 = i_29_ & new_n794;
  assign new_n796 = new_n143 & new_n158;
  assign new_n797 = new_n795 & new_n796;
  assign new_n798 = new_n541 & new_n797;
  assign new_n799 = new_n549 & new_n798;
  assign o_45_ = new_n793 & new_n799;
  assign new_n801 = i_28_ & i_29_;
  assign new_n802 = ~i_15_ & new_n801;
  assign o_10_ = ~i_37_ & new_n802;
  assign new_n804 = i_63_ & ~i_62_;
  assign new_n805 = ~i_61_ & new_n804;
  assign new_n806 = ~i_64_ & new_n805;
  assign new_n807 = new_n132 & new_n806;
  assign new_n808 = new_n181 & new_n807;
  assign new_n809 = new_n191 & new_n808;
  assign o_53_ = new_n219 & new_n809;
  assign new_n811 = new_n132 & new_n478;
  assign new_n812 = new_n293 & new_n811;
  assign new_n813 = new_n133 & new_n812;
  assign new_n814 = new_n438 & new_n606;
  assign new_n815 = i_9_ & new_n198;
  assign new_n816 = new_n213 & new_n815;
  assign new_n817 = new_n168 & new_n816;
  assign new_n818 = new_n541 & new_n814;
  assign new_n819 = new_n817 & new_n818;
  assign o_46_ = new_n813 & new_n819;
  assign new_n821 = new_n337 & new_n531;
  assign new_n822 = new_n498 & new_n821;
  assign new_n823 = ~i_25_ & new_n235;
  assign new_n824 = i_8_ & new_n198;
  assign new_n825 = new_n353 & new_n823;
  assign new_n826 = new_n824 & new_n825;
  assign new_n827 = new_n298 & new_n822;
  assign o_61_ = new_n826 & new_n827;
  assign new_n829 = new_n135 & new_n230;
  assign new_n830 = new_n179 & new_n829;
  assign new_n831 = ~i_32_ & ~i_33_;
  assign new_n832 = ~i_31_ & new_n831;
  assign new_n833 = new_n457 & new_n832;
  assign new_n834 = new_n160 & new_n833;
  assign new_n835 = new_n191 & new_n830;
  assign new_n836 = new_n834 & new_n835;
  assign new_n837 = i_23_ & ~i_22_;
  assign new_n838 = ~i_21_ & new_n837;
  assign new_n839 = new_n150 & new_n838;
  assign new_n840 = new_n257 & new_n839;
  assign new_n841 = new_n253 & new_n840;
  assign new_n842 = new_n217 & new_n841;
  assign new_n843 = new_n749 & new_n836;
  assign o_9_ = new_n842 & new_n843;
  assign new_n845 = ~i_46_ & i_47_;
  assign new_n846 = ~i_43_ & new_n845;
  assign new_n847 = new_n347 & new_n846;
  assign new_n848 = new_n189 & new_n847;
  assign new_n849 = new_n160 & new_n505;
  assign new_n850 = new_n320 & new_n849;
  assign new_n851 = ~i_60_ & new_n848;
  assign o_62_ = new_n850 & new_n851;
  assign new_n853 = i_56_ & new_n298;
  assign new_n854 = new_n492 & new_n853;
  assign new_n855 = new_n189 & new_n854;
  assign o_63_ = new_n850 & new_n855;
  assign new_n857 = i_53_ & new_n265;
  assign new_n858 = new_n272 & new_n857;
  assign new_n859 = new_n536 & new_n858;
  assign new_n860 = new_n267 & new_n859;
  assign o_49_ = new_n551 & new_n860;
  assign new_n862 = i_43_ & ~i_37_;
  assign new_n863 = ~i_15_ & new_n235;
  assign o_7_ = new_n862 & new_n863;
  assign new_n865 = new_n189 & new_n493;
  assign new_n866 = i_30_ & i_29_;
  assign new_n867 = ~i_28_ & new_n866;
  assign new_n868 = new_n505 & new_n867;
  assign new_n869 = new_n320 & new_n868;
  assign o_64_ = new_n865 & new_n869;
  assign new_n871 = ~i_39_ & i_38_;
  assign new_n872 = ~i_37_ & new_n871;
  assign new_n873 = new_n750 & new_n872;
  assign new_n874 = new_n266 & new_n399;
  assign new_n875 = new_n393 & new_n874;
  assign new_n876 = new_n873 & new_n875;
  assign new_n877 = new_n834 & new_n876;
  assign new_n878 = new_n559 & new_n877;
  assign o_8_ = new_n261 & new_n878;
  assign new_n880 = ~i_50_ & ~i_43_;
  assign new_n881 = i_40_ & new_n880;
  assign new_n882 = new_n285 & new_n881;
  assign new_n883 = new_n288 & new_n882;
  assign o_59_ = ~i_58_ & new_n883;
  assign new_n885 = i_14_ & new_n513;
  assign o_6_ = new_n512 & new_n885;
  assign new_n887 = ~i_45_ & i_44_;
  assign new_n888 = ~i_43_ & new_n887;
  assign new_n889 = ~i_39_ & ~i_38_;
  assign new_n890 = ~i_37_ & new_n889;
  assign new_n891 = new_n143 & new_n888;
  assign new_n892 = new_n890 & new_n891;
  assign new_n893 = new_n366 & new_n367;
  assign new_n894 = new_n363 & new_n893;
  assign new_n895 = new_n892 & new_n894;
  assign new_n896 = new_n834 & new_n895;
  assign new_n897 = ~i_64_ & new_n605;
  assign new_n898 = new_n896 & new_n897;
  assign o_3_ = new_n261 & new_n898;
  assign o_4_ = i_15_ & i_29_;
  assign o_5_ = i_29_;
endmodule


