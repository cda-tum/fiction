// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3, pj0,
    pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4, pl1,
    pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0, pp0,
    pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3, pq2,
    pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2, pu3,
    pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0, pz3,
    pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po,
    pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, pl4, px, ph1, pi0, pj3, pk2, pm4, py, ph2, pi3,
    pj0, pk1, pn4, pz, ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pi4,
    pl1, pm0, pn3, po2, pj4, pl2, pm3, pn0, po1, pk4, pl3, pm2, pn1, po0,
    pp0, pq1, pr2, ps3, pa, pp1, pq0, pr3, ps2, pb, pp2, pq3, ps1, pc, pp3,
    pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1, pu0, pv3, pw2, pf, pt2,
    pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0, py1, pz2, pi, px1, py0,
    pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl, pm, pn, po;
  output pe5, pf6, pg7, ph8, pi9, pd5, pf7, pg6, ph9, pi8, pd6, pe7, pg5, pj8,
    pk9, pd7, pe6, pf5, pj9, pk8, pa5, pb6, pc7, pl8, pm9, pb7, pc6, pl9,
    pm8, pa7, pc5, pn8, po9, pa6, pb5, pn9, po8, pa9, pm5, pn6, po7, pa8,
    pl5, pn7, po6, pb8, pc9, pl6, pm7, po5, pb9, pc8, pl7, pm6, pn5, po4,
    pd8, pe9, pi5, pj6, pk7, pd9, pe8, ph5, pj7, pk6, pf8, pg9, ph6, pi7,
    pk5, pf9, pg8, ph7, pi6, pj5, pt4, pu5, pv6, pw7, px8, pt5, pu4, pv7,
    pw6, py8, pt6, pu7, pv4, pw5, pz8, pt7, pu6, pv5, pw4, pp4, pq5, pr6,
    ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7, pq6, pr5, ps4, pp8,
    pq9, pp9, pq8, pr8, ps9, pr9, ps8, pt8, pu9, px4, py5, pz6, pt9, pu8,
    px5, py4, pz7, pv8, pw9, px6, py7, pz4, pv9, pw8, px7, py6, pz5;
  wire new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1459, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1516,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1524, new_n1525, new_n1526, new_n1527, new_n1528, new_n1529,
    new_n1530, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1562, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1606,
    new_n1607, new_n1608, new_n1609, new_n1610, new_n1611, new_n1612,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1706, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1723, new_n1724, new_n1725, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776, new_n1777, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1866, new_n1867, new_n1868, new_n1869, new_n1870,
    new_n1871, new_n1872, new_n1873, new_n1874, new_n1875, new_n1876,
    new_n1877, new_n1879, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1906, new_n1907, new_n1908, new_n1909,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1919, new_n1921, new_n1922, new_n1923, new_n1924,
    new_n1925, new_n1926, new_n1927, new_n1928, new_n1929, new_n1930,
    new_n1931, new_n1932, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1959, new_n1960, new_n1961, new_n1962, new_n1963, new_n1964,
    new_n1965, new_n1966, new_n1967, new_n1968, new_n1969, new_n1970,
    new_n1971, new_n1972, new_n1973, new_n1974, new_n1975, new_n1976,
    new_n1977, new_n1978, new_n1979, new_n1980, new_n1981, new_n1982,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n2000, new_n2001, new_n2002,
    new_n2003, new_n2004, new_n2005, new_n2006, new_n2007, new_n2008,
    new_n2009, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2081;
  assign pe5 = pm0 & pn3;
  assign pf6 = ~pl4 | ~pk1;
  assign new_n285 = ~pi1 & ~ph1;
  assign new_n286 = ~pj1 & new_n285;
  assign new_n287 = ~pk1 & new_n286;
  assign new_n288 = ~pl1 & new_n287;
  assign new_n289 = ~pa4 & pz3;
  assign new_n290 = ~px3 & new_n289;
  assign new_n291 = py3 & new_n290;
  assign new_n292 = ~pb4 & new_n291;
  assign new_n293 = ~pc4 & new_n292;
  assign new_n294 = pl4 & ~new_n293;
  assign new_n295 = ~new_n288 & ~new_n294;
  assign new_n296 = ~px1 & new_n295;
  assign new_n297 = po0 & ~pq0;
  assign new_n298 = pn0 & new_n297;
  assign new_n299 = ~new_n288 & new_n297;
  assign new_n300 = pq & new_n297;
  assign new_n301 = ~new_n298 & ~new_n299;
  assign new_n302 = ~new_n300 & new_n301;
  assign new_n303 = ~new_n296 & ~new_n302;
  assign new_n304 = ~pn0 & new_n303;
  assign new_n305 = new_n293 & new_n304;
  assign new_n306 = pl4 & ~py1;
  assign new_n307 = new_n304 & ~new_n306;
  assign new_n308 = px1 & new_n303;
  assign new_n309 = ~new_n306 & new_n308;
  assign new_n310 = ~pn0 & new_n288;
  assign new_n311 = new_n308 & new_n310;
  assign new_n312 = new_n293 & new_n308;
  assign new_n313 = new_n294 & new_n303;
  assign new_n314 = ~new_n306 & new_n313;
  assign new_n315 = new_n310 & new_n313;
  assign new_n316 = new_n304 & new_n310;
  assign new_n317 = new_n293 & new_n313;
  assign new_n318 = ~new_n305 & ~new_n307;
  assign new_n319 = ~new_n309 & new_n318;
  assign new_n320 = ~new_n311 & ~new_n312;
  assign new_n321 = new_n319 & new_n320;
  assign new_n322 = ~new_n316 & ~new_n317;
  assign new_n323 = ~new_n314 & ~new_n315;
  assign new_n324 = new_n322 & new_n323;
  assign pg7 = ~new_n321 | ~new_n324;
  assign new_n326 = pl4 & pz2;
  assign new_n327 = ~pk0 & pl0;
  assign new_n328 = pk0 & ~pl0;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = new_n288 & new_n329;
  assign new_n331 = ~pm0 & new_n330;
  assign new_n332 = ~pn0 & new_n331;
  assign new_n333 = py2 & ~new_n332;
  assign new_n334 = ~pl4 & new_n333;
  assign new_n335 = ~pm0 & ~pn0;
  assign new_n336 = new_n288 & new_n335;
  assign new_n337 = new_n329 & new_n336;
  assign new_n338 = po & new_n337;
  assign new_n339 = ~new_n334 & ~new_n338;
  assign new_n340 = ~new_n326 & new_n339;
  assign new_n341 = ~new_n293 & new_n340;
  assign new_n342 = new_n293 & new_n339;
  assign new_n343 = ~py2 & new_n342;
  assign new_n344 = ~py2 & new_n340;
  assign new_n345 = ~pl0 & new_n288;
  assign new_n346 = ~pk0 & new_n345;
  assign new_n347 = pl0 & new_n288;
  assign new_n348 = pk0 & new_n347;
  assign new_n349 = ~new_n346 & ~new_n348;
  assign new_n350 = ~pm0 & ~new_n349;
  assign new_n351 = ~pn0 & new_n350;
  assign new_n352 = new_n339 & new_n351;
  assign new_n353 = ~new_n341 & ~new_n343;
  assign new_n354 = ~new_n344 & ~new_n352;
  assign new_n355 = new_n353 & new_n354;
  assign new_n356 = po0 & new_n355;
  assign ph8 = ~pq0 & new_n356;
  assign new_n358 = ~px3 & ~new_n293;
  assign new_n359 = py3 & new_n358;
  assign new_n360 = ~pz3 & new_n359;
  assign new_n361 = pl4 & new_n360;
  assign new_n362 = ~pq0 & ~new_n361;
  assign new_n363 = pn0 & new_n362;
  assign new_n364 = ~new_n288 & new_n362;
  assign new_n365 = ~new_n363 & ~new_n364;
  assign new_n366 = pl4 & py3;
  assign new_n367 = ~new_n293 & new_n366;
  assign new_n368 = ~px3 & new_n367;
  assign new_n369 = pz3 & ~new_n368;
  assign new_n370 = ~new_n365 & ~new_n369;
  assign pi9 = ~po0 | ~new_n370;
  assign pd5 = pm0 & pm3;
  assign new_n373 = ~pw1 & new_n295;
  assign new_n374 = pl0 & new_n297;
  assign new_n375 = new_n301 & ~new_n374;
  assign new_n376 = ~new_n373 & ~new_n375;
  assign new_n377 = ~pn0 & new_n376;
  assign new_n378 = new_n293 & new_n377;
  assign new_n379 = pl4 & ~px1;
  assign new_n380 = new_n377 & ~new_n379;
  assign new_n381 = pw1 & new_n376;
  assign new_n382 = ~new_n379 & new_n381;
  assign new_n383 = new_n310 & new_n381;
  assign new_n384 = new_n293 & new_n381;
  assign new_n385 = new_n294 & new_n376;
  assign new_n386 = ~new_n379 & new_n385;
  assign new_n387 = new_n310 & new_n385;
  assign new_n388 = new_n310 & new_n377;
  assign new_n389 = new_n293 & new_n385;
  assign new_n390 = ~new_n378 & ~new_n380;
  assign new_n391 = ~new_n382 & new_n390;
  assign new_n392 = ~new_n383 & ~new_n384;
  assign new_n393 = new_n391 & new_n392;
  assign new_n394 = ~new_n388 & ~new_n389;
  assign new_n395 = ~new_n386 & ~new_n387;
  assign new_n396 = new_n394 & new_n395;
  assign pf7 = ~new_n393 | ~new_n396;
  assign pg6 = ~pl4 | ~pl1;
  assign new_n399 = ~py3 & new_n358;
  assign new_n400 = pl4 & new_n399;
  assign new_n401 = ~pq0 & ~new_n400;
  assign new_n402 = pn0 & new_n401;
  assign new_n403 = ~new_n288 & new_n401;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = pl4 & new_n358;
  assign new_n406 = py3 & ~new_n405;
  assign new_n407 = ~new_n404 & ~new_n406;
  assign ph9 = ~po0 | ~new_n407;
  assign new_n409 = ~pq0 & pz2;
  assign new_n410 = new_n310 & new_n329;
  assign new_n411 = ~pm0 & new_n410;
  assign new_n412 = ~new_n294 & ~new_n411;
  assign new_n413 = new_n409 & new_n412;
  assign new_n414 = po0 & new_n413;
  assign new_n415 = new_n288 & new_n297;
  assign new_n416 = pp & ~pm0;
  assign new_n417 = ~pn0 & new_n416;
  assign new_n418 = new_n329 & new_n415;
  assign new_n419 = new_n417 & new_n418;
  assign pi8 = new_n414 | new_n419;
  assign pd6 = ~pi1 | ~pl4;
  assign new_n422 = ~pv1 & new_n295;
  assign new_n423 = pk0 & new_n297;
  assign new_n424 = new_n301 & ~new_n423;
  assign new_n425 = ~new_n422 & ~new_n424;
  assign new_n426 = ~pn0 & new_n425;
  assign new_n427 = new_n293 & new_n426;
  assign new_n428 = pl4 & ~pw1;
  assign new_n429 = new_n426 & ~new_n428;
  assign new_n430 = pv1 & new_n425;
  assign new_n431 = ~new_n428 & new_n430;
  assign new_n432 = new_n310 & new_n430;
  assign new_n433 = new_n293 & new_n430;
  assign new_n434 = new_n294 & new_n425;
  assign new_n435 = ~new_n428 & new_n434;
  assign new_n436 = new_n310 & new_n434;
  assign new_n437 = new_n310 & new_n426;
  assign new_n438 = new_n293 & new_n434;
  assign new_n439 = ~new_n427 & ~new_n429;
  assign new_n440 = ~new_n431 & new_n439;
  assign new_n441 = ~new_n432 & ~new_n433;
  assign new_n442 = new_n440 & new_n441;
  assign new_n443 = ~new_n437 & ~new_n438;
  assign new_n444 = ~new_n435 & ~new_n436;
  assign new_n445 = new_n443 & new_n444;
  assign pe7 = ~new_n442 | ~new_n445;
  assign pg5 = pm0 & pp3;
  assign new_n448 = pa3 & ~pq0;
  assign new_n449 = ~pk1 & ~pj1;
  assign new_n450 = ~pl1 & new_n449;
  assign new_n451 = pe4 & pf4;
  assign new_n452 = ~pg4 & new_n451;
  assign new_n453 = ~ph4 & new_n452;
  assign new_n454 = pk1 & pj1;
  assign new_n455 = ph1 & ~px0;
  assign new_n456 = pi1 & ~py0;
  assign new_n457 = pb1 & ~pk1;
  assign new_n458 = ~pj1 & new_n457;
  assign new_n459 = pa1 & ~pl1;
  assign new_n460 = pz0 & new_n459;
  assign new_n461 = pa1 & pb1;
  assign new_n462 = ~pj1 & new_n461;
  assign new_n463 = pz0 & new_n457;
  assign new_n464 = pz0 & new_n461;
  assign new_n465 = ~pk1 & ~pl1;
  assign new_n466 = ~pj1 & new_n465;
  assign new_n467 = ~pj1 & new_n459;
  assign new_n468 = pz0 & new_n465;
  assign new_n469 = ~new_n467 & ~new_n468;
  assign new_n470 = ~new_n464 & ~new_n466;
  assign new_n471 = new_n469 & new_n470;
  assign new_n472 = ~new_n458 & ~new_n460;
  assign new_n473 = ~new_n462 & ~new_n463;
  assign new_n474 = new_n472 & new_n473;
  assign new_n475 = new_n471 & new_n474;
  assign new_n476 = ~new_n455 & ~new_n456;
  assign new_n477 = ~new_n475 & new_n476;
  assign new_n478 = ~new_n288 & ~new_n454;
  assign new_n479 = ~new_n477 & new_n478;
  assign new_n480 = ~new_n453 & new_n479;
  assign new_n481 = ~pj1 & new_n480;
  assign new_n482 = ~pl1 & new_n480;
  assign new_n483 = ~new_n481 & ~new_n482;
  assign new_n484 = pk1 & pl1;
  assign new_n485 = ~new_n483 & ~new_n484;
  assign new_n486 = pk4 & new_n485;
  assign new_n487 = ~pi1 & new_n465;
  assign new_n488 = ~pj1 & new_n487;
  assign new_n489 = new_n450 & new_n486;
  assign new_n490 = new_n488 & new_n489;
  assign new_n491 = ~pi1 & new_n486;
  assign new_n492 = new_n488 & new_n491;
  assign new_n493 = ~ph1 & new_n489;
  assign new_n494 = ~ph1 & new_n491;
  assign new_n495 = ~new_n490 & ~new_n492;
  assign new_n496 = ~new_n493 & ~new_n494;
  assign new_n497 = new_n495 & new_n496;
  assign new_n498 = new_n448 & new_n497;
  assign new_n499 = po0 & new_n498;
  assign new_n500 = pb3 & ~new_n453;
  assign new_n501 = pk4 & new_n500;
  assign new_n502 = ph1 & ~new_n488;
  assign new_n503 = pi1 & ~new_n450;
  assign new_n504 = pj1 & pl1;
  assign new_n505 = ~new_n484 & ~new_n504;
  assign new_n506 = ~new_n454 & new_n505;
  assign new_n507 = ph1 & new_n506;
  assign new_n508 = ~new_n450 & new_n506;
  assign new_n509 = pi1 & new_n506;
  assign new_n510 = ~new_n507 & ~new_n508;
  assign new_n511 = ~new_n509 & new_n510;
  assign new_n512 = ~new_n502 & ~new_n503;
  assign new_n513 = ~new_n511 & new_n512;
  assign new_n514 = new_n297 & ~new_n477;
  assign new_n515 = new_n501 & new_n513;
  assign new_n516 = new_n514 & new_n515;
  assign pj8 = new_n499 | new_n516;
  assign new_n518 = ~pq0 & ~new_n293;
  assign new_n519 = ~px3 & new_n518;
  assign new_n520 = pz3 & py3;
  assign new_n521 = ~pa4 & ~pb4;
  assign new_n522 = pl4 & new_n521;
  assign new_n523 = new_n520 & new_n522;
  assign new_n524 = po0 & new_n523;
  assign new_n525 = ~new_n310 & new_n519;
  assign new_n526 = new_n524 & new_n525;
  assign new_n527 = pb4 & ~pq0;
  assign new_n528 = py3 & ~px3;
  assign new_n529 = pl4 & new_n289;
  assign new_n530 = new_n528 & new_n529;
  assign new_n531 = ~new_n293 & new_n530;
  assign new_n532 = ~new_n310 & ~new_n531;
  assign new_n533 = new_n527 & new_n532;
  assign new_n534 = po0 & new_n533;
  assign new_n535 = pm0 & ~pn0;
  assign new_n536 = po0 & new_n535;
  assign new_n537 = ~pq0 & new_n536;
  assign new_n538 = new_n288 & new_n537;
  assign new_n539 = ~new_n526 & ~new_n534;
  assign pk9 = new_n538 | ~new_n539;
  assign new_n541 = ~pu1 & new_n295;
  assign new_n542 = pm0 & new_n297;
  assign new_n543 = new_n301 & ~new_n542;
  assign new_n544 = ~new_n541 & ~new_n543;
  assign new_n545 = ~pn0 & new_n544;
  assign new_n546 = new_n293 & new_n545;
  assign new_n547 = pl4 & ~pv1;
  assign new_n548 = new_n545 & ~new_n547;
  assign new_n549 = pu1 & new_n544;
  assign new_n550 = ~new_n547 & new_n549;
  assign new_n551 = new_n310 & new_n549;
  assign new_n552 = new_n293 & new_n549;
  assign new_n553 = new_n294 & new_n544;
  assign new_n554 = ~new_n547 & new_n553;
  assign new_n555 = new_n310 & new_n553;
  assign new_n556 = new_n310 & new_n545;
  assign new_n557 = new_n293 & new_n553;
  assign new_n558 = ~new_n546 & ~new_n548;
  assign new_n559 = ~new_n550 & new_n558;
  assign new_n560 = ~new_n551 & ~new_n552;
  assign new_n561 = new_n559 & new_n560;
  assign new_n562 = ~new_n556 & ~new_n557;
  assign new_n563 = ~new_n554 & ~new_n555;
  assign new_n564 = new_n562 & new_n563;
  assign pd7 = ~new_n561 | ~new_n564;
  assign pe6 = ~pl4 | ~pj1;
  assign pf5 = po3 & pm0;
  assign new_n568 = pl4 & new_n520;
  assign new_n569 = new_n358 & new_n568;
  assign new_n570 = ~new_n288 & new_n569;
  assign new_n571 = pn0 & new_n288;
  assign new_n572 = ~new_n570 & ~new_n571;
  assign new_n573 = new_n329 & new_n572;
  assign new_n574 = pa4 & new_n573;
  assign new_n575 = new_n288 & new_n573;
  assign new_n576 = new_n288 & new_n572;
  assign new_n577 = pm0 & new_n576;
  assign new_n578 = ~new_n288 & new_n572;
  assign new_n579 = pa4 & new_n578;
  assign new_n580 = pa4 & new_n572;
  assign new_n581 = pm0 & new_n580;
  assign new_n582 = ~new_n574 & ~new_n575;
  assign new_n583 = ~new_n577 & new_n582;
  assign new_n584 = ~new_n579 & ~new_n581;
  assign new_n585 = new_n583 & new_n584;
  assign new_n586 = ~pn0 & new_n585;
  assign new_n587 = ~new_n359 & new_n586;
  assign new_n588 = ~new_n529 & new_n586;
  assign new_n589 = ~pa4 & new_n585;
  assign new_n590 = ~new_n529 & new_n589;
  assign new_n591 = new_n310 & new_n589;
  assign new_n592 = ~new_n359 & new_n589;
  assign new_n593 = ~new_n293 & new_n568;
  assign new_n594 = ~px3 & new_n593;
  assign new_n595 = new_n585 & new_n594;
  assign new_n596 = ~new_n529 & new_n595;
  assign new_n597 = new_n310 & new_n595;
  assign new_n598 = new_n310 & new_n586;
  assign new_n599 = ~new_n359 & new_n595;
  assign new_n600 = ~new_n587 & ~new_n588;
  assign new_n601 = ~new_n590 & new_n600;
  assign new_n602 = ~new_n591 & ~new_n592;
  assign new_n603 = new_n601 & new_n602;
  assign new_n604 = ~new_n598 & ~new_n599;
  assign new_n605 = ~new_n596 & ~new_n597;
  assign new_n606 = new_n604 & new_n605;
  assign new_n607 = new_n603 & new_n606;
  assign new_n608 = po0 & new_n607;
  assign pj9 = ~pq0 & new_n608;
  assign new_n610 = pb3 & ~pq0;
  assign new_n611 = new_n497 & new_n610;
  assign new_n612 = po0 & new_n611;
  assign new_n613 = pc3 & ~new_n453;
  assign new_n614 = pk4 & new_n613;
  assign new_n615 = new_n513 & new_n614;
  assign new_n616 = new_n514 & new_n615;
  assign pk8 = new_n612 | new_n616;
  assign new_n618 = ~pj3 & pl0;
  assign new_n619 = pk0 & new_n618;
  assign new_n620 = ~pj3 & ~pl0;
  assign new_n621 = ~pk0 & new_n620;
  assign new_n622 = ~new_n619 & ~new_n621;
  assign new_n623 = pm0 & new_n622;
  assign new_n624 = pl0 & new_n623;
  assign new_n625 = pk0 & new_n624;
  assign new_n626 = ~pl0 & new_n623;
  assign new_n627 = ~pk0 & new_n626;
  assign new_n628 = pr3 & new_n623;
  assign new_n629 = ~new_n625 & ~new_n627;
  assign pa5 = new_n628 | ~new_n629;
  assign new_n631 = pm1 & pl1;
  assign pb6 = pk4 | ~new_n631;
  assign new_n633 = ~pt1 & new_n295;
  assign new_n634 = pd0 & new_n297;
  assign new_n635 = new_n301 & ~new_n634;
  assign new_n636 = ~new_n633 & ~new_n635;
  assign new_n637 = ~pn0 & new_n636;
  assign new_n638 = new_n293 & new_n637;
  assign new_n639 = pl4 & ~pu1;
  assign new_n640 = new_n637 & ~new_n639;
  assign new_n641 = pt1 & new_n636;
  assign new_n642 = ~new_n639 & new_n641;
  assign new_n643 = new_n310 & new_n641;
  assign new_n644 = new_n293 & new_n641;
  assign new_n645 = new_n294 & new_n636;
  assign new_n646 = ~new_n639 & new_n645;
  assign new_n647 = new_n310 & new_n645;
  assign new_n648 = new_n310 & new_n637;
  assign new_n649 = new_n293 & new_n645;
  assign new_n650 = ~new_n638 & ~new_n640;
  assign new_n651 = ~new_n642 & new_n650;
  assign new_n652 = ~new_n643 & ~new_n644;
  assign new_n653 = new_n651 & new_n652;
  assign new_n654 = ~new_n648 & ~new_n649;
  assign new_n655 = ~new_n646 & ~new_n647;
  assign new_n656 = new_n654 & new_n655;
  assign pc7 = ~new_n653 | ~new_n656;
  assign new_n658 = pc3 & ~pq0;
  assign new_n659 = new_n497 & new_n658;
  assign new_n660 = po0 & new_n659;
  assign new_n661 = pd3 & ~new_n453;
  assign new_n662 = pk4 & new_n661;
  assign new_n663 = new_n513 & new_n662;
  assign new_n664 = new_n514 & new_n663;
  assign pl8 = new_n660 | new_n664;
  assign new_n666 = ~pq0 & new_n288;
  assign new_n667 = po0 & new_n666;
  assign new_n668 = ~pn0 & new_n667;
  assign new_n669 = ~pg1 & ~pq0;
  assign new_n670 = pd4 & pk4;
  assign new_n671 = ~new_n477 & new_n670;
  assign new_n672 = ~new_n453 & new_n671;
  assign new_n673 = ~new_n453 & ~new_n477;
  assign new_n674 = pk4 & new_n673;
  assign new_n675 = ~pd4 & ~new_n674;
  assign new_n676 = ~new_n672 & ~new_n675;
  assign new_n677 = new_n669 & new_n676;
  assign new_n678 = po0 & new_n677;
  assign pm9 = new_n668 | new_n678;
  assign new_n680 = ~ps1 & new_n295;
  assign new_n681 = pe0 & new_n297;
  assign new_n682 = new_n301 & ~new_n681;
  assign new_n683 = ~new_n680 & ~new_n682;
  assign new_n684 = ~pn0 & new_n683;
  assign new_n685 = new_n293 & new_n684;
  assign new_n686 = pl4 & ~pt1;
  assign new_n687 = new_n684 & ~new_n686;
  assign new_n688 = ps1 & new_n683;
  assign new_n689 = ~new_n686 & new_n688;
  assign new_n690 = new_n310 & new_n688;
  assign new_n691 = new_n293 & new_n688;
  assign new_n692 = new_n294 & new_n683;
  assign new_n693 = ~new_n686 & new_n692;
  assign new_n694 = new_n310 & new_n692;
  assign new_n695 = new_n310 & new_n684;
  assign new_n696 = new_n293 & new_n692;
  assign new_n697 = ~new_n685 & ~new_n687;
  assign new_n698 = ~new_n689 & new_n697;
  assign new_n699 = ~new_n690 & ~new_n691;
  assign new_n700 = new_n698 & new_n699;
  assign new_n701 = ~new_n695 & ~new_n696;
  assign new_n702 = ~new_n693 & ~new_n694;
  assign new_n703 = new_n701 & new_n702;
  assign pb7 = ~new_n700 | ~new_n703;
  assign pc6 = ~pl4 | ~ph1;
  assign new_n706 = ~pa4 & new_n520;
  assign new_n707 = ~pb4 & ~pc4;
  assign new_n708 = pl4 & new_n707;
  assign new_n709 = new_n706 & new_n708;
  assign new_n710 = po0 & new_n709;
  assign new_n711 = new_n525 & new_n710;
  assign new_n712 = pc4 & ~pq0;
  assign new_n713 = pz3 & new_n528;
  assign new_n714 = new_n522 & new_n713;
  assign new_n715 = ~new_n293 & new_n714;
  assign new_n716 = ~new_n310 & ~new_n715;
  assign new_n717 = new_n712 & new_n716;
  assign new_n718 = po0 & new_n717;
  assign new_n719 = po0 & new_n335;
  assign new_n720 = ~pq0 & new_n719;
  assign new_n721 = new_n288 & new_n720;
  assign new_n722 = ~new_n711 & ~new_n718;
  assign pl9 = new_n721 | ~new_n722;
  assign new_n724 = pd3 & ~pq0;
  assign new_n725 = new_n497 & new_n724;
  assign new_n726 = po0 & new_n725;
  assign new_n727 = pe3 & ~new_n453;
  assign new_n728 = pk4 & new_n727;
  assign new_n729 = new_n513 & new_n728;
  assign new_n730 = new_n514 & new_n729;
  assign pm8 = new_n726 | new_n730;
  assign new_n732 = ~pr1 & new_n295;
  assign new_n733 = pf0 & new_n297;
  assign new_n734 = new_n301 & ~new_n733;
  assign new_n735 = ~new_n732 & ~new_n734;
  assign new_n736 = ~pn0 & new_n735;
  assign new_n737 = new_n293 & new_n736;
  assign new_n738 = pl4 & ~ps1;
  assign new_n739 = new_n736 & ~new_n738;
  assign new_n740 = pr1 & new_n735;
  assign new_n741 = ~new_n738 & new_n740;
  assign new_n742 = new_n310 & new_n740;
  assign new_n743 = new_n293 & new_n740;
  assign new_n744 = new_n294 & new_n735;
  assign new_n745 = ~new_n738 & new_n744;
  assign new_n746 = new_n310 & new_n744;
  assign new_n747 = new_n310 & new_n736;
  assign new_n748 = new_n293 & new_n744;
  assign new_n749 = ~new_n737 & ~new_n739;
  assign new_n750 = ~new_n741 & new_n749;
  assign new_n751 = ~new_n742 & ~new_n743;
  assign new_n752 = new_n750 & new_n751;
  assign new_n753 = ~new_n747 & ~new_n748;
  assign new_n754 = ~new_n745 & ~new_n746;
  assign new_n755 = new_n753 & new_n754;
  assign pa7 = ~new_n752 | ~new_n755;
  assign new_n757 = pl0 & ~pl3;
  assign new_n758 = pk0 & new_n757;
  assign new_n759 = ~pl0 & ~pl3;
  assign new_n760 = ~pk0 & new_n759;
  assign new_n761 = ~new_n758 & ~new_n760;
  assign new_n762 = pm0 & new_n761;
  assign new_n763 = pl0 & new_n762;
  assign new_n764 = pk0 & new_n763;
  assign new_n765 = ~pl0 & new_n762;
  assign new_n766 = ~pk0 & new_n765;
  assign new_n767 = pt3 & new_n762;
  assign new_n768 = ~new_n764 & ~new_n766;
  assign pc5 = new_n767 | ~new_n768;
  assign new_n770 = pe3 & ~pq0;
  assign new_n771 = new_n497 & new_n770;
  assign new_n772 = po0 & new_n771;
  assign new_n773 = pf3 & ~new_n453;
  assign new_n774 = pk4 & new_n773;
  assign new_n775 = new_n513 & new_n774;
  assign new_n776 = new_n514 & new_n775;
  assign pn8 = new_n772 | new_n776;
  assign new_n778 = ~pd4 & ~new_n453;
  assign new_n779 = pe4 & ~pf4;
  assign new_n780 = pk4 & new_n779;
  assign new_n781 = new_n778 & new_n780;
  assign new_n782 = ~new_n477 & new_n781;
  assign new_n783 = ~new_n310 & ~new_n782;
  assign new_n784 = ~pg1 & new_n783;
  assign new_n785 = ~pq0 & new_n784;
  assign new_n786 = ~pd4 & pe4;
  assign new_n787 = pk4 & new_n786;
  assign new_n788 = ~new_n477 & new_n787;
  assign new_n789 = ~new_n453 & new_n788;
  assign new_n790 = pf4 & ~new_n789;
  assign new_n791 = new_n785 & ~new_n790;
  assign po9 = ~po0 | ~new_n791;
  assign new_n793 = pk1 & pm1;
  assign pa6 = pk4 | ~new_n793;
  assign new_n795 = ~pk3 & pl0;
  assign new_n796 = pk0 & new_n795;
  assign new_n797 = ~pk3 & ~pl0;
  assign new_n798 = ~pk0 & new_n797;
  assign new_n799 = ~new_n796 & ~new_n798;
  assign new_n800 = pm0 & new_n799;
  assign new_n801 = pl0 & new_n800;
  assign new_n802 = pk0 & new_n801;
  assign new_n803 = ~pl0 & new_n800;
  assign new_n804 = ~pk0 & new_n803;
  assign new_n805 = ps3 & new_n800;
  assign new_n806 = ~new_n802 & ~new_n804;
  assign pb5 = new_n805 | ~new_n806;
  assign new_n808 = ~pd4 & ~pe4;
  assign new_n809 = pk4 & new_n808;
  assign new_n810 = ~new_n477 & new_n809;
  assign new_n811 = ~new_n453 & new_n810;
  assign new_n812 = ~new_n310 & ~new_n811;
  assign new_n813 = ~pg1 & new_n812;
  assign new_n814 = ~pq0 & new_n813;
  assign new_n815 = ~pd4 & pk4;
  assign new_n816 = ~new_n477 & new_n815;
  assign new_n817 = ~new_n453 & new_n816;
  assign new_n818 = pe4 & ~new_n817;
  assign new_n819 = new_n814 & ~new_n818;
  assign pn9 = ~po0 | ~new_n819;
  assign new_n821 = pf3 & ~pq0;
  assign new_n822 = new_n497 & new_n821;
  assign new_n823 = po0 & new_n822;
  assign new_n824 = pg3 & ~new_n453;
  assign new_n825 = pk4 & new_n824;
  assign new_n826 = new_n513 & new_n825;
  assign new_n827 = new_n514 & new_n826;
  assign po8 = new_n823 | new_n827;
  assign new_n829 = ~pq0 & pr3;
  assign new_n830 = new_n497 & new_n829;
  assign new_n831 = po0 & new_n830;
  assign new_n832 = ps3 & ~new_n453;
  assign new_n833 = pk4 & new_n832;
  assign new_n834 = new_n513 & new_n833;
  assign new_n835 = new_n514 & new_n834;
  assign pa9 = new_n831 | new_n835;
  assign new_n837 = ~pf1 & ~pi4;
  assign new_n838 = pf1 & pi4;
  assign pn6 = new_n837 | new_n838;
  assign new_n840 = ~pf2 & new_n295;
  assign new_n841 = py & new_n297;
  assign new_n842 = new_n301 & ~new_n841;
  assign new_n843 = ~new_n840 & ~new_n842;
  assign new_n844 = ~pn0 & new_n843;
  assign new_n845 = new_n293 & new_n844;
  assign new_n846 = ~pg2 & pl4;
  assign new_n847 = new_n844 & ~new_n846;
  assign new_n848 = pf2 & new_n843;
  assign new_n849 = ~new_n846 & new_n848;
  assign new_n850 = new_n310 & new_n848;
  assign new_n851 = new_n293 & new_n848;
  assign new_n852 = new_n294 & new_n843;
  assign new_n853 = ~new_n846 & new_n852;
  assign new_n854 = new_n310 & new_n852;
  assign new_n855 = new_n310 & new_n844;
  assign new_n856 = new_n293 & new_n852;
  assign new_n857 = ~new_n845 & ~new_n847;
  assign new_n858 = ~new_n849 & new_n857;
  assign new_n859 = ~new_n850 & ~new_n851;
  assign new_n860 = new_n858 & new_n859;
  assign new_n861 = ~new_n855 & ~new_n856;
  assign new_n862 = ~new_n853 & ~new_n854;
  assign new_n863 = new_n861 & new_n862;
  assign po7 = ~new_n860 | ~new_n863;
  assign new_n865 = pl0 & ph;
  assign new_n866 = pp & ~pl0;
  assign new_n867 = pk0 & new_n866;
  assign new_n868 = ~pk0 & ph;
  assign new_n869 = ~new_n865 & ~new_n867;
  assign new_n870 = ~new_n868 & new_n869;
  assign new_n871 = new_n310 & new_n870;
  assign new_n872 = ~pm0 & new_n871;
  assign new_n873 = pl4 & ~ps2;
  assign new_n874 = ~new_n336 & new_n873;
  assign new_n875 = ~new_n293 & new_n874;
  assign new_n876 = ~pm0 & new_n310;
  assign new_n877 = ~new_n294 & ~new_n876;
  assign new_n878 = ~pr2 & new_n877;
  assign new_n879 = ~new_n872 & ~new_n875;
  assign new_n880 = ~new_n878 & new_n879;
  assign new_n881 = po0 & new_n880;
  assign pa8 = ~pq0 & new_n881;
  assign pl5 = pg1 & ~pj4;
  assign new_n884 = ~pe2 & new_n295;
  assign new_n885 = px & new_n297;
  assign new_n886 = new_n301 & ~new_n885;
  assign new_n887 = ~new_n884 & ~new_n886;
  assign new_n888 = ~pn0 & new_n887;
  assign new_n889 = new_n293 & new_n888;
  assign new_n890 = ~pf2 & pl4;
  assign new_n891 = new_n888 & ~new_n890;
  assign new_n892 = pe2 & new_n887;
  assign new_n893 = ~new_n890 & new_n892;
  assign new_n894 = new_n310 & new_n892;
  assign new_n895 = new_n293 & new_n892;
  assign new_n896 = new_n294 & new_n887;
  assign new_n897 = ~new_n890 & new_n896;
  assign new_n898 = new_n310 & new_n896;
  assign new_n899 = new_n310 & new_n888;
  assign new_n900 = new_n293 & new_n896;
  assign new_n901 = ~new_n889 & ~new_n891;
  assign new_n902 = ~new_n893 & new_n901;
  assign new_n903 = ~new_n894 & ~new_n895;
  assign new_n904 = new_n902 & new_n903;
  assign new_n905 = ~new_n899 & ~new_n900;
  assign new_n906 = ~new_n897 & ~new_n898;
  assign new_n907 = new_n905 & new_n906;
  assign pn7 = ~new_n904 | ~new_n907;
  assign new_n909 = px3 & new_n289;
  assign new_n910 = py3 & new_n909;
  assign new_n911 = ~pb4 & new_n910;
  assign po6 = ~pc4 & new_n911;
  assign new_n913 = pl4 & pt2;
  assign new_n914 = ps2 & ~new_n332;
  assign new_n915 = ~pl4 & new_n914;
  assign new_n916 = pi & new_n337;
  assign new_n917 = ~new_n915 & ~new_n916;
  assign new_n918 = ~new_n913 & new_n917;
  assign new_n919 = ~new_n293 & new_n918;
  assign new_n920 = new_n293 & new_n917;
  assign new_n921 = ~ps2 & new_n920;
  assign new_n922 = ~ps2 & new_n918;
  assign new_n923 = new_n351 & new_n917;
  assign new_n924 = ~new_n919 & ~new_n921;
  assign new_n925 = ~new_n922 & ~new_n923;
  assign new_n926 = new_n924 & new_n925;
  assign new_n927 = po0 & new_n926;
  assign pb8 = ~pq0 & new_n927;
  assign new_n929 = ~pq0 & pt3;
  assign new_n930 = new_n497 & new_n929;
  assign new_n931 = po0 & new_n930;
  assign new_n932 = pu3 & ~new_n453;
  assign new_n933 = pk4 & new_n932;
  assign new_n934 = new_n513 & new_n933;
  assign new_n935 = new_n514 & new_n934;
  assign pc9 = new_n931 | new_n935;
  assign new_n937 = ~pd2 & new_n295;
  assign new_n938 = pw & new_n297;
  assign new_n939 = new_n301 & ~new_n938;
  assign new_n940 = ~new_n937 & ~new_n939;
  assign new_n941 = ~pn0 & new_n940;
  assign new_n942 = new_n293 & new_n941;
  assign new_n943 = ~pe2 & pl4;
  assign new_n944 = new_n941 & ~new_n943;
  assign new_n945 = pd2 & new_n940;
  assign new_n946 = ~new_n943 & new_n945;
  assign new_n947 = new_n310 & new_n945;
  assign new_n948 = new_n293 & new_n945;
  assign new_n949 = new_n294 & new_n940;
  assign new_n950 = ~new_n943 & new_n949;
  assign new_n951 = new_n310 & new_n949;
  assign new_n952 = new_n310 & new_n941;
  assign new_n953 = new_n293 & new_n949;
  assign new_n954 = ~new_n942 & ~new_n944;
  assign new_n955 = ~new_n946 & new_n954;
  assign new_n956 = ~new_n947 & ~new_n948;
  assign new_n957 = new_n955 & new_n956;
  assign new_n958 = ~new_n952 & ~new_n953;
  assign new_n959 = ~new_n950 & ~new_n951;
  assign new_n960 = new_n958 & new_n959;
  assign pm7 = ~new_n957 | ~new_n960;
  assign new_n962 = pi1 & ~pn0;
  assign po5 = pk4 | ~new_n962;
  assign new_n964 = ps3 & ~pq0;
  assign new_n965 = new_n497 & new_n964;
  assign new_n966 = po0 & new_n965;
  assign new_n967 = pt3 & ~new_n453;
  assign new_n968 = pk4 & new_n967;
  assign new_n969 = new_n513 & new_n968;
  assign new_n970 = new_n514 & new_n969;
  assign pb9 = new_n966 | new_n970;
  assign new_n972 = pl4 & pu2;
  assign new_n973 = pt2 & ~new_n332;
  assign new_n974 = ~pl4 & new_n973;
  assign new_n975 = pj & new_n337;
  assign new_n976 = ~new_n974 & ~new_n975;
  assign new_n977 = ~new_n972 & new_n976;
  assign new_n978 = ~new_n293 & new_n977;
  assign new_n979 = new_n293 & new_n976;
  assign new_n980 = ~pt2 & new_n979;
  assign new_n981 = ~pt2 & new_n977;
  assign new_n982 = new_n351 & new_n976;
  assign new_n983 = ~new_n978 & ~new_n980;
  assign new_n984 = ~new_n981 & ~new_n982;
  assign new_n985 = new_n983 & new_n984;
  assign new_n986 = po0 & new_n985;
  assign pc8 = ~pq0 & new_n986;
  assign new_n988 = ~pc2 & new_n295;
  assign new_n989 = pv & new_n297;
  assign new_n990 = new_n301 & ~new_n989;
  assign new_n991 = ~new_n988 & ~new_n990;
  assign new_n992 = ~pn0 & new_n991;
  assign new_n993 = new_n293 & new_n992;
  assign new_n994 = ~pd2 & pl4;
  assign new_n995 = new_n992 & ~new_n994;
  assign new_n996 = pc2 & new_n991;
  assign new_n997 = ~new_n994 & new_n996;
  assign new_n998 = new_n310 & new_n996;
  assign new_n999 = new_n293 & new_n996;
  assign new_n1000 = new_n294 & new_n991;
  assign new_n1001 = ~new_n994 & new_n1000;
  assign new_n1002 = new_n310 & new_n1000;
  assign new_n1003 = new_n310 & new_n992;
  assign new_n1004 = new_n293 & new_n1000;
  assign new_n1005 = ~new_n993 & ~new_n995;
  assign new_n1006 = ~new_n997 & new_n1005;
  assign new_n1007 = ~new_n998 & ~new_n999;
  assign new_n1008 = new_n1006 & new_n1007;
  assign new_n1009 = ~new_n1003 & ~new_n1004;
  assign new_n1010 = ~new_n1001 & ~new_n1002;
  assign new_n1011 = new_n1009 & new_n1010;
  assign pl7 = ~new_n1008 | ~new_n1011;
  assign new_n1013 = ph1 & ~pn0;
  assign pn5 = pk4 | ~new_n1013;
  assign new_n1015 = pl4 & pv2;
  assign new_n1016 = pu2 & ~new_n332;
  assign new_n1017 = ~pl4 & new_n1016;
  assign new_n1018 = pk & new_n337;
  assign new_n1019 = ~new_n1017 & ~new_n1018;
  assign new_n1020 = ~new_n1015 & new_n1019;
  assign new_n1021 = ~new_n293 & new_n1020;
  assign new_n1022 = new_n293 & new_n1019;
  assign new_n1023 = ~pu2 & new_n1022;
  assign new_n1024 = ~pu2 & new_n1020;
  assign new_n1025 = new_n351 & new_n1019;
  assign new_n1026 = ~new_n1021 & ~new_n1023;
  assign new_n1027 = ~new_n1024 & ~new_n1025;
  assign new_n1028 = new_n1026 & new_n1027;
  assign new_n1029 = po0 & new_n1028;
  assign pd8 = ~pq0 & new_n1029;
  assign new_n1031 = ~pq0 & pv3;
  assign new_n1032 = new_n497 & new_n1031;
  assign new_n1033 = po0 & new_n1032;
  assign new_n1034 = pw3 & ~new_n453;
  assign new_n1035 = pk4 & new_n1034;
  assign new_n1036 = new_n513 & new_n1035;
  assign new_n1037 = new_n514 & new_n1036;
  assign pe9 = new_n1033 | new_n1037;
  assign pi5 = pm0 & pr3;
  assign new_n1040 = ~pb2 & new_n295;
  assign new_n1041 = pu & new_n297;
  assign new_n1042 = new_n301 & ~new_n1041;
  assign new_n1043 = ~new_n1040 & ~new_n1042;
  assign new_n1044 = ~pn0 & new_n1043;
  assign new_n1045 = new_n293 & new_n1044;
  assign new_n1046 = ~pc2 & pl4;
  assign new_n1047 = new_n1044 & ~new_n1046;
  assign new_n1048 = pb2 & new_n1043;
  assign new_n1049 = ~new_n1046 & new_n1048;
  assign new_n1050 = new_n310 & new_n1048;
  assign new_n1051 = new_n293 & new_n1048;
  assign new_n1052 = new_n294 & new_n1043;
  assign new_n1053 = ~new_n1046 & new_n1052;
  assign new_n1054 = new_n310 & new_n1052;
  assign new_n1055 = new_n310 & new_n1044;
  assign new_n1056 = new_n293 & new_n1052;
  assign new_n1057 = ~new_n1045 & ~new_n1047;
  assign new_n1058 = ~new_n1049 & new_n1057;
  assign new_n1059 = ~new_n1050 & ~new_n1051;
  assign new_n1060 = new_n1058 & new_n1059;
  assign new_n1061 = ~new_n1055 & ~new_n1056;
  assign new_n1062 = ~new_n1053 & ~new_n1054;
  assign new_n1063 = new_n1061 & new_n1062;
  assign pk7 = ~new_n1060 | ~new_n1063;
  assign new_n1065 = ~pq0 & pu3;
  assign new_n1066 = new_n497 & new_n1065;
  assign new_n1067 = po0 & new_n1066;
  assign new_n1068 = pv3 & ~new_n453;
  assign new_n1069 = pk4 & new_n1068;
  assign new_n1070 = new_n513 & new_n1069;
  assign new_n1071 = new_n514 & new_n1070;
  assign pd9 = new_n1067 | new_n1071;
  assign new_n1073 = pl4 & pw2;
  assign new_n1074 = pv2 & ~new_n332;
  assign new_n1075 = ~pl4 & new_n1074;
  assign new_n1076 = pl & new_n337;
  assign new_n1077 = ~new_n1075 & ~new_n1076;
  assign new_n1078 = ~new_n1073 & new_n1077;
  assign new_n1079 = ~new_n293 & new_n1078;
  assign new_n1080 = new_n293 & new_n1077;
  assign new_n1081 = ~pv2 & new_n1080;
  assign new_n1082 = ~pv2 & new_n1078;
  assign new_n1083 = new_n351 & new_n1077;
  assign new_n1084 = ~new_n1079 & ~new_n1081;
  assign new_n1085 = ~new_n1082 & ~new_n1083;
  assign new_n1086 = new_n1084 & new_n1085;
  assign new_n1087 = po0 & new_n1086;
  assign pe8 = ~pq0 & new_n1087;
  assign ph5 = pm0 & pq3;
  assign new_n1090 = ~pa2 & new_n295;
  assign new_n1091 = pt & new_n297;
  assign new_n1092 = new_n301 & ~new_n1091;
  assign new_n1093 = ~new_n1090 & ~new_n1092;
  assign new_n1094 = ~pn0 & new_n1093;
  assign new_n1095 = new_n293 & new_n1094;
  assign new_n1096 = ~pb2 & pl4;
  assign new_n1097 = new_n1094 & ~new_n1096;
  assign new_n1098 = pa2 & new_n1093;
  assign new_n1099 = ~new_n1096 & new_n1098;
  assign new_n1100 = new_n310 & new_n1098;
  assign new_n1101 = new_n293 & new_n1098;
  assign new_n1102 = new_n294 & new_n1093;
  assign new_n1103 = ~new_n1096 & new_n1102;
  assign new_n1104 = new_n310 & new_n1102;
  assign new_n1105 = new_n310 & new_n1094;
  assign new_n1106 = new_n293 & new_n1102;
  assign new_n1107 = ~new_n1095 & ~new_n1097;
  assign new_n1108 = ~new_n1099 & new_n1107;
  assign new_n1109 = ~new_n1100 & ~new_n1101;
  assign new_n1110 = new_n1108 & new_n1109;
  assign new_n1111 = ~new_n1105 & ~new_n1106;
  assign new_n1112 = ~new_n1103 & ~new_n1104;
  assign new_n1113 = new_n1111 & new_n1112;
  assign pj7 = ~new_n1110 | ~new_n1113;
  assign new_n1115 = pl4 & px2;
  assign new_n1116 = pw2 & ~new_n332;
  assign new_n1117 = ~pl4 & new_n1116;
  assign new_n1118 = pm & new_n337;
  assign new_n1119 = ~new_n1117 & ~new_n1118;
  assign new_n1120 = ~new_n1115 & new_n1119;
  assign new_n1121 = ~new_n293 & new_n1120;
  assign new_n1122 = new_n293 & new_n1119;
  assign new_n1123 = ~pw2 & new_n1122;
  assign new_n1124 = ~pw2 & new_n1120;
  assign new_n1125 = new_n351 & new_n1119;
  assign new_n1126 = ~new_n1121 & ~new_n1123;
  assign new_n1127 = ~new_n1124 & ~new_n1125;
  assign new_n1128 = new_n1126 & new_n1127;
  assign new_n1129 = po0 & new_n1128;
  assign pf8 = ~pq0 & new_n1129;
  assign new_n1131 = px3 & ~new_n293;
  assign new_n1132 = pl4 & new_n1131;
  assign new_n1133 = ~new_n301 & ~new_n1132;
  assign new_n1134 = ~new_n293 & new_n1133;
  assign new_n1135 = pl4 & new_n1134;
  assign new_n1136 = px3 & new_n1133;
  assign pg9 = new_n1135 | new_n1136;
  assign new_n1138 = ~pz1 & new_n295;
  assign new_n1139 = ps & new_n297;
  assign new_n1140 = new_n301 & ~new_n1139;
  assign new_n1141 = ~new_n1138 & ~new_n1140;
  assign new_n1142 = ~pn0 & new_n1141;
  assign new_n1143 = new_n293 & new_n1142;
  assign new_n1144 = ~pa2 & pl4;
  assign new_n1145 = new_n1142 & ~new_n1144;
  assign new_n1146 = pz1 & new_n1141;
  assign new_n1147 = ~new_n1144 & new_n1146;
  assign new_n1148 = new_n310 & new_n1146;
  assign new_n1149 = new_n293 & new_n1146;
  assign new_n1150 = new_n294 & new_n1141;
  assign new_n1151 = ~new_n1144 & new_n1150;
  assign new_n1152 = new_n310 & new_n1150;
  assign new_n1153 = new_n310 & new_n1142;
  assign new_n1154 = new_n293 & new_n1150;
  assign new_n1155 = ~new_n1143 & ~new_n1145;
  assign new_n1156 = ~new_n1147 & new_n1155;
  assign new_n1157 = ~new_n1148 & ~new_n1149;
  assign new_n1158 = new_n1156 & new_n1157;
  assign new_n1159 = ~new_n1153 & ~new_n1154;
  assign new_n1160 = ~new_n1151 & ~new_n1152;
  assign new_n1161 = new_n1159 & new_n1160;
  assign pi7 = ~new_n1158 | ~new_n1161;
  assign pk5 = pm0 & pt3;
  assign new_n1164 = ~pq0 & pw3;
  assign new_n1165 = ~ph1 & new_n450;
  assign new_n1166 = ~pi1 & new_n1165;
  assign new_n1167 = pj1 & ~new_n465;
  assign new_n1168 = ~new_n1166 & ~new_n1167;
  assign new_n1169 = ~new_n477 & new_n1168;
  assign new_n1170 = ~pk1 & new_n1169;
  assign new_n1171 = ~pl1 & new_n1169;
  assign new_n1172 = ~new_n1170 & ~new_n1171;
  assign new_n1173 = ~new_n453 & ~new_n1172;
  assign new_n1174 = pk4 & new_n1173;
  assign new_n1175 = new_n450 & new_n1174;
  assign new_n1176 = new_n488 & new_n1175;
  assign new_n1177 = ~pi1 & new_n1174;
  assign new_n1178 = new_n488 & new_n1177;
  assign new_n1179 = ~ph1 & new_n1175;
  assign new_n1180 = ~ph1 & new_n1177;
  assign new_n1181 = ~new_n1176 & ~new_n1178;
  assign new_n1182 = ~new_n1179 & ~new_n1180;
  assign new_n1183 = new_n1181 & new_n1182;
  assign new_n1184 = new_n1164 & new_n1183;
  assign new_n1185 = po0 & new_n1184;
  assign new_n1186 = pt0 & new_n450;
  assign new_n1187 = pi1 & new_n1186;
  assign new_n1188 = ~pj1 & pv0;
  assign new_n1189 = pk1 & new_n1188;
  assign new_n1190 = ~pl1 & new_n1189;
  assign new_n1191 = ~new_n465 & ~new_n1190;
  assign new_n1192 = ~pw0 & new_n1191;
  assign new_n1193 = pj1 & new_n1191;
  assign new_n1194 = pj1 & ~new_n1190;
  assign new_n1195 = ~pu0 & new_n1194;
  assign new_n1196 = ~pj1 & ~new_n1190;
  assign new_n1197 = ~pw0 & new_n1196;
  assign new_n1198 = ~pw0 & ~new_n1190;
  assign new_n1199 = ~pu0 & new_n1198;
  assign new_n1200 = ~pk1 & pl1;
  assign new_n1201 = ~new_n1190 & ~new_n1200;
  assign new_n1202 = ~new_n465 & new_n1201;
  assign new_n1203 = ~pu0 & new_n1201;
  assign new_n1204 = ~pj1 & new_n1201;
  assign new_n1205 = ~new_n1203 & ~new_n1204;
  assign new_n1206 = ~new_n1199 & ~new_n1202;
  assign new_n1207 = new_n1205 & new_n1206;
  assign new_n1208 = ~new_n1192 & ~new_n1193;
  assign new_n1209 = ~new_n1195 & ~new_n1197;
  assign new_n1210 = new_n1208 & new_n1209;
  assign new_n1211 = new_n1207 & new_n1210;
  assign new_n1212 = ~pi1 & new_n1211;
  assign new_n1213 = ~new_n1187 & ~new_n1212;
  assign new_n1214 = ~ps0 & new_n1213;
  assign new_n1215 = ~pi1 & ph1;
  assign new_n1216 = new_n1213 & ~new_n1215;
  assign new_n1217 = ph1 & ~new_n1215;
  assign new_n1218 = ph1 & ~new_n450;
  assign new_n1219 = ph1 & ~ps0;
  assign new_n1220 = ~new_n450 & new_n1213;
  assign new_n1221 = ~new_n1214 & ~new_n1216;
  assign new_n1222 = ~new_n1217 & new_n1221;
  assign new_n1223 = ~new_n1218 & ~new_n1219;
  assign new_n1224 = ~new_n1220 & new_n1223;
  assign new_n1225 = new_n1222 & new_n1224;
  assign new_n1226 = new_n674 & new_n1225;
  assign new_n1227 = new_n297 & new_n1226;
  assign pf9 = new_n1185 | new_n1227;
  assign new_n1229 = pl4 & py2;
  assign new_n1230 = px2 & ~new_n332;
  assign new_n1231 = ~pl4 & new_n1230;
  assign new_n1232 = pn & new_n337;
  assign new_n1233 = ~new_n1231 & ~new_n1232;
  assign new_n1234 = ~new_n1229 & new_n1233;
  assign new_n1235 = ~new_n293 & new_n1234;
  assign new_n1236 = new_n293 & new_n1233;
  assign new_n1237 = ~px2 & new_n1236;
  assign new_n1238 = ~px2 & new_n1234;
  assign new_n1239 = new_n351 & new_n1233;
  assign new_n1240 = ~new_n1235 & ~new_n1237;
  assign new_n1241 = ~new_n1238 & ~new_n1239;
  assign new_n1242 = new_n1240 & new_n1241;
  assign new_n1243 = po0 & new_n1242;
  assign pg8 = ~pq0 & new_n1243;
  assign new_n1245 = ~py1 & new_n295;
  assign new_n1246 = pr & new_n297;
  assign new_n1247 = new_n301 & ~new_n1246;
  assign new_n1248 = ~new_n1245 & ~new_n1247;
  assign new_n1249 = ~pn0 & new_n1248;
  assign new_n1250 = new_n293 & new_n1249;
  assign new_n1251 = pl4 & ~pz1;
  assign new_n1252 = new_n1249 & ~new_n1251;
  assign new_n1253 = py1 & new_n1248;
  assign new_n1254 = ~new_n1251 & new_n1253;
  assign new_n1255 = new_n310 & new_n1253;
  assign new_n1256 = new_n293 & new_n1253;
  assign new_n1257 = new_n294 & new_n1248;
  assign new_n1258 = ~new_n1251 & new_n1257;
  assign new_n1259 = new_n310 & new_n1257;
  assign new_n1260 = new_n310 & new_n1249;
  assign new_n1261 = new_n293 & new_n1257;
  assign new_n1262 = ~new_n1250 & ~new_n1252;
  assign new_n1263 = ~new_n1254 & new_n1262;
  assign new_n1264 = ~new_n1255 & ~new_n1256;
  assign new_n1265 = new_n1263 & new_n1264;
  assign new_n1266 = ~new_n1260 & ~new_n1261;
  assign new_n1267 = ~new_n1258 & ~new_n1259;
  assign new_n1268 = new_n1266 & new_n1267;
  assign ph7 = ~new_n1265 | ~new_n1268;
  assign pj5 = pm0 & ps3;
  assign new_n1271 = ~pc4 & new_n521;
  assign new_n1272 = py3 & new_n1271;
  assign new_n1273 = pz3 & new_n1272;
  assign new_n1274 = ~new_n520 & new_n1273;
  assign new_n1275 = ~new_n1271 & new_n1273;
  assign new_n1276 = pn1 & ~new_n1271;
  assign new_n1277 = pf1 & ~pi4;
  assign new_n1278 = ~pf1 & pi4;
  assign new_n1279 = ~new_n1277 & ~new_n1278;
  assign new_n1280 = pn1 & new_n1279;
  assign new_n1281 = pn1 & ~new_n520;
  assign new_n1282 = new_n1273 & new_n1279;
  assign new_n1283 = ~new_n1274 & ~new_n1275;
  assign new_n1284 = ~new_n1276 & new_n1283;
  assign new_n1285 = ~new_n1280 & ~new_n1281;
  assign new_n1286 = ~new_n1282 & new_n1285;
  assign pu5 = ~new_n1284 | ~new_n1286;
  assign new_n1288 = ~pg4 & ~ph4;
  assign new_n1289 = pe4 & new_n1288;
  assign new_n1290 = pf4 & new_n1289;
  assign new_n1291 = ph1 & ~new_n1290;
  assign new_n1292 = ~px0 & new_n1291;
  assign new_n1293 = pi1 & ~new_n1290;
  assign new_n1294 = ~py0 & new_n1293;
  assign new_n1295 = ~pg1 & new_n451;
  assign new_n1296 = pd4 & new_n1295;
  assign new_n1297 = ~pg4 & new_n1296;
  assign new_n1298 = ~ph4 & new_n1297;
  assign new_n1299 = new_n1290 & ~new_n1298;
  assign new_n1300 = pl1 & ~new_n1298;
  assign new_n1301 = ~pb1 & new_n1300;
  assign new_n1302 = ~pn4 & ~new_n1298;
  assign new_n1303 = ~new_n1299 & ~new_n1301;
  assign new_n1304 = ~new_n1302 & new_n1303;
  assign new_n1305 = pa1 & new_n1304;
  assign new_n1306 = ~pj1 & new_n1305;
  assign new_n1307 = pz0 & new_n1305;
  assign new_n1308 = ~pk1 & new_n1304;
  assign new_n1309 = ~pj1 & new_n1308;
  assign new_n1310 = pz0 & new_n1304;
  assign new_n1311 = ~pk1 & new_n1310;
  assign new_n1312 = new_n1290 & new_n1304;
  assign new_n1313 = ~new_n1306 & ~new_n1307;
  assign new_n1314 = ~new_n1309 & new_n1313;
  assign new_n1315 = ~new_n1311 & ~new_n1312;
  assign new_n1316 = new_n1314 & new_n1315;
  assign new_n1317 = ~new_n1292 & ~new_n1294;
  assign new_n1318 = ~new_n1316 & new_n1317;
  assign new_n1319 = pm1 & new_n1318;
  assign new_n1320 = po0 & ~new_n1319;
  assign new_n1321 = ~pq0 & new_n1320;
  assign new_n1322 = pp0 & new_n1321;
  assign new_n1323 = ~pn0 & new_n1322;
  assign new_n1324 = pm1 & new_n1321;
  assign pv6 = new_n1323 | new_n1324;
  assign new_n1326 = pl0 & pd;
  assign new_n1327 = ~pl0 & pl;
  assign new_n1328 = pk0 & new_n1327;
  assign new_n1329 = ~pk0 & pd;
  assign new_n1330 = ~new_n1326 & ~new_n1328;
  assign new_n1331 = ~new_n1329 & new_n1330;
  assign new_n1332 = new_n310 & new_n1331;
  assign new_n1333 = ~pm0 & new_n1332;
  assign new_n1334 = pl4 & ~po2;
  assign new_n1335 = ~new_n336 & new_n1334;
  assign new_n1336 = ~new_n293 & new_n1335;
  assign new_n1337 = ~pn2 & new_n877;
  assign new_n1338 = ~new_n1333 & ~new_n1336;
  assign new_n1339 = ~new_n1337 & new_n1338;
  assign new_n1340 = po0 & new_n1339;
  assign pw7 = ~pq0 & new_n1340;
  assign new_n1342 = po3 & ~pq0;
  assign new_n1343 = new_n497 & new_n1342;
  assign new_n1344 = po0 & new_n1343;
  assign new_n1345 = pp3 & ~new_n453;
  assign new_n1346 = pk4 & new_n1345;
  assign new_n1347 = new_n513 & new_n1346;
  assign new_n1348 = new_n514 & new_n1347;
  assign px8 = new_n1344 | new_n1348;
  assign new_n1350 = pl0 & pc;
  assign new_n1351 = ~pl0 & pk;
  assign new_n1352 = pk0 & new_n1351;
  assign new_n1353 = ~pk0 & pc;
  assign new_n1354 = ~new_n1350 & ~new_n1352;
  assign new_n1355 = ~new_n1353 & new_n1354;
  assign new_n1356 = new_n310 & new_n1355;
  assign new_n1357 = ~pm0 & new_n1356;
  assign new_n1358 = pl4 & ~pn2;
  assign new_n1359 = ~new_n336 & new_n1358;
  assign new_n1360 = ~new_n293 & new_n1359;
  assign new_n1361 = ~pm2 & new_n877;
  assign new_n1362 = ~new_n1357 & ~new_n1360;
  assign new_n1363 = ~new_n1361 & new_n1362;
  assign new_n1364 = po0 & new_n1363;
  assign pv7 = ~pq0 & new_n1364;
  assign new_n1366 = ~pn1 & new_n295;
  assign new_n1367 = pj0 & new_n297;
  assign new_n1368 = new_n301 & ~new_n1367;
  assign new_n1369 = ~new_n1366 & ~new_n1368;
  assign new_n1370 = ~pn0 & new_n1369;
  assign new_n1371 = new_n293 & new_n1370;
  assign new_n1372 = pl4 & ~po1;
  assign new_n1373 = new_n1370 & ~new_n1372;
  assign new_n1374 = pn1 & new_n1369;
  assign new_n1375 = ~new_n1372 & new_n1374;
  assign new_n1376 = new_n310 & new_n1374;
  assign new_n1377 = new_n293 & new_n1374;
  assign new_n1378 = new_n294 & new_n1369;
  assign new_n1379 = ~new_n1372 & new_n1378;
  assign new_n1380 = new_n310 & new_n1378;
  assign new_n1381 = new_n310 & new_n1370;
  assign new_n1382 = new_n293 & new_n1378;
  assign new_n1383 = ~new_n1371 & ~new_n1373;
  assign new_n1384 = ~new_n1375 & new_n1383;
  assign new_n1385 = ~new_n1376 & ~new_n1377;
  assign new_n1386 = new_n1384 & new_n1385;
  assign new_n1387 = ~new_n1381 & ~new_n1382;
  assign new_n1388 = ~new_n1379 & ~new_n1380;
  assign new_n1389 = new_n1387 & new_n1388;
  assign pw6 = ~new_n1386 | ~new_n1389;
  assign new_n1391 = ~pq0 & pp3;
  assign new_n1392 = new_n497 & new_n1391;
  assign new_n1393 = po0 & new_n1392;
  assign new_n1394 = pq3 & ~new_n453;
  assign new_n1395 = pk4 & new_n1394;
  assign new_n1396 = new_n513 & new_n1395;
  assign new_n1397 = new_n514 & new_n1396;
  assign py8 = new_n1393 | new_n1397;
  assign new_n1399 = ~pe1 & ~pn0;
  assign new_n1400 = new_n288 & new_n1399;
  assign new_n1401 = ~pe1 & new_n288;
  assign new_n1402 = ~pn0 & new_n1401;
  assign new_n1403 = ~pk1 & ~new_n1402;
  assign new_n1404 = po0 & ~new_n1403;
  assign new_n1405 = ~pq0 & new_n1404;
  assign new_n1406 = new_n1400 & new_n1405;
  assign new_n1407 = ~new_n288 & new_n1406;
  assign new_n1408 = pn0 & new_n1406;
  assign new_n1409 = ~pg1 & new_n1405;
  assign new_n1410 = pn0 & new_n1409;
  assign new_n1411 = ~pc1 & ~pe1;
  assign new_n1412 = ~pe1 & ~pd1;
  assign new_n1413 = ~pc1 & ~pd1;
  assign new_n1414 = ~new_n1411 & ~new_n1412;
  assign new_n1415 = ~new_n1413 & new_n1414;
  assign new_n1416 = new_n1409 & new_n1415;
  assign new_n1417 = ~new_n288 & new_n1409;
  assign new_n1418 = new_n1406 & new_n1415;
  assign new_n1419 = ~new_n1407 & ~new_n1408;
  assign new_n1420 = ~new_n1410 & new_n1419;
  assign new_n1421 = ~new_n1416 & ~new_n1417;
  assign new_n1422 = ~new_n1418 & new_n1421;
  assign pt6 = ~new_n1420 | ~new_n1422;
  assign new_n1424 = pl0 & pb;
  assign new_n1425 = ~pl0 & pj;
  assign new_n1426 = pk0 & new_n1425;
  assign new_n1427 = ~pk0 & pb;
  assign new_n1428 = ~new_n1424 & ~new_n1426;
  assign new_n1429 = ~new_n1427 & new_n1428;
  assign new_n1430 = new_n310 & new_n1429;
  assign new_n1431 = ~pm0 & new_n1430;
  assign new_n1432 = pl4 & ~pm2;
  assign new_n1433 = ~new_n336 & new_n1432;
  assign new_n1434 = ~new_n293 & new_n1433;
  assign new_n1435 = ~pl2 & new_n877;
  assign new_n1436 = ~new_n1431 & ~new_n1434;
  assign new_n1437 = ~new_n1435 & new_n1436;
  assign new_n1438 = po0 & new_n1437;
  assign pu7 = ~pq0 & new_n1438;
  assign new_n1440 = ~pe3 & pl0;
  assign new_n1441 = pk0 & new_n1440;
  assign new_n1442 = ~pe3 & ~pl0;
  assign new_n1443 = ~pk0 & new_n1442;
  assign new_n1444 = ~new_n1441 & ~new_n1443;
  assign new_n1445 = pm0 & new_n1444;
  assign new_n1446 = pl0 & new_n1445;
  assign new_n1447 = pk0 & new_n1446;
  assign new_n1448 = ~pl0 & new_n1445;
  assign new_n1449 = ~pk0 & new_n1448;
  assign new_n1450 = pm3 & new_n1445;
  assign new_n1451 = ~new_n1447 & ~new_n1449;
  assign pv4 = new_n1450 | ~new_n1451;
  assign new_n1453 = ~pq0 & pq3;
  assign new_n1454 = new_n497 & new_n1453;
  assign new_n1455 = po0 & new_n1454;
  assign new_n1456 = pr3 & ~new_n453;
  assign new_n1457 = pk4 & new_n1456;
  assign new_n1458 = new_n513 & new_n1457;
  assign new_n1459 = new_n514 & new_n1458;
  assign pz8 = new_n1455 | new_n1459;
  assign new_n1461 = pl0 & pa;
  assign new_n1462 = ~pl0 & pi;
  assign new_n1463 = pk0 & new_n1462;
  assign new_n1464 = ~pk0 & pa;
  assign new_n1465 = ~new_n1461 & ~new_n1463;
  assign new_n1466 = ~new_n1464 & new_n1465;
  assign new_n1467 = new_n310 & new_n1466;
  assign new_n1468 = ~pm0 & new_n1467;
  assign new_n1469 = pl4 & ~pl2;
  assign new_n1470 = ~new_n336 & new_n1469;
  assign new_n1471 = ~new_n293 & new_n1470;
  assign new_n1472 = ~pk2 & new_n877;
  assign new_n1473 = ~new_n1468 & ~new_n1471;
  assign new_n1474 = ~new_n1472 & new_n1473;
  assign new_n1475 = po0 & new_n1474;
  assign pt7 = ~pq0 & new_n1475;
  assign new_n1477 = po0 & ~new_n1402;
  assign new_n1478 = ~pq0 & new_n1477;
  assign new_n1479 = pl1 & new_n1478;
  assign new_n1480 = ~pg1 & new_n1479;
  assign new_n1481 = ~pd1 & new_n288;
  assign new_n1482 = ~pn0 & new_n1481;
  assign new_n1483 = ~pc1 & new_n1482;
  assign new_n1484 = new_n1478 & new_n1483;
  assign pu6 = new_n1480 | new_n1484;
  assign new_n1486 = ~pf3 & pl0;
  assign new_n1487 = pk0 & new_n1486;
  assign new_n1488 = ~pf3 & ~pl0;
  assign new_n1489 = ~pk0 & new_n1488;
  assign new_n1490 = ~new_n1487 & ~new_n1489;
  assign new_n1491 = pm0 & new_n1490;
  assign new_n1492 = pl0 & new_n1491;
  assign new_n1493 = pk0 & new_n1492;
  assign new_n1494 = ~pl0 & new_n1491;
  assign new_n1495 = ~pk0 & new_n1494;
  assign new_n1496 = pn3 & new_n1491;
  assign new_n1497 = ~new_n1493 & ~new_n1495;
  assign pw4 = new_n1496 | ~new_n1497;
  assign new_n1499 = ~pd3 & ~pl3;
  assign new_n1500 = ~pd3 & pl0;
  assign new_n1501 = ~new_n759 & ~new_n1499;
  assign new_n1502 = ~new_n1500 & new_n1501;
  assign new_n1503 = ~pm0 & ~pt3;
  assign new_n1504 = ~pd3 & ~pl0;
  assign new_n1505 = ~new_n757 & ~new_n1499;
  assign new_n1506 = ~new_n1504 & new_n1505;
  assign new_n1507 = new_n1502 & ~new_n1503;
  assign new_n1508 = new_n1506 & new_n1507;
  assign new_n1509 = ~new_n1503 & new_n1506;
  assign new_n1510 = ~pk0 & new_n1509;
  assign new_n1511 = pk0 & new_n1507;
  assign new_n1512 = ~pm0 & ~new_n1503;
  assign new_n1513 = ~new_n1508 & ~new_n1510;
  assign new_n1514 = ~new_n1511 & ~new_n1512;
  assign pp4 = ~new_n1513 | ~new_n1514;
  assign new_n1516 = pk1 & ~pn0;
  assign pq5 = pk4 | ~new_n1516;
  assign new_n1518 = ~pi1 & ~new_n1402;
  assign new_n1519 = po0 & ~new_n1518;
  assign new_n1520 = ~pq0 & new_n1519;
  assign new_n1521 = new_n1400 & new_n1520;
  assign new_n1522 = ~new_n288 & new_n1521;
  assign new_n1523 = pn0 & new_n1521;
  assign new_n1524 = ~pg1 & new_n1520;
  assign new_n1525 = pn0 & new_n1524;
  assign new_n1526 = ~pe1 & pd1;
  assign new_n1527 = ~new_n1411 & ~new_n1526;
  assign new_n1528 = ~new_n1413 & new_n1527;
  assign new_n1529 = new_n1524 & new_n1528;
  assign new_n1530 = ~new_n288 & new_n1524;
  assign new_n1531 = new_n1521 & new_n1528;
  assign new_n1532 = ~new_n1522 & ~new_n1523;
  assign new_n1533 = ~new_n1525 & new_n1532;
  assign new_n1534 = ~new_n1529 & ~new_n1530;
  assign new_n1535 = ~new_n1531 & new_n1534;
  assign pr6 = ~new_n1533 | ~new_n1535;
  assign new_n1537 = ~pj2 & new_n295;
  assign new_n1538 = pc0 & new_n297;
  assign new_n1539 = new_n301 & ~new_n1538;
  assign new_n1540 = ~new_n1537 & ~new_n1539;
  assign new_n1541 = ~pn0 & new_n1540;
  assign new_n1542 = new_n293 & new_n1541;
  assign new_n1543 = pl4 & ~pk2;
  assign new_n1544 = new_n1541 & ~new_n1543;
  assign new_n1545 = pj2 & new_n1540;
  assign new_n1546 = ~new_n1543 & new_n1545;
  assign new_n1547 = new_n310 & new_n1545;
  assign new_n1548 = new_n293 & new_n1545;
  assign new_n1549 = new_n294 & new_n1540;
  assign new_n1550 = ~new_n1543 & new_n1549;
  assign new_n1551 = new_n310 & new_n1549;
  assign new_n1552 = new_n310 & new_n1541;
  assign new_n1553 = new_n293 & new_n1549;
  assign new_n1554 = ~new_n1542 & ~new_n1544;
  assign new_n1555 = ~new_n1546 & new_n1554;
  assign new_n1556 = ~new_n1547 & ~new_n1548;
  assign new_n1557 = new_n1555 & new_n1556;
  assign new_n1558 = ~new_n1552 & ~new_n1553;
  assign new_n1559 = ~new_n1550 & ~new_n1551;
  assign new_n1560 = new_n1558 & new_n1559;
  assign ps7 = ~new_n1557 | ~new_n1560;
  assign new_n1562 = pj1 & ~pn0;
  assign pp5 = pk4 | ~new_n1562;
  assign new_n1564 = ~pc3 & ~pk3;
  assign new_n1565 = ~pc3 & pl0;
  assign new_n1566 = ~new_n797 & ~new_n1564;
  assign new_n1567 = ~new_n1565 & new_n1566;
  assign new_n1568 = ~pm0 & ~ps3;
  assign new_n1569 = ~pc3 & ~pl0;
  assign new_n1570 = ~new_n795 & ~new_n1564;
  assign new_n1571 = ~new_n1569 & new_n1570;
  assign new_n1572 = new_n1567 & ~new_n1568;
  assign new_n1573 = new_n1571 & new_n1572;
  assign new_n1574 = ~new_n1568 & new_n1571;
  assign new_n1575 = ~pk0 & new_n1574;
  assign new_n1576 = pk0 & new_n1572;
  assign new_n1577 = ~pm0 & ~new_n1568;
  assign new_n1578 = ~new_n1573 & ~new_n1575;
  assign new_n1579 = ~new_n1576 & ~new_n1577;
  assign pq4 = ~new_n1578 | ~new_n1579;
  assign new_n1581 = ~pi2 & new_n295;
  assign new_n1582 = pb0 & new_n297;
  assign new_n1583 = new_n301 & ~new_n1582;
  assign new_n1584 = ~new_n1581 & ~new_n1583;
  assign new_n1585 = ~pn0 & new_n1584;
  assign new_n1586 = new_n293 & new_n1585;
  assign new_n1587 = ~pj2 & pl4;
  assign new_n1588 = new_n1585 & ~new_n1587;
  assign new_n1589 = pi2 & new_n1584;
  assign new_n1590 = ~new_n1587 & new_n1589;
  assign new_n1591 = new_n310 & new_n1589;
  assign new_n1592 = new_n293 & new_n1589;
  assign new_n1593 = new_n294 & new_n1584;
  assign new_n1594 = ~new_n1587 & new_n1593;
  assign new_n1595 = new_n310 & new_n1593;
  assign new_n1596 = new_n310 & new_n1585;
  assign new_n1597 = new_n293 & new_n1593;
  assign new_n1598 = ~new_n1586 & ~new_n1588;
  assign new_n1599 = ~new_n1590 & new_n1598;
  assign new_n1600 = ~new_n1591 & ~new_n1592;
  assign new_n1601 = new_n1599 & new_n1600;
  assign new_n1602 = ~new_n1596 & ~new_n1597;
  assign new_n1603 = ~new_n1594 & ~new_n1595;
  assign new_n1604 = new_n1602 & new_n1603;
  assign pr7 = ~new_n1601 | ~new_n1604;
  assign new_n1606 = ~pj1 & ~new_n1402;
  assign new_n1607 = po0 & ~new_n1606;
  assign new_n1608 = ~pq0 & new_n1607;
  assign new_n1609 = new_n1400 & new_n1608;
  assign new_n1610 = ~new_n288 & new_n1609;
  assign new_n1611 = pn0 & new_n1609;
  assign new_n1612 = ~pg1 & new_n1608;
  assign new_n1613 = pn0 & new_n1612;
  assign new_n1614 = pc1 & ~pe1;
  assign new_n1615 = ~new_n1412 & ~new_n1614;
  assign new_n1616 = ~new_n1413 & new_n1615;
  assign new_n1617 = new_n1612 & new_n1616;
  assign new_n1618 = ~new_n288 & new_n1612;
  assign new_n1619 = new_n1609 & new_n1616;
  assign new_n1620 = ~new_n1610 & ~new_n1611;
  assign new_n1621 = ~new_n1613 & new_n1620;
  assign new_n1622 = ~new_n1617 & ~new_n1618;
  assign new_n1623 = ~new_n1619 & new_n1622;
  assign ps6 = ~new_n1621 | ~new_n1623;
  assign pp6 = new_n297 & new_n1318;
  assign new_n1626 = ~ph2 & new_n295;
  assign new_n1627 = pa0 & new_n297;
  assign new_n1628 = new_n301 & ~new_n1627;
  assign new_n1629 = ~new_n1626 & ~new_n1628;
  assign new_n1630 = ~pn0 & new_n1629;
  assign new_n1631 = new_n293 & new_n1630;
  assign new_n1632 = pl4 & ~pi2;
  assign new_n1633 = new_n1630 & ~new_n1632;
  assign new_n1634 = ph2 & new_n1629;
  assign new_n1635 = ~new_n1632 & new_n1634;
  assign new_n1636 = new_n310 & new_n1634;
  assign new_n1637 = new_n293 & new_n1634;
  assign new_n1638 = new_n294 & new_n1629;
  assign new_n1639 = ~new_n1632 & new_n1638;
  assign new_n1640 = new_n310 & new_n1638;
  assign new_n1641 = new_n310 & new_n1630;
  assign new_n1642 = new_n293 & new_n1638;
  assign new_n1643 = ~new_n1631 & ~new_n1633;
  assign new_n1644 = ~new_n1635 & new_n1643;
  assign new_n1645 = ~new_n1636 & ~new_n1637;
  assign new_n1646 = new_n1644 & new_n1645;
  assign new_n1647 = ~new_n1641 & ~new_n1642;
  assign new_n1648 = ~new_n1639 & ~new_n1640;
  assign new_n1649 = new_n1647 & new_n1648;
  assign pq7 = ~new_n1646 | ~new_n1649;
  assign new_n1651 = ~pb3 & ~pj3;
  assign new_n1652 = ~pb3 & pl0;
  assign new_n1653 = ~new_n620 & ~new_n1651;
  assign new_n1654 = ~new_n1652 & new_n1653;
  assign new_n1655 = ~pm0 & ~pr3;
  assign new_n1656 = ~pb3 & ~pl0;
  assign new_n1657 = ~new_n618 & ~new_n1651;
  assign new_n1658 = ~new_n1656 & new_n1657;
  assign new_n1659 = new_n1654 & ~new_n1655;
  assign new_n1660 = new_n1658 & new_n1659;
  assign new_n1661 = ~new_n1655 & new_n1658;
  assign new_n1662 = ~pk0 & new_n1661;
  assign new_n1663 = pk0 & new_n1659;
  assign new_n1664 = ~pm0 & ~new_n1655;
  assign new_n1665 = ~new_n1660 & ~new_n1662;
  assign new_n1666 = ~new_n1663 & ~new_n1664;
  assign pr4 = ~new_n1665 | ~new_n1666;
  assign new_n1668 = ~pg2 & new_n295;
  assign new_n1669 = pz & new_n297;
  assign new_n1670 = new_n301 & ~new_n1669;
  assign new_n1671 = ~new_n1668 & ~new_n1670;
  assign new_n1672 = ~pn0 & new_n1671;
  assign new_n1673 = new_n293 & new_n1672;
  assign new_n1674 = pl4 & ~ph2;
  assign new_n1675 = new_n1672 & ~new_n1674;
  assign new_n1676 = pg2 & new_n1671;
  assign new_n1677 = ~new_n1674 & new_n1676;
  assign new_n1678 = new_n310 & new_n1676;
  assign new_n1679 = new_n293 & new_n1676;
  assign new_n1680 = new_n294 & new_n1671;
  assign new_n1681 = ~new_n1674 & new_n1680;
  assign new_n1682 = new_n310 & new_n1680;
  assign new_n1683 = new_n310 & new_n1672;
  assign new_n1684 = new_n293 & new_n1680;
  assign new_n1685 = ~new_n1673 & ~new_n1675;
  assign new_n1686 = ~new_n1677 & new_n1685;
  assign new_n1687 = ~new_n1678 & ~new_n1679;
  assign new_n1688 = new_n1686 & new_n1687;
  assign new_n1689 = ~new_n1683 & ~new_n1684;
  assign new_n1690 = ~new_n1681 & ~new_n1682;
  assign new_n1691 = new_n1689 & new_n1690;
  assign pp7 = ~new_n1688 | ~new_n1691;
  assign new_n1693 = ph1 & new_n669;
  assign new_n1694 = pc1 & pe1;
  assign new_n1695 = pe1 & pd1;
  assign new_n1696 = ~new_n1694 & ~new_n1695;
  assign new_n1697 = ~pn0 & new_n1696;
  assign new_n1698 = new_n288 & new_n1697;
  assign new_n1699 = new_n1693 & ~new_n1698;
  assign new_n1700 = po0 & new_n1699;
  assign new_n1701 = ~pc1 & new_n297;
  assign new_n1702 = new_n288 & new_n1412;
  assign new_n1703 = new_n1701 & new_n1702;
  assign new_n1704 = ~pn0 & new_n1703;
  assign pq6 = new_n1700 | new_n1704;
  assign new_n1706 = pl1 & ~pn0;
  assign pr5 = pk4 | ~new_n1706;
  assign new_n1708 = ~pi3 & ~pl0;
  assign new_n1709 = ~pa3 & ~pi3;
  assign new_n1710 = ~pa3 & pl0;
  assign new_n1711 = ~new_n1708 & ~new_n1709;
  assign new_n1712 = ~new_n1710 & new_n1711;
  assign new_n1713 = ~pm0 & ~pq3;
  assign new_n1714 = ~pi3 & pl0;
  assign new_n1715 = ~pa3 & ~pl0;
  assign new_n1716 = ~new_n1709 & ~new_n1714;
  assign new_n1717 = ~new_n1715 & new_n1716;
  assign new_n1718 = new_n1712 & ~new_n1713;
  assign new_n1719 = new_n1717 & new_n1718;
  assign new_n1720 = ~new_n1713 & new_n1717;
  assign new_n1721 = ~pk0 & new_n1720;
  assign new_n1722 = pk0 & new_n1718;
  assign new_n1723 = ~pm0 & ~new_n1713;
  assign new_n1724 = ~new_n1719 & ~new_n1721;
  assign new_n1725 = ~new_n1722 & ~new_n1723;
  assign ps4 = ~new_n1724 | ~new_n1725;
  assign new_n1727 = pg3 & ~pq0;
  assign new_n1728 = new_n497 & new_n1727;
  assign new_n1729 = po0 & new_n1728;
  assign new_n1730 = ph3 & ~new_n453;
  assign new_n1731 = pk4 & new_n1730;
  assign new_n1732 = new_n513 & new_n1731;
  assign new_n1733 = new_n514 & new_n1732;
  assign pp8 = new_n1729 | new_n1733;
  assign new_n1735 = pf4 & new_n786;
  assign new_n1736 = pk4 & new_n1288;
  assign new_n1737 = ~pg1 & ~new_n453;
  assign new_n1738 = new_n1735 & new_n1736;
  assign new_n1739 = new_n1737 & new_n1738;
  assign new_n1740 = ~new_n310 & new_n514;
  assign new_n1741 = new_n1739 & new_n1740;
  assign new_n1742 = ph4 & new_n669;
  assign new_n1743 = pe4 & new_n778;
  assign new_n1744 = pf4 & ~pg4;
  assign new_n1745 = pk4 & new_n1744;
  assign new_n1746 = new_n1743 & new_n1745;
  assign new_n1747 = ~new_n477 & new_n1746;
  assign new_n1748 = ~new_n310 & ~new_n1747;
  assign new_n1749 = new_n1742 & new_n1748;
  assign new_n1750 = po0 & new_n1749;
  assign new_n1751 = ~new_n1741 & ~new_n1750;
  assign pq9 = new_n538 | ~new_n1751;
  assign new_n1753 = ~pq0 & ~new_n477;
  assign new_n1754 = ~new_n453 & new_n1753;
  assign new_n1755 = ~pd4 & ~pg1;
  assign new_n1756 = pe4 & new_n1755;
  assign new_n1757 = new_n1745 & new_n1756;
  assign new_n1758 = po0 & new_n1757;
  assign new_n1759 = ~new_n310 & new_n1754;
  assign new_n1760 = new_n1758 & new_n1759;
  assign new_n1761 = pg4 & new_n669;
  assign new_n1762 = pk4 & new_n451;
  assign new_n1763 = new_n778 & new_n1762;
  assign new_n1764 = ~new_n477 & new_n1763;
  assign new_n1765 = ~new_n310 & ~new_n1764;
  assign new_n1766 = new_n1761 & new_n1765;
  assign new_n1767 = po0 & new_n1766;
  assign new_n1768 = pl0 & pm0;
  assign new_n1769 = ~pk0 & new_n1768;
  assign new_n1770 = ~pl0 & pm0;
  assign new_n1771 = pk0 & new_n1770;
  assign new_n1772 = ~new_n1769 & ~new_n1771;
  assign new_n1773 = ~pn0 & new_n1772;
  assign new_n1774 = po0 & new_n1773;
  assign new_n1775 = ~pq0 & new_n1774;
  assign new_n1776 = new_n288 & new_n1775;
  assign new_n1777 = ~new_n1760 & ~new_n1767;
  assign pp9 = new_n1776 | ~new_n1777;
  assign new_n1779 = ph3 & ~pq0;
  assign new_n1780 = new_n497 & new_n1779;
  assign new_n1781 = po0 & new_n1780;
  assign new_n1782 = pi3 & ~new_n453;
  assign new_n1783 = pk4 & new_n1782;
  assign new_n1784 = new_n513 & new_n1783;
  assign new_n1785 = new_n514 & new_n1784;
  assign pq8 = new_n1781 | new_n1785;
  assign new_n1787 = pi3 & ~pq0;
  assign new_n1788 = new_n497 & new_n1787;
  assign new_n1789 = po0 & new_n1788;
  assign new_n1790 = pj3 & ~new_n453;
  assign new_n1791 = pk4 & new_n1790;
  assign new_n1792 = new_n513 & new_n1791;
  assign new_n1793 = new_n514 & new_n1792;
  assign pr8 = new_n1789 | new_n1793;
  assign new_n1795 = pj4 & new_n669;
  assign new_n1796 = ps0 & new_n450;
  assign new_n1797 = ~pi1 & new_n1796;
  assign new_n1798 = pt0 & new_n465;
  assign new_n1799 = ~pj1 & new_n1798;
  assign new_n1800 = pi1 & ~new_n1799;
  assign new_n1801 = ~pi1 & ~pk1;
  assign new_n1802 = ~pl1 & new_n1801;
  assign new_n1803 = ~pu0 & new_n1802;
  assign new_n1804 = ~ph1 & new_n1803;
  assign new_n1805 = ~pl1 & ~new_n453;
  assign new_n1806 = ~pk1 & new_n1805;
  assign new_n1807 = ~pj1 & ~new_n453;
  assign new_n1808 = ~new_n1806 & ~new_n1807;
  assign new_n1809 = ~new_n484 & ~new_n1808;
  assign new_n1810 = ~new_n477 & new_n1809;
  assign new_n1811 = pk4 & new_n1810;
  assign new_n1812 = pn4 & new_n1811;
  assign new_n1813 = ~new_n1800 & ~new_n1804;
  assign new_n1814 = new_n1812 & new_n1813;
  assign new_n1815 = ~pi1 & ~pj1;
  assign new_n1816 = new_n1797 & new_n1814;
  assign new_n1817 = ~new_n1815 & new_n1816;
  assign new_n1818 = ~pl1 & ~pv0;
  assign new_n1819 = ~pk1 & ~pw0;
  assign new_n1820 = ~new_n465 & ~new_n1818;
  assign new_n1821 = ~new_n1819 & new_n1820;
  assign new_n1822 = new_n1816 & new_n1821;
  assign new_n1823 = new_n1814 & new_n1821;
  assign new_n1824 = ~ph1 & new_n1823;
  assign new_n1825 = ph1 & new_n1816;
  assign new_n1826 = new_n1814 & ~new_n1815;
  assign new_n1827 = ~ph1 & new_n1826;
  assign new_n1828 = ~new_n1817 & ~new_n1822;
  assign new_n1829 = ~new_n1824 & new_n1828;
  assign new_n1830 = ~new_n1825 & ~new_n1827;
  assign new_n1831 = new_n1829 & new_n1830;
  assign new_n1832 = new_n1795 & new_n1831;
  assign new_n1833 = po0 & new_n1832;
  assign new_n1834 = ~pg1 & new_n673;
  assign new_n1835 = ~pj4 & pk4;
  assign new_n1836 = pn4 & new_n1835;
  assign new_n1837 = po0 & new_n1836;
  assign new_n1838 = ~pq0 & new_n1837;
  assign new_n1839 = new_n1225 & new_n1834;
  assign new_n1840 = new_n1838 & new_n1839;
  assign ps9 = new_n1833 | new_n1840;
  assign new_n1842 = pi4 & pn1;
  assign new_n1843 = ~new_n293 & new_n297;
  assign new_n1844 = ~new_n1842 & new_n1843;
  assign new_n1845 = pl4 & new_n1844;
  assign new_n1846 = pn1 & new_n1845;
  assign new_n1847 = pi4 & new_n1845;
  assign pr9 = new_n1846 | new_n1847;
  assign new_n1849 = pj3 & ~pq0;
  assign new_n1850 = new_n497 & new_n1849;
  assign new_n1851 = po0 & new_n1850;
  assign new_n1852 = pk3 & ~new_n453;
  assign new_n1853 = pk4 & new_n1852;
  assign new_n1854 = new_n513 & new_n1853;
  assign new_n1855 = new_n514 & new_n1854;
  assign ps8 = new_n1851 | new_n1855;
  assign new_n1857 = pk3 & ~pq0;
  assign new_n1858 = new_n497 & new_n1857;
  assign new_n1859 = po0 & new_n1858;
  assign new_n1860 = pl3 & ~new_n453;
  assign new_n1861 = pk4 & new_n1860;
  assign new_n1862 = new_n513 & new_n1861;
  assign new_n1863 = new_n514 & new_n1862;
  assign pt8 = new_n1859 | new_n1863;
  assign pu9 = pm1 & new_n1843;
  assign new_n1866 = ~pg3 & pl0;
  assign new_n1867 = pk0 & new_n1866;
  assign new_n1868 = ~pg3 & ~pl0;
  assign new_n1869 = ~pk0 & new_n1868;
  assign new_n1870 = ~new_n1867 & ~new_n1869;
  assign new_n1871 = pm0 & new_n1870;
  assign new_n1872 = pl0 & new_n1871;
  assign new_n1873 = pk0 & new_n1872;
  assign new_n1874 = ~pl0 & new_n1871;
  assign new_n1875 = ~pk0 & new_n1874;
  assign new_n1876 = po3 & new_n1871;
  assign new_n1877 = ~new_n1873 & ~new_n1875;
  assign px4 = new_n1876 | ~new_n1877;
  assign new_n1879 = pi1 & pm1;
  assign py5 = pk4 | ~new_n1879;
  assign new_n1881 = ~pq1 & new_n295;
  assign new_n1882 = pg0 & new_n297;
  assign new_n1883 = new_n301 & ~new_n1882;
  assign new_n1884 = ~new_n1881 & ~new_n1883;
  assign new_n1885 = ~pn0 & new_n1884;
  assign new_n1886 = new_n293 & new_n1885;
  assign new_n1887 = pl4 & ~pr1;
  assign new_n1888 = new_n1885 & ~new_n1887;
  assign new_n1889 = pq1 & new_n1884;
  assign new_n1890 = ~new_n1887 & new_n1889;
  assign new_n1891 = new_n310 & new_n1889;
  assign new_n1892 = new_n293 & new_n1889;
  assign new_n1893 = new_n294 & new_n1884;
  assign new_n1894 = ~new_n1887 & new_n1893;
  assign new_n1895 = new_n310 & new_n1893;
  assign new_n1896 = new_n310 & new_n1885;
  assign new_n1897 = new_n293 & new_n1893;
  assign new_n1898 = ~new_n1886 & ~new_n1888;
  assign new_n1899 = ~new_n1890 & new_n1898;
  assign new_n1900 = ~new_n1891 & ~new_n1892;
  assign new_n1901 = new_n1899 & new_n1900;
  assign new_n1902 = ~new_n1896 & ~new_n1897;
  assign new_n1903 = ~new_n1894 & ~new_n1895;
  assign new_n1904 = new_n1902 & new_n1903;
  assign pz6 = ~new_n1901 | ~new_n1904;
  assign new_n1906 = pm1 & ~pq0;
  assign new_n1907 = new_n706 & new_n1906;
  assign new_n1908 = po0 & new_n1907;
  assign new_n1909 = ~pb4 & new_n1908;
  assign pt9 = ~pc4 & new_n1909;
  assign new_n1911 = pl3 & ~pq0;
  assign new_n1912 = new_n497 & new_n1911;
  assign new_n1913 = po0 & new_n1912;
  assign new_n1914 = pm3 & ~new_n453;
  assign new_n1915 = pk4 & new_n1914;
  assign new_n1916 = new_n513 & new_n1915;
  assign new_n1917 = new_n514 & new_n1916;
  assign pu8 = new_n1913 | new_n1917;
  assign new_n1919 = ph1 & pm1;
  assign px5 = pk4 | ~new_n1919;
  assign new_n1921 = ~ph3 & pl0;
  assign new_n1922 = pk0 & new_n1921;
  assign new_n1923 = ~ph3 & ~pl0;
  assign new_n1924 = ~pk0 & new_n1923;
  assign new_n1925 = ~new_n1922 & ~new_n1924;
  assign new_n1926 = pm0 & new_n1925;
  assign new_n1927 = pl0 & new_n1926;
  assign new_n1928 = pk0 & new_n1927;
  assign new_n1929 = ~pl0 & new_n1926;
  assign new_n1930 = ~pk0 & new_n1929;
  assign new_n1931 = pp3 & new_n1926;
  assign new_n1932 = ~new_n1928 & ~new_n1930;
  assign py4 = new_n1931 | ~new_n1932;
  assign new_n1934 = pl0 & pg;
  assign new_n1935 = ~pl0 & po;
  assign new_n1936 = pk0 & new_n1935;
  assign new_n1937 = ~pk0 & pg;
  assign new_n1938 = ~new_n1934 & ~new_n1936;
  assign new_n1939 = ~new_n1937 & new_n1938;
  assign new_n1940 = new_n310 & new_n1939;
  assign new_n1941 = ~pm0 & new_n1940;
  assign new_n1942 = pl4 & ~pr2;
  assign new_n1943 = ~new_n336 & new_n1942;
  assign new_n1944 = ~new_n293 & new_n1943;
  assign new_n1945 = ~pq2 & new_n877;
  assign new_n1946 = ~new_n1941 & ~new_n1944;
  assign new_n1947 = ~new_n1945 & new_n1946;
  assign new_n1948 = po0 & new_n1947;
  assign pz7 = ~pq0 & new_n1948;
  assign new_n1950 = pm3 & ~pq0;
  assign new_n1951 = new_n497 & new_n1950;
  assign new_n1952 = po0 & new_n1951;
  assign new_n1953 = pn3 & ~new_n453;
  assign new_n1954 = pk4 & new_n1953;
  assign new_n1955 = new_n513 & new_n1954;
  assign new_n1956 = new_n514 & new_n1955;
  assign pv8 = new_n1952 | new_n1956;
  assign pw9 = pk4 & new_n514;
  assign new_n1959 = ~po1 & new_n295;
  assign new_n1960 = pi0 & new_n297;
  assign new_n1961 = new_n301 & ~new_n1960;
  assign new_n1962 = ~new_n1959 & ~new_n1961;
  assign new_n1963 = ~pn0 & new_n1962;
  assign new_n1964 = new_n293 & new_n1963;
  assign new_n1965 = pl4 & ~pp1;
  assign new_n1966 = new_n1963 & ~new_n1965;
  assign new_n1967 = po1 & new_n1962;
  assign new_n1968 = ~new_n1965 & new_n1967;
  assign new_n1969 = new_n310 & new_n1967;
  assign new_n1970 = new_n293 & new_n1967;
  assign new_n1971 = new_n294 & new_n1962;
  assign new_n1972 = ~new_n1965 & new_n1971;
  assign new_n1973 = new_n310 & new_n1971;
  assign new_n1974 = new_n310 & new_n1963;
  assign new_n1975 = new_n293 & new_n1971;
  assign new_n1976 = ~new_n1964 & ~new_n1966;
  assign new_n1977 = ~new_n1968 & new_n1976;
  assign new_n1978 = ~new_n1969 & ~new_n1970;
  assign new_n1979 = new_n1977 & new_n1978;
  assign new_n1980 = ~new_n1974 & ~new_n1975;
  assign new_n1981 = ~new_n1972 & ~new_n1973;
  assign new_n1982 = new_n1980 & new_n1981;
  assign px6 = ~new_n1979 | ~new_n1982;
  assign new_n1984 = pl0 & pf;
  assign new_n1985 = ~pl0 & pn;
  assign new_n1986 = pk0 & new_n1985;
  assign new_n1987 = ~pk0 & pf;
  assign new_n1988 = ~new_n1984 & ~new_n1986;
  assign new_n1989 = ~new_n1987 & new_n1988;
  assign new_n1990 = new_n310 & new_n1989;
  assign new_n1991 = ~pm0 & new_n1990;
  assign new_n1992 = pl4 & ~pq2;
  assign new_n1993 = ~new_n336 & new_n1992;
  assign new_n1994 = ~new_n293 & new_n1993;
  assign new_n1995 = ~pp2 & new_n877;
  assign new_n1996 = ~new_n1991 & ~new_n1994;
  assign new_n1997 = ~new_n1995 & new_n1996;
  assign new_n1998 = po0 & new_n1997;
  assign py7 = ~pq0 & new_n1998;
  assign new_n2000 = pk0 & new_n1714;
  assign new_n2001 = ~pk0 & new_n1708;
  assign new_n2002 = ~new_n2000 & ~new_n2001;
  assign new_n2003 = pm0 & new_n2002;
  assign new_n2004 = pl0 & new_n2003;
  assign new_n2005 = pk0 & new_n2004;
  assign new_n2006 = ~pl0 & new_n2003;
  assign new_n2007 = ~pk0 & new_n2006;
  assign new_n2008 = pq3 & new_n2003;
  assign new_n2009 = ~new_n2005 & ~new_n2007;
  assign pz4 = new_n2008 | ~new_n2009;
  assign new_n2011 = ~pa1 & pk1;
  assign new_n2012 = ~pb1 & pl1;
  assign new_n2013 = ~new_n2011 & ~new_n2012;
  assign new_n2014 = ~new_n453 & new_n2013;
  assign new_n2015 = pz0 & new_n2014;
  assign new_n2016 = py0 & new_n2015;
  assign new_n2017 = ~pj1 & new_n2014;
  assign new_n2018 = py0 & new_n2017;
  assign new_n2019 = ~pi1 & new_n2015;
  assign new_n2020 = ~pi1 & new_n2017;
  assign new_n2021 = ~new_n2016 & ~new_n2018;
  assign new_n2022 = ~new_n2019 & ~new_n2020;
  assign new_n2023 = new_n2021 & new_n2022;
  assign new_n2024 = ~new_n455 & ~new_n2023;
  assign new_n2025 = pn4 & new_n2024;
  assign new_n2026 = new_n477 & ~new_n2025;
  assign new_n2027 = po0 & ~new_n2026;
  assign new_n2028 = ~pq0 & new_n2027;
  assign new_n2029 = new_n2025 & new_n2028;
  assign new_n2030 = new_n1318 & new_n2028;
  assign pv9 = new_n2029 | new_n2030;
  assign new_n2032 = pn3 & ~pq0;
  assign new_n2033 = new_n497 & new_n2032;
  assign new_n2034 = po0 & new_n2033;
  assign new_n2035 = po3 & ~new_n453;
  assign new_n2036 = pk4 & new_n2035;
  assign new_n2037 = new_n513 & new_n2036;
  assign new_n2038 = new_n514 & new_n2037;
  assign pw8 = new_n2034 | new_n2038;
  assign new_n2040 = pl0 & pe;
  assign new_n2041 = ~pl0 & pm;
  assign new_n2042 = pk0 & new_n2041;
  assign new_n2043 = ~pk0 & pe;
  assign new_n2044 = ~new_n2040 & ~new_n2042;
  assign new_n2045 = ~new_n2043 & new_n2044;
  assign new_n2046 = new_n310 & new_n2045;
  assign new_n2047 = ~pm0 & new_n2046;
  assign new_n2048 = pl4 & ~pp2;
  assign new_n2049 = ~new_n336 & new_n2048;
  assign new_n2050 = ~new_n293 & new_n2049;
  assign new_n2051 = ~po2 & new_n877;
  assign new_n2052 = ~new_n2047 & ~new_n2050;
  assign new_n2053 = ~new_n2051 & new_n2052;
  assign new_n2054 = po0 & new_n2053;
  assign px7 = ~pq0 & new_n2054;
  assign new_n2056 = ~pp1 & new_n295;
  assign new_n2057 = ph0 & new_n297;
  assign new_n2058 = new_n301 & ~new_n2057;
  assign new_n2059 = ~new_n2056 & ~new_n2058;
  assign new_n2060 = ~pn0 & new_n2059;
  assign new_n2061 = new_n293 & new_n2060;
  assign new_n2062 = pl4 & ~pq1;
  assign new_n2063 = new_n2060 & ~new_n2062;
  assign new_n2064 = pp1 & new_n2059;
  assign new_n2065 = ~new_n2062 & new_n2064;
  assign new_n2066 = new_n310 & new_n2064;
  assign new_n2067 = new_n293 & new_n2064;
  assign new_n2068 = new_n294 & new_n2059;
  assign new_n2069 = ~new_n2062 & new_n2068;
  assign new_n2070 = new_n310 & new_n2068;
  assign new_n2071 = new_n310 & new_n2060;
  assign new_n2072 = new_n293 & new_n2068;
  assign new_n2073 = ~new_n2061 & ~new_n2063;
  assign new_n2074 = ~new_n2065 & new_n2073;
  assign new_n2075 = ~new_n2066 & ~new_n2067;
  assign new_n2076 = new_n2074 & new_n2075;
  assign new_n2077 = ~new_n2071 & ~new_n2072;
  assign new_n2078 = ~new_n2069 & ~new_n2070;
  assign new_n2079 = new_n2077 & new_n2078;
  assign py6 = ~new_n2076 | ~new_n2079;
  assign new_n2081 = pj1 & pm1;
  assign pz5 = pk4 | ~new_n2081;
  assign pl6 = ~pl1;
  assign po4 = ~pg1;
  assign pj6 = ~pj1;
  assign pk6 = ~pk1;
  assign ph6 = ~ph1;
  assign pi6 = ~pi1;
  assign pm5 = pm4;
  assign pm6 = pk4;
  assign pt4 = pu3;
  assign pt5 = pu5;
  assign pu4 = pv3;
  assign pw5 = pu5;
  assign pv5 = pu5;
  assign ps5 = pu5;
endmodule


