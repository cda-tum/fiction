// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_  );
  input  i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17,
    new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25,
    new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33,
    new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41,
    new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49,
    new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57,
    new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157, new_n158, new_n159, new_n160,
    new_n161, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176, new_n178, new_n179, new_n180, new_n181, new_n182,
    new_n183, new_n184, new_n185, new_n186, new_n187, new_n188, new_n189,
    new_n190, new_n191, new_n192, new_n193, new_n194, new_n195, new_n196,
    new_n197, new_n198, new_n199, new_n200, new_n201, new_n202, new_n203,
    new_n204, new_n205, new_n206, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n216, new_n217,
    new_n218, new_n219, new_n220, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n255, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387;
  assign new_n11 = ~i_5_ & ~i_4_;
  assign new_n12 = i_3_ & new_n11;
  assign new_n13 = i_1_ & ~i_2_;
  assign new_n14 = i_0_ & new_n13;
  assign new_n15 = ~i_6_ & new_n12;
  assign new_n16 = new_n14 & new_n15;
  assign new_n17 = ~i_5_ & i_4_;
  assign new_n18 = i_3_ & new_n17;
  assign new_n19 = ~i_1_ & ~i_2_;
  assign new_n20 = i_0_ & new_n19;
  assign new_n21 = ~i_6_ & new_n18;
  assign new_n22 = new_n20 & new_n21;
  assign new_n23 = i_6_ & new_n18;
  assign new_n24 = new_n14 & new_n23;
  assign new_n25 = ~new_n16 & ~new_n22;
  assign new_n26 = ~new_n24 & new_n25;
  assign new_n27 = ~i_3_ & new_n11;
  assign new_n28 = i_1_ & i_2_;
  assign new_n29 = ~i_0_ & new_n28;
  assign new_n30 = i_6_ & new_n27;
  assign new_n31 = new_n29 & new_n30;
  assign new_n32 = ~i_1_ & i_2_;
  assign new_n33 = ~i_0_ & new_n32;
  assign new_n34 = ~i_6_ & new_n27;
  assign new_n35 = new_n33 & new_n34;
  assign new_n36 = i_5_ & ~i_4_;
  assign new_n37 = ~i_3_ & new_n36;
  assign new_n38 = i_6_ & new_n37;
  assign new_n39 = new_n33 & new_n38;
  assign new_n40 = ~new_n31 & ~new_n35;
  assign new_n41 = ~new_n39 & new_n40;
  assign new_n42 = ~i_0_ & new_n13;
  assign new_n43 = new_n21 & new_n42;
  assign new_n44 = i_3_ & new_n36;
  assign new_n45 = ~i_6_ & new_n44;
  assign new_n46 = new_n20 & new_n45;
  assign new_n47 = i_5_ & i_4_;
  assign new_n48 = i_3_ & new_n47;
  assign new_n49 = i_6_ & new_n48;
  assign new_n50 = new_n20 & new_n49;
  assign new_n51 = ~new_n43 & ~new_n46;
  assign new_n52 = ~new_n50 & new_n51;
  assign new_n53 = new_n26 & new_n41;
  assign new_n54 = new_n52 & new_n53;
  assign new_n55 = ~i_0_ & new_n19;
  assign new_n56 = ~i_6_ & new_n37;
  assign new_n57 = new_n55 & new_n56;
  assign new_n58 = new_n20 & new_n38;
  assign new_n59 = i_0_ & new_n32;
  assign new_n60 = new_n30 & new_n59;
  assign new_n61 = ~new_n57 & ~new_n58;
  assign new_n62 = ~new_n60 & new_n61;
  assign new_n63 = i_6_ & new_n12;
  assign new_n64 = new_n33 & new_n63;
  assign new_n65 = new_n14 & new_n30;
  assign new_n66 = ~i_3_ & new_n17;
  assign new_n67 = i_6_ & new_n66;
  assign new_n68 = new_n42 & new_n67;
  assign new_n69 = ~new_n64 & ~new_n65;
  assign new_n70 = ~new_n68 & new_n69;
  assign new_n71 = new_n38 & new_n42;
  assign new_n72 = ~i_3_ & new_n47;
  assign new_n73 = i_6_ & new_n72;
  assign new_n74 = new_n55 & new_n73;
  assign new_n75 = new_n33 & new_n67;
  assign new_n76 = ~new_n71 & ~new_n74;
  assign new_n77 = ~new_n75 & new_n76;
  assign new_n78 = new_n62 & new_n70;
  assign new_n79 = new_n77 & new_n78;
  assign new_n80 = ~i_6_ & new_n66;
  assign new_n81 = new_n14 & new_n80;
  assign new_n82 = new_n23 & new_n59;
  assign new_n83 = new_n42 & new_n45;
  assign new_n84 = ~new_n81 & ~new_n82;
  assign new_n85 = ~new_n83 & new_n84;
  assign new_n86 = i_6_ & new_n44;
  assign new_n87 = new_n14 & new_n86;
  assign new_n88 = ~i_6_ & new_n48;
  assign new_n89 = new_n55 & new_n88;
  assign new_n90 = new_n42 & new_n49;
  assign new_n91 = ~new_n87 & ~new_n89;
  assign new_n92 = ~new_n90 & new_n91;
  assign new_n93 = new_n15 & new_n59;
  assign new_n94 = ~i_6_ & new_n72;
  assign new_n95 = new_n20 & new_n94;
  assign new_n96 = new_n14 & new_n73;
  assign new_n97 = ~new_n93 & ~new_n95;
  assign new_n98 = ~new_n96 & new_n97;
  assign new_n99 = new_n85 & new_n92;
  assign new_n100 = new_n98 & new_n99;
  assign new_n101 = new_n54 & new_n79;
  assign new_n102 = new_n100 & new_n101;
  assign new_n103 = new_n30 & new_n55;
  assign new_n104 = new_n23 & new_n55;
  assign new_n105 = new_n55 & new_n80;
  assign new_n106 = new_n20 & new_n67;
  assign new_n107 = ~new_n104 & ~new_n105;
  assign new_n108 = ~new_n106 & new_n107;
  assign new_n109 = new_n20 & new_n34;
  assign new_n110 = new_n15 & new_n55;
  assign new_n111 = new_n20 & new_n63;
  assign new_n112 = ~new_n109 & ~new_n110;
  assign new_n113 = ~new_n111 & new_n112;
  assign new_n114 = new_n34 & new_n42;
  assign new_n115 = new_n42 & new_n63;
  assign new_n116 = new_n55 & new_n86;
  assign new_n117 = ~new_n114 & ~new_n115;
  assign new_n118 = ~new_n116 & new_n117;
  assign new_n119 = new_n108 & new_n113;
  assign new_n120 = new_n118 & new_n119;
  assign new_n121 = ~new_n103 & new_n120;
  assign new_n122 = new_n56 & new_n59;
  assign new_n123 = new_n33 & new_n49;
  assign new_n124 = new_n29 & new_n86;
  assign new_n125 = ~new_n122 & ~new_n123;
  assign new_n126 = ~new_n124 & new_n125;
  assign new_n127 = new_n33 & new_n45;
  assign new_n128 = i_0_ & new_n28;
  assign new_n129 = new_n67 & new_n128;
  assign new_n130 = new_n29 & new_n80;
  assign new_n131 = ~new_n127 & ~new_n129;
  assign new_n132 = ~new_n130 & new_n131;
  assign new_n133 = new_n59 & new_n73;
  assign new_n134 = new_n33 & new_n94;
  assign new_n135 = new_n29 & new_n56;
  assign new_n136 = ~new_n133 & ~new_n134;
  assign new_n137 = ~new_n135 & new_n136;
  assign new_n138 = new_n126 & new_n132;
  assign new_n139 = new_n137 & new_n138;
  assign new_n140 = new_n15 & new_n29;
  assign new_n141 = new_n59 & new_n80;
  assign new_n142 = new_n34 & new_n128;
  assign new_n143 = ~new_n140 & ~new_n141;
  assign new_n144 = ~new_n142 & new_n143;
  assign new_n145 = new_n14 & new_n56;
  assign new_n146 = new_n21 & new_n33;
  assign new_n147 = new_n63 & new_n128;
  assign new_n148 = ~new_n145 & ~new_n146;
  assign new_n149 = ~new_n147 & new_n148;
  assign new_n150 = new_n42 & new_n94;
  assign new_n151 = new_n59 & new_n86;
  assign new_n152 = new_n23 & new_n29;
  assign new_n153 = ~new_n150 & ~new_n151;
  assign new_n154 = ~new_n152 & new_n153;
  assign new_n155 = new_n144 & new_n149;
  assign new_n156 = new_n154 & new_n155;
  assign new_n157 = new_n59 & new_n88;
  assign new_n158 = new_n21 & new_n128;
  assign new_n159 = new_n45 & new_n128;
  assign new_n160 = ~new_n157 & ~new_n158;
  assign new_n161 = ~new_n159 & new_n160;
  assign new_n162 = new_n29 & new_n73;
  assign new_n163 = new_n38 & new_n128;
  assign new_n164 = new_n14 & new_n88;
  assign new_n165 = ~new_n162 & ~new_n163;
  assign new_n166 = ~new_n164 & new_n165;
  assign new_n167 = new_n94 & new_n128;
  assign new_n168 = new_n29 & new_n88;
  assign new_n169 = new_n49 & new_n128;
  assign new_n170 = ~new_n167 & ~new_n168;
  assign new_n171 = ~new_n169 & new_n170;
  assign new_n172 = new_n161 & new_n166;
  assign new_n173 = new_n171 & new_n172;
  assign new_n174 = new_n139 & new_n156;
  assign new_n175 = new_n173 & new_n174;
  assign new_n176 = new_n102 & new_n121;
  assign o_1_ = ~new_n175 | ~new_n176;
  assign new_n178 = i_3_ & i_1_;
  assign new_n179 = i_0_ & new_n178;
  assign new_n180 = i_4_ & new_n179;
  assign new_n181 = i_4_ & i_1_;
  assign new_n182 = i_0_ & new_n181;
  assign new_n183 = i_6_ & new_n182;
  assign new_n184 = i_6_ & new_n179;
  assign new_n185 = ~new_n180 & ~new_n183;
  assign new_n186 = ~new_n184 & new_n185;
  assign new_n187 = i_3_ & i_4_;
  assign new_n188 = i_0_ & new_n187;
  assign new_n189 = i_6_ & new_n188;
  assign new_n190 = i_1_ & new_n187;
  assign new_n191 = i_6_ & new_n190;
  assign new_n192 = ~new_n189 & ~new_n191;
  assign new_n193 = i_5_ & new_n190;
  assign new_n194 = i_5_ & new_n182;
  assign new_n195 = i_5_ & i_1_;
  assign new_n196 = i_0_ & new_n195;
  assign new_n197 = i_6_ & new_n196;
  assign new_n198 = ~new_n193 & ~new_n194;
  assign new_n199 = ~new_n197 & new_n198;
  assign new_n200 = new_n186 & new_n192;
  assign new_n201 = new_n199 & new_n200;
  assign new_n202 = i_2_ & new_n187;
  assign new_n203 = i_5_ & new_n202;
  assign new_n204 = i_4_ & i_2_;
  assign new_n205 = i_0_ & new_n204;
  assign new_n206 = i_5_ & new_n205;
  assign new_n207 = i_6_ & new_n128;
  assign new_n208 = ~new_n203 & ~new_n206;
  assign new_n209 = ~new_n207 & new_n208;
  assign new_n210 = i_5_ & i_3_;
  assign new_n211 = i_2_ & new_n210;
  assign new_n212 = i_6_ & new_n211;
  assign new_n213 = i_1_ & new_n204;
  assign new_n214 = i_5_ & new_n213;
  assign new_n215 = i_3_ & i_2_;
  assign new_n216 = i_1_ & new_n215;
  assign new_n217 = i_5_ & new_n216;
  assign new_n218 = ~new_n212 & ~new_n214;
  assign new_n219 = ~new_n217 & new_n218;
  assign new_n220 = i_4_ & new_n216;
  assign new_n221 = i_2_ & new_n47;
  assign new_n222 = i_6_ & new_n221;
  assign new_n223 = i_6_ & new_n213;
  assign new_n224 = ~new_n220 & ~new_n222;
  assign new_n225 = ~new_n223 & new_n224;
  assign new_n226 = new_n209 & new_n219;
  assign new_n227 = new_n225 & new_n226;
  assign new_n228 = i_0_ & new_n215;
  assign new_n229 = i_6_ & new_n228;
  assign new_n230 = i_5_ & new_n188;
  assign new_n231 = ~new_n49 & ~new_n229;
  assign new_n232 = ~new_n230 & new_n231;
  assign new_n233 = i_1_ & new_n47;
  assign new_n234 = i_6_ & new_n233;
  assign new_n235 = i_5_ & new_n179;
  assign new_n236 = i_0_ & new_n47;
  assign new_n237 = i_6_ & new_n236;
  assign new_n238 = ~new_n234 & ~new_n235;
  assign new_n239 = ~new_n237 & new_n238;
  assign new_n240 = i_5_ & new_n128;
  assign new_n241 = i_1_ & new_n210;
  assign new_n242 = i_6_ & new_n241;
  assign new_n243 = i_5_ & i_2_;
  assign new_n244 = i_1_ & new_n243;
  assign new_n245 = i_6_ & new_n244;
  assign new_n246 = ~new_n240 & ~new_n242;
  assign new_n247 = ~new_n245 & new_n246;
  assign new_n248 = new_n232 & new_n239;
  assign new_n249 = new_n247 & new_n248;
  assign new_n250 = i_5_ & new_n228;
  assign new_n251 = i_3_ & new_n128;
  assign new_n252 = i_0_ & new_n210;
  assign new_n253 = i_6_ & new_n252;
  assign new_n254 = ~new_n250 & ~new_n251;
  assign new_n255 = ~new_n253 & new_n254;
  assign new_n256 = i_4_ & new_n128;
  assign new_n257 = i_6_ & new_n202;
  assign new_n258 = i_4_ & new_n228;
  assign new_n259 = ~new_n256 & ~new_n257;
  assign new_n260 = ~new_n258 & new_n259;
  assign new_n261 = i_0_ & new_n243;
  assign new_n262 = i_6_ & new_n261;
  assign new_n263 = i_6_ & new_n216;
  assign new_n264 = i_6_ & new_n205;
  assign new_n265 = ~new_n262 & ~new_n263;
  assign new_n266 = ~new_n264 & new_n265;
  assign new_n267 = new_n255 & new_n260;
  assign new_n268 = new_n266 & new_n267;
  assign new_n269 = new_n227 & new_n249;
  assign new_n270 = new_n268 & new_n269;
  assign o_2_ = ~new_n201 | ~new_n270;
  assign new_n272 = ~i_5_ & ~i_6_;
  assign new_n273 = i_4_ & new_n272;
  assign new_n274 = new_n20 & new_n273;
  assign new_n275 = i_5_ & ~i_6_;
  assign new_n276 = i_4_ & new_n275;
  assign new_n277 = ~i_3_ & ~i_2_;
  assign new_n278 = ~i_1_ & new_n277;
  assign new_n279 = new_n276 & new_n278;
  assign new_n280 = ~i_3_ & new_n275;
  assign new_n281 = new_n42 & new_n280;
  assign new_n282 = ~new_n274 & ~new_n279;
  assign new_n283 = ~new_n281 & new_n282;
  assign new_n284 = ~i_4_ & new_n272;
  assign new_n285 = new_n14 & new_n284;
  assign new_n286 = ~i_6_ & ~i_4_;
  assign new_n287 = i_3_ & new_n286;
  assign new_n288 = new_n20 & new_n287;
  assign new_n289 = i_5_ & i_6_;
  assign new_n290 = ~i_4_ & new_n289;
  assign new_n291 = new_n55 & new_n290;
  assign new_n292 = ~new_n285 & ~new_n288;
  assign new_n293 = ~new_n291 & new_n292;
  assign new_n294 = new_n283 & new_n293;
  assign new_n295 = i_3_ & new_n272;
  assign new_n296 = new_n42 & new_n295;
  assign new_n297 = ~i_5_ & i_6_;
  assign new_n298 = ~i_4_ & new_n297;
  assign new_n299 = ~i_3_ & ~i_1_;
  assign new_n300 = i_0_ & new_n299;
  assign new_n301 = new_n298 & new_n300;
  assign new_n302 = new_n33 & new_n287;
  assign new_n303 = ~new_n296 & ~new_n301;
  assign new_n304 = ~new_n302 & new_n303;
  assign new_n305 = new_n42 & new_n298;
  assign new_n306 = new_n20 & new_n37;
  assign new_n307 = i_1_ & new_n277;
  assign new_n308 = new_n273 & new_n307;
  assign new_n309 = ~new_n305 & ~new_n306;
  assign new_n310 = ~new_n308 & new_n309;
  assign new_n311 = i_3_ & ~i_2_;
  assign new_n312 = ~i_1_ & new_n311;
  assign new_n313 = new_n298 & new_n312;
  assign new_n314 = ~i_3_ & new_n272;
  assign new_n315 = new_n29 & new_n314;
  assign new_n316 = new_n33 & new_n298;
  assign new_n317 = ~new_n313 & ~new_n315;
  assign new_n318 = ~new_n316 & new_n317;
  assign new_n319 = new_n304 & new_n310;
  assign new_n320 = new_n318 & new_n319;
  assign new_n321 = new_n294 & new_n320;
  assign new_n322 = new_n42 & new_n66;
  assign new_n323 = ~i_4_ & new_n275;
  assign new_n324 = ~i_3_ & i_2_;
  assign new_n325 = ~i_1_ & new_n324;
  assign new_n326 = new_n323 & new_n325;
  assign new_n327 = new_n33 & new_n66;
  assign new_n328 = ~new_n322 & ~new_n326;
  assign new_n329 = ~new_n327 & new_n328;
  assign new_n330 = i_3_ & new_n289;
  assign new_n331 = new_n128 & new_n330;
  assign new_n332 = new_n37 & new_n42;
  assign new_n333 = new_n20 & new_n66;
  assign new_n334 = ~new_n331 & ~new_n332;
  assign new_n335 = ~new_n333 & new_n334;
  assign new_n336 = new_n55 & new_n72;
  assign new_n337 = new_n14 & new_n27;
  assign new_n338 = i_4_ & new_n289;
  assign new_n339 = new_n128 & new_n338;
  assign new_n340 = ~new_n336 & ~new_n337;
  assign new_n341 = ~new_n339 & new_n340;
  assign new_n342 = new_n329 & new_n335;
  assign new_n343 = new_n341 & new_n342;
  assign new_n344 = new_n33 & new_n280;
  assign new_n345 = i_3_ & ~i_1_;
  assign new_n346 = ~i_0_ & new_n345;
  assign new_n347 = new_n273 & new_n346;
  assign new_n348 = i_4_ & new_n297;
  assign new_n349 = new_n55 & new_n348;
  assign new_n350 = ~new_n344 & ~new_n347;
  assign new_n351 = ~new_n349 & new_n350;
  assign new_n352 = i_3_ & new_n275;
  assign new_n353 = new_n55 & new_n352;
  assign new_n354 = new_n59 & new_n284;
  assign new_n355 = new_n228 & new_n338;
  assign new_n356 = ~new_n353 & ~new_n354;
  assign new_n357 = ~new_n355 & new_n356;
  assign new_n358 = new_n29 & new_n284;
  assign new_n359 = new_n273 & new_n325;
  assign new_n360 = i_1_ & new_n324;
  assign new_n361 = new_n284 & new_n360;
  assign new_n362 = ~new_n358 & ~new_n359;
  assign new_n363 = ~new_n361 & new_n362;
  assign new_n364 = new_n351 & new_n357;
  assign new_n365 = new_n363 & new_n364;
  assign new_n366 = new_n42 & new_n323;
  assign new_n367 = new_n216 & new_n338;
  assign new_n368 = i_6_ & i_4_;
  assign new_n369 = i_3_ & new_n368;
  assign new_n370 = new_n128 & new_n369;
  assign new_n371 = ~new_n366 & ~new_n367;
  assign new_n372 = ~new_n370 & new_n371;
  assign new_n373 = new_n27 & new_n29;
  assign new_n374 = new_n179 & new_n338;
  assign new_n375 = ~i_0_ & new_n324;
  assign new_n376 = new_n323 & new_n375;
  assign new_n377 = ~new_n373 & ~new_n374;
  assign new_n378 = ~new_n376 & new_n377;
  assign new_n379 = new_n48 & new_n128;
  assign new_n380 = new_n33 & new_n37;
  assign new_n381 = new_n307 & new_n323;
  assign new_n382 = ~new_n379 & ~new_n380;
  assign new_n383 = ~new_n381 & new_n382;
  assign new_n384 = new_n372 & new_n378;
  assign new_n385 = new_n383 & new_n384;
  assign new_n386 = new_n343 & new_n365;
  assign new_n387 = new_n385 & new_n386;
  assign o_0_ = ~new_n321 | ~new_n387;
endmodule


