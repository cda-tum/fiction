// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    _128_9_, _113_4_, _469_24_, _101_0_, _210_16_, _224_20_, _214_17_,
    _116_5_, _104_1_, _137_12_, _234_22_, _217_18_, _107_2_, _134_11_,
    _952_31_, _110_3_, _221_19_, _131_10_, _227_21_, _953_32_, _472_25_,
    _900_29_, _478_27_, _140_13_, _122_7_, _119_6_, _237_23_, _898_28_,
    _146_15_, _125_8_, _475_26_, _143_14_, _902_30_,
    _36_854_, _12_862_, _42_852_, _39_853_, _63_902_, _33_855_, _75_866_,
    _66_903_, _69_908_, _72_909_, _18_860_, _48_850_, _51_899_, _30_856_,
    _57_912_, _60_901_, _27_857_, _54_900_, _9_863_, _21_859_, _24_858_,
    _45_851_, _3_865_, _15_861_, _6_864_  );
  input  _128_9_, _113_4_, _469_24_, _101_0_, _210_16_, _224_20_,
    _214_17_, _116_5_, _104_1_, _137_12_, _234_22_, _217_18_, _107_2_,
    _134_11_, _952_31_, _110_3_, _221_19_, _131_10_, _227_21_, _953_32_,
    _472_25_, _900_29_, _478_27_, _140_13_, _122_7_, _119_6_, _237_23_,
    _898_28_, _146_15_, _125_8_, _475_26_, _143_14_, _902_30_;
  output _36_854_, _12_862_, _42_852_, _39_853_, _63_902_, _33_855_, _75_866_,
    _66_903_, _69_908_, _72_909_, _18_860_, _48_850_, _51_899_, _30_856_,
    _57_912_, _60_901_, _27_857_, _54_900_, _9_863_, _21_859_, _24_858_,
    _45_851_, _3_865_, _15_861_, _6_864_;
  wire new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157, new_n158, new_n159, new_n160,
    new_n161, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n330, new_n331, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n381, new_n382, new_n383, new_n384,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n392,
    new_n393, new_n394, new_n395, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n411, new_n412, new_n414, new_n415, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n425,
    new_n426, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n436, new_n437, new_n438, new_n439, new_n441, new_n442,
    new_n444, new_n445, new_n446, new_n447, new_n449, new_n450, new_n452,
    new_n453, new_n455, new_n456, new_n458, new_n459, new_n461, new_n462,
    new_n464, new_n465, new_n467, new_n468;
  assign new_n59 = ~_140_13_ & _125_8_;
  assign new_n60 = _140_13_ & ~_125_8_;
  assign new_n61 = ~new_n59 & ~new_n60;
  assign new_n62 = ~_146_15_ & new_n61;
  assign new_n63 = _146_15_ & ~new_n61;
  assign new_n64 = ~new_n62 & ~new_n63;
  assign new_n65 = ~_953_32_ & ~_237_23_;
  assign new_n66 = _214_17_ & new_n65;
  assign new_n67 = _143_14_ & new_n66;
  assign new_n68 = ~_143_14_ & ~new_n66;
  assign new_n69 = ~new_n67 & ~new_n68;
  assign new_n70 = ~_131_10_ & new_n69;
  assign new_n71 = _131_10_ & ~new_n69;
  assign new_n72 = ~new_n70 & ~new_n71;
  assign new_n73 = new_n64 & ~new_n72;
  assign new_n74 = ~new_n64 & new_n72;
  assign new_n75 = ~new_n73 & ~new_n74;
  assign new_n76 = ~_113_4_ & _122_7_;
  assign new_n77 = _113_4_ & ~_122_7_;
  assign new_n78 = ~new_n76 & ~new_n77;
  assign new_n79 = ~_104_1_ & new_n78;
  assign new_n80 = _104_1_ & ~new_n78;
  assign new_n81 = ~new_n79 & ~new_n80;
  assign new_n82 = new_n75 & ~new_n81;
  assign new_n83 = ~new_n75 & new_n81;
  assign new_n84 = ~new_n82 & ~new_n83;
  assign new_n85 = ~_902_30_ & ~new_n84;
  assign new_n86 = ~_475_26_ & new_n85;
  assign new_n87 = _475_26_ & ~new_n85;
  assign new_n88 = ~new_n86 & ~new_n87;
  assign new_n89 = ~_116_5_ & _122_7_;
  assign new_n90 = _116_5_ & ~_122_7_;
  assign new_n91 = ~new_n89 & ~new_n90;
  assign new_n92 = ~_107_2_ & new_n91;
  assign new_n93 = _107_2_ & ~new_n91;
  assign new_n94 = ~new_n92 & ~new_n93;
  assign new_n95 = ~_128_9_ & _143_14_;
  assign new_n96 = _128_9_ & ~_143_14_;
  assign new_n97 = ~new_n95 & ~new_n96;
  assign new_n98 = ~_134_11_ & new_n97;
  assign new_n99 = _134_11_ & ~new_n97;
  assign new_n100 = ~new_n98 & ~new_n99;
  assign new_n101 = new_n94 & ~new_n100;
  assign new_n102 = ~new_n94 & new_n100;
  assign new_n103 = ~new_n101 & ~new_n102;
  assign new_n104 = _234_22_ & ~_953_32_;
  assign new_n105 = _217_18_ & new_n104;
  assign new_n106 = new_n103 & new_n105;
  assign new_n107 = ~new_n103 & ~new_n105;
  assign new_n108 = ~new_n106 & ~new_n107;
  assign new_n109 = ~_902_30_ & ~new_n108;
  assign new_n110 = ~_478_27_ & new_n109;
  assign new_n111 = _478_27_ & ~new_n109;
  assign new_n112 = ~new_n110 & ~new_n111;
  assign new_n113 = new_n88 & ~new_n112;
  assign new_n114 = _234_22_ & _237_23_;
  assign new_n115 = ~_953_32_ & ~new_n114;
  assign new_n116 = _952_31_ & new_n115;
  assign new_n117 = _902_30_ & ~new_n114;
  assign new_n118 = _953_32_ & new_n117;
  assign new_n119 = ~_900_29_ & new_n118;
  assign new_n120 = ~new_n116 & ~new_n119;
  assign new_n121 = _110_3_ & ~_140_13_;
  assign new_n122 = ~_110_3_ & _140_13_;
  assign new_n123 = ~new_n121 & ~new_n122;
  assign new_n124 = _227_21_ & ~_953_32_;
  assign new_n125 = new_n123 & new_n124;
  assign new_n126 = ~new_n123 & ~new_n124;
  assign new_n127 = ~new_n125 & ~new_n126;
  assign new_n128 = ~_104_1_ & _107_2_;
  assign new_n129 = _104_1_ & ~_107_2_;
  assign new_n130 = ~new_n128 & ~new_n129;
  assign new_n131 = ~_101_0_ & new_n130;
  assign new_n132 = _101_0_ & ~new_n130;
  assign new_n133 = ~new_n131 & ~new_n132;
  assign new_n134 = _146_15_ & ~_143_14_;
  assign new_n135 = ~_146_15_ & _143_14_;
  assign new_n136 = ~new_n134 & ~new_n135;
  assign new_n137 = ~_128_9_ & new_n136;
  assign new_n138 = _128_9_ & ~new_n136;
  assign new_n139 = ~new_n137 & ~new_n138;
  assign new_n140 = new_n133 & new_n139;
  assign new_n141 = ~new_n133 & ~new_n139;
  assign new_n142 = ~new_n140 & ~new_n141;
  assign new_n143 = _137_12_ & ~_134_11_;
  assign new_n144 = ~_137_12_ & _134_11_;
  assign new_n145 = ~new_n143 & ~new_n144;
  assign new_n146 = ~_131_10_ & new_n145;
  assign new_n147 = _131_10_ & ~new_n145;
  assign new_n148 = ~new_n146 & ~new_n147;
  assign new_n149 = new_n142 & new_n148;
  assign new_n150 = ~new_n142 & ~new_n148;
  assign new_n151 = ~new_n149 & ~new_n150;
  assign new_n152 = new_n127 & new_n151;
  assign new_n153 = ~new_n127 & ~new_n151;
  assign new_n154 = ~new_n152 & ~new_n153;
  assign new_n155 = ~_902_30_ & ~new_n154;
  assign new_n156 = ~_469_24_ & new_n155;
  assign new_n157 = _469_24_ & ~new_n155;
  assign new_n158 = ~new_n156 & ~new_n157;
  assign new_n159 = _234_22_ & ~_902_30_;
  assign new_n160 = _221_19_ & ~new_n159;
  assign new_n161 = ~new_n158 & ~new_n160;
  assign new_n162 = _210_16_ & new_n65;
  assign new_n163 = _101_0_ & new_n162;
  assign new_n164 = ~_101_0_ & ~new_n162;
  assign new_n165 = ~new_n163 & ~new_n164;
  assign new_n166 = ~new_n139 & ~new_n148;
  assign new_n167 = new_n139 & new_n148;
  assign new_n168 = ~new_n166 & ~new_n167;
  assign new_n169 = ~_116_5_ & _119_6_;
  assign new_n170 = _116_5_ & ~_119_6_;
  assign new_n171 = ~new_n169 & ~new_n170;
  assign new_n172 = ~_113_4_ & new_n171;
  assign new_n173 = _113_4_ & ~new_n171;
  assign new_n174 = ~new_n172 & ~new_n173;
  assign new_n175 = new_n168 & new_n174;
  assign new_n176 = ~new_n168 & ~new_n174;
  assign new_n177 = ~new_n175 & ~new_n176;
  assign new_n178 = ~new_n165 & new_n177;
  assign new_n179 = new_n165 & ~new_n177;
  assign new_n180 = ~new_n178 & ~new_n179;
  assign new_n181 = ~_902_30_ & ~new_n180;
  assign new_n182 = ~_472_25_ & new_n181;
  assign new_n183 = _472_25_ & ~new_n181;
  assign new_n184 = ~new_n182 & ~new_n183;
  assign new_n185 = _128_9_ & ~_119_6_;
  assign new_n186 = ~_128_9_ & _119_6_;
  assign new_n187 = ~new_n185 & ~new_n186;
  assign new_n188 = ~_110_3_ & new_n187;
  assign new_n189 = _110_3_ & ~new_n187;
  assign new_n190 = ~new_n188 & ~new_n189;
  assign new_n191 = ~new_n64 & new_n190;
  assign new_n192 = new_n64 & ~new_n190;
  assign new_n193 = ~new_n191 & ~new_n192;
  assign new_n194 = _221_19_ & new_n104;
  assign new_n195 = ~_137_12_ & ~new_n194;
  assign new_n196 = _137_12_ & new_n194;
  assign new_n197 = ~new_n195 & ~new_n196;
  assign new_n198 = new_n193 & new_n197;
  assign new_n199 = ~new_n193 & ~new_n197;
  assign new_n200 = ~new_n198 & ~new_n199;
  assign new_n201 = ~_902_30_ & ~new_n200;
  assign new_n202 = _217_18_ & ~new_n159;
  assign new_n203 = new_n201 & ~new_n202;
  assign new_n204 = ~new_n201 & new_n202;
  assign new_n205 = ~new_n203 & ~new_n204;
  assign new_n206 = ~new_n184 & new_n205;
  assign new_n207 = ~_125_8_ & new_n139;
  assign new_n208 = _125_8_ & ~new_n139;
  assign new_n209 = ~new_n207 & ~new_n208;
  assign new_n210 = _224_20_ & ~_953_32_;
  assign new_n211 = new_n209 & new_n210;
  assign new_n212 = ~new_n209 & ~new_n210;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = ~new_n133 & ~new_n174;
  assign new_n215 = new_n133 & new_n174;
  assign new_n216 = ~new_n214 & ~new_n215;
  assign new_n217 = ~_110_3_ & _122_7_;
  assign new_n218 = _110_3_ & ~_122_7_;
  assign new_n219 = ~new_n217 & ~new_n218;
  assign new_n220 = new_n216 & new_n219;
  assign new_n221 = ~new_n216 & ~new_n219;
  assign new_n222 = ~new_n220 & ~new_n221;
  assign new_n223 = ~new_n213 & ~new_n222;
  assign new_n224 = new_n213 & new_n222;
  assign new_n225 = ~new_n223 & ~new_n224;
  assign new_n226 = ~_902_30_ & new_n225;
  assign new_n227 = ~_237_23_ & ~_902_30_;
  assign new_n228 = _210_16_ & ~new_n227;
  assign new_n229 = new_n226 & ~new_n228;
  assign new_n230 = ~new_n226 & new_n228;
  assign new_n231 = ~new_n229 & ~new_n230;
  assign new_n232 = _214_17_ & ~new_n227;
  assign new_n233 = new_n231 & ~new_n232;
  assign new_n234 = new_n113 & ~new_n120;
  assign new_n235 = new_n161 & new_n234;
  assign new_n236 = new_n206 & new_n235;
  assign new_n237 = new_n233 & new_n236;
  assign new_n238 = _134_11_ & ~new_n237;
  assign new_n239 = ~_134_11_ & new_n237;
  assign _36_854_ = new_n238 | new_n239;
  assign new_n241 = new_n88 & new_n112;
  assign new_n242 = ~_898_28_ & new_n118;
  assign new_n243 = ~new_n116 & ~new_n242;
  assign new_n244 = new_n184 & ~new_n205;
  assign new_n245 = ~new_n231 & ~new_n232;
  assign new_n246 = new_n241 & ~new_n243;
  assign new_n247 = new_n161 & new_n246;
  assign new_n248 = new_n244 & new_n247;
  assign new_n249 = new_n245 & new_n248;
  assign new_n250 = _110_3_ & ~new_n249;
  assign new_n251 = ~_110_3_ & new_n249;
  assign _12_862_ = new_n250 | new_n251;
  assign new_n253 = ~new_n88 & new_n112;
  assign new_n254 = ~new_n120 & new_n253;
  assign new_n255 = new_n161 & new_n254;
  assign new_n256 = new_n244 & new_n255;
  assign new_n257 = new_n233 & new_n256;
  assign new_n258 = _140_13_ & ~new_n257;
  assign new_n259 = ~_140_13_ & new_n257;
  assign _42_852_ = new_n258 | new_n259;
  assign new_n261 = ~new_n184 & ~new_n205;
  assign new_n262 = ~new_n120 & new_n241;
  assign new_n263 = new_n161 & new_n262;
  assign new_n264 = new_n261 & new_n263;
  assign new_n265 = new_n233 & new_n264;
  assign new_n266 = _137_12_ & ~new_n265;
  assign new_n267 = ~_137_12_ & new_n265;
  assign _39_853_ = new_n266 | new_n267;
  assign new_n269 = ~_952_31_ & _953_32_;
  assign new_n270 = new_n235 & new_n261;
  assign new_n271 = new_n245 & new_n270;
  assign new_n272 = new_n206 & new_n255;
  assign new_n273 = new_n233 & new_n272;
  assign new_n274 = new_n158 & ~new_n160;
  assign new_n275 = new_n254 & new_n274;
  assign new_n276 = new_n244 & new_n275;
  assign new_n277 = new_n245 & new_n276;
  assign new_n278 = new_n255 & new_n261;
  assign new_n279 = new_n245 & new_n278;
  assign new_n280 = ~new_n88 & ~new_n112;
  assign new_n281 = ~new_n120 & new_n280;
  assign new_n282 = new_n161 & new_n281;
  assign new_n283 = new_n206 & new_n282;
  assign new_n284 = new_n245 & new_n283;
  assign new_n285 = ~new_n237 & ~new_n265;
  assign new_n286 = ~new_n271 & new_n285;
  assign new_n287 = ~new_n273 & new_n286;
  assign new_n288 = ~new_n277 & new_n287;
  assign new_n289 = ~new_n279 & new_n288;
  assign new_n290 = ~new_n257 & new_n289;
  assign new_n291 = ~new_n284 & new_n290;
  assign new_n292 = ~new_n243 & new_n253;
  assign new_n293 = new_n274 & new_n292;
  assign new_n294 = new_n206 & new_n293;
  assign new_n295 = new_n245 & new_n294;
  assign new_n296 = new_n184 & new_n205;
  assign new_n297 = new_n161 & new_n292;
  assign new_n298 = new_n296 & new_n297;
  assign new_n299 = new_n245 & new_n298;
  assign new_n300 = new_n113 & ~new_n243;
  assign new_n301 = new_n161 & new_n300;
  assign new_n302 = new_n296 & new_n301;
  assign new_n303 = new_n245 & new_n302;
  assign new_n304 = new_n206 & new_n247;
  assign new_n305 = new_n245 & new_n304;
  assign new_n306 = ~new_n243 & new_n280;
  assign new_n307 = new_n274 & new_n306;
  assign new_n308 = new_n296 & new_n307;
  assign new_n309 = new_n245 & new_n308;
  assign new_n310 = new_n274 & new_n300;
  assign new_n311 = new_n206 & new_n310;
  assign new_n312 = new_n245 & new_n311;
  assign new_n313 = new_n246 & new_n274;
  assign new_n314 = new_n261 & new_n313;
  assign new_n315 = new_n245 & new_n314;
  assign new_n316 = ~new_n249 & ~new_n295;
  assign new_n317 = ~new_n299 & new_n316;
  assign new_n318 = ~new_n303 & new_n317;
  assign new_n319 = ~new_n305 & new_n318;
  assign new_n320 = ~new_n309 & new_n319;
  assign new_n321 = ~new_n312 & new_n320;
  assign new_n322 = ~new_n315 & new_n321;
  assign new_n323 = new_n291 & new_n322;
  assign new_n324 = _902_30_ & ~new_n323;
  assign new_n325 = _478_27_ & new_n324;
  assign new_n326 = new_n108 & new_n325;
  assign new_n327 = ~new_n108 & ~new_n325;
  assign new_n328 = ~new_n326 & ~new_n327;
  assign _63_902_ = ~new_n269 & ~new_n328;
  assign new_n330 = _131_10_ & ~new_n273;
  assign new_n331 = ~_131_10_ & new_n273;
  assign _33_855_ = new_n330 | new_n331;
  assign new_n333 = new_n116 & new_n253;
  assign new_n334 = new_n274 & new_n333;
  assign new_n335 = new_n296 & new_n334;
  assign new_n336 = new_n233 & new_n335;
  assign new_n337 = new_n113 & new_n116;
  assign new_n338 = new_n274 & new_n337;
  assign new_n339 = new_n296 & new_n338;
  assign new_n340 = new_n233 & new_n339;
  assign new_n341 = new_n116 & new_n241;
  assign new_n342 = new_n161 & new_n341;
  assign new_n343 = new_n296 & new_n342;
  assign new_n344 = new_n233 & new_n343;
  assign new_n345 = new_n274 & new_n341;
  assign new_n346 = new_n206 & new_n345;
  assign new_n347 = new_n233 & new_n346;
  assign new_n348 = new_n296 & new_n345;
  assign new_n349 = new_n245 & new_n348;
  assign new_n350 = new_n231 & new_n232;
  assign new_n351 = new_n348 & new_n350;
  assign new_n352 = new_n244 & new_n345;
  assign new_n353 = new_n233 & new_n352;
  assign new_n354 = new_n158 & new_n160;
  assign new_n355 = new_n341 & new_n354;
  assign new_n356 = new_n296 & new_n355;
  assign new_n357 = new_n233 & new_n356;
  assign new_n358 = ~new_n336 & ~new_n340;
  assign new_n359 = ~new_n344 & new_n358;
  assign new_n360 = ~new_n347 & new_n359;
  assign new_n361 = ~new_n349 & new_n360;
  assign new_n362 = ~new_n351 & new_n361;
  assign new_n363 = ~new_n353 & new_n362;
  assign new_n364 = ~new_n357 & new_n363;
  assign new_n365 = new_n291 & new_n364;
  assign new_n366 = new_n322 & new_n365;
  assign new_n367 = new_n184 & ~new_n232;
  assign new_n368 = new_n112 & new_n367;
  assign new_n369 = new_n88 & new_n368;
  assign new_n370 = new_n205 & new_n369;
  assign new_n371 = ~new_n160 & new_n370;
  assign new_n372 = new_n158 & new_n371;
  assign new_n373 = new_n231 & new_n372;
  assign new_n374 = new_n366 & ~new_n373;
  assign new_n375 = _952_31_ & new_n374;
  assign new_n376 = ~_953_32_ & new_n375;
  assign new_n377 = ~_952_31_ & ~new_n373;
  assign new_n378 = ~_952_31_ & new_n377;
  assign new_n379 = ~_953_32_ & new_n378;
  assign _75_866_ = ~new_n376 & ~new_n379;
  assign new_n381 = new_n202 & new_n324;
  assign new_n382 = new_n200 & new_n381;
  assign new_n383 = ~new_n200 & ~new_n381;
  assign new_n384 = ~new_n382 & ~new_n383;
  assign _66_903_ = ~new_n269 & ~new_n384;
  assign new_n386 = ~_953_32_ & ~new_n322;
  assign new_n387 = _953_32_ & ~_898_28_;
  assign new_n388 = new_n222 & ~new_n387;
  assign new_n389 = ~new_n386 & new_n388;
  assign new_n390 = new_n386 & ~new_n388;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = _224_20_ & _898_28_;
  assign new_n393 = _953_32_ & ~new_n392;
  assign new_n394 = new_n391 & new_n393;
  assign new_n395 = ~new_n391 & ~new_n393;
  assign _69_908_ = new_n394 | new_n395;
  assign new_n397 = ~_953_32_ & ~new_n291;
  assign new_n398 = new_n61 & new_n168;
  assign new_n399 = ~new_n61 & ~new_n168;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = _953_32_ & ~_900_29_;
  assign new_n402 = new_n400 & ~new_n401;
  assign new_n403 = ~new_n397 & new_n402;
  assign new_n404 = new_n397 & ~new_n402;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = _227_21_ & _900_29_;
  assign new_n407 = _953_32_ & ~new_n406;
  assign new_n408 = new_n405 & new_n407;
  assign new_n409 = ~new_n405 & ~new_n407;
  assign _72_909_ = new_n408 | new_n409;
  assign new_n411 = _116_5_ & ~new_n312;
  assign new_n412 = ~_116_5_ & new_n312;
  assign _18_860_ = new_n411 | new_n412;
  assign new_n414 = _146_15_ & ~new_n279;
  assign new_n415 = ~_146_15_ & new_n279;
  assign _48_850_ = new_n414 | new_n415;
  assign new_n417 = new_n213 & ~new_n222;
  assign new_n418 = ~new_n213 & new_n222;
  assign new_n419 = ~new_n417 & ~new_n418;
  assign new_n420 = new_n228 & new_n324;
  assign new_n421 = new_n419 & new_n420;
  assign new_n422 = ~new_n419 & ~new_n420;
  assign new_n423 = ~new_n421 & ~new_n422;
  assign _51_899_ = ~new_n269 & ~new_n423;
  assign new_n425 = _128_9_ & ~new_n271;
  assign new_n426 = ~_128_9_ & new_n271;
  assign _30_856_ = new_n425 | new_n426;
  assign new_n428 = _472_25_ & new_n324;
  assign new_n429 = new_n177 & new_n428;
  assign new_n430 = ~new_n177 & ~new_n428;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = ~new_n165 & new_n431;
  assign new_n433 = new_n165 & ~new_n431;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign _57_912_ = ~new_n269 & ~new_n434;
  assign new_n436 = _475_26_ & new_n324;
  assign new_n437 = new_n84 & new_n436;
  assign new_n438 = ~new_n84 & ~new_n436;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign _60_901_ = ~new_n269 & ~new_n439;
  assign new_n441 = _125_8_ & ~new_n277;
  assign new_n442 = ~_125_8_ & new_n277;
  assign _27_857_ = new_n441 | new_n442;
  assign new_n444 = _469_24_ & new_n324;
  assign new_n445 = new_n154 & new_n444;
  assign new_n446 = ~new_n154 & ~new_n444;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign _54_900_ = ~new_n269 & ~new_n447;
  assign new_n449 = _107_2_ & ~new_n303;
  assign new_n450 = ~_107_2_ & new_n303;
  assign _9_863_ = new_n449 | new_n450;
  assign new_n452 = _119_6_ & ~new_n315;
  assign new_n453 = ~_119_6_ & new_n315;
  assign _21_859_ = new_n452 | new_n453;
  assign new_n455 = _122_7_ & ~new_n309;
  assign new_n456 = ~_122_7_ & new_n309;
  assign _24_858_ = new_n455 | new_n456;
  assign new_n458 = _143_14_ & ~new_n284;
  assign new_n459 = ~_143_14_ & new_n284;
  assign _45_851_ = new_n458 | new_n459;
  assign new_n461 = _101_0_ & ~new_n305;
  assign new_n462 = ~_101_0_ & new_n305;
  assign _3_865_ = new_n461 | new_n462;
  assign new_n464 = _113_4_ & ~new_n295;
  assign new_n465 = ~_113_4_ & new_n295;
  assign _15_861_ = new_n464 | new_n465;
  assign new_n467 = _104_1_ & ~new_n299;
  assign new_n468 = ~_104_1_ & new_n299;
  assign _6_864_ = new_n467 | new_n468;
endmodule


