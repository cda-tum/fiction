// Benchmark "top" written by ABC on Mon Nov 27 17:03:31 2023

module top ( 
    count0, count1, count2, count3, count4, count5, count6, count7,
    selectp10, selectp11, selectp12, selectp13, selectp14, selectp15,
    selectp16, selectp17, selectp18, selectp19, selectp110, selectp111,
    selectp112, selectp113, selectp114, selectp115, selectp116, selectp117,
    selectp118, selectp119, selectp120, selectp121, selectp122, selectp123,
    selectp124, selectp125, selectp126, selectp127, selectp128, selectp129,
    selectp130, selectp131, selectp132, selectp133, selectp134, selectp135,
    selectp136, selectp137, selectp138, selectp139, selectp140, selectp141,
    selectp142, selectp143, selectp144, selectp145, selectp146, selectp147,
    selectp148, selectp149, selectp150, selectp151, selectp152, selectp153,
    selectp154, selectp155, selectp156, selectp157, selectp158, selectp159,
    selectp160, selectp161, selectp162, selectp163, selectp164, selectp165,
    selectp166, selectp167, selectp168, selectp169, selectp170, selectp171,
    selectp172, selectp173, selectp174, selectp175, selectp176, selectp177,
    selectp178, selectp179, selectp180, selectp181, selectp182, selectp183,
    selectp184, selectp185, selectp186, selectp187, selectp188, selectp189,
    selectp190, selectp191, selectp192, selectp193, selectp194, selectp195,
    selectp196, selectp197, selectp198, selectp199, selectp1100,
    selectp1101, selectp1102, selectp1103, selectp1104, selectp1105,
    selectp1106, selectp1107, selectp1108, selectp1109, selectp1110,
    selectp1111, selectp1112, selectp1113, selectp1114, selectp1115,
    selectp1116, selectp1117, selectp1118, selectp1119, selectp1120,
    selectp1121, selectp1122, selectp1123, selectp1124, selectp1125,
    selectp1126, selectp1127, selectp20, selectp21, selectp22, selectp23,
    selectp24, selectp25, selectp26, selectp27, selectp28, selectp29,
    selectp210, selectp211, selectp212, selectp213, selectp214, selectp215,
    selectp216, selectp217, selectp218, selectp219, selectp220, selectp221,
    selectp222, selectp223, selectp224, selectp225, selectp226, selectp227,
    selectp228, selectp229, selectp230, selectp231, selectp232, selectp233,
    selectp234, selectp235, selectp236, selectp237, selectp238, selectp239,
    selectp240, selectp241, selectp242, selectp243, selectp244, selectp245,
    selectp246, selectp247, selectp248, selectp249, selectp250, selectp251,
    selectp252, selectp253, selectp254, selectp255, selectp256, selectp257,
    selectp258, selectp259, selectp260, selectp261, selectp262, selectp263,
    selectp264, selectp265, selectp266, selectp267, selectp268, selectp269,
    selectp270, selectp271, selectp272, selectp273, selectp274, selectp275,
    selectp276, selectp277, selectp278, selectp279, selectp280, selectp281,
    selectp282, selectp283, selectp284, selectp285, selectp286, selectp287,
    selectp288, selectp289, selectp290, selectp291, selectp292, selectp293,
    selectp294, selectp295, selectp296, selectp297, selectp298, selectp299,
    selectp2100, selectp2101, selectp2102, selectp2103, selectp2104,
    selectp2105, selectp2106, selectp2107, selectp2108, selectp2109,
    selectp2110, selectp2111, selectp2112, selectp2113, selectp2114,
    selectp2115, selectp2116, selectp2117, selectp2118, selectp2119,
    selectp2120, selectp2121, selectp2122, selectp2123, selectp2124,
    selectp2125, selectp2126, selectp2127  );
  input  count0, count1, count2, count3, count4, count5, count6, count7;
  output selectp10, selectp11, selectp12, selectp13, selectp14, selectp15,
    selectp16, selectp17, selectp18, selectp19, selectp110, selectp111,
    selectp112, selectp113, selectp114, selectp115, selectp116, selectp117,
    selectp118, selectp119, selectp120, selectp121, selectp122, selectp123,
    selectp124, selectp125, selectp126, selectp127, selectp128, selectp129,
    selectp130, selectp131, selectp132, selectp133, selectp134, selectp135,
    selectp136, selectp137, selectp138, selectp139, selectp140, selectp141,
    selectp142, selectp143, selectp144, selectp145, selectp146, selectp147,
    selectp148, selectp149, selectp150, selectp151, selectp152, selectp153,
    selectp154, selectp155, selectp156, selectp157, selectp158, selectp159,
    selectp160, selectp161, selectp162, selectp163, selectp164, selectp165,
    selectp166, selectp167, selectp168, selectp169, selectp170, selectp171,
    selectp172, selectp173, selectp174, selectp175, selectp176, selectp177,
    selectp178, selectp179, selectp180, selectp181, selectp182, selectp183,
    selectp184, selectp185, selectp186, selectp187, selectp188, selectp189,
    selectp190, selectp191, selectp192, selectp193, selectp194, selectp195,
    selectp196, selectp197, selectp198, selectp199, selectp1100,
    selectp1101, selectp1102, selectp1103, selectp1104, selectp1105,
    selectp1106, selectp1107, selectp1108, selectp1109, selectp1110,
    selectp1111, selectp1112, selectp1113, selectp1114, selectp1115,
    selectp1116, selectp1117, selectp1118, selectp1119, selectp1120,
    selectp1121, selectp1122, selectp1123, selectp1124, selectp1125,
    selectp1126, selectp1127, selectp20, selectp21, selectp22, selectp23,
    selectp24, selectp25, selectp26, selectp27, selectp28, selectp29,
    selectp210, selectp211, selectp212, selectp213, selectp214, selectp215,
    selectp216, selectp217, selectp218, selectp219, selectp220, selectp221,
    selectp222, selectp223, selectp224, selectp225, selectp226, selectp227,
    selectp228, selectp229, selectp230, selectp231, selectp232, selectp233,
    selectp234, selectp235, selectp236, selectp237, selectp238, selectp239,
    selectp240, selectp241, selectp242, selectp243, selectp244, selectp245,
    selectp246, selectp247, selectp248, selectp249, selectp250, selectp251,
    selectp252, selectp253, selectp254, selectp255, selectp256, selectp257,
    selectp258, selectp259, selectp260, selectp261, selectp262, selectp263,
    selectp264, selectp265, selectp266, selectp267, selectp268, selectp269,
    selectp270, selectp271, selectp272, selectp273, selectp274, selectp275,
    selectp276, selectp277, selectp278, selectp279, selectp280, selectp281,
    selectp282, selectp283, selectp284, selectp285, selectp286, selectp287,
    selectp288, selectp289, selectp290, selectp291, selectp292, selectp293,
    selectp294, selectp295, selectp296, selectp297, selectp298, selectp299,
    selectp2100, selectp2101, selectp2102, selectp2103, selectp2104,
    selectp2105, selectp2106, selectp2107, selectp2108, selectp2109,
    selectp2110, selectp2111, selectp2112, selectp2113, selectp2114,
    selectp2115, selectp2116, selectp2117, selectp2118, selectp2119,
    selectp2120, selectp2121, selectp2122, selectp2123, selectp2124,
    selectp2125, selectp2126, selectp2127;
  wire new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n272,
    new_n273, new_n275, new_n276, new_n278, new_n280, new_n281, new_n283,
    new_n284, new_n286, new_n288, new_n290, new_n291, new_n293, new_n295,
    new_n296, new_n298, new_n300, new_n302, new_n304, new_n306, new_n308,
    new_n309, new_n326, new_n327, new_n344, new_n345, new_n362, new_n363,
    new_n380, new_n397, new_n414, new_n431, new_n432, new_n449, new_n466,
    new_n483, new_n500, new_n501, new_n518, new_n535, new_n552;
  assign new_n265 = ~count6 & count7;
  assign new_n266 = ~count4 & ~count5;
  assign new_n267 = new_n265 & new_n266;
  assign new_n268 = ~count1 & ~count3;
  assign new_n269 = ~count0 & ~count2;
  assign new_n270 = new_n268 & new_n269;
  assign selectp10 = new_n267 & new_n270;
  assign new_n272 = count0 & ~count2;
  assign new_n273 = new_n268 & new_n272;
  assign selectp11 = new_n267 & new_n273;
  assign new_n275 = count1 & ~count3;
  assign new_n276 = new_n269 & new_n275;
  assign selectp12 = new_n267 & new_n276;
  assign new_n278 = new_n272 & new_n275;
  assign selectp13 = new_n267 & new_n278;
  assign new_n280 = ~count0 & count2;
  assign new_n281 = new_n268 & new_n280;
  assign selectp14 = new_n267 & new_n281;
  assign new_n283 = count0 & count2;
  assign new_n284 = new_n268 & new_n283;
  assign selectp15 = new_n267 & new_n284;
  assign new_n286 = new_n275 & new_n280;
  assign selectp16 = new_n267 & new_n286;
  assign new_n288 = new_n275 & new_n283;
  assign selectp17 = new_n267 & new_n288;
  assign new_n290 = ~count1 & count3;
  assign new_n291 = new_n269 & new_n290;
  assign selectp18 = new_n267 & new_n291;
  assign new_n293 = new_n272 & new_n290;
  assign selectp19 = new_n267 & new_n293;
  assign new_n295 = count1 & count3;
  assign new_n296 = new_n269 & new_n295;
  assign selectp110 = new_n267 & new_n296;
  assign new_n298 = new_n272 & new_n295;
  assign selectp111 = new_n267 & new_n298;
  assign new_n300 = new_n280 & new_n290;
  assign selectp112 = new_n267 & new_n300;
  assign new_n302 = new_n283 & new_n290;
  assign selectp113 = new_n267 & new_n302;
  assign new_n304 = new_n280 & new_n295;
  assign selectp114 = new_n267 & new_n304;
  assign new_n306 = new_n283 & new_n295;
  assign selectp115 = new_n267 & new_n306;
  assign new_n308 = count4 & ~count5;
  assign new_n309 = new_n265 & new_n308;
  assign selectp116 = new_n270 & new_n309;
  assign selectp117 = new_n273 & new_n309;
  assign selectp118 = new_n276 & new_n309;
  assign selectp119 = new_n278 & new_n309;
  assign selectp120 = new_n281 & new_n309;
  assign selectp121 = new_n284 & new_n309;
  assign selectp122 = new_n286 & new_n309;
  assign selectp123 = new_n288 & new_n309;
  assign selectp124 = new_n291 & new_n309;
  assign selectp125 = new_n293 & new_n309;
  assign selectp126 = new_n296 & new_n309;
  assign selectp127 = new_n298 & new_n309;
  assign selectp128 = new_n300 & new_n309;
  assign selectp129 = new_n302 & new_n309;
  assign selectp130 = new_n304 & new_n309;
  assign selectp131 = new_n306 & new_n309;
  assign new_n326 = ~count4 & count5;
  assign new_n327 = new_n265 & new_n326;
  assign selectp132 = new_n270 & new_n327;
  assign selectp133 = new_n273 & new_n327;
  assign selectp134 = new_n276 & new_n327;
  assign selectp135 = new_n278 & new_n327;
  assign selectp136 = new_n281 & new_n327;
  assign selectp137 = new_n284 & new_n327;
  assign selectp138 = new_n286 & new_n327;
  assign selectp139 = new_n288 & new_n327;
  assign selectp140 = new_n291 & new_n327;
  assign selectp141 = new_n293 & new_n327;
  assign selectp142 = new_n296 & new_n327;
  assign selectp143 = new_n298 & new_n327;
  assign selectp144 = new_n300 & new_n327;
  assign selectp145 = new_n302 & new_n327;
  assign selectp146 = new_n304 & new_n327;
  assign selectp147 = new_n306 & new_n327;
  assign new_n344 = count4 & count5;
  assign new_n345 = new_n265 & new_n344;
  assign selectp148 = new_n270 & new_n345;
  assign selectp149 = new_n273 & new_n345;
  assign selectp150 = new_n276 & new_n345;
  assign selectp151 = new_n278 & new_n345;
  assign selectp152 = new_n281 & new_n345;
  assign selectp153 = new_n284 & new_n345;
  assign selectp154 = new_n286 & new_n345;
  assign selectp155 = new_n288 & new_n345;
  assign selectp156 = new_n291 & new_n345;
  assign selectp157 = new_n293 & new_n345;
  assign selectp158 = new_n296 & new_n345;
  assign selectp159 = new_n298 & new_n345;
  assign selectp160 = new_n300 & new_n345;
  assign selectp161 = new_n302 & new_n345;
  assign selectp162 = new_n304 & new_n345;
  assign selectp163 = new_n306 & new_n345;
  assign new_n362 = count6 & count7;
  assign new_n363 = new_n266 & new_n362;
  assign selectp164 = new_n270 & new_n363;
  assign selectp165 = new_n273 & new_n363;
  assign selectp166 = new_n276 & new_n363;
  assign selectp167 = new_n278 & new_n363;
  assign selectp168 = new_n281 & new_n363;
  assign selectp169 = new_n284 & new_n363;
  assign selectp170 = new_n286 & new_n363;
  assign selectp171 = new_n288 & new_n363;
  assign selectp172 = new_n291 & new_n363;
  assign selectp173 = new_n293 & new_n363;
  assign selectp174 = new_n296 & new_n363;
  assign selectp175 = new_n298 & new_n363;
  assign selectp176 = new_n300 & new_n363;
  assign selectp177 = new_n302 & new_n363;
  assign selectp178 = new_n304 & new_n363;
  assign selectp179 = new_n306 & new_n363;
  assign new_n380 = new_n308 & new_n362;
  assign selectp180 = new_n270 & new_n380;
  assign selectp181 = new_n273 & new_n380;
  assign selectp182 = new_n276 & new_n380;
  assign selectp183 = new_n278 & new_n380;
  assign selectp184 = new_n281 & new_n380;
  assign selectp185 = new_n284 & new_n380;
  assign selectp186 = new_n286 & new_n380;
  assign selectp187 = new_n288 & new_n380;
  assign selectp188 = new_n291 & new_n380;
  assign selectp189 = new_n293 & new_n380;
  assign selectp190 = new_n296 & new_n380;
  assign selectp191 = new_n298 & new_n380;
  assign selectp192 = new_n300 & new_n380;
  assign selectp193 = new_n302 & new_n380;
  assign selectp194 = new_n304 & new_n380;
  assign selectp195 = new_n306 & new_n380;
  assign new_n397 = new_n326 & new_n362;
  assign selectp196 = new_n270 & new_n397;
  assign selectp197 = new_n273 & new_n397;
  assign selectp198 = new_n276 & new_n397;
  assign selectp199 = new_n278 & new_n397;
  assign selectp1100 = new_n281 & new_n397;
  assign selectp1101 = new_n284 & new_n397;
  assign selectp1102 = new_n286 & new_n397;
  assign selectp1103 = new_n288 & new_n397;
  assign selectp1104 = new_n291 & new_n397;
  assign selectp1105 = new_n293 & new_n397;
  assign selectp1106 = new_n296 & new_n397;
  assign selectp1107 = new_n298 & new_n397;
  assign selectp1108 = new_n300 & new_n397;
  assign selectp1109 = new_n302 & new_n397;
  assign selectp1110 = new_n304 & new_n397;
  assign selectp1111 = new_n306 & new_n397;
  assign new_n414 = new_n344 & new_n362;
  assign selectp1112 = new_n270 & new_n414;
  assign selectp1113 = new_n273 & new_n414;
  assign selectp1114 = new_n276 & new_n414;
  assign selectp1115 = new_n278 & new_n414;
  assign selectp1116 = new_n281 & new_n414;
  assign selectp1117 = new_n284 & new_n414;
  assign selectp1118 = new_n286 & new_n414;
  assign selectp1119 = new_n288 & new_n414;
  assign selectp1120 = new_n291 & new_n414;
  assign selectp1121 = new_n293 & new_n414;
  assign selectp1122 = new_n296 & new_n414;
  assign selectp1123 = new_n298 & new_n414;
  assign selectp1124 = new_n300 & new_n414;
  assign selectp1125 = new_n302 & new_n414;
  assign selectp1126 = new_n304 & new_n414;
  assign selectp1127 = new_n306 & new_n414;
  assign new_n431 = ~count6 & ~count7;
  assign new_n432 = new_n266 & new_n431;
  assign selectp20 = new_n270 & new_n432;
  assign selectp21 = new_n273 & new_n432;
  assign selectp22 = new_n276 & new_n432;
  assign selectp23 = new_n278 & new_n432;
  assign selectp24 = new_n281 & new_n432;
  assign selectp25 = new_n284 & new_n432;
  assign selectp26 = new_n286 & new_n432;
  assign selectp27 = new_n288 & new_n432;
  assign selectp28 = new_n291 & new_n432;
  assign selectp29 = new_n293 & new_n432;
  assign selectp210 = new_n296 & new_n432;
  assign selectp211 = new_n298 & new_n432;
  assign selectp212 = new_n300 & new_n432;
  assign selectp213 = new_n302 & new_n432;
  assign selectp214 = new_n304 & new_n432;
  assign selectp215 = new_n306 & new_n432;
  assign new_n449 = new_n308 & new_n431;
  assign selectp216 = new_n270 & new_n449;
  assign selectp217 = new_n273 & new_n449;
  assign selectp218 = new_n276 & new_n449;
  assign selectp219 = new_n278 & new_n449;
  assign selectp220 = new_n281 & new_n449;
  assign selectp221 = new_n284 & new_n449;
  assign selectp222 = new_n286 & new_n449;
  assign selectp223 = new_n288 & new_n449;
  assign selectp224 = new_n291 & new_n449;
  assign selectp225 = new_n293 & new_n449;
  assign selectp226 = new_n296 & new_n449;
  assign selectp227 = new_n298 & new_n449;
  assign selectp228 = new_n300 & new_n449;
  assign selectp229 = new_n302 & new_n449;
  assign selectp230 = new_n304 & new_n449;
  assign selectp231 = new_n306 & new_n449;
  assign new_n466 = new_n326 & new_n431;
  assign selectp232 = new_n270 & new_n466;
  assign selectp233 = new_n273 & new_n466;
  assign selectp234 = new_n276 & new_n466;
  assign selectp235 = new_n278 & new_n466;
  assign selectp236 = new_n281 & new_n466;
  assign selectp237 = new_n284 & new_n466;
  assign selectp238 = new_n286 & new_n466;
  assign selectp239 = new_n288 & new_n466;
  assign selectp240 = new_n291 & new_n466;
  assign selectp241 = new_n293 & new_n466;
  assign selectp242 = new_n296 & new_n466;
  assign selectp243 = new_n298 & new_n466;
  assign selectp244 = new_n300 & new_n466;
  assign selectp245 = new_n302 & new_n466;
  assign selectp246 = new_n304 & new_n466;
  assign selectp247 = new_n306 & new_n466;
  assign new_n483 = new_n344 & new_n431;
  assign selectp248 = new_n270 & new_n483;
  assign selectp249 = new_n273 & new_n483;
  assign selectp250 = new_n276 & new_n483;
  assign selectp251 = new_n278 & new_n483;
  assign selectp252 = new_n281 & new_n483;
  assign selectp253 = new_n284 & new_n483;
  assign selectp254 = new_n286 & new_n483;
  assign selectp255 = new_n288 & new_n483;
  assign selectp256 = new_n291 & new_n483;
  assign selectp257 = new_n293 & new_n483;
  assign selectp258 = new_n296 & new_n483;
  assign selectp259 = new_n298 & new_n483;
  assign selectp260 = new_n300 & new_n483;
  assign selectp261 = new_n302 & new_n483;
  assign selectp262 = new_n304 & new_n483;
  assign selectp263 = new_n306 & new_n483;
  assign new_n500 = count6 & ~count7;
  assign new_n501 = new_n266 & new_n500;
  assign selectp264 = new_n270 & new_n501;
  assign selectp265 = new_n273 & new_n501;
  assign selectp266 = new_n276 & new_n501;
  assign selectp267 = new_n278 & new_n501;
  assign selectp268 = new_n281 & new_n501;
  assign selectp269 = new_n284 & new_n501;
  assign selectp270 = new_n286 & new_n501;
  assign selectp271 = new_n288 & new_n501;
  assign selectp272 = new_n291 & new_n501;
  assign selectp273 = new_n293 & new_n501;
  assign selectp274 = new_n296 & new_n501;
  assign selectp275 = new_n298 & new_n501;
  assign selectp276 = new_n300 & new_n501;
  assign selectp277 = new_n302 & new_n501;
  assign selectp278 = new_n304 & new_n501;
  assign selectp279 = new_n306 & new_n501;
  assign new_n518 = new_n308 & new_n500;
  assign selectp280 = new_n270 & new_n518;
  assign selectp281 = new_n273 & new_n518;
  assign selectp282 = new_n276 & new_n518;
  assign selectp283 = new_n278 & new_n518;
  assign selectp284 = new_n281 & new_n518;
  assign selectp285 = new_n284 & new_n518;
  assign selectp286 = new_n286 & new_n518;
  assign selectp287 = new_n288 & new_n518;
  assign selectp288 = new_n291 & new_n518;
  assign selectp289 = new_n293 & new_n518;
  assign selectp290 = new_n296 & new_n518;
  assign selectp291 = new_n298 & new_n518;
  assign selectp292 = new_n300 & new_n518;
  assign selectp293 = new_n302 & new_n518;
  assign selectp294 = new_n304 & new_n518;
  assign selectp295 = new_n306 & new_n518;
  assign new_n535 = new_n326 & new_n500;
  assign selectp296 = new_n270 & new_n535;
  assign selectp297 = new_n273 & new_n535;
  assign selectp298 = new_n276 & new_n535;
  assign selectp299 = new_n278 & new_n535;
  assign selectp2100 = new_n281 & new_n535;
  assign selectp2101 = new_n284 & new_n535;
  assign selectp2102 = new_n286 & new_n535;
  assign selectp2103 = new_n288 & new_n535;
  assign selectp2104 = new_n291 & new_n535;
  assign selectp2105 = new_n293 & new_n535;
  assign selectp2106 = new_n296 & new_n535;
  assign selectp2107 = new_n298 & new_n535;
  assign selectp2108 = new_n300 & new_n535;
  assign selectp2109 = new_n302 & new_n535;
  assign selectp2110 = new_n304 & new_n535;
  assign selectp2111 = new_n306 & new_n535;
  assign new_n552 = new_n344 & new_n500;
  assign selectp2112 = new_n270 & new_n552;
  assign selectp2113 = new_n273 & new_n552;
  assign selectp2114 = new_n276 & new_n552;
  assign selectp2115 = new_n278 & new_n552;
  assign selectp2116 = new_n281 & new_n552;
  assign selectp2117 = new_n284 & new_n552;
  assign selectp2118 = new_n286 & new_n552;
  assign selectp2119 = new_n288 & new_n552;
  assign selectp2120 = new_n291 & new_n552;
  assign selectp2121 = new_n293 & new_n552;
  assign selectp2122 = new_n296 & new_n552;
  assign selectp2123 = new_n298 & new_n552;
  assign selectp2124 = new_n300 & new_n552;
  assign selectp2125 = new_n302 & new_n552;
  assign selectp2126 = new_n304 & new_n552;
  assign selectp2127 = new_n306 & new_n552;
endmodule


