// Benchmark "b11" written by ABC on Wed Sep  5 10:17:20 2018

module b11 ( clock, 
    X_IN_5_, X_IN_4_, X_IN_3_, X_IN_2_, X_IN_1_, X_IN_0_, STBI,
    X_OUT_REG_5_, X_OUT_REG_4_, X_OUT_REG_3_, X_OUT_REG_2_, X_OUT_REG_1_,
    X_OUT_REG_0_  );
  input  clock;
  input  X_IN_5_, X_IN_4_, X_IN_3_, X_IN_2_, X_IN_1_, X_IN_0_, STBI;
  output X_OUT_REG_5_, X_OUT_REG_4_, X_OUT_REG_3_, X_OUT_REG_2_, X_OUT_REG_1_,
    X_OUT_REG_0_;
  reg R_IN_REG_5_, R_IN_REG_4_, R_IN_REG_3_, R_IN_REG_2_, R_IN_REG_1_,
    R_IN_REG_0_, CONT_REG_5_, CONT_REG_4_, CONT_REG_3_, CONT_REG_2_,
    CONT_REG_1_, CONT_REG_0_, CONT1_REG_8_, CONT1_REG_7_, CONT1_REG_6_,
    CONT1_REG_5_, CONT1_REG_4_, CONT1_REG_3_, CONT1_REG_2_, CONT1_REG_1_,
    CONT1_REG_0_, X_OUT_REG_5_, X_OUT_REG_4_, X_OUT_REG_3_, X_OUT_REG_2_,
    X_OUT_REG_1_, X_OUT_REG_0_, STATO_REG_3_, STATO_REG_2_, STATO_REG_1_,
    STATO_REG_0_;
  wire n107, n108_1, n109, n110, n112, n113_1, n115, n116, n118_1, n119,
    n121, n122, n124, n125, n127, n128_1, n129, n130, n131, n132, n133_1,
    n134, n135, n136, n137_1, n138, n139, n140, n141_1, n142, n143, n144,
    n145_1, n146, n147, n148, n149_1, n150, n151, n152, n153_1, n154, n155,
    n156, n157_1, n158, n159, n160, n161, n162_1, n163, n164, n165, n166,
    n167_1, n168, n169, n170, n171, n172_1, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n189, n190,
    n191, n192, n193, n195, n196, n197, n198, n199, n201, n202, n203, n204,
    n205, n207, n208, n209, n210, n211, n213, n214, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n658, n659, n660,
    n661, n662, n663, n664, n666, n667, n668, n669, n670, n672, n673, n674,
    n675, n677, n678, n679, n680, n682, n683, n684, n685, n687, n688, n689,
    n690, n692, n694, n695, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n28,
    n33, n38, n43, n48, n53, n58, n63, n68, n73, n78, n83, n88, n93, n98,
    n103, n108, n113, n118, n123, n128, n133, n137, n141, n145, n149, n153,
    n157, n162, n167, n172;
  assign n107 = ~STATO_REG_2_ & ~STATO_REG_1_;
  assign n108_1 = ~STATO_REG_3_ & n107;
  assign n109 = X_IN_5_ & n108_1;
  assign n110 = R_IN_REG_5_ & ~n108_1;
  assign n28 = n109 | n110;
  assign n112 = X_IN_4_ & n108_1;
  assign n113_1 = R_IN_REG_4_ & ~n108_1;
  assign n33 = n112 | n113_1;
  assign n115 = X_IN_3_ & n108_1;
  assign n116 = R_IN_REG_3_ & ~n108_1;
  assign n38 = n115 | n116;
  assign n118_1 = X_IN_2_ & n108_1;
  assign n119 = R_IN_REG_2_ & ~n108_1;
  assign n43 = n118_1 | n119;
  assign n121 = X_IN_1_ & n108_1;
  assign n122 = R_IN_REG_1_ & ~n108_1;
  assign n48 = n121 | n122;
  assign n124 = X_IN_0_ & n108_1;
  assign n125 = R_IN_REG_0_ & ~n108_1;
  assign n53 = n124 | n125;
  assign n127 = ~STATO_REG_2_ & STATO_REG_1_;
  assign n128_1 = ~STATO_REG_0_ & n127;
  assign n129 = ~R_IN_REG_2_ & R_IN_REG_1_;
  assign n130 = R_IN_REG_3_ & ~R_IN_REG_1_;
  assign n131 = R_IN_REG_2_ & ~R_IN_REG_0_;
  assign n132 = ~R_IN_REG_4_ & R_IN_REG_0_;
  assign n133_1 = R_IN_REG_5_ & ~R_IN_REG_3_;
  assign n134 = ~R_IN_REG_5_ & R_IN_REG_4_;
  assign n135 = ~n131 & ~n132;
  assign n136 = ~n133_1 & n135;
  assign n137_1 = ~n134 & n136;
  assign n138 = ~n129 & ~n130;
  assign n139 = n137_1 & n138;
  assign n140 = n128_1 & n139;
  assign n141_1 = ~STATO_REG_0_ & n107;
  assign n142 = ~STATO_REG_3_ & n141_1;
  assign n143 = ~n140 & ~n142;
  assign n144 = CONT_REG_5_ & n143;
  assign n145_1 = CONT_REG_1_ & CONT_REG_0_;
  assign n146 = CONT_REG_2_ & n145_1;
  assign n147 = CONT_REG_3_ & n146;
  assign n148 = CONT_REG_4_ & n147;
  assign n149_1 = ~CONT_REG_5_ & n148;
  assign n150 = CONT_REG_5_ & ~n148;
  assign n151 = ~n149_1 & ~n150;
  assign n152 = CONT_REG_5_ & n139;
  assign n153_1 = R_IN_REG_5_ & ~n139;
  assign n154 = n152 & ~n153_1;
  assign n155 = ~R_IN_REG_3_ & ~n139;
  assign n156 = ~CONT_REG_3_ & n139;
  assign n157_1 = ~n155 & n156;
  assign n158 = ~R_IN_REG_4_ & ~n139;
  assign n159 = ~CONT_REG_4_ & n139;
  assign n160 = ~n158 & n159;
  assign n161 = CONT_REG_2_ & n139;
  assign n162_1 = R_IN_REG_2_ & ~n139;
  assign n163 = n161 & ~n162_1;
  assign n164 = n155 & ~n156;
  assign n165 = R_IN_REG_1_ & ~n139;
  assign n166 = ~CONT_REG_1_ & n139;
  assign n167_1 = n165 & n166;
  assign n168 = ~n161 & n162_1;
  assign n169 = ~R_IN_REG_0_ & ~n139;
  assign n170 = CONT_REG_0_ & n139;
  assign n171 = ~n165 & ~n166;
  assign n172_1 = ~n169 & ~n170;
  assign n173 = ~n171 & n172_1;
  assign n174 = ~n167_1 & ~n168;
  assign n175 = ~n173 & n174;
  assign n176 = ~n163 & ~n164;
  assign n177 = ~n175 & n176;
  assign n178 = ~n157_1 & ~n160;
  assign n179 = ~n177 & n178;
  assign n180 = n158 & ~n159;
  assign n181 = ~n179 & ~n180;
  assign n182 = ~n152 & n153_1;
  assign n183 = ~n181 & ~n182;
  assign n184 = ~n154 & ~n183;
  assign n185 = STATO_REG_1_ & ~n143;
  assign n186 = n184 & n185;
  assign n187 = ~n151 & n186;
  assign n58 = n144 | n187;
  assign n189 = CONT_REG_4_ & n143;
  assign n190 = ~CONT_REG_4_ & n147;
  assign n191 = CONT_REG_4_ & ~n147;
  assign n192 = ~n190 & ~n191;
  assign n193 = n186 & ~n192;
  assign n63 = n189 | n193;
  assign n195 = CONT_REG_3_ & n143;
  assign n196 = ~CONT_REG_3_ & n146;
  assign n197 = CONT_REG_3_ & ~n146;
  assign n198 = ~n196 & ~n197;
  assign n199 = n186 & ~n198;
  assign n68 = n195 | n199;
  assign n201 = CONT_REG_2_ & n143;
  assign n202 = ~CONT_REG_2_ & n145_1;
  assign n203 = CONT_REG_2_ & ~n145_1;
  assign n204 = ~n202 & ~n203;
  assign n205 = n186 & ~n204;
  assign n73 = n201 | n205;
  assign n207 = CONT_REG_1_ & n143;
  assign n208 = ~CONT_REG_1_ & CONT_REG_0_;
  assign n209 = CONT_REG_1_ & ~CONT_REG_0_;
  assign n210 = ~n208 & ~n209;
  assign n211 = n186 & ~n210;
  assign n78 = n207 | n211;
  assign n213 = CONT_REG_0_ & n143;
  assign n214 = ~CONT_REG_0_ & n186;
  assign n83 = n213 | n214;
  assign n216 = CONT1_REG_2_ & CONT1_REG_1_;
  assign n217 = ~CONT1_REG_3_ & ~n216;
  assign n218 = ~CONT1_REG_4_ & n217;
  assign n219 = CONT1_REG_5_ & ~n218;
  assign n220 = CONT1_REG_6_ & n219;
  assign n221 = CONT1_REG_7_ & n220;
  assign n222 = ~CONT1_REG_8_ & n221;
  assign n223 = CONT1_REG_8_ & ~n221;
  assign n224 = ~n222 & ~n223;
  assign n225 = STATO_REG_2_ & STATO_REG_1_;
  assign n226 = STATO_REG_1_ & STATO_REG_0_;
  assign n227 = n127 & n139;
  assign n228 = ~CONT1_REG_7_ & ~CONT1_REG_6_;
  assign n229 = ~CONT1_REG_8_ & ~n228;
  assign n230 = STATO_REG_1_ & ~n229;
  assign n231 = CONT1_REG_1_ & CONT1_REG_0_;
  assign n232 = ~CONT1_REG_2_ & ~n231;
  assign n233 = CONT1_REG_4_ & CONT1_REG_3_;
  assign n234 = ~n232 & n233;
  assign n235 = ~CONT1_REG_6_ & ~n234;
  assign n236 = ~CONT1_REG_7_ & n235;
  assign n237 = ~CONT1_REG_5_ & n236;
  assign n238 = ~CONT1_REG_8_ & ~n237;
  assign n239 = STATO_REG_0_ & ~n238;
  assign n240 = STATO_REG_2_ & ~n230;
  assign n241 = ~n239 & n240;
  assign n242 = ~n226 & ~n227;
  assign n243 = ~n241 & n242;
  assign n244 = n225 & ~n243;
  assign n245 = ~STATO_REG_0_ & n244;
  assign n246 = ~n224 & n245;
  assign n247 = CONT1_REG_5_ & STATO_REG_3_;
  assign n248 = CONT1_REG_8_ & ~STATO_REG_3_;
  assign n249 = n247 & ~n248;
  assign n250 = ~n247 & n248;
  assign n251 = ~n249 & ~n250;
  assign n252 = CONT1_REG_6_ & ~STATO_REG_3_;
  assign n253 = ~n247 & n252;
  assign n254 = n247 & ~n252;
  assign n255 = CONT1_REG_5_ & ~STATO_REG_3_;
  assign n256 = ~n247 & n255;
  assign n257 = n247 & ~n255;
  assign n258 = CONT1_REG_3_ & ~STATO_REG_3_;
  assign n259 = ~CONT1_REG_3_ & STATO_REG_3_;
  assign n260 = n258 & n259;
  assign n261 = ~n258 & ~n259;
  assign n262 = CONT1_REG_1_ & ~STATO_REG_3_;
  assign n263 = ~CONT1_REG_1_ & STATO_REG_3_;
  assign n264 = n262 & n263;
  assign n265 = ~n262 & ~n263;
  assign n266 = CONT1_REG_0_ & STATO_REG_3_;
  assign n267 = CONT1_REG_0_ & ~STATO_REG_3_;
  assign n268 = n266 & ~n267;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~n264 & ~n269;
  assign n271 = CONT1_REG_2_ & STATO_REG_3_;
  assign n272 = ~n270 & ~n271;
  assign n273 = CONT1_REG_2_ & ~STATO_REG_3_;
  assign n274 = n270 & n271;
  assign n275 = n273 & ~n274;
  assign n276 = ~n272 & ~n275;
  assign n277 = ~n261 & ~n276;
  assign n278 = ~n260 & ~n277;
  assign n279 = ~CONT1_REG_4_ & STATO_REG_3_;
  assign n280 = ~n278 & n279;
  assign n281 = CONT1_REG_4_ & ~STATO_REG_3_;
  assign n282 = n278 & ~n279;
  assign n283 = n281 & ~n282;
  assign n284 = ~n280 & ~n283;
  assign n285 = ~n257 & ~n284;
  assign n286 = ~n256 & ~n285;
  assign n287 = ~n254 & ~n286;
  assign n288 = ~n253 & ~n287;
  assign n289 = ~n247 & ~n288;
  assign n290 = CONT1_REG_7_ & ~STATO_REG_3_;
  assign n291 = n247 & n288;
  assign n292 = n290 & ~n291;
  assign n293 = ~n289 & ~n292;
  assign n294 = ~n251 & ~n293;
  assign n295 = n251 & n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = ~STATO_REG_1_ & ~n243;
  assign n298 = STATO_REG_0_ & n297;
  assign n299 = ~n296 & n298;
  assign n300 = CONT1_REG_8_ & n243;
  assign n301 = R_IN_REG_1_ & CONT1_REG_8_;
  assign n302 = ~R_IN_REG_1_ & ~CONT1_REG_8_;
  assign n303 = ~n301 & ~n302;
  assign n304 = R_IN_REG_1_ & CONT1_REG_6_;
  assign n305 = ~R_IN_REG_1_ & ~CONT1_REG_6_;
  assign n306 = ~n304 & ~n305;
  assign n307 = R_IN_REG_1_ & CONT1_REG_5_;
  assign n308 = ~R_IN_REG_1_ & ~CONT1_REG_5_;
  assign n309 = ~n307 & ~n308;
  assign n310 = R_IN_REG_5_ & ~n309;
  assign n311 = ~R_IN_REG_5_ & n309;
  assign n312 = R_IN_REG_1_ & CONT1_REG_4_;
  assign n313 = ~R_IN_REG_1_ & ~CONT1_REG_4_;
  assign n314 = ~n312 & ~n313;
  assign n315 = R_IN_REG_4_ & ~n314;
  assign n316 = ~R_IN_REG_4_ & n314;
  assign n317 = R_IN_REG_1_ & CONT1_REG_3_;
  assign n318 = ~R_IN_REG_1_ & ~CONT1_REG_3_;
  assign n319 = ~n317 & ~n318;
  assign n320 = R_IN_REG_3_ & ~n319;
  assign n321 = ~R_IN_REG_3_ & n319;
  assign n322 = R_IN_REG_1_ & CONT1_REG_2_;
  assign n323 = ~R_IN_REG_1_ & ~CONT1_REG_2_;
  assign n324 = ~n322 & ~n323;
  assign n325 = R_IN_REG_2_ & ~n324;
  assign n326 = ~R_IN_REG_2_ & n324;
  assign n327 = R_IN_REG_1_ & CONT1_REG_1_;
  assign n328 = ~R_IN_REG_1_ & ~CONT1_REG_1_;
  assign n329 = ~n327 & ~n328;
  assign n330 = R_IN_REG_1_ & ~n329;
  assign n331 = ~R_IN_REG_1_ & n329;
  assign n332 = R_IN_REG_1_ & CONT1_REG_0_;
  assign n333 = ~R_IN_REG_1_ & ~CONT1_REG_0_;
  assign n334 = ~n332 & ~n333;
  assign n335 = R_IN_REG_0_ & ~n334;
  assign n336 = ~R_IN_REG_0_ & n334;
  assign n337 = ~R_IN_REG_1_ & ~n336;
  assign n338 = ~n335 & ~n337;
  assign n339 = ~n331 & ~n338;
  assign n340 = ~n330 & ~n339;
  assign n341 = ~n326 & ~n340;
  assign n342 = ~n325 & ~n341;
  assign n343 = ~n321 & ~n342;
  assign n344 = ~n320 & ~n343;
  assign n345 = ~n316 & ~n344;
  assign n346 = ~n315 & ~n345;
  assign n347 = ~n311 & ~n346;
  assign n348 = ~n310 & ~n347;
  assign n349 = ~n306 & ~n348;
  assign n350 = R_IN_REG_1_ & CONT1_REG_7_;
  assign n351 = ~R_IN_REG_1_ & ~CONT1_REG_7_;
  assign n352 = ~n350 & ~n351;
  assign n353 = n349 & ~n352;
  assign n354 = ~n303 & ~n353;
  assign n355 = n303 & n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~STATO_REG_0_ & n297;
  assign n358 = ~n356 & n357;
  assign n359 = R_IN_REG_3_ & CONT1_REG_8_;
  assign n360 = ~R_IN_REG_3_ & ~CONT1_REG_8_;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~R_IN_REG_3_ & R_IN_REG_2_;
  assign n363 = R_IN_REG_3_ & ~R_IN_REG_2_;
  assign n364 = ~n362 & ~n363;
  assign n365 = R_IN_REG_3_ & ~n364;
  assign n366 = ~R_IN_REG_3_ & n364;
  assign n367 = ~n365 & ~n366;
  assign n368 = CONT1_REG_4_ & n367;
  assign n369 = ~CONT1_REG_4_ & ~n367;
  assign n370 = R_IN_REG_3_ & R_IN_REG_2_;
  assign n371 = ~R_IN_REG_3_ & ~R_IN_REG_2_;
  assign n372 = ~n370 & ~n371;
  assign n373 = CONT1_REG_3_ & ~n372;
  assign n374 = ~CONT1_REG_3_ & n372;
  assign n375 = R_IN_REG_3_ & n362;
  assign n376 = ~R_IN_REG_3_ & ~n362;
  assign n377 = ~n375 & ~n376;
  assign n378 = CONT1_REG_2_ & n377;
  assign n379 = ~CONT1_REG_2_ & ~n377;
  assign n380 = CONT1_REG_0_ & n372;
  assign n381 = ~CONT1_REG_0_ & ~n372;
  assign n382 = ~R_IN_REG_3_ & ~n381;
  assign n383 = ~n380 & ~n382;
  assign n384 = ~n367 & ~n383;
  assign n385 = n367 & n383;
  assign n386 = CONT1_REG_1_ & ~n385;
  assign n387 = ~n384 & ~n386;
  assign n388 = ~n379 & ~n387;
  assign n389 = ~n378 & ~n388;
  assign n390 = ~n374 & ~n389;
  assign n391 = ~n373 & ~n390;
  assign n392 = ~n369 & ~n391;
  assign n393 = ~n368 & ~n392;
  assign n394 = CONT1_REG_5_ & ~n393;
  assign n395 = ~CONT1_REG_5_ & n393;
  assign n396 = ~n377 & ~n395;
  assign n397 = ~n394 & ~n396;
  assign n398 = CONT1_REG_6_ & ~n397;
  assign n399 = ~CONT1_REG_6_ & n397;
  assign n400 = ~R_IN_REG_3_ & ~n399;
  assign n401 = ~n398 & ~n400;
  assign n402 = CONT1_REG_7_ & ~n401;
  assign n403 = ~CONT1_REG_7_ & n401;
  assign n404 = ~R_IN_REG_3_ & ~n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = ~n361 & ~n405;
  assign n407 = n361 & n405;
  assign n408 = ~n406 & ~n407;
  assign n409 = STATO_REG_0_ & n244;
  assign n410 = n408 & n409;
  assign n411 = ~n246 & ~n299;
  assign n412 = ~n300 & n411;
  assign n413 = ~n358 & n412;
  assign n88 = n410 | ~n413;
  assign n415 = ~CONT1_REG_7_ & n220;
  assign n416 = CONT1_REG_7_ & ~n220;
  assign n417 = ~n415 & ~n416;
  assign n418 = n245 & ~n417;
  assign n419 = n247 & ~n290;
  assign n420 = ~n247 & n290;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n288 & ~n421;
  assign n423 = n288 & n421;
  assign n424 = ~n422 & ~n423;
  assign n425 = n298 & ~n424;
  assign n426 = CONT1_REG_7_ & n243;
  assign n427 = ~n349 & ~n352;
  assign n428 = n349 & n352;
  assign n429 = ~n427 & ~n428;
  assign n430 = n357 & ~n429;
  assign n431 = R_IN_REG_3_ & CONT1_REG_7_;
  assign n432 = ~R_IN_REG_3_ & ~CONT1_REG_7_;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n401 & ~n433;
  assign n435 = n401 & n433;
  assign n436 = ~n434 & ~n435;
  assign n437 = n409 & n436;
  assign n438 = ~n418 & ~n425;
  assign n439 = ~n426 & n438;
  assign n440 = ~n430 & n439;
  assign n93 = n437 | ~n440;
  assign n442 = ~CONT1_REG_6_ & n219;
  assign n443 = CONT1_REG_6_ & ~n219;
  assign n444 = ~n442 & ~n443;
  assign n445 = n245 & ~n444;
  assign n446 = ~STATO_REG_2_ & ~n243;
  assign n447 = STATO_REG_0_ & n446;
  assign n448 = R_IN_REG_0_ & n447;
  assign n449 = CONT_REG_5_ & n448;
  assign n450 = n306 & n348;
  assign n451 = ~n349 & ~n450;
  assign n452 = n357 & n451;
  assign n453 = CONT1_REG_6_ & n243;
  assign n454 = ~n253 & ~n254;
  assign n455 = ~n286 & ~n454;
  assign n456 = n286 & n454;
  assign n457 = ~n455 & ~n456;
  assign n458 = n298 & ~n457;
  assign n459 = R_IN_REG_3_ & CONT1_REG_6_;
  assign n460 = ~R_IN_REG_3_ & ~CONT1_REG_6_;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n397 & ~n461;
  assign n463 = n397 & n461;
  assign n464 = ~n462 & ~n463;
  assign n465 = n409 & n464;
  assign n466 = ~n453 & ~n458;
  assign n467 = ~n465 & n466;
  assign n468 = ~n445 & ~n449;
  assign n469 = ~n452 & n468;
  assign n98 = ~n467 | ~n469;
  assign n471 = CONT_REG_4_ & n448;
  assign n472 = ~R_IN_REG_0_ & n447;
  assign n473 = CONT_REG_5_ & n472;
  assign n474 = ~n256 & ~n257;
  assign n475 = ~n284 & ~n474;
  assign n476 = n284 & n474;
  assign n477 = ~n475 & ~n476;
  assign n478 = n298 & ~n477;
  assign n479 = CONT1_REG_5_ & n243;
  assign n480 = ~CONT1_REG_5_ & ~n377;
  assign n481 = CONT1_REG_5_ & n377;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n393 & ~n482;
  assign n484 = n393 & n482;
  assign n485 = ~n483 & ~n484;
  assign n486 = n409 & n485;
  assign n487 = ~n479 & ~n486;
  assign n488 = ~CONT1_REG_5_ & ~CONT1_REG_4_;
  assign n489 = n217 & n488;
  assign n490 = ~n219 & ~n489;
  assign n491 = n244 & n490;
  assign n492 = R_IN_REG_5_ & n446;
  assign n493 = ~n310 & ~n311;
  assign n494 = n346 & n493;
  assign n495 = ~n346 & ~n493;
  assign n496 = ~n494 & ~n495;
  assign n497 = n297 & ~n496;
  assign n498 = ~n491 & ~n492;
  assign n499 = ~n497 & n498;
  assign n500 = ~STATO_REG_0_ & ~n499;
  assign n501 = ~n471 & ~n473;
  assign n502 = ~n478 & n501;
  assign n503 = n487 & n502;
  assign n103 = n500 | ~n503;
  assign n505 = CONT_REG_3_ & n448;
  assign n506 = CONT_REG_4_ & n472;
  assign n507 = ~n279 & ~n281;
  assign n508 = n279 & n281;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~n278 & ~n509;
  assign n511 = n278 & n509;
  assign n512 = ~n510 & ~n511;
  assign n513 = n298 & ~n512;
  assign n514 = CONT1_REG_4_ & n243;
  assign n515 = ~n368 & ~n369;
  assign n516 = ~n391 & ~n515;
  assign n517 = n391 & n515;
  assign n518 = ~n516 & ~n517;
  assign n519 = n409 & ~n518;
  assign n520 = ~n514 & ~n519;
  assign n521 = CONT1_REG_4_ & ~n217;
  assign n522 = ~n218 & ~n521;
  assign n523 = n244 & ~n522;
  assign n524 = R_IN_REG_4_ & n446;
  assign n525 = ~n315 & ~n316;
  assign n526 = n344 & n525;
  assign n527 = ~n344 & ~n525;
  assign n528 = ~n526 & ~n527;
  assign n529 = n297 & ~n528;
  assign n530 = ~n523 & ~n524;
  assign n531 = ~n529 & n530;
  assign n532 = ~STATO_REG_0_ & ~n531;
  assign n533 = ~n505 & ~n506;
  assign n534 = ~n513 & n533;
  assign n535 = n520 & n534;
  assign n108 = n532 | ~n535;
  assign n537 = CONT_REG_2_ & n448;
  assign n538 = CONT_REG_3_ & n472;
  assign n539 = ~n260 & ~n261;
  assign n540 = ~n276 & ~n539;
  assign n541 = n276 & n539;
  assign n542 = ~n540 & ~n541;
  assign n543 = n298 & ~n542;
  assign n544 = CONT1_REG_3_ & n243;
  assign n545 = ~CONT1_REG_3_ & ~n372;
  assign n546 = CONT1_REG_3_ & n372;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n389 & ~n547;
  assign n549 = n389 & n547;
  assign n550 = ~n548 & ~n549;
  assign n551 = n409 & n550;
  assign n552 = ~n544 & ~n551;
  assign n553 = CONT1_REG_3_ & n216;
  assign n554 = ~n217 & ~n553;
  assign n555 = n244 & ~n554;
  assign n556 = R_IN_REG_3_ & n446;
  assign n557 = ~n320 & ~n321;
  assign n558 = n342 & n557;
  assign n559 = ~n342 & ~n557;
  assign n560 = ~n558 & ~n559;
  assign n561 = n297 & ~n560;
  assign n562 = ~n555 & ~n556;
  assign n563 = ~n561 & n562;
  assign n564 = ~STATO_REG_0_ & ~n563;
  assign n565 = ~n537 & ~n538;
  assign n566 = ~n543 & n565;
  assign n567 = n552 & n566;
  assign n113 = n564 | ~n567;
  assign n569 = CONT_REG_1_ & n448;
  assign n570 = CONT_REG_2_ & n472;
  assign n571 = n271 & ~n273;
  assign n572 = ~n271 & n273;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n270 & ~n573;
  assign n575 = n270 & n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = n298 & ~n576;
  assign n578 = CONT1_REG_2_ & n243;
  assign n579 = ~n378 & ~n379;
  assign n580 = ~n387 & ~n579;
  assign n581 = n387 & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = n409 & ~n582;
  assign n584 = ~n578 & ~n583;
  assign n585 = CONT1_REG_2_ & ~CONT1_REG_1_;
  assign n586 = ~CONT1_REG_2_ & CONT1_REG_1_;
  assign n587 = ~n585 & ~n586;
  assign n588 = n244 & ~n587;
  assign n589 = R_IN_REG_2_ & n446;
  assign n590 = ~n325 & ~n326;
  assign n591 = n340 & n590;
  assign n592 = ~n340 & ~n590;
  assign n593 = ~n591 & ~n592;
  assign n594 = n297 & ~n593;
  assign n595 = ~n588 & ~n589;
  assign n596 = ~n594 & n595;
  assign n597 = ~STATO_REG_0_ & ~n596;
  assign n598 = ~n569 & ~n570;
  assign n599 = ~n577 & n598;
  assign n600 = n584 & n599;
  assign n118 = n597 | ~n600;
  assign n602 = CONT_REG_0_ & n448;
  assign n603 = CONT_REG_1_ & n472;
  assign n604 = ~n264 & ~n265;
  assign n605 = ~n268 & ~n604;
  assign n606 = n268 & n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = n298 & ~n607;
  assign n609 = CONT1_REG_1_ & n243;
  assign n610 = ~CONT1_REG_1_ & ~n367;
  assign n611 = CONT1_REG_1_ & n367;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n383 & ~n612;
  assign n614 = n383 & n612;
  assign n615 = ~n613 & ~n614;
  assign n616 = n409 & n615;
  assign n617 = ~n609 & ~n616;
  assign n618 = ~n330 & ~n331;
  assign n619 = n338 & n618;
  assign n620 = ~n338 & ~n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = n297 & ~n621;
  assign n623 = R_IN_REG_1_ & n446;
  assign n624 = ~CONT1_REG_1_ & n244;
  assign n625 = ~n622 & ~n623;
  assign n626 = ~n624 & n625;
  assign n627 = ~STATO_REG_0_ & ~n626;
  assign n628 = ~n602 & ~n603;
  assign n629 = ~n608 & n628;
  assign n630 = n617 & n629;
  assign n123 = n627 | ~n630;
  assign n632 = ~n266 & n267;
  assign n633 = ~n268 & ~n632;
  assign n634 = n298 & ~n633;
  assign n635 = R_IN_REG_3_ & CONT1_REG_0_;
  assign n636 = ~R_IN_REG_3_ & ~CONT1_REG_0_;
  assign n637 = ~n635 & ~n636;
  assign n638 = n372 & ~n637;
  assign n639 = ~n372 & n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = n409 & n640;
  assign n642 = CONT_REG_0_ & n472;
  assign n643 = CONT1_REG_0_ & n243;
  assign n644 = ~n335 & ~n336;
  assign n645 = R_IN_REG_1_ & n644;
  assign n646 = ~R_IN_REG_1_ & ~n644;
  assign n647 = ~n645 & ~n646;
  assign n648 = n297 & ~n647;
  assign n649 = R_IN_REG_0_ & n446;
  assign n650 = CONT1_REG_0_ & n244;
  assign n651 = ~n648 & ~n649;
  assign n652 = ~n650 & n651;
  assign n653 = ~STATO_REG_0_ & ~n652;
  assign n654 = ~n634 & ~n641;
  assign n655 = ~n642 & n654;
  assign n656 = ~n643 & n655;
  assign n128 = n653 | ~n656;
  assign n658 = X_OUT_REG_5_ & ~n141_1;
  assign n659 = ~CONT1_REG_8_ & n141_1;
  assign n660 = n247 & n659;
  assign n661 = STATO_REG_3_ & n141_1;
  assign n662 = CONT1_REG_8_ & n661;
  assign n663 = ~n477 & n662;
  assign n664 = ~n658 & ~n660;
  assign n133 = n663 | ~n664;
  assign n666 = X_OUT_REG_4_ & ~n141_1;
  assign n667 = ~CONT1_REG_8_ & n661;
  assign n668 = CONT1_REG_4_ & n667;
  assign n669 = ~n512 & n662;
  assign n670 = ~n666 & ~n668;
  assign n137 = n669 | ~n670;
  assign n672 = X_OUT_REG_3_ & ~n141_1;
  assign n673 = CONT1_REG_3_ & n667;
  assign n674 = ~n542 & n662;
  assign n675 = ~n672 & ~n673;
  assign n141 = n674 | ~n675;
  assign n677 = X_OUT_REG_2_ & ~n141_1;
  assign n678 = n271 & n659;
  assign n679 = ~n576 & n662;
  assign n680 = ~n677 & ~n678;
  assign n145 = n679 | ~n680;
  assign n682 = X_OUT_REG_1_ & ~n141_1;
  assign n683 = CONT1_REG_1_ & n667;
  assign n684 = ~n607 & n662;
  assign n685 = ~n682 & ~n683;
  assign n149 = n684 | ~n685;
  assign n687 = X_OUT_REG_0_ & ~n141_1;
  assign n688 = n266 & n659;
  assign n689 = ~n633 & n662;
  assign n690 = ~n687 & ~n688;
  assign n153 = n689 | ~n690;
  assign n692 = STATO_REG_0_ & n225;
  assign n157 = n140 | n692;
  assign n694 = STATO_REG_0_ & n127;
  assign n695 = STATO_REG_2_ & ~n226;
  assign n162 = n694 | n695;
  assign n697 = R_IN_REG_1_ & ~STATO_REG_1_;
  assign n698 = ~STATO_REG_0_ & n697;
  assign n699 = ~STATO_REG_1_ & ~n238;
  assign n700 = STATO_REG_0_ & ~n699;
  assign n701 = ~n698 & ~n700;
  assign n702 = STATO_REG_2_ & n701;
  assign n703 = ~STBI & STATO_REG_0_;
  assign n704 = n107 & n703;
  assign n705 = n128_1 & ~n139;
  assign n706 = ~n184 & n705;
  assign n707 = ~n702 & ~n704;
  assign n167 = n706 | ~n707;
  assign n709 = ~STBI & ~STATO_REG_2_;
  assign n710 = ~R_IN_REG_1_ & ~STATO_REG_0_;
  assign n711 = ~STATO_REG_1_ & ~n709;
  assign n712 = ~n710 & n711;
  assign n713 = ~STATO_REG_0_ & n225;
  assign n714 = ~n229 & n713;
  assign n715 = ~n705 & ~n712;
  assign n716 = ~n714 & n715;
  assign n172 = n141_1 | ~n716;
  always @ (posedge clock) begin
    R_IN_REG_5_ <= n28;
    R_IN_REG_4_ <= n33;
    R_IN_REG_3_ <= n38;
    R_IN_REG_2_ <= n43;
    R_IN_REG_1_ <= n48;
    R_IN_REG_0_ <= n53;
    CONT_REG_5_ <= n58;
    CONT_REG_4_ <= n63;
    CONT_REG_3_ <= n68;
    CONT_REG_2_ <= n73;
    CONT_REG_1_ <= n78;
    CONT_REG_0_ <= n83;
    CONT1_REG_8_ <= n88;
    CONT1_REG_7_ <= n93;
    CONT1_REG_6_ <= n98;
    CONT1_REG_5_ <= n103;
    CONT1_REG_4_ <= n108;
    CONT1_REG_3_ <= n113;
    CONT1_REG_2_ <= n118;
    CONT1_REG_1_ <= n123;
    CONT1_REG_0_ <= n128;
    X_OUT_REG_5_ <= n133;
    X_OUT_REG_4_ <= n137;
    X_OUT_REG_3_ <= n141;
    X_OUT_REG_2_ <= n145;
    X_OUT_REG_1_ <= n149;
    X_OUT_REG_0_ <= n153;
    STATO_REG_3_ <= n157;
    STATO_REG_2_ <= n162;
    STATO_REG_1_ <= n167;
    STATO_REG_0_ <= n172;
  end
endmodule


