// Benchmark "top" written by ABC on Mon Nov 27 16:51:57 2023

module top ( 
    \1 , \5 , \9 , \12 , \15 , \18 , \23 , \26 , \29 , \32 , \35 , \38 ,
    \41 , \44 , \47 , \50 , \53 , \54 , \55 , \56 , \57 , \58 , \59 , \60 ,
    \61 , \62 , \63 , \64 , \65 , \66 , \69 , \70 , \73 , \74 , \75 , \76 ,
    \77 , \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86 , \87 , \88 ,
    \89 , \94 , \97 , \100 , \103 , \106 , \109 , \110 , \111 , \112 ,
    \113 , \114 , \115 , \118 , \121 , \124 , \127 , \130 , \133 , \134 ,
    \135 , \138 , \141 , \144 , \147 , \150 , \151 , \152 , \153 , \154 ,
    \155 , \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 , \164 ,
    \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 , \174 ,
    \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 , \184 ,
    \185 , \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 , \194 ,
    \195 , \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 , \204 ,
    \205 , \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 , \214 ,
    \215 , \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 , \224 ,
    \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 , \234 ,
    \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \245 , \248 ,
    \251 , \254 , \257 , \260 , \263 , \267 , \271 , \274 , \277 , \280 ,
    \283 , \286 , \289 , \293 , \296 , \299 , \303 , \307 , \310 , \313 ,
    \316 , \319 , \322 , \325 , \328 , \331 , \334 , \337 , \340 , \343 ,
    \346 , \349 , \352 , \355 , \358 , \361 , \364 , \367 , \382 ,
    \387 , \388 , \478 , \482 , \484 , \486 , \489 , \492 , \501 , \505 ,
    \507 , \509 , \511 , \513 , \515 , \517 , \519 , \535 , \537 , \539 ,
    \541 , \543 , \545 , \547 , \549 , \551 , \553 , \556 , \559 , \561 ,
    \563 , \565 , \567 , \569 , \571 , \573 , \582 , \643 , \707 , \813 ,
    \881 , \882 , \883 , \884 , \885 , \889 , \945 , \1110 , \1111 ,
    \1112 , \1113 , \1114 , \1489 , \1490 , \1781 , \10025 , \10101 ,
    \10102 , \10103 , \10104 , \10109 , \10110 , \10111 , \10112 , \10350 ,
    \10351 , \10352 , \10353 , \10574 , \10575 , \10576 , \10628 , \10632 ,
    \10641 , \10704 , \10706 , \10711 , \10712 , \10713 , \10714 , \10715 ,
    \10716 , \10717 , \10718 , \10729 , \10759 , \10760 , \10761 , \10762 ,
    \10763 , \10827 , \10837 , \10838 , \10839 , \10840 , \10868 , \10869 ,
    \10870 , \10871 , \10905 , \10906 , \10907 , \10908 , \11333 , \11334 ,
    \11340 , \11342   );
  input  \1 , \5 , \9 , \12 , \15 , \18 , \23 , \26 , \29 , \32 , \35 ,
    \38 , \41 , \44 , \47 , \50 , \53 , \54 , \55 , \56 , \57 , \58 , \59 ,
    \60 , \61 , \62 , \63 , \64 , \65 , \66 , \69 , \70 , \73 , \74 , \75 ,
    \76 , \77 , \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86 , \87 ,
    \88 , \89 , \94 , \97 , \100 , \103 , \106 , \109 , \110 , \111 ,
    \112 , \113 , \114 , \115 , \118 , \121 , \124 , \127 , \130 , \133 ,
    \134 , \135 , \138 , \141 , \144 , \147 , \150 , \151 , \152 , \153 ,
    \154 , \155 , \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 ,
    \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 ,
    \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 ,
    \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 ,
    \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 ,
    \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 ,
    \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 ,
    \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ,
    \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \245 ,
    \248 , \251 , \254 , \257 , \260 , \263 , \267 , \271 , \274 , \277 ,
    \280 , \283 , \286 , \289 , \293 , \296 , \299 , \303 , \307 , \310 ,
    \313 , \316 , \319 , \322 , \325 , \328 , \331 , \334 , \337 , \340 ,
    \343 , \346 , \349 , \352 , \355 , \358 , \361 , \364 , \367 , \382 ;
  output \387 , \388 , \478 , \482 , \484 , \486 , \489 , \492 , \501 , \505 ,
    \507 , \509 , \511 , \513 , \515 , \517 , \519 , \535 , \537 , \539 ,
    \541 , \543 , \545 , \547 , \549 , \551 , \553 , \556 , \559 , \561 ,
    \563 , \565 , \567 , \569 , \571 , \573 , \582 , \643 , \707 , \813 ,
    \881 , \882 , \883 , \884 , \885 , \889 , \945 , \1110 , \1111 ,
    \1112 , \1113 , \1114 , \1489 , \1490 , \1781 , \10025 , \10101 ,
    \10102 , \10103 , \10104 , \10109 , \10110 , \10111 , \10112 , \10350 ,
    \10351 , \10352 , \10353 , \10574 , \10575 , \10576 , \10628 , \10632 ,
    \10641 , \10704 , \10706 , \10711 , \10712 , \10713 , \10714 , \10715 ,
    \10716 , \10717 , \10718 , \10729 , \10759 , \10760 , \10761 , \10762 ,
    \10763 , \10827 , \10837 , \10838 , \10839 , \10840 , \10868 , \10869 ,
    \10870 , \10871 , \10905 , \10906 , \10907 , \10908 , \11333 , \11334 ,
    \11340 , \11342 ;
  wire new_n316, new_n317, new_n319, new_n320, new_n322, new_n323, new_n325,
    new_n326, new_n329, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n917, new_n919, new_n921, new_n923, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1408, new_n1409,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1422, new_n1423, new_n1424, new_n1425, new_n1426, new_n1427,
    new_n1428, new_n1429, new_n1430, new_n1431, new_n1432, new_n1433,
    new_n1434, new_n1436, new_n1437, new_n1438, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1445, new_n1446, new_n1447, new_n1449,
    new_n1451, new_n1452, new_n1453, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1460, new_n1462, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1470, new_n1471, new_n1472, new_n1474,
    new_n1475, new_n1476, new_n1477, new_n1478, new_n1480, new_n1482,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1489, new_n1490,
    new_n1492, new_n1494, new_n1495, new_n1496, new_n1497, new_n1498,
    new_n1499, new_n1500, new_n1501, new_n1502, new_n1503, new_n1504,
    new_n1505, new_n1507, new_n1508, new_n1510, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1523, new_n1525, new_n1526, new_n1527, new_n1529,
    new_n1530, new_n1531, new_n1533, new_n1535, new_n1536, new_n1537,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1657, new_n1658, new_n1659, new_n1660,
    new_n1661, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1677, new_n1678,
    new_n1679, new_n1680, new_n1681, new_n1682, new_n1683, new_n1684,
    new_n1685, new_n1686, new_n1687, new_n1688, new_n1689, new_n1690,
    new_n1691, new_n1692, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1698, new_n1699, new_n1700, new_n1701, new_n1702,
    new_n1703, new_n1704, new_n1705, new_n1706, new_n1707, new_n1708,
    new_n1709, new_n1710, new_n1711, new_n1712, new_n1713, new_n1714,
    new_n1715, new_n1716, new_n1717, new_n1718, new_n1719, new_n1720,
    new_n1721, new_n1723, new_n1724, new_n1725, new_n1726, new_n1727,
    new_n1728, new_n1729, new_n1730, new_n1731, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1737, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799;
  assign \881  = \5  | \57 ;
  assign new_n316 = \150  & \184 ;
  assign new_n317 = \228  & \240 ;
  assign \882  = ~new_n316 | ~new_n317;
  assign new_n319 = \152  & \210 ;
  assign new_n320 = \218  & \230 ;
  assign \883  = ~new_n319 | ~new_n320;
  assign new_n322 = \182  & \183 ;
  assign new_n323 = \185  & \186 ;
  assign \884  = ~new_n322 | ~new_n323;
  assign new_n325 = \162  & \172 ;
  assign new_n326 = \188  & \199 ;
  assign \885  = ~new_n325 | ~new_n326;
  assign \1110  = \5  | ~\242 ;
  assign new_n329 = ~\5  & \133 ;
  assign \1113  = ~\134  | ~new_n329;
  assign \1781  = \1  & \163 ;
  assign new_n332 = ~\18  & ~\41 ;
  assign new_n333 = \310  & new_n332;
  assign new_n334 = ~\18  & \41 ;
  assign new_n335 = ~\310  & new_n334;
  assign new_n336 = ~new_n333 & ~new_n335;
  assign new_n337 = ~\367  & ~new_n336;
  assign new_n338 = \367  & new_n336;
  assign \10025  = ~new_n337 & ~new_n338;
  assign new_n340 = ~\263  & ~\267 ;
  assign new_n341 = \382  & ~new_n340;
  assign new_n342 = ~\38  & new_n341;
  assign new_n343 = \9  & \12 ;
  assign new_n344 = ~\18  & ~new_n343;
  assign new_n345 = \213  & ~new_n343;
  assign new_n346 = ~new_n344 & ~new_n345;
  assign new_n347 = ~\260  & ~new_n346;
  assign new_n348 = \260  & new_n346;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = \214  & ~new_n343;
  assign new_n351 = ~new_n344 & ~new_n350;
  assign new_n352 = ~\257  & ~new_n351;
  assign new_n353 = \257  & new_n351;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = \215  & ~new_n343;
  assign new_n356 = ~new_n344 & ~new_n355;
  assign new_n357 = \106  & new_n356;
  assign new_n358 = ~\106  & ~new_n356;
  assign new_n359 = \216  & ~new_n343;
  assign new_n360 = ~new_n344 & ~new_n359;
  assign new_n361 = \254  & new_n360;
  assign new_n362 = ~\254  & ~new_n360;
  assign new_n363 = \209  & ~new_n343;
  assign new_n364 = ~new_n344 & ~new_n363;
  assign new_n365 = ~\251  & ~new_n364;
  assign new_n366 = ~new_n362 & ~new_n365;
  assign new_n367 = ~new_n361 & ~new_n366;
  assign new_n368 = ~new_n358 & ~new_n367;
  assign new_n369 = ~new_n357 & ~new_n368;
  assign new_n370 = \18  & ~new_n343;
  assign new_n371 = ~\209  & ~\216 ;
  assign new_n372 = \209  & \216 ;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = new_n370 & new_n373;
  assign new_n375 = \251  & \254 ;
  assign new_n376 = ~\251  & ~\254 ;
  assign new_n377 = ~new_n375 & ~new_n376;
  assign new_n378 = ~new_n374 & new_n377;
  assign new_n379 = new_n374 & ~new_n377;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = ~new_n361 & ~new_n362;
  assign new_n382 = new_n380 & new_n381;
  assign new_n383 = ~new_n357 & new_n382;
  assign new_n384 = \153  & ~new_n343;
  assign new_n385 = ~new_n344 & ~new_n384;
  assign new_n386 = \303  & new_n385;
  assign new_n387 = \154  & ~new_n343;
  assign new_n388 = ~new_n344 & ~new_n387;
  assign new_n389 = \299  & new_n388;
  assign new_n390 = ~\299  & ~new_n388;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = \155  & ~new_n343;
  assign new_n393 = ~new_n344 & ~new_n392;
  assign new_n394 = ~\296  & ~new_n393;
  assign new_n395 = \18  & ~\156 ;
  assign new_n396 = ~new_n343 & ~new_n395;
  assign new_n397 = \293  & ~new_n396;
  assign new_n398 = \296  & new_n393;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = ~new_n394 & ~new_n399;
  assign new_n401 = \157  & ~new_n343;
  assign new_n402 = ~new_n344 & ~new_n401;
  assign new_n403 = ~\289  & ~new_n402;
  assign new_n404 = \289  & new_n402;
  assign new_n405 = ~\18  & \135 ;
  assign new_n406 = \18  & \158 ;
  assign new_n407 = ~new_n405 & ~new_n406;
  assign new_n408 = ~\286  & ~new_n407;
  assign new_n409 = \286  & new_n407;
  assign new_n410 = ~new_n408 & ~new_n409;
  assign new_n411 = ~\18  & \144 ;
  assign new_n412 = \18  & \159 ;
  assign new_n413 = ~new_n411 & ~new_n412;
  assign new_n414 = ~\283  & ~new_n413;
  assign new_n415 = \283  & new_n413;
  assign new_n416 = ~\18  & ~\138 ;
  assign new_n417 = \18  & ~\160 ;
  assign new_n418 = ~new_n416 & ~new_n417;
  assign new_n419 = ~\280  & new_n418;
  assign new_n420 = \280  & ~new_n418;
  assign new_n421 = ~new_n419 & ~new_n420;
  assign new_n422 = ~\18  & \147 ;
  assign new_n423 = \18  & \151 ;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = \277  & new_n424;
  assign new_n426 = new_n421 & ~new_n425;
  assign new_n427 = ~\18  & ~\66 ;
  assign new_n428 = \18  & ~\219 ;
  assign new_n429 = ~new_n427 & ~new_n428;
  assign new_n430 = \364  & ~new_n429;
  assign new_n431 = ~\364  & new_n429;
  assign new_n432 = ~\18  & \50 ;
  assign new_n433 = \18  & \220 ;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign new_n435 = ~\361  & ~new_n434;
  assign new_n436 = \361  & new_n434;
  assign new_n437 = ~\18  & \32 ;
  assign new_n438 = \18  & \221 ;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = \358  & new_n439;
  assign new_n441 = ~\358  & ~new_n439;
  assign new_n442 = ~new_n440 & ~new_n441;
  assign new_n443 = ~\18  & \35 ;
  assign new_n444 = \18  & \222 ;
  assign new_n445 = ~new_n443 & ~new_n444;
  assign new_n446 = ~\355  & ~new_n445;
  assign new_n447 = \355  & new_n445;
  assign new_n448 = ~\18  & ~\47 ;
  assign new_n449 = \18  & ~\223 ;
  assign new_n450 = ~new_n448 & ~new_n449;
  assign new_n451 = ~\352  & new_n450;
  assign new_n452 = \352  & ~new_n450;
  assign new_n453 = ~new_n451 & ~new_n452;
  assign new_n454 = ~\18  & \118 ;
  assign new_n455 = \18  & \217 ;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457 = ~\340  & ~new_n456;
  assign new_n458 = \340  & new_n456;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = ~\18  & \100 ;
  assign new_n461 = \18  & \231 ;
  assign new_n462 = ~new_n460 & ~new_n461;
  assign new_n463 = ~\334  & ~new_n462;
  assign new_n464 = \334  & new_n462;
  assign new_n465 = ~new_n463 & ~new_n464;
  assign new_n466 = ~\18  & \124 ;
  assign new_n467 = \18  & \232 ;
  assign new_n468 = ~new_n466 & ~new_n467;
  assign new_n469 = ~\331  & ~new_n468;
  assign new_n470 = ~\18  & \127 ;
  assign new_n471 = \18  & \233 ;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = ~\328  & ~new_n472;
  assign new_n474 = \328  & new_n472;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = ~\18  & \130 ;
  assign new_n477 = \18  & \234 ;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = ~\325  & ~new_n478;
  assign new_n480 = new_n475 & ~new_n479;
  assign new_n481 = ~\18  & \103 ;
  assign new_n482 = \18  & \235 ;
  assign new_n483 = ~new_n481 & ~new_n482;
  assign new_n484 = ~\322  & ~new_n483;
  assign new_n485 = ~\18  & \23 ;
  assign new_n486 = \18  & \236 ;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = ~\319  & ~new_n487;
  assign new_n489 = ~\18  & ~\29 ;
  assign new_n490 = \18  & ~\238 ;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = ~\313  & new_n491;
  assign new_n493 = \313  & ~new_n491;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = ~new_n335 & ~new_n338;
  assign new_n496 = new_n494 & ~new_n495;
  assign new_n497 = ~new_n492 & ~new_n496;
  assign new_n498 = ~\18  & \26 ;
  assign new_n499 = \18  & \237 ;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = \316  & new_n500;
  assign new_n502 = ~\316  & ~new_n500;
  assign new_n503 = ~new_n501 & ~new_n502;
  assign new_n504 = ~new_n497 & new_n503;
  assign new_n505 = ~new_n335 & ~new_n492;
  assign new_n506 = ~new_n493 & ~new_n501;
  assign new_n507 = ~new_n505 & new_n506;
  assign new_n508 = ~new_n502 & ~new_n507;
  assign new_n509 = ~new_n504 & new_n508;
  assign new_n510 = \319  & new_n487;
  assign new_n511 = ~new_n488 & ~new_n510;
  assign new_n512 = ~new_n509 & new_n511;
  assign new_n513 = ~new_n488 & ~new_n512;
  assign new_n514 = \322  & new_n483;
  assign new_n515 = ~new_n484 & ~new_n514;
  assign new_n516 = ~new_n513 & new_n515;
  assign new_n517 = ~new_n484 & ~new_n516;
  assign new_n518 = new_n480 & new_n517;
  assign new_n519 = \325  & new_n478;
  assign new_n520 = new_n475 & new_n519;
  assign new_n521 = ~new_n474 & ~new_n520;
  assign new_n522 = ~new_n518 & new_n521;
  assign new_n523 = \331  & new_n468;
  assign new_n524 = ~new_n469 & ~new_n523;
  assign new_n525 = new_n522 & new_n524;
  assign new_n526 = ~new_n469 & ~new_n525;
  assign new_n527 = new_n465 & ~new_n526;
  assign new_n528 = ~new_n463 & ~new_n527;
  assign new_n529 = new_n459 & ~new_n528;
  assign new_n530 = ~new_n457 & ~new_n529;
  assign new_n531 = ~\18  & \121 ;
  assign new_n532 = \18  & \224 ;
  assign new_n533 = ~new_n531 & ~new_n532;
  assign new_n534 = \349  & new_n533;
  assign new_n535 = ~\349  & ~new_n533;
  assign new_n536 = ~\18  & ~\94 ;
  assign new_n537 = \18  & ~\225 ;
  assign new_n538 = ~new_n536 & ~new_n537;
  assign new_n539 = ~\346  & new_n538;
  assign new_n540 = \18  & ~\226 ;
  assign new_n541 = ~\18  & ~\97 ;
  assign new_n542 = ~new_n540 & ~new_n541;
  assign new_n543 = ~\343  & new_n542;
  assign new_n544 = new_n459 & ~new_n543;
  assign new_n545 = ~new_n539 & new_n544;
  assign new_n546 = \346  & ~new_n538;
  assign new_n547 = \343  & ~new_n542;
  assign new_n548 = ~new_n458 & ~new_n547;
  assign new_n549 = ~new_n539 & ~new_n543;
  assign new_n550 = ~new_n548 & new_n549;
  assign new_n551 = ~new_n546 & ~new_n550;
  assign new_n552 = ~new_n545 & new_n551;
  assign new_n553 = ~new_n535 & ~new_n552;
  assign new_n554 = ~new_n534 & ~new_n553;
  assign new_n555 = new_n530 & ~new_n554;
  assign new_n556 = ~new_n539 & ~new_n546;
  assign new_n557 = ~new_n543 & ~new_n547;
  assign new_n558 = new_n556 & new_n557;
  assign new_n559 = new_n553 & ~new_n558;
  assign new_n560 = ~new_n534 & ~new_n559;
  assign new_n561 = ~new_n555 & new_n560;
  assign new_n562 = new_n453 & new_n561;
  assign new_n563 = ~new_n451 & ~new_n562;
  assign new_n564 = ~new_n447 & ~new_n563;
  assign new_n565 = ~new_n446 & ~new_n564;
  assign new_n566 = new_n442 & new_n565;
  assign new_n567 = ~new_n440 & ~new_n566;
  assign new_n568 = ~new_n436 & new_n567;
  assign new_n569 = ~new_n435 & ~new_n568;
  assign new_n570 = ~new_n431 & new_n569;
  assign new_n571 = ~new_n430 & ~new_n570;
  assign new_n572 = new_n426 & new_n571;
  assign new_n573 = ~\277  & ~new_n424;
  assign new_n574 = ~new_n419 & ~new_n573;
  assign new_n575 = ~new_n420 & ~new_n574;
  assign new_n576 = ~new_n572 & ~new_n575;
  assign new_n577 = ~new_n415 & ~new_n576;
  assign new_n578 = ~new_n414 & ~new_n577;
  assign new_n579 = new_n410 & ~new_n578;
  assign new_n580 = ~new_n408 & ~new_n579;
  assign new_n581 = ~new_n404 & ~new_n580;
  assign new_n582 = ~new_n403 & ~new_n581;
  assign new_n583 = ~new_n397 & ~new_n582;
  assign new_n584 = ~new_n394 & ~new_n398;
  assign new_n585 = ~\293  & new_n396;
  assign new_n586 = new_n584 & ~new_n585;
  assign new_n587 = ~new_n583 & new_n586;
  assign new_n588 = ~new_n400 & ~new_n587;
  assign new_n589 = new_n391 & ~new_n588;
  assign new_n590 = ~new_n389 & ~new_n589;
  assign new_n591 = ~\303  & ~new_n385;
  assign new_n592 = ~new_n386 & ~new_n591;
  assign new_n593 = ~new_n590 & new_n592;
  assign new_n594 = ~new_n386 & ~new_n593;
  assign new_n595 = new_n383 & new_n594;
  assign new_n596 = ~new_n369 & ~new_n595;
  assign new_n597 = new_n354 & ~new_n596;
  assign new_n598 = ~new_n352 & ~new_n597;
  assign new_n599 = new_n349 & ~new_n598;
  assign new_n600 = ~new_n347 & ~new_n599;
  assign new_n601 = \263  & \382 ;
  assign new_n602 = \267  & new_n601;
  assign new_n603 = \38  & ~new_n602;
  assign new_n604 = new_n600 & ~new_n603;
  assign \10101  = ~new_n342 & ~new_n604;
  assign new_n606 = \85  & new_n405;
  assign new_n607 = ~\179  & \283 ;
  assign new_n608 = ~\178  & \286 ;
  assign new_n609 = ~new_n607 & ~new_n608;
  assign new_n610 = \18  & ~new_n609;
  assign new_n611 = ~\85  & ~\135 ;
  assign new_n612 = ~\84  & ~\144 ;
  assign new_n613 = ~new_n611 & ~new_n612;
  assign new_n614 = ~\18  & ~new_n613;
  assign new_n615 = \84  & new_n411;
  assign new_n616 = ~\83  & new_n416;
  assign new_n617 = \65  & new_n422;
  assign new_n618 = ~\18  & ~\65 ;
  assign new_n619 = ~\147  & new_n618;
  assign new_n620 = \18  & ~\171 ;
  assign new_n621 = \277  & new_n620;
  assign new_n622 = ~\62  & new_n427;
  assign new_n623 = \61  & new_n432;
  assign new_n624 = ~\190  & \361 ;
  assign new_n625 = ~\191  & \358 ;
  assign new_n626 = ~new_n624 & ~new_n625;
  assign new_n627 = \18  & ~new_n626;
  assign new_n628 = ~\50  & ~\61 ;
  assign new_n629 = ~\32  & ~\60 ;
  assign new_n630 = ~new_n628 & ~new_n629;
  assign new_n631 = ~\18  & ~new_n630;
  assign new_n632 = \79  & new_n443;
  assign new_n633 = ~\18  & ~\35 ;
  assign new_n634 = ~\79  & new_n633;
  assign new_n635 = \18  & ~\192 ;
  assign new_n636 = \355  & new_n635;
  assign new_n637 = \77  & new_n454;
  assign new_n638 = \18  & \200 ;
  assign new_n639 = ~new_n460 & ~new_n638;
  assign new_n640 = \18  & ~\334 ;
  assign new_n641 = ~\18  & \56 ;
  assign new_n642 = ~new_n640 & ~new_n641;
  assign new_n643 = new_n639 & new_n642;
  assign new_n644 = \55  & new_n466;
  assign new_n645 = ~\201  & \331 ;
  assign new_n646 = ~\202  & \328 ;
  assign new_n647 = ~new_n645 & ~new_n646;
  assign new_n648 = \18  & ~new_n647;
  assign new_n649 = ~\54  & ~\127 ;
  assign new_n650 = ~\55  & ~\124 ;
  assign new_n651 = ~new_n649 & ~new_n650;
  assign new_n652 = ~\18  & ~new_n651;
  assign new_n653 = \53  & new_n476;
  assign new_n654 = \202  & ~\328 ;
  assign new_n655 = \203  & ~\325 ;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = \18  & ~new_n656;
  assign new_n658 = \54  & new_n470;
  assign new_n659 = ~\18  & ~\130 ;
  assign new_n660 = ~\53  & new_n659;
  assign new_n661 = \18  & ~\203 ;
  assign new_n662 = \325  & new_n661;
  assign new_n663 = \18  & \204 ;
  assign new_n664 = ~new_n481 & ~new_n663;
  assign new_n665 = \18  & ~\322 ;
  assign new_n666 = ~\18  & \73 ;
  assign new_n667 = ~new_n665 & ~new_n666;
  assign new_n668 = new_n664 & new_n667;
  assign new_n669 = ~new_n664 & ~new_n667;
  assign new_n670 = \18  & \205 ;
  assign new_n671 = ~new_n485 & ~new_n670;
  assign new_n672 = \18  & ~\319 ;
  assign new_n673 = ~\18  & \75 ;
  assign new_n674 = ~new_n672 & ~new_n673;
  assign new_n675 = ~new_n671 & ~new_n674;
  assign new_n676 = \18  & \206 ;
  assign new_n677 = ~new_n498 & ~new_n676;
  assign new_n678 = \18  & ~\316 ;
  assign new_n679 = ~\18  & \76 ;
  assign new_n680 = ~new_n678 & ~new_n679;
  assign new_n681 = new_n677 & new_n680;
  assign new_n682 = new_n671 & new_n674;
  assign new_n683 = ~new_n677 & ~new_n680;
  assign new_n684 = ~\18  & \29 ;
  assign new_n685 = ~\70  & new_n332;
  assign new_n686 = \89  & ~new_n685;
  assign new_n687 = \70  & new_n334;
  assign new_n688 = ~new_n686 & ~new_n687;
  assign new_n689 = \18  & ~\207 ;
  assign new_n690 = \313  & new_n689;
  assign new_n691 = ~new_n688 & ~new_n690;
  assign new_n692 = ~new_n684 & ~new_n691;
  assign new_n693 = \74  & ~new_n692;
  assign new_n694 = ~new_n489 & new_n691;
  assign new_n695 = \18  & \207 ;
  assign new_n696 = ~\313  & new_n695;
  assign new_n697 = ~new_n683 & ~new_n696;
  assign new_n698 = ~new_n694 & new_n697;
  assign new_n699 = ~new_n693 & new_n698;
  assign new_n700 = ~new_n681 & ~new_n682;
  assign new_n701 = ~new_n699 & new_n700;
  assign new_n702 = ~new_n669 & ~new_n675;
  assign new_n703 = ~new_n701 & new_n702;
  assign new_n704 = ~new_n660 & ~new_n662;
  assign new_n705 = ~new_n668 & new_n704;
  assign new_n706 = ~new_n703 & new_n705;
  assign new_n707 = ~new_n653 & ~new_n658;
  assign new_n708 = ~new_n657 & new_n707;
  assign new_n709 = ~new_n706 & new_n708;
  assign new_n710 = ~new_n648 & ~new_n652;
  assign new_n711 = ~new_n709 & new_n710;
  assign new_n712 = ~new_n639 & ~new_n642;
  assign new_n713 = \18  & \201 ;
  assign new_n714 = ~\331  & new_n713;
  assign new_n715 = ~new_n644 & ~new_n714;
  assign new_n716 = ~new_n712 & new_n715;
  assign new_n717 = ~new_n711 & new_n716;
  assign new_n718 = ~new_n643 & ~new_n717;
  assign new_n719 = \18  & \187 ;
  assign new_n720 = ~\340  & new_n719;
  assign new_n721 = ~new_n637 & ~new_n720;
  assign new_n722 = ~new_n718 & new_n721;
  assign new_n723 = ~\194  & \349 ;
  assign new_n724 = ~\195  & \346 ;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = \18  & ~new_n725;
  assign new_n727 = ~\81  & ~\121 ;
  assign new_n728 = ~\59  & ~\94 ;
  assign new_n729 = ~new_n727 & ~new_n728;
  assign new_n730 = ~\18  & ~new_n729;
  assign new_n731 = ~new_n726 & ~new_n730;
  assign new_n732 = ~\77  & ~\118 ;
  assign new_n733 = ~\78  & ~\97 ;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = ~\18  & ~new_n734;
  assign new_n736 = ~\196  & \343 ;
  assign new_n737 = ~\187  & \340 ;
  assign new_n738 = ~new_n736 & ~new_n737;
  assign new_n739 = \18  & ~new_n738;
  assign new_n740 = ~\80  & new_n448;
  assign new_n741 = \18  & ~\193 ;
  assign new_n742 = \352  & new_n741;
  assign new_n743 = ~new_n740 & ~new_n742;
  assign new_n744 = ~new_n735 & ~new_n739;
  assign new_n745 = new_n743 & new_n744;
  assign new_n746 = new_n731 & new_n745;
  assign new_n747 = ~new_n722 & new_n746;
  assign new_n748 = ~\18  & \47 ;
  assign new_n749 = \80  & new_n748;
  assign new_n750 = \18  & \194 ;
  assign new_n751 = ~\349  & new_n750;
  assign new_n752 = \81  & new_n531;
  assign new_n753 = \59  & \94 ;
  assign new_n754 = \78  & \97 ;
  assign new_n755 = ~\18  & ~new_n753;
  assign new_n756 = ~new_n754 & new_n755;
  assign new_n757 = \195  & ~\346 ;
  assign new_n758 = \196  & ~\343 ;
  assign new_n759 = \18  & ~new_n757;
  assign new_n760 = ~new_n758 & new_n759;
  assign new_n761 = ~new_n756 & ~new_n760;
  assign new_n762 = new_n731 & new_n761;
  assign new_n763 = ~new_n751 & ~new_n752;
  assign new_n764 = ~new_n762 & new_n763;
  assign new_n765 = new_n743 & ~new_n764;
  assign new_n766 = \18  & \193 ;
  assign new_n767 = ~\352  & new_n766;
  assign new_n768 = ~new_n749 & ~new_n767;
  assign new_n769 = ~new_n765 & new_n768;
  assign new_n770 = ~new_n747 & new_n769;
  assign new_n771 = ~new_n634 & ~new_n636;
  assign new_n772 = ~new_n770 & new_n771;
  assign new_n773 = \192  & ~\355 ;
  assign new_n774 = \191  & ~\358 ;
  assign new_n775 = ~new_n773 & ~new_n774;
  assign new_n776 = \18  & ~new_n775;
  assign new_n777 = \60  & new_n437;
  assign new_n778 = ~new_n632 & ~new_n777;
  assign new_n779 = ~new_n776 & new_n778;
  assign new_n780 = ~new_n772 & new_n779;
  assign new_n781 = ~new_n627 & ~new_n631;
  assign new_n782 = ~new_n780 & new_n781;
  assign new_n783 = \189  & ~\364 ;
  assign new_n784 = \190  & ~\361 ;
  assign new_n785 = ~new_n783 & ~new_n784;
  assign new_n786 = \18  & ~new_n785;
  assign new_n787 = ~\18  & \66 ;
  assign new_n788 = \62  & new_n787;
  assign new_n789 = ~new_n623 & ~new_n788;
  assign new_n790 = ~new_n786 & new_n789;
  assign new_n791 = ~new_n782 & new_n790;
  assign new_n792 = \18  & ~\189 ;
  assign new_n793 = \364  & new_n792;
  assign new_n794 = ~new_n622 & ~new_n793;
  assign \10704  = ~new_n791 & new_n794;
  assign new_n796 = ~new_n619 & ~new_n621;
  assign new_n797 = \10704  & new_n796;
  assign new_n798 = \18  & \171 ;
  assign new_n799 = ~\277  & new_n798;
  assign new_n800 = ~new_n617 & ~new_n799;
  assign new_n801 = ~new_n797 & new_n800;
  assign new_n802 = \18  & ~\180 ;
  assign new_n803 = \280  & new_n802;
  assign new_n804 = ~new_n616 & ~new_n803;
  assign new_n805 = ~new_n801 & new_n804;
  assign new_n806 = \179  & ~\283 ;
  assign new_n807 = \180  & ~\280 ;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = \18  & ~new_n808;
  assign new_n810 = ~\18  & \138 ;
  assign new_n811 = \83  & new_n810;
  assign new_n812 = ~new_n615 & ~new_n811;
  assign new_n813 = ~new_n809 & new_n812;
  assign new_n814 = ~new_n805 & new_n813;
  assign new_n815 = ~new_n610 & ~new_n614;
  assign new_n816 = ~new_n814 & new_n815;
  assign new_n817 = \178  & ~\286 ;
  assign new_n818 = \177  & ~new_n343;
  assign new_n819 = ~\289  & new_n818;
  assign new_n820 = ~new_n817 & ~new_n819;
  assign new_n821 = \18  & ~new_n820;
  assign new_n822 = \64  & new_n344;
  assign new_n823 = ~new_n606 & ~new_n822;
  assign new_n824 = ~new_n821 & new_n823;
  assign new_n825 = ~new_n816 & new_n824;
  assign new_n826 = \63  & \110 ;
  assign new_n827 = ~\18  & \64 ;
  assign new_n828 = \86  & new_n827;
  assign new_n829 = \109  & new_n826;
  assign new_n830 = new_n828 & new_n829;
  assign new_n831 = \289  & ~new_n818;
  assign new_n832 = ~\174  & \299 ;
  assign new_n833 = ~\175  & \296 ;
  assign new_n834 = ~new_n832 & ~new_n833;
  assign new_n835 = ~\173  & \303 ;
  assign new_n836 = ~\176  & \293 ;
  assign new_n837 = ~new_n343 & ~new_n836;
  assign new_n838 = ~\293  & ~\303 ;
  assign new_n839 = ~\296  & ~\299 ;
  assign new_n840 = new_n838 & new_n839;
  assign new_n841 = ~new_n837 & ~new_n840;
  assign new_n842 = \18  & ~new_n835;
  assign new_n843 = new_n834 & new_n842;
  assign new_n844 = ~new_n831 & new_n843;
  assign new_n845 = ~new_n841 & new_n844;
  assign new_n846 = ~new_n344 & ~new_n830;
  assign new_n847 = ~new_n845 & new_n846;
  assign new_n848 = ~new_n825 & ~new_n847;
  assign new_n849 = ~\63  & ~\110 ;
  assign new_n850 = ~\86  & ~\109 ;
  assign new_n851 = new_n849 & new_n850;
  assign new_n852 = new_n344 & ~new_n851;
  assign new_n853 = \173  & ~\303 ;
  assign new_n854 = \175  & ~\296 ;
  assign new_n855 = \176  & ~\293 ;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = new_n834 & ~new_n856;
  assign new_n858 = \174  & ~\299 ;
  assign new_n859 = ~new_n853 & ~new_n858;
  assign new_n860 = ~new_n857 & new_n859;
  assign new_n861 = new_n370 & ~new_n835;
  assign new_n862 = ~new_n860 & new_n861;
  assign new_n863 = ~new_n852 & ~new_n862;
  assign new_n864 = ~new_n848 & new_n863;
  assign new_n865 = \18  & ~\169 ;
  assign new_n866 = \254  & new_n865;
  assign new_n867 = ~new_n343 & ~new_n866;
  assign new_n868 = ~\106  & ~\260 ;
  assign new_n869 = \18  & new_n376;
  assign new_n870 = new_n868 & new_n869;
  assign new_n871 = \88  & \112 ;
  assign new_n872 = ~\18  & \87 ;
  assign new_n873 = \111  & new_n872;
  assign new_n874 = \113  & new_n871;
  assign new_n875 = new_n873 & new_n874;
  assign new_n876 = ~new_n867 & ~new_n870;
  assign new_n877 = ~new_n875 & new_n876;
  assign new_n878 = ~new_n864 & ~new_n877;
  assign new_n879 = ~\87  & ~\111 ;
  assign new_n880 = ~\18  & ~\113 ;
  assign new_n881 = new_n879 & new_n880;
  assign new_n882 = ~\106  & \168 ;
  assign new_n883 = \169  & ~new_n375;
  assign new_n884 = \18  & ~new_n376;
  assign new_n885 = ~new_n882 & new_n884;
  assign new_n886 = ~new_n883 & new_n885;
  assign new_n887 = ~new_n343 & ~new_n881;
  assign new_n888 = ~new_n886 & new_n887;
  assign new_n889 = ~new_n878 & ~new_n888;
  assign new_n890 = ~\166  & \260 ;
  assign new_n891 = \167  & ~new_n343;
  assign new_n892 = \257  & ~new_n891;
  assign new_n893 = \106  & ~\168 ;
  assign new_n894 = ~new_n890 & ~new_n893;
  assign new_n895 = ~new_n892 & new_n894;
  assign new_n896 = \18  & ~new_n895;
  assign new_n897 = ~new_n889 & ~new_n896;
  assign new_n898 = \166  & ~\260 ;
  assign new_n899 = \167  & ~\257 ;
  assign new_n900 = ~new_n890 & new_n899;
  assign new_n901 = ~new_n898 & ~new_n900;
  assign new_n902 = new_n370 & ~new_n901;
  assign new_n903 = ~\88  & ~\112 ;
  assign new_n904 = new_n344 & ~new_n903;
  assign new_n905 = ~\245  & ~\271 ;
  assign new_n906 = \382  & new_n905;
  assign new_n907 = \38  & ~new_n906;
  assign new_n908 = ~new_n904 & ~new_n907;
  assign new_n909 = ~new_n902 & new_n908;
  assign new_n910 = ~new_n897 & new_n909;
  assign new_n911 = \245  & \271 ;
  assign new_n912 = ~\38  & \382 ;
  assign new_n913 = ~new_n911 & new_n912;
  assign \10102  = ~new_n910 & ~new_n913;
  assign new_n915 = new_n513 & ~new_n515;
  assign \10109  = ~new_n516 & ~new_n915;
  assign new_n917 = new_n509 & ~new_n511;
  assign \10110  = ~new_n512 & ~new_n917;
  assign new_n919 = new_n497 & ~new_n503;
  assign \10111  = ~new_n504 & ~new_n919;
  assign new_n921 = ~new_n494 & new_n495;
  assign \10112  = ~new_n496 & ~new_n921;
  assign new_n923 = ~new_n465 & new_n526;
  assign \10350  = ~new_n527 & ~new_n923;
  assign new_n925 = ~new_n522 & ~new_n524;
  assign \10351  = ~new_n525 & ~new_n925;
  assign new_n927 = ~new_n475 & new_n479;
  assign new_n928 = ~new_n475 & ~new_n519;
  assign new_n929 = ~new_n517 & new_n928;
  assign new_n930 = ~new_n520 & ~new_n927;
  assign new_n931 = ~new_n518 & new_n930;
  assign \10352  = new_n929 | ~new_n931;
  assign new_n933 = ~new_n479 & ~new_n519;
  assign new_n934 = new_n517 & ~new_n933;
  assign new_n935 = ~new_n517 & new_n933;
  assign \10353  = ~new_n934 & ~new_n935;
  assign new_n937 = \29  & new_n470;
  assign new_n938 = \233  & ~\238 ;
  assign new_n939 = ~new_n471 & ~new_n490;
  assign new_n940 = ~new_n938 & ~new_n939;
  assign new_n941 = ~\127  & new_n489;
  assign new_n942 = ~new_n937 & ~new_n941;
  assign new_n943 = ~new_n940 & new_n942;
  assign new_n944 = ~\100  & new_n466;
  assign new_n945 = ~\124  & new_n460;
  assign new_n946 = ~\231  & ~\232 ;
  assign new_n947 = \231  & \232 ;
  assign new_n948 = \18  & ~new_n946;
  assign new_n949 = ~new_n947 & new_n948;
  assign new_n950 = ~new_n944 & ~new_n945;
  assign new_n951 = ~new_n949 & new_n950;
  assign new_n952 = new_n500 & ~new_n951;
  assign new_n953 = ~new_n500 & new_n951;
  assign new_n954 = ~new_n952 & ~new_n953;
  assign new_n955 = \44  & ~new_n478;
  assign new_n956 = ~\44  & new_n478;
  assign new_n957 = ~new_n955 & ~new_n956;
  assign new_n958 = new_n334 & new_n957;
  assign new_n959 = new_n332 & ~new_n957;
  assign new_n960 = ~\229  & ~\239 ;
  assign new_n961 = \229  & \239 ;
  assign new_n962 = ~new_n960 & ~new_n961;
  assign new_n963 = \234  & ~new_n962;
  assign new_n964 = ~\234  & new_n962;
  assign new_n965 = \18  & ~new_n963;
  assign new_n966 = ~new_n964 & new_n965;
  assign new_n967 = ~new_n958 & ~new_n959;
  assign new_n968 = ~new_n966 & new_n967;
  assign new_n969 = ~\23  & new_n481;
  assign new_n970 = ~\103  & new_n485;
  assign new_n971 = ~\235  & ~\236 ;
  assign new_n972 = \235  & \236 ;
  assign new_n973 = \18  & ~new_n971;
  assign new_n974 = ~new_n972 & new_n973;
  assign new_n975 = ~new_n969 & ~new_n970;
  assign new_n976 = ~new_n974 & new_n975;
  assign new_n977 = ~new_n968 & new_n976;
  assign new_n978 = new_n968 & ~new_n976;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980 = new_n954 & ~new_n979;
  assign new_n981 = ~new_n954 & new_n979;
  assign new_n982 = ~new_n980 & ~new_n981;
  assign new_n983 = new_n943 & new_n982;
  assign new_n984 = ~new_n943 & ~new_n982;
  assign new_n985 = ~\213  & ~\215 ;
  assign new_n986 = \213  & \215 ;
  assign new_n987 = ~new_n985 & ~new_n986;
  assign new_n988 = ~\212  & ~\214 ;
  assign new_n989 = \212  & \214 ;
  assign new_n990 = ~new_n988 & ~new_n989;
  assign new_n991 = \211  & ~new_n990;
  assign new_n992 = ~\211  & new_n990;
  assign new_n993 = ~new_n991 & ~new_n992;
  assign new_n994 = new_n373 & new_n993;
  assign new_n995 = ~new_n373 & ~new_n993;
  assign new_n996 = ~new_n994 & ~new_n995;
  assign new_n997 = new_n987 & new_n996;
  assign new_n998 = ~new_n987 & ~new_n996;
  assign new_n999 = new_n370 & ~new_n997;
  assign new_n1000 = ~new_n998 & new_n999;
  assign new_n1001 = \18  & ~\161 ;
  assign new_n1002 = ~\18  & ~\141 ;
  assign new_n1003 = ~new_n1001 & ~new_n1002;
  assign new_n1004 = new_n413 & ~new_n1003;
  assign new_n1005 = ~new_n413 & new_n1003;
  assign new_n1006 = ~new_n1004 & ~new_n1005;
  assign new_n1007 = \153  & ~\154 ;
  assign new_n1008 = ~\153  & \154 ;
  assign new_n1009 = ~new_n1007 & ~new_n1008;
  assign new_n1010 = new_n370 & ~new_n1009;
  assign new_n1011 = \155  & ~\157 ;
  assign new_n1012 = ~\155  & \157 ;
  assign new_n1013 = ~new_n1011 & ~new_n1012;
  assign new_n1014 = new_n396 & new_n1013;
  assign new_n1015 = new_n370 & ~new_n395;
  assign new_n1016 = ~new_n343 & ~new_n1013;
  assign new_n1017 = ~new_n1015 & new_n1016;
  assign new_n1018 = ~new_n1014 & ~new_n1017;
  assign new_n1019 = new_n1010 & ~new_n1018;
  assign new_n1020 = ~new_n1010 & new_n1018;
  assign new_n1021 = ~new_n1019 & ~new_n1020;
  assign new_n1022 = new_n1006 & new_n1021;
  assign new_n1023 = ~new_n1006 & ~new_n1021;
  assign new_n1024 = ~new_n1022 & ~new_n1023;
  assign new_n1025 = new_n407 & ~new_n424;
  assign new_n1026 = ~new_n407 & new_n424;
  assign new_n1027 = ~new_n1025 & ~new_n1026;
  assign new_n1028 = new_n418 & new_n1027;
  assign new_n1029 = ~new_n418 & ~new_n1027;
  assign new_n1030 = ~new_n1028 & ~new_n1029;
  assign new_n1031 = ~new_n1024 & ~new_n1030;
  assign new_n1032 = new_n1024 & new_n1030;
  assign new_n1033 = ~new_n1031 & ~new_n1032;
  assign new_n1034 = new_n445 & ~new_n456;
  assign new_n1035 = ~new_n445 & new_n456;
  assign new_n1036 = ~new_n1034 & ~new_n1035;
  assign new_n1037 = ~new_n429 & new_n533;
  assign new_n1038 = new_n429 & ~new_n533;
  assign new_n1039 = ~new_n1037 & ~new_n1038;
  assign new_n1040 = \220  & ~\227 ;
  assign new_n1041 = ~\220  & \227 ;
  assign new_n1042 = ~new_n1040 & ~new_n1041;
  assign new_n1043 = \18  & ~new_n1042;
  assign new_n1044 = ~\50  & ~\115 ;
  assign new_n1045 = \50  & \115 ;
  assign new_n1046 = ~\18  & ~new_n1044;
  assign new_n1047 = ~new_n1045 & new_n1046;
  assign new_n1048 = ~new_n1043 & ~new_n1047;
  assign new_n1049 = ~\32  & new_n748;
  assign new_n1050 = ~\47  & new_n437;
  assign new_n1051 = ~\221  & ~\223 ;
  assign new_n1052 = \221  & \223 ;
  assign new_n1053 = \18  & ~new_n1051;
  assign new_n1054 = ~new_n1052 & new_n1053;
  assign new_n1055 = ~new_n1049 & ~new_n1050;
  assign new_n1056 = ~new_n1054 & new_n1055;
  assign new_n1057 = new_n538 & ~new_n1056;
  assign new_n1058 = ~new_n538 & new_n1056;
  assign new_n1059 = ~new_n1057 & ~new_n1058;
  assign new_n1060 = new_n1048 & new_n1059;
  assign new_n1061 = ~new_n1048 & ~new_n1059;
  assign new_n1062 = ~new_n1060 & ~new_n1061;
  assign new_n1063 = new_n542 & ~new_n1062;
  assign new_n1064 = ~new_n542 & new_n1062;
  assign new_n1065 = ~new_n1063 & ~new_n1064;
  assign new_n1066 = new_n1039 & ~new_n1065;
  assign new_n1067 = ~new_n1039 & new_n1065;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n1036 & ~new_n1068;
  assign new_n1070 = ~new_n1036 & new_n1068;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = ~new_n1000 & ~new_n1033;
  assign new_n1073 = ~new_n983 & new_n1072;
  assign new_n1074 = ~new_n984 & new_n1073;
  assign \10574  = new_n1071 | ~new_n1074;
  assign new_n1076 = \277  & ~\299 ;
  assign new_n1077 = ~\277  & \299 ;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = \18  & ~new_n1078;
  assign new_n1080 = ~\65  & ~\109 ;
  assign new_n1081 = \65  & \109 ;
  assign new_n1082 = ~\18  & ~new_n1080;
  assign new_n1083 = ~new_n1081 & new_n1082;
  assign new_n1084 = ~new_n1079 & ~new_n1083;
  assign new_n1085 = ~\289  & ~\296 ;
  assign new_n1086 = \289  & \296 ;
  assign new_n1087 = ~new_n1085 & ~new_n1086;
  assign new_n1088 = \18  & ~new_n1087;
  assign new_n1089 = ~\18  & ~\64 ;
  assign new_n1090 = ~\86  & new_n1089;
  assign new_n1091 = ~new_n828 & ~new_n1090;
  assign new_n1092 = ~new_n1088 & new_n1091;
  assign new_n1093 = \280  & ~\286 ;
  assign new_n1094 = ~\280  & \286 ;
  assign new_n1095 = ~new_n1093 & ~new_n1094;
  assign new_n1096 = \18  & ~new_n1095;
  assign new_n1097 = ~\83  & ~\85 ;
  assign new_n1098 = \83  & \85 ;
  assign new_n1099 = ~\18  & ~new_n1097;
  assign new_n1100 = ~new_n1098 & new_n1099;
  assign new_n1101 = ~new_n1096 & ~new_n1100;
  assign new_n1102 = ~new_n1092 & new_n1101;
  assign new_n1103 = new_n1092 & ~new_n1101;
  assign new_n1104 = ~new_n1102 & ~new_n1103;
  assign new_n1105 = \274  & ~\283 ;
  assign new_n1106 = ~\274  & \283 ;
  assign new_n1107 = ~new_n1105 & ~new_n1106;
  assign new_n1108 = \18  & ~new_n1107;
  assign new_n1109 = ~\82  & ~\84 ;
  assign new_n1110 = \82  & \84 ;
  assign new_n1111 = ~\18  & ~new_n1109;
  assign new_n1112 = ~new_n1110 & new_n1111;
  assign new_n1113 = ~new_n1108 & ~new_n1112;
  assign new_n1114 = new_n1104 & ~new_n1113;
  assign new_n1115 = ~new_n1104 & new_n1113;
  assign new_n1116 = ~new_n1114 & ~new_n1115;
  assign new_n1117 = \293  & \303 ;
  assign new_n1118 = ~new_n838 & ~new_n1117;
  assign new_n1119 = \18  & ~new_n1118;
  assign new_n1120 = ~new_n826 & ~new_n849;
  assign new_n1121 = ~\18  & ~new_n1120;
  assign new_n1122 = ~new_n1119 & ~new_n1121;
  assign new_n1123 = ~new_n1116 & new_n1122;
  assign new_n1124 = new_n1116 & ~new_n1122;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = new_n1084 & ~new_n1125;
  assign new_n1127 = ~new_n1084 & new_n1125;
  assign new_n1128 = ~new_n1126 & ~new_n1127;
  assign new_n1129 = \307  & ~\313 ;
  assign new_n1130 = ~\307  & \313 ;
  assign new_n1131 = ~new_n1129 & ~new_n1130;
  assign new_n1132 = \18  & ~new_n1131;
  assign new_n1133 = ~\69  & ~\74 ;
  assign new_n1134 = \69  & \74 ;
  assign new_n1135 = ~\18  & ~new_n1133;
  assign new_n1136 = ~new_n1134 & new_n1135;
  assign new_n1137 = ~new_n1132 & ~new_n1136;
  assign new_n1138 = ~new_n667 & new_n1137;
  assign new_n1139 = new_n667 & ~new_n1137;
  assign new_n1140 = ~new_n1138 & ~new_n1139;
  assign new_n1141 = ~\310  & ~\328 ;
  assign new_n1142 = \310  & \328 ;
  assign new_n1143 = ~new_n1141 & ~new_n1142;
  assign new_n1144 = \18  & ~new_n1143;
  assign new_n1145 = ~\54  & \70 ;
  assign new_n1146 = \54  & ~\70 ;
  assign new_n1147 = ~\18  & ~new_n1145;
  assign new_n1148 = ~new_n1146 & new_n1147;
  assign new_n1149 = ~new_n1144 & ~new_n1148;
  assign new_n1150 = new_n1140 & ~new_n1149;
  assign new_n1151 = ~new_n1140 & new_n1149;
  assign new_n1152 = ~new_n1150 & ~new_n1151;
  assign new_n1153 = new_n642 & ~new_n680;
  assign new_n1154 = ~new_n642 & new_n680;
  assign new_n1155 = ~new_n1153 & ~new_n1154;
  assign new_n1156 = new_n674 & new_n1155;
  assign new_n1157 = ~new_n674 & ~new_n1155;
  assign new_n1158 = ~new_n1156 & ~new_n1157;
  assign new_n1159 = \325  & ~\331 ;
  assign new_n1160 = ~\325  & \331 ;
  assign new_n1161 = ~new_n1159 & ~new_n1160;
  assign new_n1162 = \18  & ~new_n1161;
  assign new_n1163 = ~\53  & ~\55 ;
  assign new_n1164 = \53  & \55 ;
  assign new_n1165 = ~\18  & ~new_n1163;
  assign new_n1166 = ~new_n1164 & new_n1165;
  assign new_n1167 = ~new_n1162 & ~new_n1166;
  assign new_n1168 = new_n1158 & ~new_n1167;
  assign new_n1169 = ~new_n1158 & new_n1167;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = new_n1152 & new_n1170;
  assign new_n1172 = ~new_n1152 & ~new_n1170;
  assign new_n1173 = ~\352  & ~\355 ;
  assign new_n1174 = \352  & \355 ;
  assign new_n1175 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = \18  & ~new_n1175;
  assign new_n1177 = ~\79  & \80 ;
  assign new_n1178 = \79  & ~\80 ;
  assign new_n1179 = ~\18  & ~new_n1177;
  assign new_n1180 = ~new_n1178 & new_n1179;
  assign new_n1181 = ~new_n1176 & ~new_n1180;
  assign new_n1182 = \337  & ~\361 ;
  assign new_n1183 = ~\337  & \361 ;
  assign new_n1184 = ~new_n1182 & ~new_n1183;
  assign new_n1185 = \18  & ~new_n1184;
  assign new_n1186 = ~\58  & ~\61 ;
  assign new_n1187 = \58  & \61 ;
  assign new_n1188 = ~\18  & ~new_n1186;
  assign new_n1189 = ~new_n1187 & new_n1188;
  assign new_n1190 = ~new_n1185 & ~new_n1189;
  assign new_n1191 = ~\340  & ~\358 ;
  assign new_n1192 = \340  & \358 ;
  assign new_n1193 = ~new_n1191 & ~new_n1192;
  assign new_n1194 = \18  & ~new_n1193;
  assign new_n1195 = ~\60  & \77 ;
  assign new_n1196 = \60  & ~\77 ;
  assign new_n1197 = ~\18  & ~new_n1195;
  assign new_n1198 = ~new_n1196 & new_n1197;
  assign new_n1199 = ~new_n1194 & ~new_n1198;
  assign new_n1200 = ~new_n1190 & new_n1199;
  assign new_n1201 = new_n1190 & ~new_n1199;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign new_n1203 = \343  & ~\346 ;
  assign new_n1204 = ~\343  & \346 ;
  assign new_n1205 = ~new_n1203 & ~new_n1204;
  assign new_n1206 = \18  & ~new_n1205;
  assign new_n1207 = ~\59  & ~\78 ;
  assign new_n1208 = \59  & \78 ;
  assign new_n1209 = ~\18  & ~new_n1207;
  assign new_n1210 = ~new_n1208 & new_n1209;
  assign new_n1211 = ~new_n1206 & ~new_n1210;
  assign new_n1212 = new_n1202 & ~new_n1211;
  assign new_n1213 = ~new_n1202 & new_n1211;
  assign new_n1214 = ~new_n1212 & ~new_n1213;
  assign new_n1215 = new_n1181 & new_n1214;
  assign new_n1216 = ~new_n1181 & ~new_n1214;
  assign new_n1217 = ~new_n1215 & ~new_n1216;
  assign new_n1218 = \349  & ~\364 ;
  assign new_n1219 = ~\349  & \364 ;
  assign new_n1220 = ~new_n1218 & ~new_n1219;
  assign new_n1221 = \18  & ~new_n1220;
  assign new_n1222 = ~\62  & ~\81 ;
  assign new_n1223 = \62  & \81 ;
  assign new_n1224 = ~\18  & ~new_n1222;
  assign new_n1225 = ~new_n1223 & new_n1224;
  assign new_n1226 = ~new_n1221 & ~new_n1225;
  assign new_n1227 = new_n1217 & ~new_n1226;
  assign new_n1228 = ~new_n1217 & new_n1226;
  assign new_n1229 = ~\106  & ~\254 ;
  assign new_n1230 = \106  & \254 ;
  assign new_n1231 = ~new_n1229 & ~new_n1230;
  assign new_n1232 = \18  & ~new_n1231;
  assign new_n1233 = ~\18  & new_n879;
  assign new_n1234 = ~new_n873 & ~new_n1233;
  assign new_n1235 = ~new_n1232 & new_n1234;
  assign new_n1236 = \263  & \267 ;
  assign new_n1237 = ~new_n340 & ~new_n1236;
  assign new_n1238 = ~\248  & ~\251 ;
  assign new_n1239 = \248  & \251 ;
  assign new_n1240 = ~new_n1238 & ~new_n1239;
  assign new_n1241 = ~new_n1237 & ~new_n1240;
  assign new_n1242 = new_n1237 & new_n1240;
  assign new_n1243 = ~new_n1241 & ~new_n1242;
  assign new_n1244 = \18  & ~new_n1243;
  assign new_n1245 = ~new_n905 & ~new_n911;
  assign new_n1246 = ~\113  & ~\114 ;
  assign new_n1247 = \113  & \114 ;
  assign new_n1248 = ~new_n1246 & ~new_n1247;
  assign new_n1249 = ~new_n1245 & ~new_n1248;
  assign new_n1250 = new_n1245 & new_n1248;
  assign new_n1251 = ~new_n1249 & ~new_n1250;
  assign new_n1252 = ~\18  & ~new_n1251;
  assign new_n1253 = ~new_n1244 & ~new_n1252;
  assign new_n1254 = new_n1235 & ~new_n1253;
  assign new_n1255 = ~new_n1235 & new_n1253;
  assign new_n1256 = ~new_n1254 & ~new_n1255;
  assign new_n1257 = ~\257  & ~\260 ;
  assign new_n1258 = \257  & \260 ;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = \18  & ~new_n1259;
  assign new_n1261 = ~new_n871 & ~new_n903;
  assign new_n1262 = ~\18  & ~new_n1261;
  assign new_n1263 = ~new_n1260 & ~new_n1262;
  assign new_n1264 = new_n1256 & ~new_n1263;
  assign new_n1265 = ~new_n1256 & new_n1263;
  assign new_n1266 = ~new_n1171 & ~new_n1172;
  assign new_n1267 = ~new_n1264 & ~new_n1265;
  assign new_n1268 = new_n1266 & new_n1267;
  assign new_n1269 = ~new_n1227 & new_n1268;
  assign new_n1270 = ~new_n1228 & new_n1269;
  assign \10575  = new_n1128 | ~new_n1270;
  assign new_n1272 = ~\115  & new_n427;
  assign new_n1273 = \115  & new_n787;
  assign new_n1274 = ~\189  & \197 ;
  assign new_n1275 = \189  & ~\197 ;
  assign new_n1276 = \18  & ~new_n1274;
  assign new_n1277 = ~new_n1275 & new_n1276;
  assign new_n1278 = ~new_n1272 & ~new_n1273;
  assign new_n1279 = ~new_n1277 & new_n1278;
  assign new_n1280 = ~\118  & new_n536;
  assign new_n1281 = \94  & new_n454;
  assign new_n1282 = ~\187  & \195 ;
  assign new_n1283 = \187  & ~\195 ;
  assign new_n1284 = \18  & ~new_n1282;
  assign new_n1285 = ~new_n1283 & new_n1284;
  assign new_n1286 = ~new_n1280 & ~new_n1281;
  assign new_n1287 = ~new_n1285 & new_n1286;
  assign new_n1288 = ~\47  & new_n531;
  assign new_n1289 = ~\121  & new_n748;
  assign new_n1290 = ~\193  & ~\194 ;
  assign new_n1291 = \193  & \194 ;
  assign new_n1292 = \18  & ~new_n1290;
  assign new_n1293 = ~new_n1291 & new_n1292;
  assign new_n1294 = ~new_n1288 & ~new_n1289;
  assign new_n1295 = ~new_n1293 & new_n1294;
  assign new_n1296 = new_n1287 & ~new_n1295;
  assign new_n1297 = ~new_n1287 & new_n1295;
  assign new_n1298 = ~new_n1296 & ~new_n1297;
  assign new_n1299 = \97  & new_n443;
  assign new_n1300 = ~\97  & new_n633;
  assign new_n1301 = ~\192  & \196 ;
  assign new_n1302 = \192  & ~\196 ;
  assign new_n1303 = \18  & ~new_n1301;
  assign new_n1304 = ~new_n1302 & new_n1303;
  assign new_n1305 = ~new_n1299 & ~new_n1300;
  assign new_n1306 = ~new_n1304 & new_n1305;
  assign new_n1307 = ~\32  & new_n432;
  assign new_n1308 = ~\50  & new_n437;
  assign new_n1309 = ~\190  & ~\191 ;
  assign new_n1310 = \190  & \191 ;
  assign new_n1311 = \18  & ~new_n1309;
  assign new_n1312 = ~new_n1310 & new_n1311;
  assign new_n1313 = ~new_n1307 & ~new_n1308;
  assign new_n1314 = ~new_n1312 & new_n1313;
  assign new_n1315 = new_n1306 & ~new_n1314;
  assign new_n1316 = ~new_n1306 & new_n1314;
  assign new_n1317 = ~new_n1315 & ~new_n1316;
  assign new_n1318 = ~new_n1298 & ~new_n1317;
  assign new_n1319 = new_n1298 & new_n1317;
  assign new_n1320 = ~new_n1318 & ~new_n1319;
  assign new_n1321 = new_n1279 & ~new_n1320;
  assign new_n1322 = ~new_n1279 & new_n1320;
  assign new_n1323 = ~new_n1321 & ~new_n1322;
  assign new_n1324 = ~\166  & ~\167 ;
  assign new_n1325 = \166  & \167 ;
  assign new_n1326 = ~new_n1324 & ~new_n1325;
  assign new_n1327 = ~\165  & ~\168 ;
  assign new_n1328 = \165  & \168 ;
  assign new_n1329 = ~new_n1327 & ~new_n1328;
  assign new_n1330 = \164  & new_n1329;
  assign new_n1331 = ~\164  & ~new_n1329;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = \169  & ~\170 ;
  assign new_n1334 = ~\169  & \170 ;
  assign new_n1335 = ~new_n1333 & ~new_n1334;
  assign new_n1336 = new_n1332 & new_n1335;
  assign new_n1337 = ~new_n1332 & ~new_n1335;
  assign new_n1338 = ~new_n1336 & ~new_n1337;
  assign new_n1339 = new_n1326 & new_n1338;
  assign new_n1340 = ~new_n1326 & ~new_n1338;
  assign new_n1341 = new_n370 & ~new_n1339;
  assign new_n1342 = ~new_n1340 & new_n1341;
  assign new_n1343 = ~new_n466 & ~new_n713;
  assign new_n1344 = new_n664 & ~new_n1343;
  assign new_n1345 = ~new_n664 & new_n1343;
  assign new_n1346 = ~new_n1344 & ~new_n1345;
  assign new_n1347 = ~\26  & new_n470;
  assign new_n1348 = ~\127  & new_n498;
  assign new_n1349 = ~\202  & ~\206 ;
  assign new_n1350 = \202  & \206 ;
  assign new_n1351 = \18  & ~new_n1349;
  assign new_n1352 = ~new_n1350 & new_n1351;
  assign new_n1353 = ~new_n1347 & ~new_n1348;
  assign new_n1354 = ~new_n1352 & new_n1353;
  assign new_n1355 = ~\200  & ~\207 ;
  assign new_n1356 = \200  & \207 ;
  assign new_n1357 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = \198  & ~new_n1357;
  assign new_n1359 = ~\198  & new_n1357;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = \18  & ~new_n1360;
  assign new_n1362 = ~\41  & ~\100 ;
  assign new_n1363 = \41  & \100 ;
  assign new_n1364 = ~new_n1362 & ~new_n1363;
  assign new_n1365 = \29  & ~new_n1364;
  assign new_n1366 = ~\29  & new_n1364;
  assign new_n1367 = ~new_n1365 & ~new_n1366;
  assign new_n1368 = ~\18  & ~new_n1367;
  assign new_n1369 = ~new_n1361 & ~new_n1368;
  assign new_n1370 = new_n1354 & ~new_n1369;
  assign new_n1371 = ~new_n1354 & new_n1369;
  assign new_n1372 = ~new_n1370 & ~new_n1371;
  assign new_n1373 = \44  & new_n476;
  assign new_n1374 = ~\44  & new_n659;
  assign new_n1375 = ~\203  & \208 ;
  assign new_n1376 = \203  & ~\208 ;
  assign new_n1377 = \18  & ~new_n1375;
  assign new_n1378 = ~new_n1376 & new_n1377;
  assign new_n1379 = ~new_n1373 & ~new_n1374;
  assign new_n1380 = ~new_n1378 & new_n1379;
  assign new_n1381 = new_n671 & ~new_n1380;
  assign new_n1382 = ~new_n671 & new_n1380;
  assign new_n1383 = ~new_n1381 & ~new_n1382;
  assign new_n1384 = ~new_n1372 & ~new_n1383;
  assign new_n1385 = new_n1372 & new_n1383;
  assign new_n1386 = ~new_n1384 & ~new_n1385;
  assign new_n1387 = new_n1346 & new_n1386;
  assign new_n1388 = ~new_n1346 & ~new_n1386;
  assign new_n1389 = ~\175  & ~\176 ;
  assign new_n1390 = \175  & \176 ;
  assign new_n1391 = ~new_n1389 & ~new_n1390;
  assign new_n1392 = \173  & new_n1391;
  assign new_n1393 = ~\173  & ~new_n1391;
  assign new_n1394 = ~new_n1392 & ~new_n1393;
  assign new_n1395 = ~\174  & ~new_n1394;
  assign new_n1396 = \174  & new_n1394;
  assign new_n1397 = new_n370 & ~new_n1395;
  assign new_n1398 = ~new_n1396 & new_n1397;
  assign new_n1399 = new_n343 & new_n411;
  assign new_n1400 = ~\144  & new_n344;
  assign new_n1401 = ~\179  & ~new_n818;
  assign new_n1402 = \179  & new_n818;
  assign new_n1403 = \18  & ~new_n1401;
  assign new_n1404 = ~new_n1402 & new_n1403;
  assign new_n1405 = ~new_n1399 & ~new_n1400;
  assign new_n1406 = ~new_n1404 & new_n1405;
  assign new_n1407 = ~new_n1398 & new_n1406;
  assign new_n1408 = new_n1398 & ~new_n1406;
  assign new_n1409 = ~new_n1407 & ~new_n1408;
  assign new_n1410 = ~\141  & \147 ;
  assign new_n1411 = ~new_n422 & ~new_n1002;
  assign new_n1412 = ~new_n1410 & ~new_n1411;
  assign new_n1413 = ~\171  & \181 ;
  assign new_n1414 = \171  & ~\181 ;
  assign new_n1415 = \18  & ~new_n1413;
  assign new_n1416 = ~new_n1414 & new_n1415;
  assign new_n1417 = ~new_n1412 & ~new_n1416;
  assign new_n1418 = ~\135  & new_n416;
  assign new_n1419 = \135  & new_n810;
  assign new_n1420 = ~\178  & \180 ;
  assign new_n1421 = \178  & ~\180 ;
  assign new_n1422 = \18  & ~new_n1420;
  assign new_n1423 = ~new_n1421 & new_n1422;
  assign new_n1424 = ~new_n1418 & ~new_n1419;
  assign new_n1425 = ~new_n1423 & new_n1424;
  assign new_n1426 = new_n1417 & ~new_n1425;
  assign new_n1427 = ~new_n1417 & new_n1425;
  assign new_n1428 = ~new_n1426 & ~new_n1427;
  assign new_n1429 = new_n1409 & ~new_n1428;
  assign new_n1430 = ~new_n1409 & new_n1428;
  assign new_n1431 = ~new_n1323 & ~new_n1342;
  assign new_n1432 = ~new_n1429 & ~new_n1430;
  assign new_n1433 = new_n1431 & new_n1432;
  assign new_n1434 = ~new_n1387 & ~new_n1388;
  assign \10576  = ~new_n1433 | ~new_n1434;
  assign new_n1436 = ~new_n425 & ~new_n573;
  assign new_n1437 = ~new_n571 & new_n1436;
  assign new_n1438 = new_n571 & ~new_n1436;
  assign \10632  = new_n1437 | new_n1438;
  assign new_n1440 = \251  & new_n364;
  assign new_n1441 = ~new_n365 & ~new_n1440;
  assign new_n1442 = ~new_n594 & new_n1441;
  assign new_n1443 = new_n594 & ~new_n1441;
  assign \10641  = new_n1442 | new_n1443;
  assign new_n1445 = ~new_n403 & ~new_n404;
  assign new_n1446 = new_n580 & ~new_n1445;
  assign new_n1447 = ~new_n580 & new_n1445;
  assign \10711  = ~new_n1446 & ~new_n1447;
  assign new_n1449 = ~new_n410 & new_n578;
  assign \10712  = ~new_n579 & ~new_n1449;
  assign new_n1451 = ~new_n414 & ~new_n415;
  assign new_n1452 = new_n576 & ~new_n1451;
  assign new_n1453 = ~new_n576 & new_n1451;
  assign \10713  = ~new_n1452 & ~new_n1453;
  assign new_n1455 = ~new_n421 & new_n1437;
  assign new_n1456 = ~new_n421 & new_n425;
  assign new_n1457 = ~new_n426 & ~new_n1456;
  assign new_n1458 = ~new_n1437 & ~new_n1457;
  assign \10714  = ~new_n1455 & ~new_n1458;
  assign new_n1460 = ~new_n349 & new_n598;
  assign \10715  = ~new_n599 & ~new_n1460;
  assign new_n1462 = ~new_n354 & new_n596;
  assign \10716  = ~new_n597 & ~new_n1462;
  assign new_n1464 = new_n382 & new_n594;
  assign new_n1465 = ~new_n367 & ~new_n1464;
  assign new_n1466 = ~new_n357 & ~new_n358;
  assign new_n1467 = ~new_n1465 & new_n1466;
  assign new_n1468 = new_n1465 & ~new_n1466;
  assign \10717  = ~new_n1467 & ~new_n1468;
  assign new_n1470 = ~new_n1440 & ~new_n1442;
  assign new_n1471 = new_n381 & ~new_n1470;
  assign new_n1472 = ~new_n381 & new_n1470;
  assign \10718  = new_n1471 | new_n1472;
  assign new_n1474 = ~\882  & ~\883 ;
  assign new_n1475 = ~\884  & ~\885 ;
  assign new_n1476 = new_n1474 & new_n1475;
  assign new_n1477 = ~\10576  & new_n1476;
  assign new_n1478 = ~\10575  & new_n1477;
  assign \10729  = \10574  | ~new_n1478;
  assign new_n1480 = new_n590 & ~new_n592;
  assign \10760  = new_n593 | new_n1480;
  assign new_n1482 = ~new_n391 & new_n588;
  assign \10761  = new_n589 | new_n1482;
  assign new_n1484 = ~new_n584 & new_n585;
  assign new_n1485 = new_n583 & ~new_n585;
  assign new_n1486 = ~new_n1484 & ~new_n1485;
  assign new_n1487 = ~new_n586 & ~new_n1486;
  assign \10762  = new_n587 | new_n1487;
  assign new_n1489 = ~new_n397 & ~new_n585;
  assign new_n1490 = new_n582 & ~new_n1489;
  assign \10763  = ~new_n1485 & ~new_n1490;
  assign new_n1492 = ~new_n459 & new_n528;
  assign \10827  = ~new_n529 & ~new_n1492;
  assign new_n1494 = \263  & ~new_n603;
  assign new_n1495 = new_n341 & ~new_n1494;
  assign new_n1496 = new_n600 & ~new_n1495;
  assign new_n1497 = ~\38  & ~new_n341;
  assign new_n1498 = ~new_n602 & ~new_n1497;
  assign new_n1499 = ~new_n600 & new_n1498;
  assign new_n1500 = ~new_n1496 & ~new_n1499;
  assign new_n1501 = ~\38  & ~new_n600;
  assign new_n1502 = \38  & new_n600;
  assign new_n1503 = ~new_n1501 & ~new_n1502;
  assign new_n1504 = \267  & \382 ;
  assign new_n1505 = new_n1503 & new_n1504;
  assign \10837  = ~new_n1500 & ~new_n1505;
  assign new_n1507 = new_n601 & ~new_n1503;
  assign new_n1508 = ~new_n601 & new_n1503;
  assign \10839  = new_n1507 | new_n1508;
  assign new_n1510 = ~new_n453 & ~new_n561;
  assign \10868  = ~new_n562 & ~new_n1510;
  assign new_n1512 = ~new_n534 & ~new_n535;
  assign new_n1513 = ~new_n528 & new_n551;
  assign new_n1514 = ~new_n552 & ~new_n1513;
  assign new_n1515 = new_n1512 & ~new_n1514;
  assign new_n1516 = ~new_n1512 & new_n1514;
  assign \10869  = ~new_n1515 & ~new_n1516;
  assign new_n1518 = ~new_n530 & new_n557;
  assign new_n1519 = ~new_n543 & ~new_n1518;
  assign new_n1520 = new_n556 & ~new_n1519;
  assign new_n1521 = ~new_n556 & new_n1519;
  assign \10870  = ~new_n1520 & ~new_n1521;
  assign new_n1523 = new_n530 & ~new_n557;
  assign \10871  = ~new_n1518 & ~new_n1523;
  assign new_n1525 = ~new_n430 & ~new_n431;
  assign new_n1526 = new_n569 & new_n1525;
  assign new_n1527 = ~new_n569 & ~new_n1525;
  assign \10905  = new_n1526 | new_n1527;
  assign new_n1529 = ~new_n435 & ~new_n436;
  assign new_n1530 = ~new_n567 & new_n1529;
  assign new_n1531 = new_n567 & ~new_n1529;
  assign \10906  = new_n1530 | new_n1531;
  assign new_n1533 = ~new_n442 & ~new_n565;
  assign \10907  = new_n566 | new_n1533;
  assign new_n1535 = ~new_n446 & ~new_n447;
  assign new_n1536 = ~new_n563 & new_n1535;
  assign new_n1537 = new_n563 & ~new_n1535;
  assign \10908  = ~new_n1536 & ~new_n1537;
  assign new_n1539 = ~new_n390 & ~new_n400;
  assign new_n1540 = ~new_n586 & new_n1539;
  assign new_n1541 = ~new_n389 & ~new_n1540;
  assign new_n1542 = new_n397 & ~new_n398;
  assign new_n1543 = ~new_n394 & ~new_n397;
  assign new_n1544 = ~new_n586 & new_n1543;
  assign new_n1545 = ~new_n1542 & ~new_n1544;
  assign new_n1546 = new_n592 & ~new_n1545;
  assign new_n1547 = ~new_n592 & new_n1545;
  assign new_n1548 = ~new_n1546 & ~new_n1547;
  assign new_n1549 = new_n1541 & ~new_n1548;
  assign new_n1550 = ~new_n1541 & new_n1548;
  assign new_n1551 = ~new_n1549 & ~new_n1550;
  assign new_n1552 = new_n582 & new_n1551;
  assign new_n1553 = ~new_n586 & ~new_n1484;
  assign new_n1554 = ~new_n389 & new_n400;
  assign new_n1555 = ~new_n1539 & ~new_n1554;
  assign new_n1556 = new_n592 & ~new_n1555;
  assign new_n1557 = ~new_n592 & new_n1555;
  assign new_n1558 = ~new_n1556 & ~new_n1557;
  assign new_n1559 = new_n1553 & ~new_n1558;
  assign new_n1560 = ~new_n1553 & new_n1558;
  assign new_n1561 = ~new_n1559 & ~new_n1560;
  assign new_n1562 = ~new_n582 & new_n1561;
  assign new_n1563 = ~new_n1552 & ~new_n1562;
  assign new_n1564 = ~new_n415 & ~new_n426;
  assign new_n1565 = ~new_n575 & new_n1564;
  assign new_n1566 = ~new_n414 & ~new_n1565;
  assign new_n1567 = ~new_n409 & ~new_n579;
  assign new_n1568 = ~new_n419 & new_n573;
  assign new_n1569 = ~new_n420 & ~new_n573;
  assign new_n1570 = ~new_n426 & new_n1569;
  assign new_n1571 = ~new_n1568 & ~new_n1570;
  assign new_n1572 = new_n1445 & ~new_n1571;
  assign new_n1573 = ~new_n1445 & new_n1571;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = new_n1567 & ~new_n1574;
  assign new_n1576 = ~new_n1567 & new_n1574;
  assign new_n1577 = ~new_n1575 & ~new_n1576;
  assign new_n1578 = new_n1566 & ~new_n1577;
  assign new_n1579 = ~new_n1566 & new_n1577;
  assign new_n1580 = ~new_n1578 & ~new_n1579;
  assign new_n1581 = new_n571 & ~new_n1580;
  assign new_n1582 = new_n413 & ~new_n575;
  assign new_n1583 = \283  & ~new_n409;
  assign new_n1584 = ~new_n575 & new_n1583;
  assign new_n1585 = ~\283  & new_n409;
  assign new_n1586 = ~new_n1584 & ~new_n1585;
  assign new_n1587 = new_n1582 & new_n1586;
  assign new_n1588 = ~\283  & new_n575;
  assign new_n1589 = ~new_n408 & ~new_n1588;
  assign new_n1590 = ~\283  & new_n408;
  assign new_n1591 = ~new_n1589 & ~new_n1590;
  assign new_n1592 = ~new_n413 & new_n1591;
  assign new_n1593 = ~new_n1445 & ~new_n1587;
  assign new_n1594 = ~new_n1592 & new_n1593;
  assign new_n1595 = new_n413 & ~new_n1586;
  assign new_n1596 = ~new_n413 & new_n575;
  assign new_n1597 = ~new_n1591 & new_n1596;
  assign new_n1598 = new_n1445 & ~new_n1595;
  assign new_n1599 = ~new_n1597 & new_n1598;
  assign new_n1600 = ~new_n1594 & ~new_n1599;
  assign new_n1601 = ~new_n408 & ~new_n1583;
  assign new_n1602 = new_n1445 & ~new_n1601;
  assign new_n1603 = ~new_n1445 & new_n1601;
  assign new_n1604 = ~new_n1582 & ~new_n1596;
  assign new_n1605 = ~new_n1602 & ~new_n1603;
  assign new_n1606 = new_n1604 & new_n1605;
  assign new_n1607 = ~new_n1600 & ~new_n1606;
  assign new_n1608 = ~new_n1457 & ~new_n1607;
  assign new_n1609 = new_n1457 & new_n1607;
  assign new_n1610 = ~new_n1608 & ~new_n1609;
  assign new_n1611 = ~new_n571 & ~new_n1610;
  assign new_n1612 = ~new_n1581 & ~new_n1611;
  assign new_n1613 = new_n1563 & ~new_n1612;
  assign new_n1614 = ~new_n1563 & new_n1612;
  assign \11333  = ~new_n1613 & ~new_n1614;
  assign new_n1616 = ~new_n353 & new_n383;
  assign new_n1617 = ~new_n352 & ~new_n369;
  assign new_n1618 = ~new_n383 & new_n1617;
  assign new_n1619 = ~new_n353 & new_n369;
  assign new_n1620 = ~new_n1616 & ~new_n1619;
  assign new_n1621 = ~new_n1618 & new_n1620;
  assign new_n1622 = new_n380 & ~new_n1621;
  assign new_n1623 = ~new_n380 & new_n1621;
  assign new_n1624 = ~new_n1622 & ~new_n1623;
  assign new_n1625 = new_n594 & new_n1624;
  assign new_n1626 = ~new_n380 & new_n381;
  assign new_n1627 = ~new_n1617 & ~new_n1619;
  assign new_n1628 = new_n1626 & ~new_n1627;
  assign new_n1629 = ~new_n1626 & new_n1627;
  assign new_n1630 = ~new_n1628 & ~new_n1629;
  assign new_n1631 = ~new_n594 & new_n1630;
  assign new_n1632 = ~new_n1625 & ~new_n1631;
  assign new_n1633 = new_n354 & \10839 ;
  assign new_n1634 = ~new_n354 & ~\10839 ;
  assign new_n1635 = ~new_n1633 & ~new_n1634;
  assign new_n1636 = new_n1632 & ~new_n1635;
  assign new_n1637 = ~new_n1632 & new_n1635;
  assign new_n1638 = ~new_n1636 & ~new_n1637;
  assign new_n1639 = new_n370 & new_n987;
  assign new_n1640 = \106  & \260 ;
  assign new_n1641 = ~new_n868 & ~new_n1640;
  assign new_n1642 = new_n1639 & ~new_n1641;
  assign new_n1643 = ~new_n1639 & new_n1641;
  assign new_n1644 = ~new_n1642 & ~new_n1643;
  assign new_n1645 = \10837  & ~new_n1644;
  assign new_n1646 = ~\10837  & new_n1644;
  assign new_n1647 = ~new_n1645 & ~new_n1646;
  assign new_n1648 = new_n1638 & new_n1647;
  assign new_n1649 = ~new_n1638 & ~new_n1647;
  assign new_n1650 = ~new_n1648 & ~new_n1649;
  assign new_n1651 = ~new_n362 & new_n1440;
  assign new_n1652 = ~new_n361 & ~new_n1440;
  assign new_n1653 = ~new_n1651 & ~new_n1652;
  assign new_n1654 = new_n1650 & ~new_n1653;
  assign new_n1655 = ~new_n1650 & new_n1653;
  assign \11334  = new_n1654 | new_n1655;
  assign new_n1657 = new_n456 & ~new_n543;
  assign new_n1658 = ~new_n548 & ~new_n1657;
  assign new_n1659 = ~new_n544 & ~new_n1658;
  assign new_n1660 = ~new_n453 & new_n1512;
  assign new_n1661 = new_n453 & ~new_n1512;
  assign new_n1662 = ~new_n1660 & ~new_n1661;
  assign new_n1663 = ~new_n1659 & ~new_n1662;
  assign new_n1664 = new_n1659 & new_n1662;
  assign new_n1665 = ~new_n1663 & ~new_n1664;
  assign new_n1666 = ~new_n557 & ~new_n1665;
  assign new_n1667 = new_n557 & ~new_n1662;
  assign new_n1668 = ~new_n1666 & ~new_n1667;
  assign new_n1669 = new_n551 & ~new_n1668;
  assign new_n1670 = ~new_n551 & new_n1668;
  assign new_n1671 = ~new_n1669 & ~new_n1670;
  assign new_n1672 = ~new_n459 & new_n556;
  assign new_n1673 = new_n459 & ~new_n556;
  assign new_n1674 = ~new_n1672 & ~new_n1673;
  assign new_n1675 = new_n554 & ~new_n1674;
  assign new_n1676 = ~new_n560 & new_n1674;
  assign new_n1677 = ~new_n1675 & ~new_n1676;
  assign new_n1678 = new_n1671 & ~new_n1677;
  assign new_n1679 = ~new_n1671 & new_n1677;
  assign new_n1680 = ~new_n1678 & ~new_n1679;
  assign new_n1681 = ~new_n528 & new_n1680;
  assign new_n1682 = ~new_n556 & ~new_n557;
  assign new_n1683 = ~new_n558 & ~new_n1682;
  assign new_n1684 = ~new_n534 & new_n552;
  assign new_n1685 = ~new_n553 & ~new_n1684;
  assign new_n1686 = ~new_n1665 & new_n1685;
  assign new_n1687 = new_n1665 & ~new_n1685;
  assign new_n1688 = ~new_n1686 & ~new_n1687;
  assign new_n1689 = new_n1683 & new_n1688;
  assign new_n1690 = ~new_n1683 & ~new_n1688;
  assign new_n1691 = ~new_n1689 & ~new_n1690;
  assign new_n1692 = new_n528 & new_n1691;
  assign new_n1693 = ~new_n1681 & ~new_n1692;
  assign new_n1694 = new_n442 & new_n446;
  assign new_n1695 = ~new_n440 & ~new_n447;
  assign new_n1696 = new_n440 & new_n447;
  assign new_n1697 = ~new_n1695 & ~new_n1696;
  assign new_n1698 = ~new_n1694 & ~new_n1697;
  assign new_n1699 = ~\10905  & ~new_n1529;
  assign new_n1700 = \10905  & new_n1529;
  assign new_n1701 = ~new_n1699 & ~new_n1700;
  assign new_n1702 = new_n1698 & new_n1701;
  assign new_n1703 = ~new_n1698 & ~new_n1701;
  assign new_n1704 = ~new_n1702 & ~new_n1703;
  assign new_n1705 = new_n563 & ~new_n1704;
  assign new_n1706 = ~new_n442 & ~new_n446;
  assign new_n1707 = ~new_n1694 & ~new_n1706;
  assign new_n1708 = ~new_n441 & ~new_n1695;
  assign new_n1709 = ~new_n436 & new_n1708;
  assign new_n1710 = ~new_n435 & ~new_n1708;
  assign new_n1711 = ~new_n1709 & ~new_n1710;
  assign new_n1712 = ~new_n1525 & new_n1711;
  assign new_n1713 = new_n1525 & ~new_n1711;
  assign new_n1714 = ~new_n1712 & ~new_n1713;
  assign new_n1715 = new_n1707 & new_n1714;
  assign new_n1716 = ~new_n1707 & ~new_n1714;
  assign new_n1717 = ~new_n1715 & ~new_n1716;
  assign new_n1718 = ~new_n563 & ~new_n1717;
  assign new_n1719 = ~new_n1705 & ~new_n1718;
  assign new_n1720 = new_n1693 & ~new_n1719;
  assign new_n1721 = ~new_n1693 & new_n1719;
  assign \11340  = new_n1720 | new_n1721;
  assign new_n1723 = new_n333 & ~new_n493;
  assign new_n1724 = new_n335 & new_n492;
  assign new_n1725 = ~new_n505 & ~new_n1724;
  assign new_n1726 = ~new_n1723 & ~new_n1725;
  assign new_n1727 = new_n515 & ~new_n1726;
  assign new_n1728 = ~new_n515 & new_n1726;
  assign new_n1729 = ~new_n1727 & ~new_n1728;
  assign new_n1730 = new_n488 & ~new_n1729;
  assign new_n1731 = new_n497 & new_n503;
  assign new_n1732 = ~new_n502 & new_n510;
  assign new_n1733 = new_n502 & ~new_n510;
  assign new_n1734 = ~new_n1732 & ~new_n1733;
  assign new_n1735 = ~new_n1731 & new_n1734;
  assign new_n1736 = new_n1730 & new_n1735;
  assign new_n1737 = ~new_n509 & ~new_n1734;
  assign new_n1738 = ~new_n501 & ~new_n1737;
  assign new_n1739 = ~new_n488 & new_n1729;
  assign new_n1740 = ~new_n1738 & new_n1739;
  assign new_n1741 = new_n488 & ~new_n504;
  assign new_n1742 = ~new_n1729 & ~new_n1737;
  assign new_n1743 = ~new_n1741 & ~new_n1742;
  assign new_n1744 = ~new_n501 & ~new_n1730;
  assign new_n1745 = ~new_n1743 & new_n1744;
  assign new_n1746 = \367  & ~new_n1736;
  assign new_n1747 = ~new_n1740 & new_n1746;
  assign new_n1748 = ~new_n1745 & new_n1747;
  assign new_n1749 = ~new_n493 & new_n500;
  assign new_n1750 = new_n493 & ~new_n500;
  assign new_n1751 = ~new_n1749 & ~new_n1750;
  assign new_n1752 = ~new_n333 & new_n1751;
  assign new_n1753 = ~new_n336 & ~new_n1751;
  assign new_n1754 = ~new_n1752 & ~new_n1753;
  assign new_n1755 = ~new_n492 & new_n500;
  assign new_n1756 = new_n492 & ~new_n500;
  assign new_n1757 = new_n335 & ~new_n1755;
  assign new_n1758 = ~new_n1756 & new_n1757;
  assign new_n1759 = ~new_n1754 & ~new_n1758;
  assign new_n1760 = ~\316  & ~new_n515;
  assign new_n1761 = \316  & new_n515;
  assign new_n1762 = ~new_n1760 & ~new_n1761;
  assign new_n1763 = ~new_n488 & new_n508;
  assign new_n1764 = ~new_n508 & ~new_n510;
  assign new_n1765 = ~new_n1763 & ~new_n1764;
  assign new_n1766 = new_n1762 & ~new_n1765;
  assign new_n1767 = ~new_n1762 & new_n1765;
  assign new_n1768 = ~new_n1766 & ~new_n1767;
  assign new_n1769 = ~new_n1759 & ~new_n1768;
  assign new_n1770 = new_n1759 & new_n1768;
  assign new_n1771 = ~\367  & ~new_n1769;
  assign new_n1772 = ~new_n1770 & new_n1771;
  assign new_n1773 = ~new_n1748 & ~new_n1772;
  assign new_n1774 = new_n465 & ~new_n511;
  assign new_n1775 = ~new_n465 & new_n511;
  assign new_n1776 = ~new_n1774 & ~new_n1775;
  assign new_n1777 = new_n1773 & new_n1776;
  assign new_n1778 = ~new_n1773 & ~new_n1776;
  assign new_n1779 = ~new_n1777 & ~new_n1778;
  assign new_n1780 = ~new_n520 & ~new_n928;
  assign new_n1781 = ~new_n474 & ~new_n480;
  assign new_n1782 = ~new_n469 & new_n1781;
  assign new_n1783 = ~new_n523 & ~new_n1781;
  assign new_n1784 = ~new_n1782 & ~new_n1783;
  assign new_n1785 = ~new_n1780 & ~new_n1784;
  assign new_n1786 = new_n1780 & new_n1784;
  assign new_n1787 = ~new_n1785 & ~new_n1786;
  assign new_n1788 = new_n517 & ~new_n1787;
  assign new_n1789 = ~new_n480 & ~new_n927;
  assign new_n1790 = ~new_n469 & new_n521;
  assign new_n1791 = ~new_n521 & ~new_n523;
  assign new_n1792 = ~new_n1790 & ~new_n1791;
  assign new_n1793 = new_n1789 & ~new_n1792;
  assign new_n1794 = ~new_n1789 & new_n1792;
  assign new_n1795 = ~new_n1793 & ~new_n1794;
  assign new_n1796 = ~new_n517 & ~new_n1795;
  assign new_n1797 = ~new_n1788 & ~new_n1796;
  assign new_n1798 = new_n1779 & ~new_n1797;
  assign new_n1799 = ~new_n1779 & new_n1797;
  assign \11342  = ~new_n1798 & ~new_n1799;
  assign \582  = ~\15 ;
  assign \387  = \1 ;
  assign \388  = \1 ;
  assign \478  = \248 ;
  assign \482  = \254 ;
  assign \484  = \257 ;
  assign \486  = \260 ;
  assign \489  = \263 ;
  assign \492  = \267 ;
  assign \501  = \274 ;
  assign \505  = \280 ;
  assign \507  = \283 ;
  assign \509  = \286 ;
  assign \511  = \289 ;
  assign \513  = \293 ;
  assign \515  = \296 ;
  assign \517  = \299 ;
  assign \519  = \303 ;
  assign \535  = \307 ;
  assign \537  = \310 ;
  assign \539  = \313 ;
  assign \541  = \316 ;
  assign \543  = \319 ;
  assign \545  = \322 ;
  assign \547  = \325 ;
  assign \549  = \328 ;
  assign \551  = \331 ;
  assign \553  = \334 ;
  assign \556  = \337 ;
  assign \559  = \343 ;
  assign \561  = \346 ;
  assign \563  = \349 ;
  assign \565  = \352 ;
  assign \567  = \355 ;
  assign \569  = \358 ;
  assign \571  = \361 ;
  assign \573  = \364 ;
  assign \643  = \251 ;
  assign \707  = \277 ;
  assign \813  = \340 ;
  assign \889  = \1 ;
  assign \945  = \106 ;
  assign \1111  = \582 ;
  assign \1112  = \1110 ;
  assign \1114  = \582 ;
  assign \1489  = \1113 ;
  assign \1490  = \1 ;
  assign \10103  = \10102 ;
  assign \10104  = \10101 ;
  assign \10628  = \10102 ;
  assign \10706  = \10101 ;
  assign \10759  = \10101 ;
  assign \10838  = \10837 ;
  assign \10840  = \10839 ;
endmodule


