// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    p_193_130_, p_257_171_, p_2435_225_, p_79_60_, p_135_106_, p_142_113_,
    p_192_129_, p_209_146_, p_2096_218_, p_2454_230_, p_4_3_, p_51_36_,
    p_52_37_, p_112_87_, p_126_99_, p_179_118_, p_189_126_, p_21_14_,
    p_25_18_, p_90_69_, p_206_143_, p_253_167_, p_277_187_, p_60_43_,
    p_61_44_, p_66_49_, p_202_139_, p_22_15_, p_24_17_, p_119_94_,
    p_132_105_, p_203_140_, p_250_164_, p_267_177_, p_270_180_, p_559_193_,
    p_2443_227_, p_3_2_, p_53_38_, p_54_39_, p_102_79_, p_182_121_,
    p_212_149_, p_1961_204_, p_1986_209_, p_2090_217_, p_2430_224_,
    p_23_16_, p_169_114_, p_213_150_, p_242_156_, p_28_21_, p_29_22_,
    p_93_72_, p_94_73_, p_95_74_, p_96_75_, p_128_101_, p_651_195_,
    p_661_196_, p_14_9_, p_32_23_, p_34_25_, p_36_27_, p_67_50_, p_69_52_,
    p_104_81_, p_106_83_, p_252_166_, p_269_179_, p_276_186_, p_2_1_,
    p_72_53_, p_99_76_, p_100_77_, p_113_88_, p_125_98_, p_2451_229_,
    p_35_26_, p_116_91_, p_136_107_, p_240_154_, p_273_183_, p_62_45_,
    p_63_46_, p_64_47_, p_65_48_, p_183_122_, p_199_136_, p_1981_208_,
    p_1996_211_, p_11_8_, p_26_19_, p_140_111_, p_207_144_, p_214_151_,
    p_243_157_, p_263_173_, p_1_0_, p_186_125_, p_196_133_, p_247_161_,
    p_33_24_, p_68_51_, p_204_141_, p_266_176_, p_279_189_, p_2678_232_,
    p_19_12_, p_85_64_, p_86_65_, p_87_66_, p_88_67_, p_89_68_, p_120_95_,
    p_181_120_, p_200_137_, p_2100_219_, p_130_103_, p_180_119_,
    p_241_155_, p_265_175_, p_272_182_, p_567_194_, p_8_7_, p_15_10_,
    p_16_11_, p_80_61_, p_81_62_, p_127_100_, p_174_115_, p_184_123_,
    p_198_135_, p_210_147_, p_56_41_, p_103_80_, p_107_84_, p_244_158_,
    p_268_178_, p_1976_207_, p_195_132_, p_248_162_, p_2066_212_,
    p_2106_222_, p_2474_231_, p_43_30_, p_57_42_, p_117_92_, p_137_108_,
    p_278_188_, p_483_191_, p_1384_202_, p_1971_206_, p_7_6_, p_73_54_,
    p_74_55_, p_123_96_, p_177_116_, p_256_170_, p_1083_199_, p_1341_200_,
    p_1991_210_, p_2067_213_, p_2078_215_, p_2105_221_, p_37_28_, p_44_31_,
    p_191_128_, p_208_145_, p_255_169_, p_262_172_, p_275_185_, p_868_198_,
    p_27_20_, p_91_70_, p_92_71_, p_178_117_, p_185_124_, p_197_134_,
    p_211_148_, p_239_153_, p_246_160_, p_2084_216_, p_2104_220_,
    p_108_85_, p_205_142_, p_245_159_, p_2446_228_, p_6_5_, p_40_29_,
    p_75_56_, p_76_57_, p_194_131_, p_201_138_, p_249_163_, p_452_190_,
    p_47_32_, p_131_104_, p_141_112_, p_215_152_, p_264_174_, p_2427_223_,
    p_1966_205_, p_2438_226_, p_20_13_, p_48_33_, p_55_40_, p_115_90_,
    p_190_127_, p_254_168_, p_274_184_, p_543_192_, p_1956_203_, p_5_4_,
    p_50_35_, p_77_58_, p_78_59_, p_82_63_, p_101_78_, p_111_86_,
    p_114_89_, p_124_97_, p_129_102_, p_139_110_, p_860_197_, p_1348_201_,
    p_49_34_, p_105_82_, p_118_93_, p_138_109_, p_251_165_, p_271_181_,
    p_2072_214_,
    p_284_847_, p_171_621_, p_145_1358_, p_150_1277_, p_188_761_,
    p_221_305_, p_311_1278_, p_158_349_, p_235_307_, p_259_414_,
    p_299_692_, p_160_609_, p_367_288_, p_288_700_, p_301_694_, p_384_262_,
    p_218_311_, p_261_506_, p_236_303_, p_319_656_, p_321_848_, p_350_301_,
    p_397_1406_, p_148_851_, p_220_306_, p_369_289_, p_164_607_,
    p_411_264_, p_231_1422_, p_297_849_, p_168_623_, p_156_1046_,
    p_337_263_, p_153_671_, p_223_413_, p_303_698_, p_331_1401_,
    p_391_379_, p_395_1392_, p_282_922_, p_173_389_, p_217_423_,
    p_229_1180_, p_280_850_, p_335_299_, p_162_612_, p_227_1179_,
    p_237_309_, p_176_803_, p_305_702_, p_290_704_, p_329_1414_,
    p_286_696_, p_295_1400_, p_401_1276_, p_238_304_, p_323_923_,
    p_325_507_, p_219_302_, p_166_625_, p_409_298_, p_234_376_,
    p_308_1425_, p_225_1424_  );
  input  p_193_130_, p_257_171_, p_2435_225_, p_79_60_, p_135_106_,
    p_142_113_, p_192_129_, p_209_146_, p_2096_218_, p_2454_230_, p_4_3_,
    p_51_36_, p_52_37_, p_112_87_, p_126_99_, p_179_118_, p_189_126_,
    p_21_14_, p_25_18_, p_90_69_, p_206_143_, p_253_167_, p_277_187_,
    p_60_43_, p_61_44_, p_66_49_, p_202_139_, p_22_15_, p_24_17_,
    p_119_94_, p_132_105_, p_203_140_, p_250_164_, p_267_177_, p_270_180_,
    p_559_193_, p_2443_227_, p_3_2_, p_53_38_, p_54_39_, p_102_79_,
    p_182_121_, p_212_149_, p_1961_204_, p_1986_209_, p_2090_217_,
    p_2430_224_, p_23_16_, p_169_114_, p_213_150_, p_242_156_, p_28_21_,
    p_29_22_, p_93_72_, p_94_73_, p_95_74_, p_96_75_, p_128_101_,
    p_651_195_, p_661_196_, p_14_9_, p_32_23_, p_34_25_, p_36_27_,
    p_67_50_, p_69_52_, p_104_81_, p_106_83_, p_252_166_, p_269_179_,
    p_276_186_, p_2_1_, p_72_53_, p_99_76_, p_100_77_, p_113_88_,
    p_125_98_, p_2451_229_, p_35_26_, p_116_91_, p_136_107_, p_240_154_,
    p_273_183_, p_62_45_, p_63_46_, p_64_47_, p_65_48_, p_183_122_,
    p_199_136_, p_1981_208_, p_1996_211_, p_11_8_, p_26_19_, p_140_111_,
    p_207_144_, p_214_151_, p_243_157_, p_263_173_, p_1_0_, p_186_125_,
    p_196_133_, p_247_161_, p_33_24_, p_68_51_, p_204_141_, p_266_176_,
    p_279_189_, p_2678_232_, p_19_12_, p_85_64_, p_86_65_, p_87_66_,
    p_88_67_, p_89_68_, p_120_95_, p_181_120_, p_200_137_, p_2100_219_,
    p_130_103_, p_180_119_, p_241_155_, p_265_175_, p_272_182_, p_567_194_,
    p_8_7_, p_15_10_, p_16_11_, p_80_61_, p_81_62_, p_127_100_, p_174_115_,
    p_184_123_, p_198_135_, p_210_147_, p_56_41_, p_103_80_, p_107_84_,
    p_244_158_, p_268_178_, p_1976_207_, p_195_132_, p_248_162_,
    p_2066_212_, p_2106_222_, p_2474_231_, p_43_30_, p_57_42_, p_117_92_,
    p_137_108_, p_278_188_, p_483_191_, p_1384_202_, p_1971_206_, p_7_6_,
    p_73_54_, p_74_55_, p_123_96_, p_177_116_, p_256_170_, p_1083_199_,
    p_1341_200_, p_1991_210_, p_2067_213_, p_2078_215_, p_2105_221_,
    p_37_28_, p_44_31_, p_191_128_, p_208_145_, p_255_169_, p_262_172_,
    p_275_185_, p_868_198_, p_27_20_, p_91_70_, p_92_71_, p_178_117_,
    p_185_124_, p_197_134_, p_211_148_, p_239_153_, p_246_160_,
    p_2084_216_, p_2104_220_, p_108_85_, p_205_142_, p_245_159_,
    p_2446_228_, p_6_5_, p_40_29_, p_75_56_, p_76_57_, p_194_131_,
    p_201_138_, p_249_163_, p_452_190_, p_47_32_, p_131_104_, p_141_112_,
    p_215_152_, p_264_174_, p_2427_223_, p_1966_205_, p_2438_226_,
    p_20_13_, p_48_33_, p_55_40_, p_115_90_, p_190_127_, p_254_168_,
    p_274_184_, p_543_192_, p_1956_203_, p_5_4_, p_50_35_, p_77_58_,
    p_78_59_, p_82_63_, p_101_78_, p_111_86_, p_114_89_, p_124_97_,
    p_129_102_, p_139_110_, p_860_197_, p_1348_201_, p_49_34_, p_105_82_,
    p_118_93_, p_138_109_, p_251_165_, p_271_181_, p_2072_214_;
  output p_284_847_, p_171_621_, p_145_1358_, p_150_1277_, p_188_761_,
    p_221_305_, p_311_1278_, p_158_349_, p_235_307_, p_259_414_,
    p_299_692_, p_160_609_, p_367_288_, p_288_700_, p_301_694_, p_384_262_,
    p_218_311_, p_261_506_, p_236_303_, p_319_656_, p_321_848_, p_350_301_,
    p_397_1406_, p_148_851_, p_220_306_, p_369_289_, p_164_607_,
    p_411_264_, p_231_1422_, p_297_849_, p_168_623_, p_156_1046_,
    p_337_263_, p_153_671_, p_223_413_, p_303_698_, p_331_1401_,
    p_391_379_, p_395_1392_, p_282_922_, p_173_389_, p_217_423_,
    p_229_1180_, p_280_850_, p_335_299_, p_162_612_, p_227_1179_,
    p_237_309_, p_176_803_, p_305_702_, p_290_704_, p_329_1414_,
    p_286_696_, p_295_1400_, p_401_1276_, p_238_304_, p_323_923_,
    p_325_507_, p_219_302_, p_166_625_, p_409_298_, p_234_376_,
    p_308_1425_, p_225_1424_;
  wire new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372, new_n373, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n580, new_n581, new_n583, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n940, new_n941, new_n942,
    new_n943;
  assign new_n299 = p_651_195_ & p_543_192_;
  assign new_n300 = p_77_58_ & new_n299;
  assign new_n301 = ~p_651_195_ & p_543_192_;
  assign new_n302 = p_52_37_ & new_n301;
  assign new_n303 = p_651_195_ & ~p_543_192_;
  assign new_n304 = p_64_47_ & new_n303;
  assign new_n305 = ~p_651_195_ & ~p_543_192_;
  assign new_n306 = p_90_69_ & new_n305;
  assign new_n307 = ~new_n300 & ~new_n302;
  assign new_n308 = ~new_n304 & new_n307;
  assign p_171_621_ = ~new_n306 & new_n308;
  assign new_n310 = p_868_198_ & ~p_171_621_;
  assign new_n311 = p_79_60_ & new_n299;
  assign new_n312 = p_54_39_ & new_n301;
  assign new_n313 = p_66_49_ & new_n303;
  assign new_n314 = p_92_71_ & new_n305;
  assign new_n315 = ~new_n311 & ~new_n312;
  assign new_n316 = ~new_n313 & new_n315;
  assign new_n317 = ~new_n314 & new_n316;
  assign new_n318 = ~p_868_198_ & ~new_n317;
  assign p_284_847_ = new_n310 | new_n318;
  assign new_n320 = p_80_61_ & new_n299;
  assign new_n321 = p_55_40_ & new_n301;
  assign new_n322 = p_67_50_ & new_n303;
  assign new_n323 = p_93_72_ & new_n305;
  assign new_n324 = ~new_n320 & ~new_n321;
  assign new_n325 = ~new_n322 & new_n324;
  assign new_n326 = ~new_n323 & new_n325;
  assign new_n327 = p_860_197_ & ~new_n326;
  assign new_n328 = p_68_51_ & new_n299;
  assign new_n329 = p_43_30_ & new_n301;
  assign new_n330 = p_56_41_ & new_n303;
  assign new_n331 = p_81_62_ & new_n305;
  assign new_n332 = ~new_n328 & ~new_n329;
  assign new_n333 = ~new_n330 & new_n332;
  assign new_n334 = ~new_n331 & new_n333;
  assign new_n335 = ~new_n317 & new_n334;
  assign new_n336 = new_n317 & ~new_n334;
  assign new_n337 = ~new_n335 & ~new_n336;
  assign new_n338 = ~p_559_193_ & new_n317;
  assign new_n339 = new_n337 & new_n338;
  assign new_n340 = ~new_n337 & ~new_n338;
  assign new_n341 = ~new_n339 & ~new_n340;
  assign new_n342 = ~new_n326 & new_n341;
  assign new_n343 = new_n326 & ~new_n341;
  assign new_n344 = ~new_n342 & ~new_n343;
  assign new_n345 = ~p_860_197_ & ~new_n344;
  assign p_145_1358_ = new_n327 | new_n345;
  assign new_n347 = p_2105_221_ & p_2104_220_;
  assign new_n348 = p_116_91_ & new_n347;
  assign new_n349 = ~p_2105_221_ & p_2104_220_;
  assign new_n350 = p_104_81_ & new_n349;
  assign new_n351 = p_2105_221_ & ~p_2104_220_;
  assign new_n352 = p_128_101_ & new_n351;
  assign new_n353 = ~p_2105_221_ & ~p_2104_220_;
  assign new_n354 = p_140_111_ & new_n353;
  assign new_n355 = ~new_n348 & ~new_n350;
  assign new_n356 = ~new_n352 & new_n355;
  assign new_n357 = ~new_n354 & new_n356;
  assign new_n358 = p_29_22_ & ~new_n357;
  assign new_n359 = ~p_29_22_ & p_26_19_;
  assign new_n360 = ~new_n358 & ~new_n359;
  assign new_n361 = ~p_2067_213_ & new_n360;
  assign new_n362 = p_2067_213_ & ~new_n360;
  assign new_n363 = ~new_n361 & ~new_n362;
  assign new_n364 = p_117_92_ & new_n347;
  assign new_n365 = p_105_82_ & new_n349;
  assign new_n366 = p_129_102_ & new_n351;
  assign new_n367 = p_141_112_ & new_n353;
  assign new_n368 = ~new_n364 & ~new_n365;
  assign new_n369 = ~new_n366 & new_n368;
  assign new_n370 = ~new_n367 & new_n369;
  assign new_n371 = p_29_22_ & ~new_n370;
  assign new_n372 = ~p_29_22_ & p_32_23_;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = ~p_1996_211_ & new_n373;
  assign new_n375 = p_1996_211_ & ~new_n373;
  assign new_n376 = ~new_n374 & ~new_n375;
  assign new_n377 = p_114_89_ & new_n347;
  assign new_n378 = p_102_79_ & new_n349;
  assign new_n379 = p_126_99_ & new_n351;
  assign new_n380 = p_138_109_ & new_n353;
  assign new_n381 = ~new_n377 & ~new_n378;
  assign new_n382 = ~new_n379 & new_n381;
  assign p_164_607_ = ~new_n380 & new_n382;
  assign new_n384 = p_29_22_ & ~p_164_607_;
  assign new_n385 = ~p_29_22_ & p_27_20_;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = ~p_2078_215_ & new_n386;
  assign new_n388 = p_2078_215_ & ~new_n386;
  assign new_n389 = ~new_n387 & ~new_n388;
  assign new_n390 = p_115_90_ & new_n347;
  assign new_n391 = p_103_80_ & new_n349;
  assign new_n392 = p_127_100_ & new_n351;
  assign new_n393 = p_139_110_ & new_n353;
  assign new_n394 = ~new_n390 & ~new_n391;
  assign new_n395 = ~new_n392 & new_n394;
  assign new_n396 = ~new_n393 & new_n395;
  assign new_n397 = p_29_22_ & ~new_n396;
  assign new_n398 = ~p_29_22_ & p_33_24_;
  assign new_n399 = ~new_n397 & ~new_n398;
  assign new_n400 = ~p_2072_214_ & new_n399;
  assign new_n401 = p_2072_214_ & ~new_n399;
  assign new_n402 = ~new_n400 & ~new_n401;
  assign new_n403 = p_113_88_ & new_n347;
  assign new_n404 = p_101_78_ & new_n349;
  assign new_n405 = p_125_98_ & new_n351;
  assign new_n406 = p_137_108_ & new_n353;
  assign new_n407 = ~new_n403 & ~new_n404;
  assign new_n408 = ~new_n405 & new_n407;
  assign p_160_609_ = ~new_n406 & new_n408;
  assign new_n410 = p_29_22_ & ~p_160_609_;
  assign new_n411 = ~p_29_22_ & p_34_25_;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign new_n413 = ~p_2084_216_ & new_n412;
  assign new_n414 = p_2084_216_ & ~new_n412;
  assign new_n415 = ~new_n413 & ~new_n414;
  assign new_n416 = new_n363 & new_n376;
  assign new_n417 = new_n389 & new_n416;
  assign new_n418 = new_n402 & new_n417;
  assign new_n419 = new_n415 & new_n418;
  assign new_n420 = p_112_87_ & new_n347;
  assign new_n421 = p_100_77_ & new_n349;
  assign new_n422 = p_124_97_ & new_n351;
  assign new_n423 = p_136_107_ & new_n353;
  assign new_n424 = ~new_n420 & ~new_n421;
  assign new_n425 = ~new_n422 & new_n424;
  assign p_162_612_ = ~new_n423 & new_n425;
  assign new_n427 = p_29_22_ & ~p_162_612_;
  assign new_n428 = ~p_29_22_ & p_35_26_;
  assign new_n429 = ~new_n427 & ~new_n428;
  assign new_n430 = ~p_2090_217_ & new_n429;
  assign new_n431 = p_2090_217_ & ~new_n429;
  assign new_n432 = ~new_n430 & ~new_n431;
  assign new_n433 = p_111_86_ & new_n347;
  assign new_n434 = p_99_76_ & new_n349;
  assign new_n435 = p_123_96_ & new_n351;
  assign new_n436 = p_135_106_ & new_n353;
  assign new_n437 = ~new_n433 & ~new_n434;
  assign new_n438 = ~new_n435 & new_n437;
  assign new_n439 = ~new_n436 & new_n438;
  assign new_n440 = p_29_22_ & ~new_n439;
  assign new_n441 = p_28_21_ & ~p_29_22_;
  assign new_n442 = ~new_n440 & ~new_n441;
  assign new_n443 = new_n432 & ~new_n442;
  assign new_n444 = new_n419 & new_n443;
  assign new_n445 = p_11_8_ & p_868_198_;
  assign new_n446 = p_11_8_ & ~p_868_198_;
  assign new_n447 = ~new_n445 & ~new_n446;
  assign new_n448 = p_16_11_ & ~new_n317;
  assign new_n449 = p_4_3_ & ~p_16_11_;
  assign new_n450 = ~new_n448 & ~new_n449;
  assign new_n451 = ~p_1348_201_ & new_n450;
  assign new_n452 = p_1348_201_ & ~new_n450;
  assign new_n453 = ~new_n451 & ~new_n452;
  assign new_n454 = p_16_11_ & ~new_n334;
  assign new_n455 = p_19_12_ & ~p_16_11_;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457 = ~p_1341_200_ & new_n456;
  assign new_n458 = p_1341_200_ & ~new_n456;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = p_16_11_ & ~p_171_621_;
  assign new_n461 = ~p_16_11_ & p_5_4_;
  assign new_n462 = ~new_n460 & ~new_n461;
  assign new_n463 = ~p_1961_204_ & new_n462;
  assign new_n464 = p_1961_204_ & ~new_n462;
  assign new_n465 = ~new_n463 & ~new_n464;
  assign new_n466 = p_78_59_ & new_n299;
  assign new_n467 = p_53_38_ & new_n301;
  assign new_n468 = p_65_48_ & new_n303;
  assign new_n469 = p_91_70_ & new_n305;
  assign new_n470 = ~new_n466 & ~new_n467;
  assign new_n471 = ~new_n468 & new_n470;
  assign p_299_692_ = new_n469 | ~new_n471;
  assign new_n473 = p_16_11_ & p_299_692_;
  assign new_n474 = ~p_16_11_ & p_20_13_;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = ~p_1956_203_ & new_n475;
  assign new_n477 = p_1956_203_ & ~new_n475;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = p_76_57_ & new_n299;
  assign new_n480 = p_51_36_ & new_n301;
  assign new_n481 = p_63_46_ & new_n303;
  assign new_n482 = p_89_68_ & new_n305;
  assign new_n483 = ~new_n479 & ~new_n480;
  assign new_n484 = ~new_n481 & new_n483;
  assign p_168_623_ = ~new_n482 & new_n484;
  assign new_n486 = p_16_11_ & ~p_168_623_;
  assign new_n487 = p_21_14_ & ~p_16_11_;
  assign new_n488 = ~new_n486 & ~new_n487;
  assign new_n489 = ~p_1966_205_ & new_n488;
  assign new_n490 = p_1966_205_ & ~new_n488;
  assign new_n491 = ~new_n489 & ~new_n490;
  assign new_n492 = new_n453 & new_n459;
  assign new_n493 = new_n465 & new_n492;
  assign new_n494 = new_n478 & new_n493;
  assign new_n495 = new_n491 & new_n494;
  assign new_n496 = p_74_55_ & new_n299;
  assign new_n497 = p_49_34_ & new_n301;
  assign new_n498 = p_87_66_ & new_n305;
  assign new_n499 = ~new_n496 & ~new_n497;
  assign new_n500 = ~new_n303 & new_n499;
  assign p_288_700_ = new_n498 | ~new_n500;
  assign new_n502 = p_16_11_ & p_288_700_;
  assign new_n503 = p_23_16_ & ~p_16_11_;
  assign new_n504 = ~new_n502 & ~new_n503;
  assign new_n505 = ~p_1976_207_ & new_n504;
  assign new_n506 = p_1976_207_ & ~new_n504;
  assign new_n507 = ~new_n505 & ~new_n506;
  assign new_n508 = p_75_56_ & new_n299;
  assign new_n509 = p_50_35_ & new_n301;
  assign new_n510 = p_62_45_ & new_n303;
  assign new_n511 = p_88_67_ & new_n305;
  assign new_n512 = ~new_n508 & ~new_n509;
  assign new_n513 = ~new_n510 & new_n512;
  assign p_166_625_ = ~new_n511 & new_n513;
  assign new_n515 = p_16_11_ & ~p_166_625_;
  assign new_n516 = p_22_15_ & ~p_16_11_;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = ~p_1971_206_ & new_n517;
  assign new_n519 = p_1971_206_ & ~new_n517;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = p_72_53_ & new_n299;
  assign new_n522 = p_47_32_ & new_n301;
  assign new_n523 = p_60_43_ & new_n303;
  assign new_n524 = p_85_64_ & new_n305;
  assign new_n525 = ~new_n521 & ~new_n522;
  assign new_n526 = ~new_n523 & new_n525;
  assign p_290_704_ = new_n524 | ~new_n526;
  assign new_n528 = p_16_11_ & p_290_704_;
  assign new_n529 = p_24_17_ & ~p_16_11_;
  assign new_n530 = ~new_n528 & ~new_n529;
  assign new_n531 = ~p_1986_209_ & new_n530;
  assign new_n532 = p_1986_209_ & ~new_n530;
  assign new_n533 = ~new_n531 & ~new_n532;
  assign new_n534 = p_73_54_ & new_n299;
  assign new_n535 = p_48_33_ & new_n301;
  assign new_n536 = p_61_44_ & new_n303;
  assign new_n537 = p_86_65_ & new_n305;
  assign new_n538 = ~new_n534 & ~new_n535;
  assign new_n539 = ~new_n536 & new_n538;
  assign p_305_702_ = new_n537 | ~new_n539;
  assign new_n541 = p_16_11_ & p_305_702_;
  assign new_n542 = ~p_16_11_ & p_6_5_;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign new_n544 = ~p_1981_208_ & new_n543;
  assign new_n545 = p_1981_208_ & ~new_n543;
  assign new_n546 = ~new_n544 & ~new_n545;
  assign new_n547 = p_107_84_ & new_n347;
  assign new_n548 = p_95_74_ & new_n349;
  assign new_n549 = p_119_94_ & new_n351;
  assign new_n550 = p_131_104_ & new_n353;
  assign new_n551 = ~new_n547 & ~new_n548;
  assign new_n552 = ~new_n549 & new_n551;
  assign new_n553 = ~new_n550 & new_n552;
  assign new_n554 = p_29_22_ & ~new_n553;
  assign new_n555 = p_25_18_ & ~p_29_22_;
  assign new_n556 = ~new_n554 & ~new_n555;
  assign new_n557 = ~p_1991_210_ & new_n556;
  assign new_n558 = p_1991_210_ & ~new_n556;
  assign new_n559 = ~new_n557 & ~new_n558;
  assign new_n560 = new_n507 & new_n520;
  assign new_n561 = new_n533 & new_n560;
  assign new_n562 = new_n546 & new_n561;
  assign new_n563 = new_n559 & new_n562;
  assign new_n564 = new_n495 & new_n563;
  assign new_n565 = new_n444 & ~new_n447;
  assign p_311_1278_ = new_n564 & new_n565;
  assign new_n567 = p_3_2_ & p_1_0_;
  assign new_n568 = p_69_52_ & p_57_42_;
  assign new_n569 = p_108_85_ & new_n568;
  assign new_n570 = p_120_95_ & new_n569;
  assign new_n571 = p_567_194_ & ~new_n570;
  assign new_n572 = p_44_31_ & p_82_63_;
  assign new_n573 = p_96_75_ & new_n572;
  assign new_n574 = p_132_105_ & new_n573;
  assign new_n575 = p_2106_222_ & ~new_n574;
  assign p_319_656_ = ~new_n571 & ~new_n575;
  assign new_n577 = p_483_191_ & ~new_n567;
  assign new_n578 = p_319_656_ & new_n577;
  assign p_188_761_ = ~p_661_196_ | ~new_n578;
  assign new_n580 = p_2084_216_ & p_2072_214_;
  assign new_n581 = p_2078_215_ & new_n580;
  assign p_158_349_ = ~p_2090_217_ | ~new_n581;
  assign new_n583 = p_661_196_ & p_15_10_;
  assign p_259_414_ = ~p_2_1_ | ~new_n583;
  assign p_325_507_ = new_n570 & new_n574;
  assign new_n586 = ~p_288_700_ & ~p_166_625_;
  assign new_n587 = p_288_700_ & p_166_625_;
  assign new_n588 = ~new_n586 & ~new_n587;
  assign new_n589 = ~p_290_704_ & p_305_702_;
  assign new_n590 = p_290_704_ & ~p_305_702_;
  assign new_n591 = ~new_n589 & ~new_n590;
  assign new_n592 = new_n588 & ~new_n591;
  assign new_n593 = ~new_n588 & new_n591;
  assign new_n594 = ~new_n592 & ~new_n593;
  assign new_n595 = ~new_n326 & new_n334;
  assign new_n596 = new_n326 & ~new_n334;
  assign new_n597 = ~new_n595 & ~new_n596;
  assign new_n598 = ~p_171_621_ & p_168_623_;
  assign new_n599 = p_171_621_ & ~p_168_623_;
  assign new_n600 = ~new_n598 & ~new_n599;
  assign new_n601 = ~new_n317 & ~p_299_692_;
  assign new_n602 = new_n317 & p_299_692_;
  assign new_n603 = ~new_n601 & ~new_n602;
  assign new_n604 = ~new_n597 & ~new_n600;
  assign new_n605 = ~new_n603 & new_n604;
  assign new_n606 = new_n600 & ~new_n603;
  assign new_n607 = new_n597 & new_n606;
  assign new_n608 = ~new_n605 & ~new_n607;
  assign new_n609 = new_n597 & ~new_n600;
  assign new_n610 = new_n603 & new_n609;
  assign new_n611 = new_n600 & new_n603;
  assign new_n612 = ~new_n597 & new_n611;
  assign new_n613 = ~new_n610 & ~new_n612;
  assign new_n614 = new_n608 & new_n613;
  assign new_n615 = new_n594 & ~new_n614;
  assign new_n616 = ~new_n594 & new_n614;
  assign new_n617 = ~new_n615 & ~new_n616;
  assign p_397_1406_ = ~p_37_28_ & new_n617;
  assign new_n619 = p_860_197_ & ~new_n317;
  assign new_n620 = ~p_860_197_ & ~new_n338;
  assign p_148_851_ = new_n619 | new_n620;
  assign new_n622 = ~p_1384_202_ & ~p_164_607_;
  assign new_n623 = p_40_29_ & new_n622;
  assign new_n624 = p_160_609_ & new_n623;
  assign new_n625 = ~p_1348_201_ & ~new_n624;
  assign new_n626 = ~p_2067_213_ & new_n624;
  assign new_n627 = ~new_n625 & ~new_n626;
  assign new_n628 = new_n317 & ~new_n627;
  assign new_n629 = ~p_1956_203_ & ~new_n624;
  assign new_n630 = ~p_2072_214_ & new_n624;
  assign new_n631 = ~new_n629 & ~new_n630;
  assign new_n632 = p_299_692_ & ~new_n631;
  assign new_n633 = ~p_299_692_ & new_n631;
  assign new_n634 = ~new_n632 & ~new_n633;
  assign new_n635 = new_n628 & ~new_n634;
  assign new_n636 = ~p_1341_200_ & ~new_n624;
  assign new_n637 = ~p_1996_211_ & new_n624;
  assign new_n638 = ~new_n636 & ~new_n637;
  assign new_n639 = new_n334 & ~new_n638;
  assign new_n640 = ~new_n317 & ~new_n627;
  assign new_n641 = new_n317 & new_n627;
  assign new_n642 = ~new_n640 & ~new_n641;
  assign new_n643 = ~new_n634 & new_n639;
  assign new_n644 = ~new_n642 & new_n643;
  assign new_n645 = ~p_299_692_ & ~new_n631;
  assign new_n646 = ~new_n635 & ~new_n644;
  assign new_n647 = ~new_n645 & new_n646;
  assign new_n648 = p_305_702_ & ~new_n624;
  assign new_n649 = p_8_7_ & new_n648;
  assign new_n650 = ~p_1981_208_ & ~new_n624;
  assign new_n651 = p_8_7_ & new_n650;
  assign new_n652 = new_n649 & new_n651;
  assign new_n653 = ~new_n649 & ~new_n651;
  assign new_n654 = ~new_n652 & ~new_n653;
  assign new_n655 = ~p_168_623_ & new_n624;
  assign new_n656 = ~p_168_623_ & ~new_n624;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign new_n658 = p_8_7_ & ~new_n657;
  assign new_n659 = ~p_1966_205_ & ~new_n624;
  assign new_n660 = ~p_2084_216_ & new_n624;
  assign new_n661 = ~new_n659 & ~new_n660;
  assign new_n662 = p_8_7_ & ~new_n661;
  assign new_n663 = new_n658 & new_n662;
  assign new_n664 = ~new_n658 & ~new_n662;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = ~p_1961_204_ & ~new_n624;
  assign new_n667 = ~p_2078_215_ & new_n624;
  assign new_n668 = ~new_n666 & ~new_n667;
  assign new_n669 = ~p_171_621_ & ~new_n668;
  assign new_n670 = p_171_621_ & new_n668;
  assign new_n671 = ~new_n669 & ~new_n670;
  assign new_n672 = ~p_166_625_ & new_n624;
  assign new_n673 = ~p_166_625_ & ~new_n624;
  assign new_n674 = ~new_n672 & ~new_n673;
  assign new_n675 = p_8_7_ & ~new_n674;
  assign new_n676 = ~p_1971_206_ & ~new_n624;
  assign new_n677 = ~p_2090_217_ & new_n624;
  assign new_n678 = ~new_n676 & ~new_n677;
  assign new_n679 = p_8_7_ & ~new_n678;
  assign new_n680 = new_n675 & new_n679;
  assign new_n681 = ~new_n675 & ~new_n679;
  assign new_n682 = ~new_n680 & ~new_n681;
  assign new_n683 = p_288_700_ & ~new_n624;
  assign new_n684 = p_8_7_ & new_n683;
  assign new_n685 = ~p_1976_207_ & ~new_n624;
  assign new_n686 = p_8_7_ & new_n685;
  assign new_n687 = new_n684 & new_n686;
  assign new_n688 = ~new_n684 & ~new_n686;
  assign new_n689 = ~new_n687 & ~new_n688;
  assign new_n690 = ~new_n654 & ~new_n665;
  assign new_n691 = ~new_n671 & new_n690;
  assign new_n692 = ~new_n682 & new_n691;
  assign new_n693 = ~new_n689 & new_n692;
  assign new_n694 = ~new_n647 & new_n693;
  assign new_n695 = ~new_n658 & new_n662;
  assign new_n696 = ~new_n654 & ~new_n689;
  assign new_n697 = new_n695 & new_n696;
  assign new_n698 = ~new_n682 & new_n697;
  assign new_n699 = p_171_621_ & ~new_n668;
  assign new_n700 = ~new_n689 & new_n699;
  assign new_n701 = ~new_n682 & new_n700;
  assign new_n702 = ~new_n654 & new_n701;
  assign new_n703 = ~new_n665 & new_n702;
  assign new_n704 = ~new_n684 & new_n686;
  assign new_n705 = ~new_n654 & new_n704;
  assign new_n706 = ~new_n675 & new_n679;
  assign new_n707 = ~new_n654 & new_n706;
  assign new_n708 = ~new_n689 & new_n707;
  assign new_n709 = ~new_n649 & new_n651;
  assign new_n710 = ~new_n698 & ~new_n703;
  assign new_n711 = ~new_n705 & new_n710;
  assign new_n712 = ~new_n708 & new_n711;
  assign new_n713 = ~new_n709 & new_n712;
  assign new_n714 = ~new_n694 & new_n713;
  assign new_n715 = p_160_609_ & ~new_n622;
  assign new_n716 = p_40_29_ & new_n715;
  assign new_n717 = ~new_n357 & ~new_n624;
  assign new_n718 = new_n716 & new_n717;
  assign new_n719 = ~p_2067_213_ & ~new_n624;
  assign new_n720 = new_n716 & new_n719;
  assign new_n721 = new_n718 & new_n720;
  assign new_n722 = ~new_n718 & ~new_n720;
  assign new_n723 = ~new_n721 & ~new_n722;
  assign new_n724 = p_290_704_ & ~new_n624;
  assign new_n725 = new_n716 & new_n724;
  assign new_n726 = ~p_1986_209_ & ~new_n624;
  assign new_n727 = new_n716 & new_n726;
  assign new_n728 = new_n725 & new_n727;
  assign new_n729 = ~new_n725 & ~new_n727;
  assign new_n730 = ~new_n728 & ~new_n729;
  assign new_n731 = ~new_n553 & ~new_n624;
  assign new_n732 = new_n716 & new_n731;
  assign new_n733 = ~p_1991_210_ & ~new_n624;
  assign new_n734 = new_n716 & new_n733;
  assign new_n735 = new_n732 & new_n734;
  assign new_n736 = ~new_n732 & ~new_n734;
  assign new_n737 = ~new_n735 & ~new_n736;
  assign new_n738 = ~new_n370 & ~new_n624;
  assign new_n739 = new_n716 & new_n738;
  assign new_n740 = ~p_1996_211_ & ~new_n624;
  assign new_n741 = new_n716 & new_n740;
  assign new_n742 = new_n739 & new_n741;
  assign new_n743 = ~new_n739 & ~new_n741;
  assign new_n744 = ~new_n742 & ~new_n743;
  assign new_n745 = ~new_n723 & ~new_n730;
  assign new_n746 = ~new_n737 & new_n745;
  assign new_n747 = ~new_n744 & new_n746;
  assign new_n748 = ~new_n725 & new_n727;
  assign new_n749 = ~new_n723 & ~new_n744;
  assign new_n750 = new_n748 & new_n749;
  assign new_n751 = ~new_n737 & new_n750;
  assign new_n752 = ~new_n739 & new_n741;
  assign new_n753 = ~new_n723 & new_n752;
  assign new_n754 = ~new_n732 & new_n734;
  assign new_n755 = ~new_n723 & new_n754;
  assign new_n756 = ~new_n744 & new_n755;
  assign new_n757 = ~new_n718 & new_n720;
  assign new_n758 = ~new_n751 & ~new_n753;
  assign new_n759 = ~new_n756 & new_n758;
  assign new_n760 = ~new_n757 & new_n759;
  assign new_n761 = ~new_n747 & new_n760;
  assign new_n762 = ~new_n714 & ~new_n761;
  assign new_n763 = new_n714 & ~new_n760;
  assign p_329_1414_ = new_n762 | new_n763;
  assign new_n765 = p_868_198_ & ~p_168_623_;
  assign new_n766 = ~p_868_198_ & p_299_692_;
  assign p_297_849_ = new_n765 | new_n766;
  assign new_n768 = ~p_2096_218_ & ~new_n439;
  assign new_n769 = ~new_n439 & ~new_n768;
  assign new_n770 = ~p_2096_218_ & ~new_n768;
  assign new_n771 = ~new_n769 & ~new_n770;
  assign new_n772 = ~new_n347 & ~new_n349;
  assign new_n773 = ~new_n351 & new_n772;
  assign new_n774 = ~new_n353 & new_n773;
  assign new_n775 = ~p_2100_219_ & ~new_n774;
  assign new_n776 = ~new_n774 & ~new_n775;
  assign new_n777 = ~p_2100_219_ & ~new_n775;
  assign new_n778 = ~new_n776 & ~new_n777;
  assign p_156_1046_ = ~new_n771 | ~new_n778;
  assign new_n780 = p_860_197_ & ~new_n334;
  assign p_153_671_ = ~p_860_197_ | new_n780;
  assign p_223_413_ = ~p_661_196_ | ~p_7_6_;
  assign new_n783 = ~new_n338 & ~new_n603;
  assign new_n784 = ~new_n597 & new_n783;
  assign new_n785 = ~new_n597 & new_n603;
  assign new_n786 = new_n338 & new_n785;
  assign new_n787 = ~new_n784 & ~new_n786;
  assign new_n788 = new_n338 & ~new_n603;
  assign new_n789 = new_n597 & new_n788;
  assign new_n790 = new_n597 & new_n603;
  assign new_n791 = ~new_n338 & new_n790;
  assign new_n792 = ~new_n789 & ~new_n791;
  assign new_n793 = new_n787 & new_n792;
  assign new_n794 = new_n594 & ~new_n793;
  assign new_n795 = ~new_n594 & new_n793;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = p_868_198_ & ~new_n796;
  assign new_n798 = ~p_868_198_ & ~new_n326;
  assign p_331_1401_ = new_n797 | new_n798;
  assign new_n800 = p_160_609_ & ~p_162_612_;
  assign new_n801 = ~p_160_609_ & p_162_612_;
  assign new_n802 = ~new_n800 & ~new_n801;
  assign new_n803 = new_n439 & ~new_n774;
  assign new_n804 = ~new_n439 & new_n774;
  assign new_n805 = ~new_n803 & ~new_n804;
  assign new_n806 = new_n802 & ~new_n805;
  assign new_n807 = ~new_n802 & new_n805;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = p_118_93_ & new_n347;
  assign new_n810 = p_106_83_ & new_n349;
  assign new_n811 = p_130_103_ & new_n351;
  assign new_n812 = p_142_113_ & new_n353;
  assign new_n813 = ~new_n809 & ~new_n810;
  assign new_n814 = ~new_n811 & new_n813;
  assign new_n815 = ~new_n812 & new_n814;
  assign new_n816 = ~new_n553 & new_n815;
  assign new_n817 = new_n553 & ~new_n815;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = ~p_164_607_ & new_n396;
  assign new_n820 = p_164_607_ & ~new_n396;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = ~new_n357 & new_n370;
  assign new_n823 = new_n357 & ~new_n370;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = ~new_n818 & ~new_n821;
  assign new_n826 = ~new_n824 & new_n825;
  assign new_n827 = new_n821 & ~new_n824;
  assign new_n828 = new_n818 & new_n827;
  assign new_n829 = ~new_n826 & ~new_n828;
  assign new_n830 = new_n818 & ~new_n821;
  assign new_n831 = new_n824 & new_n830;
  assign new_n832 = new_n821 & new_n824;
  assign new_n833 = ~new_n818 & new_n832;
  assign new_n834 = ~new_n831 & ~new_n833;
  assign new_n835 = new_n829 & new_n834;
  assign new_n836 = new_n808 & ~new_n835;
  assign new_n837 = ~new_n808 & new_n835;
  assign new_n838 = ~new_n836 & ~new_n837;
  assign p_395_1392_ = ~p_37_28_ & new_n838;
  assign new_n840 = p_868_198_ & ~new_n338;
  assign new_n841 = ~p_868_198_ & ~new_n334;
  assign p_282_922_ = new_n840 | new_n841;
  assign p_173_389_ = p_94_73_ & p_452_190_;
  assign p_217_423_ = ~p_2106_222_ | p_223_413_;
  assign new_n845 = p_1986_209_ & ~p_1981_208_;
  assign new_n846 = ~p_1986_209_ & p_1981_208_;
  assign new_n847 = ~new_n845 & ~new_n846;
  assign new_n848 = p_1996_211_ & ~p_1991_210_;
  assign new_n849 = ~p_1996_211_ & p_1991_210_;
  assign new_n850 = ~new_n848 & ~new_n849;
  assign new_n851 = new_n847 & ~new_n850;
  assign new_n852 = ~new_n847 & new_n850;
  assign new_n853 = ~new_n851 & ~new_n852;
  assign new_n854 = ~p_2474_231_ & p_1956_203_;
  assign new_n855 = p_2474_231_ & ~p_1956_203_;
  assign new_n856 = ~new_n854 & ~new_n855;
  assign new_n857 = p_1976_207_ & ~p_1971_206_;
  assign new_n858 = ~p_1976_207_ & p_1971_206_;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = ~p_1961_204_ & p_1966_205_;
  assign new_n861 = p_1961_204_ & ~p_1966_205_;
  assign new_n862 = ~new_n860 & ~new_n861;
  assign new_n863 = ~new_n856 & ~new_n859;
  assign new_n864 = ~new_n862 & new_n863;
  assign new_n865 = new_n859 & ~new_n862;
  assign new_n866 = new_n856 & new_n865;
  assign new_n867 = ~new_n864 & ~new_n866;
  assign new_n868 = new_n856 & ~new_n859;
  assign new_n869 = new_n862 & new_n868;
  assign new_n870 = new_n859 & new_n862;
  assign new_n871 = ~new_n856 & new_n870;
  assign new_n872 = ~new_n869 & ~new_n871;
  assign new_n873 = new_n867 & new_n872;
  assign new_n874 = new_n853 & ~new_n873;
  assign new_n875 = ~new_n853 & new_n873;
  assign p_229_1180_ = ~new_n874 & ~new_n875;
  assign new_n877 = ~p_2096_218_ & p_2100_219_;
  assign new_n878 = p_2096_218_ & ~p_2100_219_;
  assign new_n879 = ~new_n877 & ~new_n878;
  assign new_n880 = ~p_2678_232_ & p_2067_213_;
  assign new_n881 = p_2678_232_ & ~p_2067_213_;
  assign new_n882 = ~new_n880 & ~new_n881;
  assign new_n883 = p_2090_217_ & ~p_2084_216_;
  assign new_n884 = ~p_2090_217_ & p_2084_216_;
  assign new_n885 = ~new_n883 & ~new_n884;
  assign new_n886 = p_2078_215_ & ~p_2072_214_;
  assign new_n887 = ~p_2078_215_ & p_2072_214_;
  assign new_n888 = ~new_n886 & ~new_n887;
  assign new_n889 = ~new_n882 & ~new_n885;
  assign new_n890 = ~new_n888 & new_n889;
  assign new_n891 = new_n885 & ~new_n888;
  assign new_n892 = new_n882 & new_n891;
  assign new_n893 = ~new_n890 & ~new_n892;
  assign new_n894 = new_n882 & ~new_n885;
  assign new_n895 = new_n888 & new_n894;
  assign new_n896 = new_n885 & new_n888;
  assign new_n897 = ~new_n882 & new_n896;
  assign new_n898 = ~new_n895 & ~new_n897;
  assign new_n899 = new_n893 & new_n898;
  assign new_n900 = new_n879 & ~new_n899;
  assign new_n901 = ~new_n879 & new_n899;
  assign p_227_1179_ = ~new_n900 & ~new_n901;
  assign new_n903 = p_483_191_ & p_319_656_;
  assign new_n904 = p_36_27_ & new_n903;
  assign p_176_803_ = ~p_661_196_ | ~new_n904;
  assign new_n906 = ~p_2454_230_ & p_2451_229_;
  assign new_n907 = p_2454_230_ & ~p_2451_229_;
  assign new_n908 = ~new_n906 & ~new_n907;
  assign new_n909 = ~p_1341_200_ & p_1348_201_;
  assign new_n910 = p_1341_200_ & ~p_1348_201_;
  assign new_n911 = ~new_n909 & ~new_n910;
  assign new_n912 = new_n908 & ~new_n911;
  assign new_n913 = ~new_n908 & new_n911;
  assign new_n914 = ~new_n912 & ~new_n913;
  assign new_n915 = ~p_2430_224_ & p_2427_223_;
  assign new_n916 = p_2430_224_ & ~p_2427_223_;
  assign new_n917 = ~new_n915 & ~new_n916;
  assign new_n918 = p_2443_227_ & ~p_2446_228_;
  assign new_n919 = ~p_2443_227_ & p_2446_228_;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = p_2435_225_ & ~p_2438_226_;
  assign new_n922 = ~p_2435_225_ & p_2438_226_;
  assign new_n923 = ~new_n921 & ~new_n922;
  assign new_n924 = ~new_n917 & ~new_n920;
  assign new_n925 = ~new_n923 & new_n924;
  assign new_n926 = new_n920 & ~new_n923;
  assign new_n927 = new_n917 & new_n926;
  assign new_n928 = ~new_n925 & ~new_n927;
  assign new_n929 = new_n917 & ~new_n920;
  assign new_n930 = new_n923 & new_n929;
  assign new_n931 = new_n920 & new_n923;
  assign new_n932 = ~new_n917 & new_n931;
  assign new_n933 = ~new_n930 & ~new_n932;
  assign new_n934 = new_n928 & new_n933;
  assign new_n935 = new_n914 & ~new_n934;
  assign new_n936 = ~new_n914 & new_n934;
  assign new_n937 = ~new_n935 & ~new_n936;
  assign p_401_1276_ = p_14_9_ & new_n937;
  assign p_234_376_ = ~p_567_194_ | p_223_413_;
  assign new_n940 = ~p_229_1180_ & ~p_401_1276_;
  assign new_n941 = ~p_397_1406_ & ~p_227_1179_;
  assign new_n942 = ~p_395_1392_ & new_n941;
  assign new_n943 = p_319_656_ & new_n940;
  assign p_308_1425_ = new_n942 & new_n943;
  assign p_231_1422_ = 1'b0;
  assign p_150_1277_ = ~p_311_1278_;
  assign p_221_305_ = ~p_96_75_;
  assign p_235_307_ = ~p_69_52_;
  assign p_301_694_ = ~p_171_621_;
  assign p_218_311_ = ~p_44_31_;
  assign p_261_506_ = ~p_325_507_;
  assign p_236_303_ = ~p_120_95_;
  assign p_220_306_ = ~p_82_63_;
  assign p_303_698_ = ~p_166_625_;
  assign p_237_309_ = ~p_57_42_;
  assign p_286_696_ = ~p_168_623_;
  assign p_238_304_ = ~p_108_85_;
  assign p_219_302_ = ~p_132_105_;
  assign p_225_1424_ = ~p_308_1425_;
  assign p_367_288_ = p_1083_199_;
  assign p_384_262_ = p_2066_212_;
  assign p_321_848_ = p_284_847_;
  assign p_350_301_ = p_452_190_;
  assign p_369_289_ = p_1083_199_;
  assign p_411_264_ = p_2066_212_;
  assign p_337_263_ = p_2066_212_;
  assign p_391_379_ = p_452_190_;
  assign p_280_850_ = p_297_849_;
  assign p_335_299_ = p_452_190_;
  assign p_295_1400_ = p_331_1401_;
  assign p_323_923_ = p_282_922_;
  assign p_409_298_ = p_452_190_;
endmodule


