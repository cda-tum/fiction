// Benchmark "b05" written by ABC on Wed Sep  5 10:17:19 2018

module b05 ( clock, 
    START,
    U646, U792, U590, U589, U589, U590, U590, U590, U661, U662, U663, U664,
    U665, U666, U667, U647, U648, U649, U650, U651, U652, U653, U792, U591,
    U589, U589, U591, U591, U591, U654, U655, U656, U657, U658, U659, U660  );
  input  clock;
  input  START;
  output U646, U792, U590, U589, U589, U590, U590, U590, U661, U662, U663,
    U664, U665, U666, U667, U647, U648, U649, U650, U651, U652, U653, U792,
    U591, U589, U589, U591, U591, U591, U654, U655, U656, U657, U658, U659,
    U660;
  reg NUM_REG_4_, NUM_REG_3_, NUM_REG_2_, NUM_REG_1_, NUM_REG_0_,
    MAR_REG_4_, MAR_REG_3_, MAR_REG_2_, MAR_REG_1_, MAR_REG_0_,
    TEMP_REG_8_, TEMP_REG_7_, TEMP_REG_6_, TEMP_REG_5_, TEMP_REG_4_,
    TEMP_REG_3_, TEMP_REG_2_, TEMP_REG_1_, TEMP_REG_0_, MAX_REG_8_,
    MAX_REG_7_, MAX_REG_6_, MAX_REG_5_, MAX_REG_4_, MAX_REG_3_, MAX_REG_2_,
    MAX_REG_1_, MAX_REG_0_, EN_DISP_REG, RES_DISP_REG, FLAG_REG,
    STATO_REG_0_, STATO_REG_1_, STATO_REG_2_;
  wire n141_1, n144, n145, n146_1, n147, n148, n149, n150, n151_1, n152,
    n153, n154, n155, n156_1, n157, n158, n159, n160, n161_1, n162, n163,
    n164, n165, n166_1, n167, n168, n170, n171_1, n172, n173, n174, n175,
    n176_1, n177, n178, n179, n180, n181_1, n182, n183, n184, n185, n186_1,
    n187, n188, n189, n190, n191_1, n192, n193, n194, n195, n196_1, n197,
    n198, n199, n200, n201_1, n202, n203, n204, n205, n206_1, n207, n208,
    n209, n210, n211_1, n212, n213, n214, n215, n216_1, n217, n218, n219,
    n220, n221_1, n222, n223, n224, n225, n226_1, n227, n228, n229, n230,
    n231_1, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n283, n284, n285, n286, n287, n289, n291, n292, n294,
    n295, n296, n297, n299, n300, n301, n302, n303, n304, n305, n306, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n485, n486, n487, n488, n489, n491,
    n493, n494, n496, n497, n498, n499, n501, n502, n503, n504, n505, n506,
    n507, n508, n510, n511, n512, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n569,
    n570, n571, n572, n573, n574, n575, n576, n578, n579, n580, n581, n582,
    n584, n586, n587, n588, n590, n591, n592, n593, n595, n596, n597, n598,
    n599, n600, n601, n602, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n752, n753, n754, n755, n756,
    n758, n759, n760, n761, n762, n764, n765, n766, n767, n768, n770, n771,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n786, n787, n788, n789, n790, n792, n793, n794, n795, n796, n798, n799,
    n800, n801, n802, n804, n805, n807, n808, n810, n811, n813, n814, n816,
    n817, n818, n819, n820, n821, n823, n824, n826, n827, n828, n830, n831,
    n833, n834, n836, n837, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n923, n924, n926, n927, n929, n930, n932, n933, n935,
    n936, n938, n939, n941, n942, n944, n945, n947, n948, n949, n950, n951,
    n952, n953, n955, n956, n957, n959, n960, n961, n963, n964, n965, n966,
    n967, n970, n66, n71, n76, n81, n86, n91, n96, n101, n106, n111, n116,
    n121, n126, n131, n136, n141, n146, n151, n156, n161, n166, n171, n176,
    n181, n186, n191, n196, n201, n206, n211, n216, n221, n226, n231;
  assign U792 = ~EN_DISP_REG & ~RES_DISP_REG;
  assign n141_1 = MAX_REG_8_ & ~EN_DISP_REG;
  assign U646 = U792 | n141_1;
  assign U589 = ~EN_DISP_REG & RES_DISP_REG;
  assign n144 = ~MAX_REG_1_ & ~MAX_REG_0_;
  assign n145 = ~MAX_REG_2_ & n144;
  assign n146_1 = ~MAX_REG_3_ & n145;
  assign n147 = ~MAX_REG_4_ & n146_1;
  assign n148 = MAX_REG_8_ & ~n147;
  assign n149 = MAX_REG_2_ & ~n144;
  assign n150 = ~n145 & ~n149;
  assign n151_1 = MAX_REG_8_ & n150;
  assign n152 = ~MAX_REG_8_ & MAX_REG_2_;
  assign n153 = ~n151_1 & ~n152;
  assign n154 = MAX_REG_3_ & ~n145;
  assign n155 = ~n146_1 & ~n154;
  assign n156_1 = MAX_REG_8_ & n155;
  assign n157 = ~MAX_REG_8_ & MAX_REG_3_;
  assign n158 = ~n156_1 & ~n157;
  assign n159 = MAX_REG_4_ & ~n146_1;
  assign n160 = ~n147 & ~n159;
  assign n161_1 = MAX_REG_8_ & n160;
  assign n162 = ~MAX_REG_8_ & MAX_REG_4_;
  assign n163 = ~n161_1 & ~n162;
  assign n164 = n153 & n158;
  assign n165 = n163 & n164;
  assign n166_1 = n148 & ~n165;
  assign n167 = ~n148 & ~n166_1;
  assign n168 = ~n148 & ~n167;
  assign U590 = U589 & ~n168;
  assign n170 = n148 & ~n168;
  assign n171_1 = n148 & n166_1;
  assign n172 = ~n148 & ~n171_1;
  assign n173 = ~n148 & n172;
  assign n174 = n148 & ~n172;
  assign n175 = ~n173 & ~n174;
  assign n176_1 = n168 & ~n175;
  assign n177 = ~n170 & ~n176_1;
  assign n178 = ~n148 & n166_1;
  assign n179 = n148 & ~n166_1;
  assign n180 = ~n178 & ~n179;
  assign n181_1 = n168 & ~n180;
  assign n182 = ~n170 & ~n181_1;
  assign n183 = ~n153 & ~n158;
  assign n184 = ~n164 & ~n183;
  assign n185 = n168 & ~n184;
  assign n186_1 = ~n158 & ~n168;
  assign n187 = ~n185 & ~n186_1;
  assign n188 = ~n163 & ~n164;
  assign n189 = ~n165 & ~n188;
  assign n190 = n168 & ~n189;
  assign n191_1 = ~n163 & ~n168;
  assign n192 = ~n190 & ~n191_1;
  assign n193 = n153 & n168;
  assign n194 = ~n153 & ~n168;
  assign n195 = ~n193 & ~n194;
  assign n196_1 = ~MAX_REG_1_ & MAX_REG_0_;
  assign n197 = MAX_REG_1_ & ~MAX_REG_0_;
  assign n198 = ~n196_1 & ~n197;
  assign n199 = MAX_REG_8_ & ~n198;
  assign n200 = ~MAX_REG_8_ & MAX_REG_1_;
  assign n201_1 = ~n199 & ~n200;
  assign n202 = n168 & ~n201_1;
  assign n203 = ~n168 & ~n201_1;
  assign n204 = ~n202 & ~n203;
  assign n205 = n195 & n204;
  assign n206_1 = ~n187 & ~n192;
  assign n207 = ~n205 & n206_1;
  assign n208 = ~n148 & n165;
  assign n209 = ~n166_1 & ~n208;
  assign n210 = n168 & n209;
  assign n211_1 = ~n170 & ~n210;
  assign n212 = ~n207 & n211_1;
  assign n213 = ~n182 & ~n212;
  assign n214 = ~n148 & n171_1;
  assign n215 = n148 & ~n171_1;
  assign n216_1 = ~n214 & ~n215;
  assign n217 = n168 & n216_1;
  assign n218 = ~n170 & ~n217;
  assign n219 = ~n213 & n218;
  assign n220 = n177 & ~n219;
  assign n221_1 = n192 & n211_1;
  assign n222 = ~n182 & ~n221_1;
  assign n223 = n218 & ~n222;
  assign n224 = n177 & ~n223;
  assign n225 = ~n220 & ~n224;
  assign n226_1 = n187 & n195;
  assign n227 = n204 & n226_1;
  assign n228 = ~n192 & ~n211_1;
  assign n229 = ~n227 & n228;
  assign n230 = n218 & ~n229;
  assign n231_1 = n182 & n230;
  assign n232 = n177 & ~n231_1;
  assign n233 = ~n195 & ~n211_1;
  assign n234 = ~n187 & n233;
  assign n235 = ~n192 & n234;
  assign n236 = n218 & ~n235;
  assign n237 = n182 & n236;
  assign n238 = n177 & ~n237;
  assign n239 = ~n232 & ~n238;
  assign n240 = ~n195 & ~n204;
  assign n241 = n187 & ~n240;
  assign n242 = n192 & n241;
  assign n243 = n211_1 & n242;
  assign n244 = ~n182 & ~n243;
  assign n245 = n218 & ~n244;
  assign n246 = n177 & ~n245;
  assign n247 = ~n239 & ~n246;
  assign n248 = n225 & ~n247;
  assign n249 = ~n187 & ~n195;
  assign n250 = ~n192 & n249;
  assign n251 = ~n204 & n250;
  assign n252 = n211_1 & n218;
  assign n253 = n182 & n252;
  assign n254 = ~n251 & n253;
  assign n255 = n177 & ~n254;
  assign n256 = ~n192 & ~n226_1;
  assign n257 = n182 & n218;
  assign n258 = n211_1 & n257;
  assign n259 = ~n256 & n258;
  assign n260 = n177 & ~n259;
  assign n261 = n187 & n192;
  assign n262 = ~n211_1 & ~n261;
  assign n263 = n218 & ~n262;
  assign n264 = n182 & n263;
  assign n265 = n177 & ~n264;
  assign n266 = ~n255 & ~n260;
  assign n267 = ~n265 & n266;
  assign n268 = ~n246 & ~n267;
  assign n269 = RES_DISP_REG & n248;
  assign n270 = ~n268 & n269;
  assign U661 = ~EN_DISP_REG & ~n270;
  assign n272 = ~n187 & ~n205;
  assign n273 = n257 & ~n272;
  assign n274 = n211_1 & n273;
  assign n275 = n192 & n274;
  assign n276 = n177 & ~n275;
  assign n277 = ~n260 & n276;
  assign n278 = ~n255 & n277;
  assign n279 = ~n246 & ~n265;
  assign n280 = ~n278 & n279;
  assign n281 = n248 & ~n280;
  assign U662 = U589 & ~n281;
  assign n283 = n225 & ~n246;
  assign n284 = n239 & n283;
  assign n285 = ~n255 & ~n265;
  assign n286 = n260 & n285;
  assign n287 = n284 & n286;
  assign U663 = U589 & ~n287;
  assign n289 = ~n239 & n283;
  assign U664 = U589 & ~n289;
  assign n291 = ~n277 & n285;
  assign n292 = n284 & ~n291;
  assign U665 = U589 & ~n292;
  assign n294 = n266 & ~n276;
  assign n295 = ~n265 & ~n294;
  assign n296 = ~n246 & ~n295;
  assign n297 = n248 & ~n296;
  assign U666 = U589 & ~n297;
  assign n299 = ~n260 & ~n276;
  assign n300 = ~n255 & ~n299;
  assign n301 = ~n232 & ~n265;
  assign n302 = ~n300 & n301;
  assign n303 = ~n238 & ~n302;
  assign n304 = ~n246 & ~n303;
  assign n305 = ~n224 & ~n304;
  assign n306 = U589 & ~n220;
  assign U667 = ~n305 & n306;
  assign n308 = ~n182 & n283;
  assign n309 = n182 & ~n283;
  assign n310 = n238 & n283;
  assign n311 = n232 & ~n238;
  assign n312 = n283 & n311;
  assign n313 = n265 & n284;
  assign n314 = ~n310 & ~n312;
  assign n315 = ~n313 & n314;
  assign n316 = ~n211_1 & n315;
  assign n317 = n211_1 & ~n315;
  assign n318 = n255 & ~n265;
  assign n319 = n284 & n318;
  assign n320 = ~n287 & ~n310;
  assign n321 = ~n319 & n320;
  assign n322 = n225 & ~n312;
  assign n323 = n321 & n322;
  assign n324 = ~n192 & n323;
  assign n325 = n192 & ~n323;
  assign n326 = ~n224 & ~n246;
  assign n327 = n265 & n326;
  assign n328 = n239 & n327;
  assign n329 = n267 & n284;
  assign n330 = ~n220 & ~n319;
  assign n331 = ~n329 & n330;
  assign n332 = ~n310 & ~n328;
  assign n333 = n331 & n332;
  assign n334 = ~n187 & n333;
  assign n335 = n187 & ~n333;
  assign n336 = n225 & n246;
  assign n337 = n321 & ~n336;
  assign n338 = ~n195 & n337;
  assign n339 = n195 & ~n337;
  assign n340 = ~n224 & n246;
  assign n341 = ~n312 & ~n340;
  assign n342 = n331 & n341;
  assign n343 = n204 & ~n342;
  assign n344 = ~n339 & ~n343;
  assign n345 = ~n338 & ~n344;
  assign n346 = ~n335 & ~n345;
  assign n347 = ~n334 & ~n346;
  assign n348 = ~n325 & ~n347;
  assign n349 = ~n324 & ~n348;
  assign n350 = ~n317 & ~n349;
  assign n351 = ~n316 & ~n350;
  assign n352 = ~n309 & ~n351;
  assign n353 = ~n308 & ~n352;
  assign n354 = n218 & n353;
  assign n355 = n177 & n354;
  assign n356 = ~n177 & ~n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = n239 & ~n276;
  assign n359 = n267 & n358;
  assign n360 = n283 & n359;
  assign n361 = ~n357 & ~n360;
  assign n362 = ~n177 & n360;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n218 & ~n353;
  assign n365 = ~n354 & ~n364;
  assign n366 = ~n360 & ~n365;
  assign n367 = ~n218 & n360;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n308 & ~n309;
  assign n370 = ~n351 & ~n369;
  assign n371 = n351 & n369;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n360 & ~n372;
  assign n374 = ~n182 & n360;
  assign n375 = ~n373 & ~n374;
  assign n376 = MAX_REG_8_ & MAX_REG_0_;
  assign n377 = ~MAX_REG_8_ & MAX_REG_0_;
  assign n378 = ~n376 & ~n377;
  assign n379 = n168 & ~n378;
  assign n380 = ~n168 & ~n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = n360 & ~n381;
  assign n383 = ~n360 & ~n381;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n204 & n360;
  assign n386 = ~n204 & n342;
  assign n387 = ~n343 & ~n386;
  assign n388 = ~n360 & ~n387;
  assign n389 = ~n385 & ~n388;
  assign n390 = ~n384 & ~n389;
  assign n391 = ~n187 & n360;
  assign n392 = ~n334 & ~n335;
  assign n393 = ~n345 & ~n392;
  assign n394 = n345 & n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~n360 & ~n395;
  assign n397 = ~n391 & ~n396;
  assign n398 = ~n195 & n360;
  assign n399 = ~n338 & ~n339;
  assign n400 = ~n343 & ~n399;
  assign n401 = n343 & n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n360 & ~n402;
  assign n404 = ~n398 & ~n403;
  assign n405 = ~n192 & n360;
  assign n406 = ~n324 & ~n325;
  assign n407 = ~n347 & ~n406;
  assign n408 = n347 & n406;
  assign n409 = ~n407 & ~n408;
  assign n410 = ~n360 & ~n409;
  assign n411 = ~n405 & ~n410;
  assign n412 = ~n316 & ~n317;
  assign n413 = ~n349 & ~n412;
  assign n414 = n349 & n412;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~n360 & ~n415;
  assign n417 = ~n211_1 & n360;
  assign n418 = ~n416 & ~n417;
  assign n419 = n397 & n404;
  assign n420 = n411 & n419;
  assign n421 = n418 & n420;
  assign n422 = n368 & n375;
  assign n423 = ~n390 & n422;
  assign n424 = n421 & n423;
  assign n425 = n363 & ~n424;
  assign n426 = n389 & n397;
  assign n427 = n411 & n426;
  assign n428 = n404 & n427;
  assign n429 = n418 & n428;
  assign n430 = n368 & n429;
  assign n431 = n375 & n430;
  assign n432 = n363 & ~n431;
  assign n433 = ~n425 & ~n432;
  assign n434 = n390 & ~n404;
  assign n435 = n397 & n411;
  assign n436 = n418 & n435;
  assign n437 = n422 & ~n434;
  assign n438 = n436 & n437;
  assign n439 = n363 & ~n438;
  assign n440 = ~n433 & ~n439;
  assign n441 = n418 & n422;
  assign n442 = n411 & n441;
  assign n443 = n397 & n442;
  assign n444 = n363 & ~n443;
  assign n445 = n384 & n389;
  assign n446 = n404 & n445;
  assign n447 = ~n397 & ~n446;
  assign n448 = n422 & ~n447;
  assign n449 = n418 & n448;
  assign n450 = n411 & n449;
  assign n451 = n363 & ~n450;
  assign n452 = ~n389 & ~n404;
  assign n453 = n422 & ~n452;
  assign n454 = n436 & n453;
  assign n455 = n363 & ~n454;
  assign n456 = ~n404 & ~n445;
  assign n457 = n422 & ~n456;
  assign n458 = n436 & n457;
  assign n459 = n363 & ~n458;
  assign n460 = ~n455 & ~n459;
  assign n461 = ~n439 & ~n460;
  assign n462 = ~n444 & ~n451;
  assign n463 = ~n461 & n462;
  assign n464 = n404 & n435;
  assign n465 = n418 & n464;
  assign n466 = n375 & n465;
  assign n467 = n368 & n466;
  assign n468 = n363 & ~n467;
  assign n469 = ~n439 & n468;
  assign n470 = n463 & ~n469;
  assign n471 = RES_DISP_REG & ~n440;
  assign n472 = n470 & n471;
  assign U647 = ~EN_DISP_REG & ~n472;
  assign n474 = n397 & n446;
  assign n475 = n422 & n474;
  assign n476 = n411 & n475;
  assign n477 = n418 & n476;
  assign n478 = n363 & ~n477;
  assign n479 = ~n432 & n478;
  assign n480 = ~n425 & n479;
  assign n481 = ~n439 & ~n468;
  assign n482 = ~n480 & n481;
  assign n483 = n463 & ~n482;
  assign U648 = U589 & ~n483;
  assign n485 = ~n439 & n462;
  assign n486 = n460 & n485;
  assign n487 = ~n425 & ~n468;
  assign n488 = n432 & n487;
  assign n489 = n486 & n488;
  assign U649 = U589 & ~n489;
  assign n491 = ~n460 & n485;
  assign U650 = U589 & ~n491;
  assign n493 = ~n479 & n487;
  assign n494 = n486 & ~n493;
  assign U651 = U589 & ~n494;
  assign n496 = ~n439 & ~n478;
  assign n497 = ~n432 & n496;
  assign n498 = ~n425 & n497;
  assign n499 = n470 & ~n498;
  assign U652 = U589 & ~n499;
  assign n501 = ~n432 & ~n478;
  assign n502 = ~n425 & ~n501;
  assign n503 = ~n459 & ~n468;
  assign n504 = ~n502 & n503;
  assign n505 = ~n455 & ~n504;
  assign n506 = ~n439 & ~n505;
  assign n507 = ~n444 & ~n506;
  assign n508 = U589 & ~n451;
  assign U653 = ~n507 & n508;
  assign n510 = ~NUM_REG_2_ & ~NUM_REG_1_;
  assign n511 = NUM_REG_3_ & ~n510;
  assign n512 = ~NUM_REG_4_ & ~n511;
  assign U591 = U589 & n512;
  assign n514 = ~NUM_REG_3_ & ~NUM_REG_2_;
  assign n515 = ~NUM_REG_1_ & n514;
  assign n516 = ~n511 & ~n515;
  assign n517 = ~n512 & n516;
  assign n518 = NUM_REG_3_ & n512;
  assign n519 = ~n517 & ~n518;
  assign n520 = NUM_REG_4_ & n511;
  assign n521 = ~n512 & ~n520;
  assign n522 = ~n512 & ~n521;
  assign n523 = NUM_REG_4_ & n512;
  assign n524 = ~n522 & ~n523;
  assign n525 = n519 & n524;
  assign n526 = NUM_REG_0_ & ~n512;
  assign n527 = NUM_REG_0_ & n512;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~NUM_REG_1_ & ~n512;
  assign n530 = NUM_REG_1_ & n512;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n528 & ~n531;
  assign n533 = ~NUM_REG_2_ & NUM_REG_1_;
  assign n534 = NUM_REG_2_ & ~NUM_REG_1_;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~n512 & n535;
  assign n537 = NUM_REG_2_ & n512;
  assign n538 = ~n536 & ~n537;
  assign n539 = n525 & ~n532;
  assign n540 = n538 & n539;
  assign n541 = n524 & n531;
  assign n542 = n538 & n541;
  assign n543 = n519 & n542;
  assign n544 = n540 & n543;
  assign n545 = ~n531 & ~n538;
  assign n546 = ~n528 & n545;
  assign n547 = n525 & ~n546;
  assign n548 = ~n544 & n547;
  assign n549 = n528 & n538;
  assign n550 = n531 & n549;
  assign n551 = ~n519 & ~n550;
  assign n552 = n524 & ~n551;
  assign n553 = n525 & n552;
  assign n554 = n524 & ~n545;
  assign n555 = n519 & n554;
  assign n556 = n528 & n531;
  assign n557 = ~n538 & ~n556;
  assign n558 = n525 & ~n557;
  assign n559 = n555 & n558;
  assign n560 = n547 & ~n559;
  assign n561 = n553 & ~n560;
  assign n562 = n524 & n538;
  assign n563 = n519 & n562;
  assign n564 = n547 & ~n563;
  assign n565 = n561 & ~n564;
  assign n566 = RES_DISP_REG & ~n548;
  assign n567 = n565 & n566;
  assign U654 = ~EN_DISP_REG & ~n567;
  assign n569 = n538 & n556;
  assign n570 = n519 & n569;
  assign n571 = n524 & n570;
  assign n572 = n543 & ~n571;
  assign n573 = n540 & n572;
  assign n574 = n547 & n563;
  assign n575 = ~n573 & n574;
  assign n576 = n561 & ~n575;
  assign U655 = U589 & ~n576;
  assign n578 = n547 & n553;
  assign n579 = n559 & n578;
  assign n580 = ~n543 & n563;
  assign n581 = n540 & n580;
  assign n582 = n579 & n581;
  assign U656 = U589 & ~n582;
  assign n584 = ~n559 & n578;
  assign U657 = U589 & ~n584;
  assign n586 = n540 & n563;
  assign n587 = ~n572 & n586;
  assign n588 = n579 & ~n587;
  assign U658 = U589 & ~n588;
  assign n590 = n540 & n571;
  assign n591 = n543 & n590;
  assign n592 = n547 & n591;
  assign n593 = n565 & ~n592;
  assign U659 = U589 & ~n593;
  assign n595 = n543 & n571;
  assign n596 = n540 & ~n595;
  assign n597 = n558 & n563;
  assign n598 = ~n596 & n597;
  assign n599 = n555 & ~n598;
  assign n600 = n547 & ~n599;
  assign n601 = n525 & ~n600;
  assign n602 = U589 & n552;
  assign U660 = ~n601 & n602;
  assign n604 = ~START & ~STATO_REG_1_;
  assign n605 = ~MAR_REG_4_ & ~MAR_REG_0_;
  assign n606 = ~MAR_REG_2_ & n605;
  assign n607 = MAR_REG_3_ & MAR_REG_1_;
  assign n608 = MAR_REG_3_ & ~MAR_REG_1_;
  assign n609 = ~n607 & ~n608;
  assign n610 = n606 & ~n609;
  assign n611 = ~MAR_REG_3_ & MAR_REG_1_;
  assign n612 = ~MAR_REG_2_ & MAR_REG_0_;
  assign n613 = MAR_REG_4_ & n612;
  assign n614 = n611 & n613;
  assign n615 = ~MAR_REG_3_ & ~MAR_REG_1_;
  assign n616 = MAR_REG_2_ & n605;
  assign n617 = n615 & n616;
  assign n618 = ~MAR_REG_4_ & ~MAR_REG_2_;
  assign n619 = MAR_REG_0_ & n618;
  assign n620 = n607 & n619;
  assign n621 = ~MAR_REG_4_ & MAR_REG_2_;
  assign n622 = MAR_REG_0_ & n621;
  assign n623 = n607 & n622;
  assign n624 = MAR_REG_4_ & ~MAR_REG_0_;
  assign n625 = ~MAR_REG_2_ & n624;
  assign n626 = n615 & n625;
  assign n627 = n608 & n613;
  assign n628 = n607 & n613;
  assign n629 = ~n623 & ~n626;
  assign n630 = ~n627 & n629;
  assign n631 = ~n628 & n630;
  assign n632 = ~n617 & ~n620;
  assign n633 = n631 & n632;
  assign n634 = n608 & n619;
  assign n635 = MAR_REG_2_ & n624;
  assign n636 = ~n613 & ~n635;
  assign n637 = n615 & ~n636;
  assign n638 = ~n616 & ~n619;
  assign n639 = ~n625 & n638;
  assign n640 = n611 & ~n639;
  assign n641 = ~n634 & ~n637;
  assign n642 = ~n640 & n641;
  assign n643 = n611 & n622;
  assign n644 = ~n610 & ~n614;
  assign n645 = n633 & n644;
  assign n646 = n642 & n645;
  assign n647 = ~n643 & n646;
  assign n648 = TEMP_REG_7_ & n647;
  assign n649 = ~TEMP_REG_8_ & ~n633;
  assign n650 = TEMP_REG_8_ & n633;
  assign n651 = ~n649 & ~n650;
  assign n652 = n615 & n622;
  assign n653 = n608 & n625;
  assign n654 = ~n652 & ~n653;
  assign n655 = MAR_REG_2_ & MAR_REG_0_;
  assign n656 = MAR_REG_4_ & n655;
  assign n657 = n615 & n656;
  assign n658 = n642 & ~n657;
  assign n659 = n611 & n635;
  assign n660 = n654 & n658;
  assign n661 = ~n659 & n660;
  assign n662 = n633 & n661;
  assign n663 = ~TEMP_REG_6_ & ~n662;
  assign n664 = TEMP_REG_6_ & n662;
  assign n665 = n615 & n619;
  assign n666 = ~n659 & ~n665;
  assign n667 = ~n626 & n666;
  assign n668 = ~n628 & n667;
  assign n669 = n608 & n655;
  assign n670 = n668 & ~n669;
  assign n671 = n607 & n656;
  assign n672 = n606 & n615;
  assign n673 = ~n616 & ~n635;
  assign n674 = n607 & ~n673;
  assign n675 = ~n610 & ~n617;
  assign n676 = ~n671 & n675;
  assign n677 = ~n672 & n676;
  assign n678 = ~n674 & n677;
  assign n679 = ~n620 & ~n623;
  assign n680 = ~n643 & n679;
  assign n681 = n678 & n680;
  assign n682 = n658 & n681;
  assign n683 = n670 & n682;
  assign n684 = ~TEMP_REG_5_ & ~n683;
  assign n685 = TEMP_REG_5_ & n683;
  assign n686 = ~n643 & ~n659;
  assign n687 = ~n614 & n686;
  assign n688 = ~n620 & n687;
  assign n689 = n678 & n688;
  assign n690 = ~TEMP_REG_4_ & ~n689;
  assign n691 = TEMP_REG_4_ & n689;
  assign n692 = n611 & n656;
  assign n693 = n654 & ~n692;
  assign n694 = ~n627 & n693;
  assign n695 = ~n610 & n694;
  assign n696 = n670 & n695;
  assign n697 = ~TEMP_REG_3_ & ~n696;
  assign n698 = TEMP_REG_3_ & n696;
  assign n699 = ~n617 & ~n627;
  assign n700 = ~n626 & n699;
  assign n701 = n688 & n700;
  assign n702 = n658 & n701;
  assign n703 = ~TEMP_REG_2_ & ~n702;
  assign n704 = TEMP_REG_2_ & n702;
  assign n705 = ~n614 & ~n692;
  assign n706 = n631 & n705;
  assign n707 = n678 & n706;
  assign n708 = n654 & n707;
  assign n709 = n654 & n688;
  assign n710 = n642 & n709;
  assign n711 = ~n623 & n710;
  assign n712 = TEMP_REG_0_ & n711;
  assign n713 = ~n708 & ~n712;
  assign n714 = n708 & n712;
  assign n715 = ~TEMP_REG_1_ & ~n714;
  assign n716 = ~n713 & ~n715;
  assign n717 = ~n704 & ~n716;
  assign n718 = ~n703 & ~n717;
  assign n719 = ~n698 & ~n718;
  assign n720 = ~n697 & ~n719;
  assign n721 = ~n691 & ~n720;
  assign n722 = ~n690 & ~n721;
  assign n723 = ~n685 & ~n722;
  assign n724 = ~n684 & ~n723;
  assign n725 = ~n664 & ~n724;
  assign n726 = ~n663 & ~n725;
  assign n727 = ~TEMP_REG_7_ & ~n647;
  assign n728 = n726 & ~n727;
  assign n729 = ~n648 & ~n651;
  assign n730 = ~n728 & n729;
  assign n731 = ~n648 & ~n726;
  assign n732 = n651 & ~n727;
  assign n733 = ~n731 & n732;
  assign n734 = ~n730 & ~n733;
  assign n735 = STATO_REG_1_ & n734;
  assign n736 = STATO_REG_0_ & ~n604;
  assign n737 = ~n735 & n736;
  assign n738 = ~FLAG_REG & STATO_REG_1_;
  assign n739 = n737 & ~n738;
  assign n740 = NUM_REG_4_ & ~n739;
  assign n741 = NUM_REG_1_ & NUM_REG_0_;
  assign n742 = NUM_REG_2_ & n741;
  assign n743 = NUM_REG_3_ & n742;
  assign n744 = ~NUM_REG_4_ & n743;
  assign n745 = NUM_REG_4_ & ~n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = STATO_REG_0_ & STATO_REG_1_;
  assign n748 = FLAG_REG & n747;
  assign n749 = ~n734 & n748;
  assign n750 = ~n746 & n749;
  assign n66 = n740 | n750;
  assign n752 = NUM_REG_3_ & ~n739;
  assign n753 = ~NUM_REG_3_ & n742;
  assign n754 = NUM_REG_3_ & ~n742;
  assign n755 = ~n753 & ~n754;
  assign n756 = n749 & ~n755;
  assign n71 = n752 | n756;
  assign n758 = NUM_REG_2_ & ~n739;
  assign n759 = ~NUM_REG_2_ & n741;
  assign n760 = NUM_REG_2_ & ~n741;
  assign n761 = ~n759 & ~n760;
  assign n762 = n749 & ~n761;
  assign n76 = n758 | n762;
  assign n764 = NUM_REG_1_ & ~n739;
  assign n765 = ~NUM_REG_1_ & NUM_REG_0_;
  assign n766 = NUM_REG_1_ & ~NUM_REG_0_;
  assign n767 = ~n765 & ~n766;
  assign n768 = n749 & ~n767;
  assign n81 = n764 | n768;
  assign n770 = NUM_REG_0_ & ~n739;
  assign n771 = ~NUM_REG_0_ & n749;
  assign n86 = n770 | n771;
  assign n773 = STATO_REG_0_ & ~STATO_REG_1_;
  assign n774 = START & n773;
  assign n775 = STATO_REG_2_ & ~n671;
  assign n776 = ~n774 & ~n775;
  assign n777 = MAR_REG_4_ & n776;
  assign n778 = MAR_REG_1_ & MAR_REG_0_;
  assign n779 = MAR_REG_2_ & n778;
  assign n780 = MAR_REG_3_ & n779;
  assign n781 = ~MAR_REG_4_ & n780;
  assign n782 = MAR_REG_4_ & ~n780;
  assign n783 = ~n781 & ~n782;
  assign n784 = STATO_REG_2_ & ~n783;
  assign n91 = n777 | n784;
  assign n786 = MAR_REG_3_ & n776;
  assign n787 = ~MAR_REG_3_ & n779;
  assign n788 = MAR_REG_3_ & ~n779;
  assign n789 = ~n787 & ~n788;
  assign n790 = STATO_REG_2_ & ~n789;
  assign n96 = n786 | n790;
  assign n792 = MAR_REG_2_ & n776;
  assign n793 = ~MAR_REG_2_ & n778;
  assign n794 = MAR_REG_2_ & ~n778;
  assign n795 = ~n793 & ~n794;
  assign n796 = STATO_REG_2_ & ~n795;
  assign n101 = n792 | n796;
  assign n798 = MAR_REG_1_ & n776;
  assign n799 = ~MAR_REG_1_ & MAR_REG_0_;
  assign n800 = MAR_REG_1_ & ~MAR_REG_0_;
  assign n801 = ~n799 & ~n800;
  assign n802 = STATO_REG_2_ & ~n801;
  assign n106 = n798 | n802;
  assign n804 = MAR_REG_0_ & n776;
  assign n805 = ~MAR_REG_0_ & STATO_REG_2_;
  assign n111 = n804 | n805;
  assign n807 = STATO_REG_1_ & ~n633;
  assign n808 = TEMP_REG_8_ & ~STATO_REG_1_;
  assign n116 = n807 | n808;
  assign n810 = STATO_REG_1_ & ~n647;
  assign n811 = TEMP_REG_7_ & ~STATO_REG_1_;
  assign n121 = n810 | n811;
  assign n813 = STATO_REG_1_ & ~n662;
  assign n814 = TEMP_REG_6_ & ~STATO_REG_1_;
  assign n126 = n813 | n814;
  assign n816 = ~n622 & ~n656;
  assign n817 = n608 & ~n816;
  assign n818 = n668 & ~n817;
  assign n819 = n682 & n818;
  assign n820 = STATO_REG_1_ & ~n819;
  assign n821 = TEMP_REG_5_ & ~STATO_REG_1_;
  assign n131 = n820 | n821;
  assign n823 = STATO_REG_1_ & ~n689;
  assign n824 = TEMP_REG_4_ & ~STATO_REG_1_;
  assign n136 = n823 | n824;
  assign n826 = n695 & n818;
  assign n827 = STATO_REG_1_ & ~n826;
  assign n828 = TEMP_REG_3_ & ~STATO_REG_1_;
  assign n141 = n827 | n828;
  assign n830 = STATO_REG_1_ & ~n702;
  assign n831 = TEMP_REG_2_ & ~STATO_REG_1_;
  assign n146 = n830 | n831;
  assign n833 = STATO_REG_1_ & ~n708;
  assign n834 = TEMP_REG_1_ & ~STATO_REG_1_;
  assign n151 = n833 | n834;
  assign n836 = STATO_REG_1_ & ~n711;
  assign n837 = TEMP_REG_0_ & ~STATO_REG_1_;
  assign n156 = n836 | n837;
  assign n839 = ~STATO_REG_0_ & STATO_REG_1_;
  assign n840 = MAX_REG_7_ & n647;
  assign n841 = ~MAX_REG_8_ & ~n633;
  assign n842 = MAX_REG_8_ & n633;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~MAX_REG_6_ & ~n662;
  assign n845 = MAX_REG_4_ & n689;
  assign n846 = MAX_REG_5_ & n683;
  assign n847 = ~MAX_REG_4_ & ~n689;
  assign n848 = ~MAX_REG_3_ & ~n696;
  assign n849 = MAX_REG_2_ & n702;
  assign n850 = MAX_REG_3_ & n696;
  assign n851 = ~MAX_REG_1_ & ~n708;
  assign n852 = MAX_REG_0_ & n711;
  assign n853 = MAX_REG_1_ & n708;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~MAX_REG_2_ & ~n702;
  assign n856 = ~n851 & ~n854;
  assign n857 = ~n855 & n856;
  assign n858 = ~n849 & ~n850;
  assign n859 = ~n857 & n858;
  assign n860 = ~n847 & ~n848;
  assign n861 = ~n859 & n860;
  assign n862 = ~n845 & ~n846;
  assign n863 = ~n861 & n862;
  assign n864 = ~MAX_REG_5_ & ~n683;
  assign n865 = ~n863 & ~n864;
  assign n866 = MAX_REG_6_ & n662;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n844 & ~n867;
  assign n869 = ~MAX_REG_7_ & ~n647;
  assign n870 = n868 & ~n869;
  assign n871 = ~n840 & ~n843;
  assign n872 = ~n870 & n871;
  assign n873 = ~n840 & ~n868;
  assign n874 = n843 & ~n869;
  assign n875 = ~n873 & n874;
  assign n876 = ~n872 & ~n875;
  assign n877 = ~n684 & ~n685;
  assign n878 = ~n722 & ~n877;
  assign n879 = n722 & n877;
  assign n880 = ~n878 & ~n879;
  assign n881 = ~n690 & ~n691;
  assign n882 = ~n720 & ~n881;
  assign n883 = n720 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n648 & ~n727;
  assign n886 = ~n726 & ~n885;
  assign n887 = n726 & n885;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~TEMP_REG_1_ & ~n708;
  assign n890 = TEMP_REG_1_ & n708;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n712 & ~n891;
  assign n893 = n712 & n891;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~TEMP_REG_0_ & ~n711;
  assign n896 = ~n712 & ~n895;
  assign n897 = ~n703 & ~n704;
  assign n898 = ~n716 & ~n897;
  assign n899 = n716 & n897;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n697 & ~n698;
  assign n902 = ~n718 & ~n901;
  assign n903 = n718 & n901;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n663 & ~n664;
  assign n906 = ~n724 & ~n905;
  assign n907 = n724 & n905;
  assign n908 = ~n906 & ~n907;
  assign n909 = n894 & n896;
  assign n910 = n900 & n909;
  assign n911 = n904 & n910;
  assign n912 = n908 & n911;
  assign n913 = n880 & n884;
  assign n914 = n734 & n913;
  assign n915 = n888 & n914;
  assign n916 = n912 & n915;
  assign n917 = n735 & ~n876;
  assign n918 = ~n916 & n917;
  assign n919 = ~n839 & ~n918;
  assign n920 = ~n633 & ~n919;
  assign n921 = MAX_REG_8_ & n919;
  assign n161 = n920 | n921;
  assign n923 = ~n647 & ~n919;
  assign n924 = MAX_REG_7_ & n919;
  assign n166 = n923 | n924;
  assign n926 = ~n662 & ~n919;
  assign n927 = MAX_REG_6_ & n919;
  assign n171 = n926 | n927;
  assign n929 = ~n819 & ~n919;
  assign n930 = MAX_REG_5_ & n919;
  assign n176 = n929 | n930;
  assign n932 = ~n689 & ~n919;
  assign n933 = MAX_REG_4_ & n919;
  assign n181 = n932 | n933;
  assign n935 = ~n826 & ~n919;
  assign n936 = MAX_REG_3_ & n919;
  assign n186 = n935 | n936;
  assign n938 = ~n702 & ~n919;
  assign n939 = MAX_REG_2_ & n919;
  assign n191 = n938 | n939;
  assign n941 = ~n708 & ~n919;
  assign n942 = MAX_REG_1_ & n919;
  assign n196 = n941 | n942;
  assign n944 = ~n711 & ~n919;
  assign n945 = MAX_REG_0_ & n919;
  assign n201 = n944 | n945;
  assign n947 = STATO_REG_1_ & ~STATO_REG_2_;
  assign n948 = ~STATO_REG_0_ & ~n947;
  assign n949 = ~n775 & n948;
  assign n950 = EN_DISP_REG & ~n949;
  assign n951 = STATO_REG_2_ & n671;
  assign n952 = STATO_REG_0_ & n951;
  assign n953 = ~n774 & ~n950;
  assign n206 = n952 | ~n953;
  assign n955 = ~STATO_REG_1_ & ~STATO_REG_2_;
  assign n956 = ~STATO_REG_0_ & n955;
  assign n957 = RES_DISP_REG & ~n956;
  assign n211 = n774 | n957;
  assign n959 = FLAG_REG & ~n737;
  assign n960 = STATO_REG_0_ & n735;
  assign n961 = ~n916 & n960;
  assign n216 = n959 | n961;
  assign n963 = ~STATO_REG_0_ & ~STATO_REG_2_;
  assign n964 = STATO_REG_1_ & ~n951;
  assign n965 = ~START & ~n964;
  assign n966 = ~n839 & ~n963;
  assign n967 = ~n775 & n966;
  assign n221 = n965 | ~n967;
  assign n226 = ~n776 | n839;
  assign n970 = START & n951;
  assign n231 = n747 | n970;
  always @ (posedge clock) begin
    NUM_REG_4_ <= n66;
    NUM_REG_3_ <= n71;
    NUM_REG_2_ <= n76;
    NUM_REG_1_ <= n81;
    NUM_REG_0_ <= n86;
    MAR_REG_4_ <= n91;
    MAR_REG_3_ <= n96;
    MAR_REG_2_ <= n101;
    MAR_REG_1_ <= n106;
    MAR_REG_0_ <= n111;
    TEMP_REG_8_ <= n116;
    TEMP_REG_7_ <= n121;
    TEMP_REG_6_ <= n126;
    TEMP_REG_5_ <= n131;
    TEMP_REG_4_ <= n136;
    TEMP_REG_3_ <= n141;
    TEMP_REG_2_ <= n146;
    TEMP_REG_1_ <= n151;
    TEMP_REG_0_ <= n156;
    MAX_REG_8_ <= n161;
    MAX_REG_7_ <= n166;
    MAX_REG_6_ <= n171;
    MAX_REG_5_ <= n176;
    MAX_REG_4_ <= n181;
    MAX_REG_3_ <= n186;
    MAX_REG_2_ <= n191;
    MAX_REG_1_ <= n196;
    MAX_REG_0_ <= n201;
    EN_DISP_REG <= n206;
    RES_DISP_REG <= n211;
    FLAG_REG <= n216;
    STATO_REG_0_ <= n221;
    STATO_REG_1_ <= n226;
    STATO_REG_2_ <= n231;
  end
endmodule


