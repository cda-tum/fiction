// Benchmark "top" written by ABC on Mon Feb 19 11:52:45 2024

module top ( 
    pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1, pf4, pr,
    pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0, pf3,
    pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw, ph0,
    pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz, ph3,
    pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2, pm3,
    pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb, pp2,
    pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe, pt1,
    pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph, px0,
    py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1, pl,
    pm, pn, po,
    pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5  );
  input  pa1, pb2, pc3, pd4, pp, pa0, pb3, pc2, pe4, pq, pa3, pb0, pc1,
    pf4, pr, pa2, pb1, pc0, pg4, ps, pd0, pe1, pf2, pg3, pt, pa4, pd1, pe0,
    pf3, pg2, pu, pb4, pd2, pe3, pf0, pg1, pv, pc4, pd3, pe2, pf1, pg0, pw,
    ph0, pi1, pj2, pk3, px, ph1, pi0, pj3, pk2, py, ph2, pi3, pj0, pk1, pz,
    ph3, pi2, pj1, pk0, ph4, pl0, pm1, pn2, po3, pl1, pm0, pn3, po2, pl2,
    pm3, pn0, po1, pl3, pm2, pn1, po0, pq1, pr2, ps3, pp1, pr3, ps2, pb,
    pp2, pq3, pr0, ps1, pc, pp3, pq2, pr1, ps0, pd, pt0, pu1, pv2, pw3, pe,
    pt1, pu0, pv3, pw2, pf, pt2, pu3, pv0, pw1, pg, pt3, pu2, pv1, pw0, ph,
    px0, py1, pz2, pi, px1, py0, pz3, pj, px2, py3, pz0, pk, px3, py2, pz1,
    pl, pm, pn, po;
  output pe5, pf6, pg7, pd5, pf7, pg6, pd6, pe7, pg5, pd7, pe6, pf5, pa5, pb6,
    pc7, pb7, pc6, pa7, pc5, pa6, pb5, pl4, pm5, pn6, po7, pa8, pl5, pm4,
    pn7, po6, pb8, pl6, pm7, pn4, po5, pc8, pl7, pm6, pn5, po4, pi5, pj6,
    pk7, ph5, pi4, pj7, pk6, ph6, pi7, pj4, pk5, ph7, pi6, pj5, pk4, pt4,
    pu5, pv6, pw7, pt5, pu4, pv7, pw6, pt6, pu7, pv4, pw5, pt7, pu6, pv5,
    pw4, pp4, pq5, pr6, ps7, pp5, pq4, pr7, ps6, pp6, pq7, pr4, ps5, pp7,
    pq6, pr5, ps4, px4, py5, pz6, px5, py4, pz7, px6, py7, pz4, px7, py6,
    pz5;
  wire new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n391,
    new_n392, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n409, new_n410, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n525, new_n526, new_n527, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1389, new_n1390,
    new_n1391, new_n1392, new_n1393, new_n1394, new_n1395, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1410, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1451, new_n1452, new_n1453, new_n1454, new_n1455, new_n1456,
    new_n1457, new_n1459, new_n1460, new_n1461, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1516,
    new_n1517, new_n1518, new_n1519, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1525, new_n1526, new_n1527, new_n1528, new_n1529,
    new_n1530, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552;
  assign new_n235 = ~pb0 & ~pv;
  assign new_n236 = ps & new_n235;
  assign new_n237 = ~pv & ~pj1;
  assign new_n238 = pb0 & ~pj1;
  assign new_n239 = ~ps & ~pj1;
  assign new_n240 = ~new_n236 & ~new_n237;
  assign new_n241 = ~new_n238 & ~new_n239;
  assign new_n242 = new_n240 & new_n241;
  assign pe5 = ~py1 & new_n242;
  assign new_n244 = pl2 & ~pm2;
  assign new_n245 = pn2 & new_n244;
  assign new_n246 = ~pe0 & ~pf0;
  assign new_n247 = pg0 & new_n246;
  assign new_n248 = ~po2 & new_n245;
  assign new_n249 = new_n247 & new_n248;
  assign new_n250 = pp2 & new_n248;
  assign new_n251 = ~new_n249 & ~new_n250;
  assign new_n252 = ~pk2 & new_n251;
  assign new_n253 = pk2 & ~new_n251;
  assign new_n254 = ~px1 & new_n253;
  assign new_n255 = ~new_n252 & ~new_n254;
  assign new_n256 = ~py1 & new_n255;
  assign new_n257 = ~px1 & new_n256;
  assign new_n258 = pk2 & new_n256;
  assign pf6 = new_n257 | new_n258;
  assign new_n260 = ~pk1 & pe;
  assign new_n261 = ~pe & ~pu0;
  assign new_n262 = pd & new_n261;
  assign new_n263 = pc & ~pd;
  assign new_n264 = ~pe & new_n263;
  assign new_n265 = ~pv2 & new_n264;
  assign new_n266 = ~new_n260 & ~new_n262;
  assign new_n267 = ~new_n265 & new_n266;
  assign new_n268 = ~pd & ~pe;
  assign new_n269 = ~py1 & new_n267;
  assign new_n270 = ~new_n268 & new_n269;
  assign new_n271 = ~pk2 & pl3;
  assign new_n272 = ~pj2 & new_n271;
  assign new_n273 = pl3 & px1;
  assign new_n274 = ~new_n272 & ~new_n273;
  assign new_n275 = px1 & new_n274;
  assign new_n276 = ~pj2 & ~pk2;
  assign new_n277 = new_n274 & new_n276;
  assign new_n278 = ~pm3 & new_n274;
  assign new_n279 = ~new_n275 & ~new_n277;
  assign new_n280 = ~new_n278 & new_n279;
  assign new_n281 = new_n269 & new_n280;
  assign new_n282 = pc & new_n269;
  assign new_n283 = ~new_n270 & ~new_n281;
  assign pg7 = new_n282 | ~new_n283;
  assign new_n285 = ~pb0 & ~pu;
  assign new_n286 = ps & new_n285;
  assign new_n287 = ~pu & ~pi1;
  assign new_n288 = pb0 & ~pi1;
  assign new_n289 = ~ps & ~pi1;
  assign new_n290 = ~new_n286 & ~new_n287;
  assign new_n291 = ~new_n288 & ~new_n289;
  assign new_n292 = new_n290 & new_n291;
  assign pd5 = ~py1 & new_n292;
  assign new_n294 = ~pj1 & pe;
  assign new_n295 = ~pt0 & ~pe;
  assign new_n296 = pd & new_n295;
  assign new_n297 = ~pu2 & new_n264;
  assign new_n298 = ~new_n294 & ~new_n296;
  assign new_n299 = ~new_n297 & new_n298;
  assign new_n300 = ~py1 & new_n299;
  assign new_n301 = ~new_n268 & new_n300;
  assign new_n302 = pk3 & ~pk2;
  assign new_n303 = ~pj2 & new_n302;
  assign new_n304 = pk3 & px1;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = px1 & new_n305;
  assign new_n307 = new_n276 & new_n305;
  assign new_n308 = ~pl3 & new_n305;
  assign new_n309 = ~new_n306 & ~new_n307;
  assign new_n310 = ~new_n308 & new_n309;
  assign new_n311 = new_n300 & new_n310;
  assign new_n312 = pc & new_n300;
  assign new_n313 = ~new_n301 & ~new_n311;
  assign pf7 = new_n312 | ~new_n313;
  assign new_n315 = ~pc & ~pd;
  assign new_n316 = ~pe & new_n315;
  assign new_n317 = px1 & new_n316;
  assign new_n318 = ~pl2 & new_n317;
  assign new_n319 = ~pe & px1;
  assign new_n320 = ~pc & new_n319;
  assign new_n321 = ~pd & new_n320;
  assign new_n322 = ~py1 & ~new_n318;
  assign new_n323 = new_n321 & new_n322;
  assign new_n324 = ~pl2 & new_n322;
  assign pg6 = new_n323 | new_n324;
  assign new_n326 = po2 & new_n244;
  assign new_n327 = pp2 & new_n244;
  assign new_n328 = ~pg0 & new_n244;
  assign new_n329 = ~new_n326 & ~new_n327;
  assign new_n330 = ~new_n328 & new_n329;
  assign new_n331 = pn2 & ~new_n330;
  assign new_n332 = pj2 & new_n331;
  assign new_n333 = ~pp2 & new_n332;
  assign new_n334 = ~po2 & new_n331;
  assign new_n335 = ~new_n333 & ~new_n334;
  assign new_n336 = ~py1 & ~new_n335;
  assign new_n337 = ~px1 & new_n336;
  assign new_n338 = pi2 & ~py1;
  assign pd6 = new_n337 | new_n338;
  assign new_n340 = ~pi1 & pe;
  assign new_n341 = ~ps0 & ~pe;
  assign new_n342 = pd & new_n341;
  assign new_n343 = ~pt2 & new_n264;
  assign new_n344 = ~new_n340 & ~new_n342;
  assign new_n345 = ~new_n343 & new_n344;
  assign new_n346 = ~py1 & new_n345;
  assign new_n347 = ~new_n268 & new_n346;
  assign new_n348 = pj3 & ~pk2;
  assign new_n349 = ~pj2 & new_n348;
  assign new_n350 = pj3 & px1;
  assign new_n351 = ~new_n349 & ~new_n350;
  assign new_n352 = px1 & new_n351;
  assign new_n353 = new_n276 & new_n351;
  assign new_n354 = ~pk3 & new_n351;
  assign new_n355 = ~new_n352 & ~new_n353;
  assign new_n356 = ~new_n354 & new_n355;
  assign new_n357 = new_n346 & new_n356;
  assign new_n358 = pc & new_n346;
  assign new_n359 = ~new_n347 & ~new_n357;
  assign pe7 = new_n358 | ~new_n359;
  assign new_n361 = ~pb0 & ~px;
  assign new_n362 = ps & new_n361;
  assign new_n363 = ~px & ~pl1;
  assign new_n364 = pb0 & ~pl1;
  assign new_n365 = ~ps & ~pl1;
  assign new_n366 = ~new_n362 & ~new_n363;
  assign new_n367 = ~new_n364 & ~new_n365;
  assign new_n368 = new_n366 & new_n367;
  assign pg5 = ~py1 & new_n368;
  assign new_n370 = ~ph1 & pe;
  assign new_n371 = ~pr0 & ~pe;
  assign new_n372 = pd & new_n371;
  assign new_n373 = ~ps2 & new_n264;
  assign new_n374 = ~new_n370 & ~new_n372;
  assign new_n375 = ~new_n373 & new_n374;
  assign new_n376 = ~py1 & new_n375;
  assign new_n377 = ~new_n268 & new_n376;
  assign new_n378 = ~pk2 & pi3;
  assign new_n379 = ~pj2 & new_n378;
  assign new_n380 = pi3 & px1;
  assign new_n381 = ~new_n379 & ~new_n380;
  assign new_n382 = px1 & new_n381;
  assign new_n383 = new_n276 & new_n381;
  assign new_n384 = ~pj3 & new_n381;
  assign new_n385 = ~new_n382 & ~new_n383;
  assign new_n386 = ~new_n384 & new_n385;
  assign new_n387 = new_n376 & new_n386;
  assign new_n388 = pc & new_n376;
  assign new_n389 = ~new_n377 & ~new_n387;
  assign pd7 = new_n388 | ~new_n389;
  assign new_n391 = ~po2 & new_n244;
  assign new_n392 = pj2 & new_n244;
  assign new_n393 = ~new_n391 & ~new_n392;
  assign new_n394 = ~po2 & new_n246;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396 = pn2 & new_n395;
  assign new_n397 = ~pp2 & new_n396;
  assign new_n398 = pg0 & new_n397;
  assign new_n399 = po2 & new_n397;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = ~pj2 & new_n400;
  assign new_n402 = pj2 & ~new_n400;
  assign new_n403 = ~px1 & new_n402;
  assign new_n404 = ~new_n401 & ~new_n403;
  assign new_n405 = ~py1 & new_n404;
  assign new_n406 = ~px1 & new_n405;
  assign new_n407 = pj2 & new_n405;
  assign pe6 = new_n406 | new_n407;
  assign new_n409 = ~pb0 & ~pw;
  assign new_n410 = ps & new_n409;
  assign new_n411 = ~pw & ~pk1;
  assign new_n412 = pb0 & ~pk1;
  assign new_n413 = ~ps & ~pk1;
  assign new_n414 = ~new_n410 & ~new_n411;
  assign new_n415 = ~new_n412 & ~new_n413;
  assign new_n416 = new_n414 & new_n415;
  assign pf5 = ~py1 & new_n416;
  assign new_n418 = ~pp & pr;
  assign new_n419 = pi & new_n418;
  assign new_n420 = ~pp & ~pf1;
  assign new_n421 = ~pr & ~pf1;
  assign new_n422 = ~pf1 & ~pi;
  assign new_n423 = ~new_n419 & ~new_n420;
  assign new_n424 = ~new_n421 & ~new_n422;
  assign new_n425 = new_n423 & new_n424;
  assign pa5 = ~py1 & new_n425;
  assign pb6 = ph2 & ~pn0;
  assign new_n428 = ~ph3 & ~pf;
  assign new_n429 = ~pg & ph;
  assign new_n430 = pf & new_n429;
  assign new_n431 = ~new_n428 & ~new_n430;
  assign new_n432 = ~py1 & new_n431;
  assign new_n433 = ph & new_n432;
  assign new_n434 = ph3 & new_n432;
  assign pc7 = new_n433 | new_n434;
  assign new_n436 = ~pg3 & ~pf;
  assign new_n437 = ~ph3 & ph;
  assign new_n438 = pf & new_n437;
  assign new_n439 = ~new_n436 & ~new_n438;
  assign new_n440 = ~py1 & new_n439;
  assign new_n441 = ph & new_n440;
  assign new_n442 = pg3 & new_n440;
  assign pb7 = new_n441 | new_n442;
  assign pc6 = pl0 & ~pn0;
  assign new_n445 = ~pf3 & ~pf;
  assign new_n446 = ~pg3 & ph;
  assign new_n447 = pf & new_n446;
  assign new_n448 = ~new_n445 & ~new_n447;
  assign new_n449 = ~py1 & new_n448;
  assign new_n450 = ph & new_n449;
  assign new_n451 = pf3 & new_n449;
  assign pa7 = new_n450 | new_n451;
  assign new_n453 = ~pb0 & ~pt;
  assign new_n454 = ps & new_n453;
  assign new_n455 = ~pt & ~ph1;
  assign new_n456 = pb0 & ~ph1;
  assign new_n457 = ~ps & ~ph1;
  assign new_n458 = ~new_n454 & ~new_n455;
  assign new_n459 = ~new_n456 & ~new_n457;
  assign new_n460 = new_n458 & new_n459;
  assign pc5 = ~py1 & new_n460;
  assign new_n462 = ~pi0 & ~pj0;
  assign new_n463 = ~pk0 & pl0;
  assign new_n464 = pd2 & new_n463;
  assign new_n465 = new_n462 & new_n464;
  assign new_n466 = ~ph0 & new_n465;
  assign new_n467 = ~pe4 & pi0;
  assign new_n468 = pf4 & ~pj0;
  assign new_n469 = pf4 & ~pg4;
  assign new_n470 = ~pk0 & new_n469;
  assign new_n471 = pf4 & pg4;
  assign new_n472 = pk0 & new_n471;
  assign new_n473 = ~pg4 & ~pk0;
  assign new_n474 = ~pj0 & new_n473;
  assign new_n475 = pg4 & pk0;
  assign new_n476 = ~pj0 & new_n475;
  assign new_n477 = ~new_n470 & ~new_n472;
  assign new_n478 = ~new_n474 & ~new_n476;
  assign new_n479 = new_n477 & new_n478;
  assign new_n480 = ~new_n467 & ~new_n468;
  assign new_n481 = ~new_n479 & new_n480;
  assign new_n482 = pi0 & new_n481;
  assign new_n483 = ~ph0 & new_n482;
  assign new_n484 = ~pe4 & new_n481;
  assign new_n485 = ~ph0 & new_n484;
  assign new_n486 = ~pd4 & new_n482;
  assign new_n487 = ~pd4 & new_n484;
  assign new_n488 = ~new_n483 & ~new_n485;
  assign new_n489 = ~new_n486 & ~new_n487;
  assign new_n490 = new_n488 & new_n489;
  assign new_n491 = ~pd4 & ~ph0;
  assign new_n492 = ~new_n490 & ~new_n491;
  assign new_n493 = pc4 & new_n492;
  assign new_n494 = pb4 & new_n493;
  assign new_n495 = pa4 & new_n494;
  assign new_n496 = pz3 & new_n495;
  assign new_n497 = py3 & new_n496;
  assign new_n498 = ph4 & new_n497;
  assign new_n499 = ~new_n466 & ~new_n498;
  assign new_n500 = ~pa2 & pf2;
  assign new_n501 = new_n499 & new_n500;
  assign new_n502 = ~pn0 & new_n501;
  assign new_n503 = ~pf2 & pe2;
  assign new_n504 = ~pa2 & ~new_n498;
  assign new_n505 = ~new_n462 & new_n504;
  assign new_n506 = ~new_n464 & new_n504;
  assign new_n507 = ph0 & new_n504;
  assign new_n508 = ~new_n505 & ~new_n506;
  assign new_n509 = ~new_n507 & new_n508;
  assign new_n510 = new_n503 & new_n509;
  assign new_n511 = ~pn0 & new_n510;
  assign new_n512 = ~pe2 & ~pn0;
  assign new_n513 = pf2 & new_n512;
  assign new_n514 = ~new_n502 & ~new_n511;
  assign pa6 = new_n513 | ~new_n514;
  assign new_n516 = ~pq & pr;
  assign new_n517 = pi & new_n516;
  assign new_n518 = ~pq & ~pg1;
  assign new_n519 = ~pr & ~pg1;
  assign new_n520 = ~pg1 & ~pi;
  assign new_n521 = ~new_n517 & ~new_n518;
  assign new_n522 = ~new_n519 & ~new_n520;
  assign new_n523 = new_n521 & new_n522;
  assign pb5 = ~py1 & new_n523;
  assign new_n525 = pg2 & ph2;
  assign new_n526 = ~pn0 & new_n525;
  assign new_n527 = pc2 & ~pn0;
  assign pl4 = new_n526 | new_n527;
  assign new_n529 = pb0 & ~pv;
  assign new_n530 = ps & new_n529;
  assign new_n531 = ~pv & ~pr1;
  assign new_n532 = ~pb0 & ~pr1;
  assign new_n533 = ~ps & ~pr1;
  assign new_n534 = ~new_n530 & ~new_n531;
  assign new_n535 = ~new_n532 & ~new_n533;
  assign new_n536 = new_n534 & new_n535;
  assign pm5 = ~py1 & new_n536;
  assign new_n538 = ~ps2 & ~pf;
  assign new_n539 = ~pt2 & ~ph;
  assign new_n540 = pf & new_n539;
  assign new_n541 = ~new_n538 & ~new_n540;
  assign new_n542 = ~py1 & new_n541;
  assign new_n543 = ~ph & new_n542;
  assign new_n544 = ps2 & new_n542;
  assign pn6 = new_n543 | new_n544;
  assign new_n546 = ~ps1 & pe;
  assign new_n547 = ~pc1 & ~pe;
  assign new_n548 = pd & new_n547;
  assign new_n549 = ~pd3 & new_n264;
  assign new_n550 = ~new_n546 & ~new_n548;
  assign new_n551 = ~new_n549 & new_n550;
  assign new_n552 = ~py1 & new_n551;
  assign new_n553 = ~new_n268 & new_n552;
  assign new_n554 = ~pk2 & pt3;
  assign new_n555 = ~pj2 & new_n554;
  assign new_n556 = pt3 & px1;
  assign new_n557 = ~new_n555 & ~new_n556;
  assign new_n558 = px1 & new_n557;
  assign new_n559 = new_n276 & new_n557;
  assign new_n560 = ~pu3 & new_n557;
  assign new_n561 = ~new_n558 & ~new_n559;
  assign new_n562 = ~new_n560 & new_n561;
  assign new_n563 = new_n552 & new_n562;
  assign new_n564 = pc & new_n552;
  assign new_n565 = ~new_n553 & ~new_n563;
  assign po7 = new_n564 | ~new_n565;
  assign new_n567 = pa4 & pz3;
  assign new_n568 = pb4 & new_n567;
  assign new_n569 = ~pd4 & pc4;
  assign new_n570 = pe4 & new_n569;
  assign new_n571 = new_n568 & new_n570;
  assign new_n572 = py3 & new_n571;
  assign new_n573 = ~pl0 & ~pn0;
  assign new_n574 = pz3 & py3;
  assign new_n575 = new_n572 & new_n573;
  assign new_n576 = ~new_n574 & new_n575;
  assign new_n577 = pa4 & pb4;
  assign new_n578 = pc4 & new_n577;
  assign new_n579 = new_n575 & ~new_n578;
  assign new_n580 = pf4 & new_n573;
  assign new_n581 = ~new_n578 & new_n580;
  assign new_n582 = ~pd4 & pe4;
  assign new_n583 = pf4 & new_n582;
  assign new_n584 = new_n580 & ~new_n583;
  assign new_n585 = ~new_n574 & new_n580;
  assign new_n586 = new_n575 & ~new_n583;
  assign new_n587 = ~new_n576 & ~new_n579;
  assign new_n588 = ~new_n581 & new_n587;
  assign new_n589 = ~new_n584 & ~new_n585;
  assign new_n590 = ~new_n586 & new_n589;
  assign pa8 = ~new_n588 | ~new_n590;
  assign new_n592 = pb0 & ~pu;
  assign new_n593 = ps & new_n592;
  assign new_n594 = ~pu & ~pq1;
  assign new_n595 = ~pb0 & ~pq1;
  assign new_n596 = ~ps & ~pq1;
  assign new_n597 = ~new_n593 & ~new_n594;
  assign new_n598 = ~new_n595 & ~new_n596;
  assign new_n599 = new_n597 & new_n598;
  assign pl5 = ~py1 & new_n599;
  assign new_n601 = ~pr & ~pj;
  assign new_n602 = pi & new_n601;
  assign new_n603 = ~pr0 & ~pj;
  assign new_n604 = pr & ~pr0;
  assign new_n605 = ~pr0 & ~pi;
  assign new_n606 = ~new_n602 & ~new_n603;
  assign new_n607 = ~new_n604 & ~new_n605;
  assign new_n608 = new_n606 & new_n607;
  assign pm4 = ~py1 & new_n608;
  assign new_n610 = ~pr1 & pe;
  assign new_n611 = ~pb1 & ~pe;
  assign new_n612 = pd & new_n611;
  assign new_n613 = ~pc3 & new_n264;
  assign new_n614 = ~new_n610 & ~new_n612;
  assign new_n615 = ~new_n613 & new_n614;
  assign new_n616 = ~py1 & new_n615;
  assign new_n617 = ~new_n268 & new_n616;
  assign new_n618 = ~pk2 & ps3;
  assign new_n619 = ~pj2 & new_n618;
  assign new_n620 = ps3 & px1;
  assign new_n621 = ~new_n619 & ~new_n620;
  assign new_n622 = px1 & new_n621;
  assign new_n623 = new_n276 & new_n621;
  assign new_n624 = ~pt3 & new_n621;
  assign new_n625 = ~new_n622 & ~new_n623;
  assign new_n626 = ~new_n624 & new_n625;
  assign new_n627 = new_n616 & new_n626;
  assign new_n628 = pc & new_n616;
  assign new_n629 = ~new_n617 & ~new_n627;
  assign pn7 = new_n628 | ~new_n629;
  assign new_n631 = ~pf & ~pt2;
  assign new_n632 = ~pu2 & ~ph;
  assign new_n633 = pf & new_n632;
  assign new_n634 = ~new_n631 & ~new_n633;
  assign new_n635 = ~py1 & new_n634;
  assign new_n636 = ~ph & new_n635;
  assign new_n637 = pt2 & new_n635;
  assign po6 = new_n636 | new_n637;
  assign new_n639 = new_n578 & new_n583;
  assign new_n640 = new_n574 & new_n639;
  assign new_n641 = pa4 & new_n574;
  assign new_n642 = new_n573 & new_n640;
  assign new_n643 = ~new_n641 & new_n642;
  assign new_n644 = pb4 & pc4;
  assign new_n645 = ~pd4 & new_n644;
  assign new_n646 = new_n642 & ~new_n645;
  assign new_n647 = pg4 & new_n573;
  assign new_n648 = ~new_n645 & new_n647;
  assign new_n649 = pe4 & pf4;
  assign new_n650 = pg4 & new_n649;
  assign new_n651 = new_n647 & ~new_n650;
  assign new_n652 = ~new_n641 & new_n647;
  assign new_n653 = new_n642 & ~new_n650;
  assign new_n654 = ~new_n643 & ~new_n646;
  assign new_n655 = ~new_n648 & new_n654;
  assign new_n656 = ~new_n651 & ~new_n652;
  assign new_n657 = ~new_n653 & new_n656;
  assign pb8 = ~new_n655 | ~new_n657;
  assign new_n659 = ~pq2 & px1;
  assign new_n660 = ~pq2 & new_n335;
  assign new_n661 = ~pi2 & new_n660;
  assign new_n662 = ~new_n659 & ~new_n661;
  assign new_n663 = ~py1 & new_n662;
  assign new_n664 = px1 & new_n663;
  assign new_n665 = ~pi2 & new_n335;
  assign new_n666 = new_n663 & new_n665;
  assign new_n667 = ~pq2 & new_n663;
  assign new_n668 = ~new_n664 & ~new_n666;
  assign pl6 = new_n667 | ~new_n668;
  assign new_n670 = ~pq1 & pe;
  assign new_n671 = ~pa1 & ~pe;
  assign new_n672 = pd & new_n671;
  assign new_n673 = ~pb3 & new_n264;
  assign new_n674 = ~new_n670 & ~new_n672;
  assign new_n675 = ~new_n673 & new_n674;
  assign new_n676 = ~py1 & new_n675;
  assign new_n677 = ~new_n268 & new_n676;
  assign new_n678 = ~pk2 & pr3;
  assign new_n679 = ~pj2 & new_n678;
  assign new_n680 = pr3 & px1;
  assign new_n681 = ~new_n679 & ~new_n680;
  assign new_n682 = px1 & new_n681;
  assign new_n683 = new_n276 & new_n681;
  assign new_n684 = ~ps3 & new_n681;
  assign new_n685 = ~new_n682 & ~new_n683;
  assign new_n686 = ~new_n684 & new_n685;
  assign new_n687 = new_n676 & new_n686;
  assign new_n688 = pc & new_n676;
  assign new_n689 = ~new_n677 & ~new_n687;
  assign pm7 = new_n688 | ~new_n689;
  assign new_n691 = ~pr & ~pk;
  assign new_n692 = pi & new_n691;
  assign new_n693 = ~ps0 & ~pk;
  assign new_n694 = pr & ~ps0;
  assign new_n695 = ~ps0 & ~pi;
  assign new_n696 = ~new_n692 & ~new_n693;
  assign new_n697 = ~new_n694 & ~new_n695;
  assign new_n698 = new_n696 & new_n697;
  assign pn4 = ~py1 & new_n698;
  assign new_n700 = pb0 & ~px;
  assign new_n701 = ps & new_n700;
  assign new_n702 = ~px & ~pt1;
  assign new_n703 = ~pb0 & ~pt1;
  assign new_n704 = ~ps & ~pt1;
  assign new_n705 = ~new_n701 & ~new_n702;
  assign new_n706 = ~new_n703 & ~new_n704;
  assign new_n707 = new_n705 & new_n706;
  assign po5 = ~py1 & new_n707;
  assign new_n709 = pb & ~new_n525;
  assign new_n710 = ~pn0 & new_n709;
  assign new_n711 = pl0 & new_n710;
  assign new_n712 = pd2 & new_n711;
  assign new_n713 = ph4 & new_n710;
  assign pc8 = new_n712 | new_n713;
  assign new_n715 = ~pp1 & pe;
  assign new_n716 = ~pe & ~pz0;
  assign new_n717 = pd & new_n716;
  assign new_n718 = ~pa3 & new_n264;
  assign new_n719 = ~new_n715 & ~new_n717;
  assign new_n720 = ~new_n718 & new_n719;
  assign new_n721 = ~py1 & new_n720;
  assign new_n722 = ~new_n268 & new_n721;
  assign new_n723 = ~pk2 & pq3;
  assign new_n724 = ~pj2 & new_n723;
  assign new_n725 = pq3 & px1;
  assign new_n726 = ~new_n724 & ~new_n725;
  assign new_n727 = px1 & new_n726;
  assign new_n728 = new_n276 & new_n726;
  assign new_n729 = ~pr3 & new_n726;
  assign new_n730 = ~new_n727 & ~new_n728;
  assign new_n731 = ~new_n729 & new_n730;
  assign new_n732 = new_n721 & new_n731;
  assign new_n733 = pc & new_n721;
  assign new_n734 = ~new_n722 & ~new_n732;
  assign pl7 = new_n733 | ~new_n734;
  assign new_n736 = pq2 & ~new_n665;
  assign new_n737 = ~px1 & new_n736;
  assign new_n738 = ~py1 & new_n737;
  assign new_n739 = px1 & new_n738;
  assign new_n740 = pr2 & pq2;
  assign new_n741 = new_n738 & ~new_n740;
  assign new_n742 = pr2 & ~py1;
  assign new_n743 = ~new_n740 & new_n742;
  assign new_n744 = new_n665 & new_n742;
  assign new_n745 = px1 & new_n742;
  assign new_n746 = new_n665 & new_n738;
  assign new_n747 = ~new_n739 & ~new_n741;
  assign new_n748 = ~new_n743 & new_n747;
  assign new_n749 = ~new_n744 & ~new_n745;
  assign new_n750 = ~new_n746 & new_n749;
  assign pm6 = ~new_n748 | ~new_n750;
  assign new_n752 = pb0 & ~pw;
  assign new_n753 = ps & new_n752;
  assign new_n754 = ~pw & ~ps1;
  assign new_n755 = ~pb0 & ~ps1;
  assign new_n756 = ~ps & ~ps1;
  assign new_n757 = ~new_n753 & ~new_n754;
  assign new_n758 = ~new_n755 & ~new_n756;
  assign new_n759 = new_n757 & new_n758;
  assign pn5 = ~py1 & new_n759;
  assign new_n761 = ~pr & ~pl;
  assign new_n762 = pi & new_n761;
  assign new_n763 = ~pt0 & ~pl;
  assign new_n764 = pr & ~pt0;
  assign new_n765 = ~pt0 & ~pi;
  assign new_n766 = ~new_n762 & ~new_n763;
  assign new_n767 = ~new_n764 & ~new_n765;
  assign new_n768 = new_n766 & new_n767;
  assign po4 = ~py1 & new_n768;
  assign new_n770 = ~pb0 & ~pz;
  assign new_n771 = ps & new_n770;
  assign new_n772 = ~pz & ~pn1;
  assign new_n773 = pb0 & ~pn1;
  assign new_n774 = ~ps & ~pn1;
  assign new_n775 = ~new_n771 & ~new_n772;
  assign new_n776 = ~new_n773 & ~new_n774;
  assign new_n777 = new_n775 & new_n776;
  assign pi5 = ~py1 & new_n777;
  assign new_n779 = pl2 & pm2;
  assign new_n780 = pn2 & new_n779;
  assign new_n781 = ~new_n321 & new_n780;
  assign new_n782 = ~py1 & new_n781;
  assign new_n783 = ~pl2 & new_n782;
  assign new_n784 = pn2 & pm2;
  assign new_n785 = po2 & new_n784;
  assign new_n786 = new_n782 & ~new_n785;
  assign new_n787 = po2 & ~py1;
  assign new_n788 = ~new_n785 & new_n787;
  assign new_n789 = new_n321 & new_n787;
  assign new_n790 = ~pl2 & new_n787;
  assign new_n791 = new_n321 & new_n782;
  assign new_n792 = ~new_n783 & ~new_n786;
  assign new_n793 = ~new_n788 & new_n792;
  assign new_n794 = ~new_n789 & ~new_n790;
  assign new_n795 = ~new_n791 & new_n794;
  assign pj6 = ~new_n793 | ~new_n795;
  assign new_n797 = ~po1 & pe;
  assign new_n798 = ~pe & ~py0;
  assign new_n799 = pd & new_n798;
  assign new_n800 = ~pz2 & new_n264;
  assign new_n801 = ~new_n797 & ~new_n799;
  assign new_n802 = ~new_n800 & new_n801;
  assign new_n803 = ~py1 & new_n802;
  assign new_n804 = ~new_n268 & new_n803;
  assign new_n805 = ~pk2 & pp3;
  assign new_n806 = ~pj2 & new_n805;
  assign new_n807 = pp3 & px1;
  assign new_n808 = ~new_n806 & ~new_n807;
  assign new_n809 = px1 & new_n808;
  assign new_n810 = new_n276 & new_n808;
  assign new_n811 = ~pq3 & new_n808;
  assign new_n812 = ~new_n809 & ~new_n810;
  assign new_n813 = ~new_n811 & new_n812;
  assign new_n814 = new_n803 & new_n813;
  assign new_n815 = pc & new_n803;
  assign new_n816 = ~new_n804 & ~new_n814;
  assign pk7 = new_n815 | ~new_n816;
  assign new_n818 = ~pb0 & ~py;
  assign new_n819 = ps & new_n818;
  assign new_n820 = ~py & ~pm1;
  assign new_n821 = pb0 & ~pm1;
  assign new_n822 = ~ps & ~pm1;
  assign new_n823 = ~new_n819 & ~new_n820;
  assign new_n824 = ~new_n821 & ~new_n822;
  assign new_n825 = new_n823 & new_n824;
  assign ph5 = ~py1 & new_n825;
  assign pi4 = pa2 | ~px1;
  assign new_n828 = ~pn1 & pe;
  assign new_n829 = ~pe & ~px0;
  assign new_n830 = pd & new_n829;
  assign new_n831 = ~py2 & new_n264;
  assign new_n832 = ~new_n828 & ~new_n830;
  assign new_n833 = ~new_n831 & new_n832;
  assign new_n834 = ~py1 & new_n833;
  assign new_n835 = ~new_n268 & new_n834;
  assign new_n836 = ~pk2 & po3;
  assign new_n837 = ~pj2 & new_n836;
  assign new_n838 = po3 & px1;
  assign new_n839 = ~new_n837 & ~new_n838;
  assign new_n840 = px1 & new_n839;
  assign new_n841 = new_n276 & new_n839;
  assign new_n842 = ~pp3 & new_n839;
  assign new_n843 = ~new_n840 & ~new_n841;
  assign new_n844 = ~new_n842 & new_n843;
  assign new_n845 = new_n834 & new_n844;
  assign new_n846 = pc & new_n834;
  assign new_n847 = ~new_n835 & ~new_n845;
  assign pj7 = new_n846 | ~new_n847;
  assign new_n849 = ~new_n321 & new_n785;
  assign new_n850 = pl2 & new_n849;
  assign new_n851 = ~py1 & new_n850;
  assign new_n852 = ~new_n779 & new_n851;
  assign new_n853 = pn2 & po2;
  assign new_n854 = pp2 & new_n853;
  assign new_n855 = new_n851 & ~new_n854;
  assign new_n856 = pp2 & ~py1;
  assign new_n857 = ~new_n854 & new_n856;
  assign new_n858 = new_n321 & new_n856;
  assign new_n859 = ~new_n779 & new_n856;
  assign new_n860 = new_n321 & new_n851;
  assign new_n861 = ~new_n852 & ~new_n855;
  assign new_n862 = ~new_n857 & new_n861;
  assign new_n863 = ~new_n858 & ~new_n859;
  assign new_n864 = ~new_n860 & new_n863;
  assign pk6 = ~new_n862 | ~new_n864;
  assign new_n866 = ~pm2 & new_n319;
  assign new_n867 = ~pc & new_n866;
  assign new_n868 = ~pd & new_n867;
  assign new_n869 = ~py1 & ~new_n868;
  assign new_n870 = new_n321 & new_n869;
  assign new_n871 = pm2 & new_n870;
  assign new_n872 = ~pm2 & new_n869;
  assign new_n873 = pl2 & new_n872;
  assign new_n874 = pl2 & new_n870;
  assign new_n875 = pm2 & new_n869;
  assign new_n876 = ~pl2 & new_n875;
  assign new_n877 = ~new_n871 & ~new_n873;
  assign new_n878 = ~new_n874 & ~new_n876;
  assign ph6 = ~new_n877 | ~new_n878;
  assign new_n880 = ~pm1 & pe;
  assign new_n881 = ~pe & ~pw0;
  assign new_n882 = pd & new_n881;
  assign new_n883 = ~px2 & new_n264;
  assign new_n884 = ~new_n880 & ~new_n882;
  assign new_n885 = ~new_n883 & new_n884;
  assign new_n886 = ~py1 & new_n885;
  assign new_n887 = ~new_n268 & new_n886;
  assign new_n888 = ~pk2 & pn3;
  assign new_n889 = ~pj2 & new_n888;
  assign new_n890 = pn3 & px1;
  assign new_n891 = ~new_n889 & ~new_n890;
  assign new_n892 = px1 & new_n891;
  assign new_n893 = new_n276 & new_n891;
  assign new_n894 = ~po3 & new_n891;
  assign new_n895 = ~new_n892 & ~new_n893;
  assign new_n896 = ~new_n894 & new_n895;
  assign new_n897 = new_n886 & new_n896;
  assign new_n898 = pc & new_n886;
  assign new_n899 = ~new_n887 & ~new_n897;
  assign pi7 = new_n898 | ~new_n899;
  assign new_n901 = ~po0 & px1;
  assign new_n902 = ~po0 & ~new_n740;
  assign new_n903 = ~pi2 & ~po0;
  assign new_n904 = ~new_n901 & ~new_n902;
  assign new_n905 = ~new_n903 & new_n904;
  assign new_n906 = new_n268 & new_n905;
  assign new_n907 = ~pc & new_n906;
  assign pj4 = py1 | new_n907;
  assign new_n909 = pb0 & ~pt;
  assign new_n910 = ps & new_n909;
  assign new_n911 = ~pt & ~pp1;
  assign new_n912 = ~pb0 & ~pp1;
  assign new_n913 = ~ps & ~pp1;
  assign new_n914 = ~new_n910 & ~new_n911;
  assign new_n915 = ~new_n912 & ~new_n913;
  assign new_n916 = new_n914 & new_n915;
  assign pk5 = ~py1 & new_n916;
  assign new_n918 = ~pl1 & pe;
  assign new_n919 = ~pe & ~pv0;
  assign new_n920 = pd & new_n919;
  assign new_n921 = ~pw2 & new_n264;
  assign new_n922 = ~new_n918 & ~new_n920;
  assign new_n923 = ~new_n921 & new_n922;
  assign new_n924 = ~py1 & new_n923;
  assign new_n925 = ~new_n268 & new_n924;
  assign new_n926 = ~pk2 & pm3;
  assign new_n927 = ~pj2 & new_n926;
  assign new_n928 = pm3 & px1;
  assign new_n929 = ~new_n927 & ~new_n928;
  assign new_n930 = px1 & new_n929;
  assign new_n931 = new_n276 & new_n929;
  assign new_n932 = ~pn3 & new_n929;
  assign new_n933 = ~new_n930 & ~new_n931;
  assign new_n934 = ~new_n932 & new_n933;
  assign new_n935 = new_n924 & new_n934;
  assign new_n936 = pc & new_n924;
  assign new_n937 = ~new_n925 & ~new_n935;
  assign ph7 = new_n936 | ~new_n937;
  assign new_n939 = ~new_n321 & new_n779;
  assign new_n940 = ~py1 & new_n939;
  assign new_n941 = ~pl2 & new_n940;
  assign new_n942 = ~new_n784 & new_n940;
  assign new_n943 = pn2 & ~py1;
  assign new_n944 = ~new_n784 & new_n943;
  assign new_n945 = new_n321 & new_n943;
  assign new_n946 = ~pl2 & new_n943;
  assign new_n947 = new_n321 & new_n940;
  assign new_n948 = ~new_n941 & ~new_n942;
  assign new_n949 = ~new_n944 & new_n948;
  assign new_n950 = ~new_n945 & ~new_n946;
  assign new_n951 = ~new_n947 & new_n950;
  assign pi6 = ~new_n949 | ~new_n951;
  assign new_n953 = ~pa0 & ~pb0;
  assign new_n954 = ps & new_n953;
  assign new_n955 = ~pa0 & ~po1;
  assign new_n956 = pb0 & ~po1;
  assign new_n957 = ~ps & ~po1;
  assign new_n958 = ~new_n954 & ~new_n955;
  assign new_n959 = ~new_n956 & ~new_n957;
  assign new_n960 = new_n958 & new_n959;
  assign pj5 = ~py1 & new_n960;
  assign new_n962 = ~pa2 & ~pj2;
  assign new_n963 = ~pk2 & new_n962;
  assign new_n964 = pi2 & pq2;
  assign new_n965 = pi2 & pr2;
  assign new_n966 = ~new_n964 & ~new_n965;
  assign new_n967 = ~pk0 & ~pl2;
  assign new_n968 = ~pj0 & ~pk0;
  assign new_n969 = ~pj0 & pl2;
  assign new_n970 = ~new_n967 & ~new_n968;
  assign new_n971 = ~pn2 & ~new_n969;
  assign new_n972 = new_n970 & new_n971;
  assign new_n973 = ~po2 & ~pp2;
  assign new_n974 = new_n972 & new_n973;
  assign new_n975 = pm2 & new_n974;
  assign new_n976 = ~pi0 & ~pl2;
  assign new_n977 = ~ph0 & ~pi0;
  assign new_n978 = ~ph0 & pl2;
  assign new_n979 = ~new_n976 & ~new_n977;
  assign new_n980 = pn2 & ~new_n978;
  assign new_n981 = new_n979 & new_n980;
  assign new_n982 = new_n974 & new_n981;
  assign new_n983 = new_n973 & new_n981;
  assign new_n984 = ~pm2 & new_n983;
  assign new_n985 = ~new_n975 & ~new_n982;
  assign new_n986 = ~new_n984 & new_n985;
  assign new_n987 = ~py1 & ~new_n986;
  assign new_n988 = new_n963 & new_n966;
  assign new_n989 = new_n987 & new_n988;
  assign new_n990 = ~pa2 & ~py1;
  assign new_n991 = pd0 & new_n965;
  assign new_n992 = pi3 & pr2;
  assign new_n993 = pd0 & new_n992;
  assign new_n994 = pi3 & ~pi2;
  assign new_n995 = pi3 & pq2;
  assign new_n996 = ~new_n991 & ~new_n993;
  assign new_n997 = ~new_n994 & new_n996;
  assign new_n998 = ~new_n964 & ~new_n995;
  assign new_n999 = new_n997 & new_n998;
  assign new_n1000 = pr2 & new_n999;
  assign new_n1001 = ~pi3 & new_n999;
  assign new_n1002 = ~new_n1000 & ~new_n1001;
  assign new_n1003 = ~pi2 & new_n1002;
  assign new_n1004 = pk2 & new_n1003;
  assign new_n1005 = pj2 & new_n1003;
  assign new_n1006 = ~pq2 & new_n1002;
  assign new_n1007 = pj2 & new_n1006;
  assign new_n1008 = ~pr2 & ~pq2;
  assign new_n1009 = pi2 & ~new_n1008;
  assign new_n1010 = new_n1006 & new_n1009;
  assign new_n1011 = pk2 & new_n1006;
  assign new_n1012 = pr2 & pz1;
  assign new_n1013 = pc0 & ~pr2;
  assign new_n1014 = pc0 & pz1;
  assign new_n1015 = ~new_n1012 & ~new_n1013;
  assign new_n1016 = ~new_n1014 & new_n1015;
  assign new_n1017 = new_n1002 & new_n1016;
  assign new_n1018 = pj2 & new_n1017;
  assign new_n1019 = new_n1009 & new_n1017;
  assign new_n1020 = new_n1003 & new_n1009;
  assign new_n1021 = pk2 & new_n1017;
  assign new_n1022 = ~new_n1004 & ~new_n1005;
  assign new_n1023 = ~new_n1007 & new_n1022;
  assign new_n1024 = ~new_n1010 & ~new_n1011;
  assign new_n1025 = new_n1023 & new_n1024;
  assign new_n1026 = ~new_n1020 & ~new_n1021;
  assign new_n1027 = ~new_n1018 & ~new_n1019;
  assign new_n1028 = new_n1026 & new_n1027;
  assign new_n1029 = new_n1025 & new_n1028;
  assign new_n1030 = new_n990 & ~new_n1029;
  assign new_n1031 = ~px1 & new_n1030;
  assign new_n1032 = ~pm0 & new_n986;
  assign new_n1033 = pa2 & ~py1;
  assign new_n1034 = new_n986 & ~new_n1033;
  assign new_n1035 = ~px1 & ~new_n1033;
  assign new_n1036 = ~pd0 & new_n503;
  assign new_n1037 = pf2 & ~pe2;
  assign new_n1038 = pd0 & new_n1037;
  assign new_n1039 = ~new_n1036 & ~new_n1038;
  assign new_n1040 = ~px1 & new_n1039;
  assign new_n1041 = ~pm0 & ~px1;
  assign new_n1042 = ~new_n990 & ~new_n1033;
  assign new_n1043 = ~new_n990 & new_n1039;
  assign new_n1044 = new_n986 & new_n1039;
  assign new_n1045 = ~pm0 & ~new_n990;
  assign new_n1046 = ~new_n1032 & ~new_n1034;
  assign new_n1047 = ~new_n1035 & new_n1046;
  assign new_n1048 = ~new_n1040 & ~new_n1041;
  assign new_n1049 = new_n1047 & new_n1048;
  assign new_n1050 = ~new_n1044 & ~new_n1045;
  assign new_n1051 = ~new_n1042 & ~new_n1043;
  assign new_n1052 = new_n1050 & new_n1051;
  assign new_n1053 = new_n1049 & new_n1052;
  assign new_n1054 = ~new_n989 & ~new_n1031;
  assign pk4 = new_n1053 | ~new_n1054;
  assign new_n1056 = ~pq & ~pr;
  assign new_n1057 = pi & new_n1056;
  assign new_n1058 = ~pq & ~py0;
  assign new_n1059 = pr & ~py0;
  assign new_n1060 = ~pi & ~py0;
  assign new_n1061 = ~new_n1057 & ~new_n1058;
  assign new_n1062 = ~new_n1059 & ~new_n1060;
  assign new_n1063 = new_n1061 & new_n1062;
  assign pt4 = ~py1 & new_n1063;
  assign new_n1065 = ~py1 & ~pz1;
  assign new_n1066 = pi3 & ~pr2;
  assign new_n1067 = ~pi2 & ~new_n276;
  assign new_n1068 = pi3 & new_n1067;
  assign new_n1069 = pc0 & ~pd0;
  assign new_n1070 = ~pd0 & ~pq2;
  assign new_n1071 = ~new_n1013 & ~new_n1069;
  assign new_n1072 = ~new_n1070 & new_n1071;
  assign new_n1073 = new_n1009 & new_n1072;
  assign new_n1074 = ~new_n1068 & ~new_n1073;
  assign new_n1075 = ~new_n1066 & new_n1074;
  assign new_n1076 = new_n986 & new_n1075;
  assign new_n1077 = ~new_n276 & new_n1075;
  assign new_n1078 = pq2 & new_n1074;
  assign new_n1079 = ~new_n276 & new_n1078;
  assign new_n1080 = new_n1009 & new_n1078;
  assign new_n1081 = new_n986 & new_n1078;
  assign new_n1082 = new_n276 & new_n1074;
  assign new_n1083 = ~new_n276 & new_n1082;
  assign new_n1084 = new_n1009 & new_n1082;
  assign new_n1085 = new_n1009 & new_n1075;
  assign new_n1086 = new_n986 & new_n1082;
  assign new_n1087 = ~new_n1076 & ~new_n1077;
  assign new_n1088 = ~new_n1079 & new_n1087;
  assign new_n1089 = ~new_n1080 & ~new_n1081;
  assign new_n1090 = new_n1088 & new_n1089;
  assign new_n1091 = ~new_n1085 & ~new_n1086;
  assign new_n1092 = ~new_n1083 & ~new_n1084;
  assign new_n1093 = new_n1091 & new_n1092;
  assign new_n1094 = new_n1090 & new_n1093;
  assign new_n1095 = new_n1065 & new_n1094;
  assign new_n1096 = ~px1 & new_n1095;
  assign new_n1097 = ~pi3 & ~pr2;
  assign new_n1098 = ~pi3 & new_n1067;
  assign new_n1099 = pd0 & ~px1;
  assign new_n1100 = ~pc0 & new_n1099;
  assign new_n1101 = pd0 & ~pq2;
  assign new_n1102 = ~px1 & new_n1101;
  assign new_n1103 = ~pr2 & ~px1;
  assign new_n1104 = ~pc0 & new_n1103;
  assign new_n1105 = ~px1 & new_n1008;
  assign new_n1106 = ~pi2 & ~px1;
  assign new_n1107 = ~new_n1100 & ~new_n1102;
  assign new_n1108 = ~new_n1104 & new_n1107;
  assign new_n1109 = ~new_n1105 & ~new_n1106;
  assign new_n1110 = new_n1108 & new_n1109;
  assign new_n1111 = ~new_n1098 & ~new_n1110;
  assign new_n1112 = ~new_n1097 & new_n1111;
  assign new_n1113 = ~new_n986 & new_n1112;
  assign new_n1114 = ~new_n276 & new_n1112;
  assign new_n1115 = pq2 & new_n1111;
  assign new_n1116 = ~new_n276 & new_n1115;
  assign new_n1117 = new_n1009 & new_n1115;
  assign new_n1118 = ~new_n986 & new_n1115;
  assign new_n1119 = new_n276 & new_n1111;
  assign new_n1120 = ~new_n276 & new_n1119;
  assign new_n1121 = new_n1009 & new_n1119;
  assign new_n1122 = new_n1009 & new_n1112;
  assign new_n1123 = ~new_n986 & new_n1119;
  assign new_n1124 = ~new_n1113 & ~new_n1114;
  assign new_n1125 = ~new_n1116 & new_n1124;
  assign new_n1126 = ~new_n1117 & ~new_n1118;
  assign new_n1127 = new_n1125 & new_n1126;
  assign new_n1128 = ~new_n1122 & ~new_n1123;
  assign new_n1129 = ~new_n1120 & ~new_n1121;
  assign new_n1130 = new_n1128 & new_n1129;
  assign new_n1131 = new_n1127 & new_n1130;
  assign new_n1132 = ~py1 & new_n1131;
  assign new_n1133 = pz1 & new_n1132;
  assign new_n1134 = ~py1 & ~px1;
  assign new_n1135 = pi2 & new_n1134;
  assign new_n1136 = pq2 & new_n1135;
  assign new_n1137 = pr2 & new_n1136;
  assign new_n1138 = ~new_n1096 & ~new_n1133;
  assign pu5 = new_n1137 | ~new_n1138;
  assign new_n1140 = ~pa3 & ~pf;
  assign new_n1141 = ~pb3 & ph;
  assign new_n1142 = pf & new_n1141;
  assign new_n1143 = ~new_n1140 & ~new_n1142;
  assign new_n1144 = ~py1 & new_n1143;
  assign new_n1145 = ph & new_n1144;
  assign new_n1146 = pa3 & new_n1144;
  assign pv6 = new_n1145 | new_n1146;
  assign new_n1148 = new_n573 & new_n641;
  assign new_n1149 = ~pz3 & new_n1148;
  assign new_n1150 = ~py3 & new_n1148;
  assign new_n1151 = pb4 & new_n573;
  assign new_n1152 = ~py3 & new_n1151;
  assign new_n1153 = ~new_n577 & new_n1151;
  assign new_n1154 = ~pz3 & new_n1151;
  assign new_n1155 = ~new_n577 & new_n1148;
  assign new_n1156 = ~new_n1149 & ~new_n1150;
  assign new_n1157 = ~new_n1152 & new_n1156;
  assign new_n1158 = ~new_n1153 & ~new_n1154;
  assign new_n1159 = ~new_n1155 & new_n1158;
  assign pw7 = ~new_n1157 | ~new_n1159;
  assign new_n1161 = ~px1 & new_n740;
  assign new_n1162 = pi2 & new_n1161;
  assign pt5 = pn0 | new_n1162;
  assign new_n1164 = pr & ~pj;
  assign new_n1165 = pi & new_n1164;
  assign new_n1166 = ~pj & ~pz0;
  assign new_n1167 = ~pr & ~pz0;
  assign new_n1168 = ~pi & ~pz0;
  assign new_n1169 = ~new_n1165 & ~new_n1166;
  assign new_n1170 = ~new_n1167 & ~new_n1168;
  assign new_n1171 = new_n1169 & new_n1170;
  assign pu4 = ~py1 & new_n1171;
  assign new_n1173 = py3 & new_n567;
  assign new_n1174 = ~pl0 & ~new_n1173;
  assign new_n1175 = ~pn0 & new_n1174;
  assign new_n1176 = py3 & new_n1175;
  assign new_n1177 = pz3 & new_n1176;
  assign new_n1178 = pa4 & new_n1175;
  assign pv7 = new_n1177 | new_n1178;
  assign new_n1180 = ~pb3 & ~pf;
  assign new_n1181 = ~pc3 & ph;
  assign new_n1182 = pf & new_n1181;
  assign new_n1183 = ~new_n1180 & ~new_n1182;
  assign new_n1184 = ~py1 & new_n1183;
  assign new_n1185 = ph & new_n1184;
  assign new_n1186 = pb3 & new_n1184;
  assign pw6 = new_n1185 | new_n1186;
  assign new_n1188 = ~pf & ~py2;
  assign new_n1189 = ~ph & ~pz2;
  assign new_n1190 = pf & new_n1189;
  assign new_n1191 = ~new_n1188 & ~new_n1190;
  assign new_n1192 = ~py1 & new_n1191;
  assign new_n1193 = ~ph & new_n1192;
  assign new_n1194 = py2 & new_n1192;
  assign pt6 = new_n1193 | new_n1194;
  assign new_n1196 = ~pl0 & ~new_n574;
  assign new_n1197 = ~pn0 & new_n1196;
  assign new_n1198 = py3 & new_n1197;
  assign new_n1199 = pz3 & new_n1197;
  assign pu7 = new_n1198 | new_n1199;
  assign new_n1201 = pr & ~pk;
  assign new_n1202 = pi & new_n1201;
  assign new_n1203 = ~pa1 & ~pk;
  assign new_n1204 = ~pa1 & ~pr;
  assign new_n1205 = ~pa1 & ~pi;
  assign new_n1206 = ~new_n1202 & ~new_n1203;
  assign new_n1207 = ~new_n1204 & ~new_n1205;
  assign new_n1208 = new_n1206 & new_n1207;
  assign pv4 = ~py1 & new_n1208;
  assign new_n1210 = pd4 & new_n644;
  assign new_n1211 = ~pe4 & ~pf4;
  assign new_n1212 = ~pg4 & new_n1211;
  assign new_n1213 = new_n1210 & new_n1212;
  assign new_n1214 = new_n641 & new_n1213;
  assign new_n1215 = ~pf4 & ~pg4;
  assign new_n1216 = pb2 & new_n1215;
  assign new_n1217 = py3 & new_n1216;
  assign new_n1218 = new_n573 & new_n1214;
  assign new_n1219 = ~new_n1217 & new_n1218;
  assign new_n1220 = ~new_n568 & new_n1218;
  assign new_n1221 = pb2 & new_n573;
  assign new_n1222 = ~new_n568 & new_n1221;
  assign new_n1223 = pd4 & pc4;
  assign new_n1224 = ~pe4 & new_n1223;
  assign new_n1225 = new_n1221 & ~new_n1224;
  assign new_n1226 = ~new_n1217 & new_n1221;
  assign new_n1227 = new_n1218 & ~new_n1224;
  assign new_n1228 = ~new_n1219 & ~new_n1220;
  assign new_n1229 = ~new_n1222 & new_n1228;
  assign new_n1230 = ~new_n1225 & ~new_n1226;
  assign new_n1231 = ~new_n1227 & new_n1230;
  assign pw5 = ~new_n1229 | ~new_n1231;
  assign pt7 = ~py3 & new_n573;
  assign new_n1234 = ~pf & ~pz2;
  assign new_n1235 = ~pg & ~ph;
  assign new_n1236 = pf & new_n1235;
  assign new_n1237 = ~new_n1234 & ~new_n1236;
  assign new_n1238 = ~py1 & new_n1237;
  assign new_n1239 = ~ph & new_n1238;
  assign new_n1240 = pz2 & new_n1238;
  assign pu6 = new_n1239 | new_n1240;
  assign new_n1242 = pa2 & ~pf2;
  assign new_n1243 = pa2 & ~pe2;
  assign new_n1244 = ~new_n498 & ~new_n1242;
  assign new_n1245 = ~new_n1243 & new_n1244;
  assign new_n1246 = ~new_n462 & new_n1245;
  assign new_n1247 = ~new_n464 & new_n1245;
  assign new_n1248 = ph0 & new_n1245;
  assign new_n1249 = ~new_n1246 & ~new_n1247;
  assign new_n1250 = ~new_n1248 & new_n1249;
  assign pv5 = ~py1 & new_n1250;
  assign new_n1252 = pr & ~pl;
  assign new_n1253 = pi & new_n1252;
  assign new_n1254 = ~pb1 & ~pl;
  assign new_n1255 = ~pr & ~pb1;
  assign new_n1256 = ~pb1 & ~pi;
  assign new_n1257 = ~new_n1253 & ~new_n1254;
  assign new_n1258 = ~new_n1255 & ~new_n1256;
  assign new_n1259 = new_n1257 & new_n1258;
  assign pw4 = ~py1 & new_n1259;
  assign new_n1261 = ~pr & ~pm;
  assign new_n1262 = pi & new_n1261;
  assign new_n1263 = ~pu0 & ~pm;
  assign new_n1264 = pr & ~pu0;
  assign new_n1265 = ~pu0 & ~pi;
  assign new_n1266 = ~new_n1262 & ~new_n1263;
  assign new_n1267 = ~new_n1264 & ~new_n1265;
  assign new_n1268 = new_n1266 & new_n1267;
  assign pp4 = ~py1 & new_n1268;
  assign new_n1270 = pb0 & ~pz;
  assign new_n1271 = ps & new_n1270;
  assign new_n1272 = ~pz & ~pv1;
  assign new_n1273 = ~pb0 & ~pv1;
  assign new_n1274 = ~ps & ~pv1;
  assign new_n1275 = ~new_n1271 & ~new_n1272;
  assign new_n1276 = ~new_n1273 & ~new_n1274;
  assign new_n1277 = new_n1275 & new_n1276;
  assign pq5 = ~py1 & new_n1277;
  assign new_n1279 = ~pw2 & ~pf;
  assign new_n1280 = ~ph & ~px2;
  assign new_n1281 = pf & new_n1280;
  assign new_n1282 = ~new_n1279 & ~new_n1281;
  assign new_n1283 = ~py1 & new_n1282;
  assign new_n1284 = ~ph & new_n1283;
  assign new_n1285 = pw2 & new_n1283;
  assign pr6 = new_n1284 | new_n1285;
  assign new_n1287 = pe & ~pw1;
  assign new_n1288 = ~pg1 & ~pe;
  assign new_n1289 = pd & new_n1288;
  assign new_n1290 = ~ph3 & new_n264;
  assign new_n1291 = ~new_n1287 & ~new_n1289;
  assign new_n1292 = ~new_n1290 & new_n1291;
  assign new_n1293 = ~py1 & new_n1292;
  assign new_n1294 = ~new_n268 & new_n1293;
  assign new_n1295 = pk2 & ~px1;
  assign new_n1296 = pj2 & ~px1;
  assign new_n1297 = ~new_n1295 & ~new_n1296;
  assign new_n1298 = px3 & new_n1297;
  assign new_n1299 = new_n1293 & new_n1298;
  assign new_n1300 = pc & new_n1293;
  assign new_n1301 = ~new_n1294 & ~new_n1299;
  assign ps7 = new_n1300 | ~new_n1301;
  assign new_n1303 = pb0 & ~py;
  assign new_n1304 = ps & new_n1303;
  assign new_n1305 = ~py & ~pu1;
  assign new_n1306 = ~pb0 & ~pu1;
  assign new_n1307 = ~ps & ~pu1;
  assign new_n1308 = ~new_n1304 & ~new_n1305;
  assign new_n1309 = ~new_n1306 & ~new_n1307;
  assign new_n1310 = new_n1308 & new_n1309;
  assign pp5 = ~py1 & new_n1310;
  assign new_n1312 = ~pr & ~pn;
  assign new_n1313 = pi & new_n1312;
  assign new_n1314 = ~pv0 & ~pn;
  assign new_n1315 = pr & ~pv0;
  assign new_n1316 = ~pv0 & ~pi;
  assign new_n1317 = ~new_n1313 & ~new_n1314;
  assign new_n1318 = ~new_n1315 & ~new_n1316;
  assign new_n1319 = new_n1317 & new_n1318;
  assign pq4 = ~py1 & new_n1319;
  assign new_n1321 = pe & ~pv1;
  assign new_n1322 = ~pf1 & ~pe;
  assign new_n1323 = pd & new_n1322;
  assign new_n1324 = ~pg3 & new_n264;
  assign new_n1325 = ~new_n1321 & ~new_n1323;
  assign new_n1326 = ~new_n1324 & new_n1325;
  assign new_n1327 = ~py1 & new_n1326;
  assign new_n1328 = ~new_n268 & new_n1327;
  assign new_n1329 = ~pk2 & pw3;
  assign new_n1330 = ~pj2 & new_n1329;
  assign new_n1331 = pw3 & px1;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = px1 & new_n1332;
  assign new_n1334 = new_n276 & new_n1332;
  assign new_n1335 = ~px3 & new_n1332;
  assign new_n1336 = ~new_n1333 & ~new_n1334;
  assign new_n1337 = ~new_n1335 & new_n1336;
  assign new_n1338 = new_n1327 & new_n1337;
  assign new_n1339 = pc & new_n1327;
  assign new_n1340 = ~new_n1328 & ~new_n1338;
  assign pr7 = new_n1339 | ~new_n1340;
  assign new_n1342 = ~pf & ~px2;
  assign new_n1343 = ~ph & ~py2;
  assign new_n1344 = pf & new_n1343;
  assign new_n1345 = ~new_n1342 & ~new_n1344;
  assign new_n1346 = ~py1 & new_n1345;
  assign new_n1347 = ~ph & new_n1346;
  assign new_n1348 = px2 & new_n1346;
  assign ps6 = new_n1347 | new_n1348;
  assign new_n1350 = ~pf & ~pu2;
  assign new_n1351 = ~pv2 & ~ph;
  assign new_n1352 = pf & new_n1351;
  assign new_n1353 = ~new_n1350 & ~new_n1352;
  assign new_n1354 = ~py1 & new_n1353;
  assign new_n1355 = ~ph & new_n1354;
  assign new_n1356 = pu2 & new_n1354;
  assign pp6 = new_n1355 | new_n1356;
  assign new_n1358 = ~pu1 & pe;
  assign new_n1359 = ~pe1 & ~pe;
  assign new_n1360 = pd & new_n1359;
  assign new_n1361 = ~pf3 & new_n264;
  assign new_n1362 = ~new_n1358 & ~new_n1360;
  assign new_n1363 = ~new_n1361 & new_n1362;
  assign new_n1364 = ~py1 & new_n1363;
  assign new_n1365 = ~new_n268 & new_n1364;
  assign new_n1366 = ~pk2 & pv3;
  assign new_n1367 = ~pj2 & new_n1366;
  assign new_n1368 = pv3 & px1;
  assign new_n1369 = ~new_n1367 & ~new_n1368;
  assign new_n1370 = px1 & new_n1369;
  assign new_n1371 = new_n276 & new_n1369;
  assign new_n1372 = ~pw3 & new_n1369;
  assign new_n1373 = ~new_n1370 & ~new_n1371;
  assign new_n1374 = ~new_n1372 & new_n1373;
  assign new_n1375 = new_n1364 & new_n1374;
  assign new_n1376 = pc & new_n1364;
  assign new_n1377 = ~new_n1365 & ~new_n1375;
  assign pq7 = new_n1376 | ~new_n1377;
  assign new_n1379 = ~pr & ~po;
  assign new_n1380 = pi & new_n1379;
  assign new_n1381 = ~pw0 & ~po;
  assign new_n1382 = pr & ~pw0;
  assign new_n1383 = ~pw0 & ~pi;
  assign new_n1384 = ~new_n1380 & ~new_n1381;
  assign new_n1385 = ~new_n1382 & ~new_n1383;
  assign new_n1386 = new_n1384 & new_n1385;
  assign pr4 = ~py1 & new_n1386;
  assign ps5 = py1 | new_n321;
  assign new_n1389 = pe & ~pt1;
  assign new_n1390 = ~pd1 & ~pe;
  assign new_n1391 = pd & new_n1390;
  assign new_n1392 = ~pe3 & new_n264;
  assign new_n1393 = ~new_n1389 & ~new_n1391;
  assign new_n1394 = ~new_n1392 & new_n1393;
  assign new_n1395 = ~py1 & new_n1394;
  assign new_n1396 = ~new_n268 & new_n1395;
  assign new_n1397 = ~pk2 & pu3;
  assign new_n1398 = ~pj2 & new_n1397;
  assign new_n1399 = pu3 & px1;
  assign new_n1400 = ~new_n1398 & ~new_n1399;
  assign new_n1401 = px1 & new_n1400;
  assign new_n1402 = new_n276 & new_n1400;
  assign new_n1403 = ~pv3 & new_n1400;
  assign new_n1404 = ~new_n1401 & ~new_n1402;
  assign new_n1405 = ~new_n1403 & new_n1404;
  assign new_n1406 = new_n1395 & new_n1405;
  assign new_n1407 = pc & new_n1395;
  assign new_n1408 = ~new_n1396 & ~new_n1406;
  assign pp7 = new_n1407 | ~new_n1408;
  assign new_n1410 = ~pv2 & ~pf;
  assign new_n1411 = ~pw2 & ~ph;
  assign new_n1412 = pf & new_n1411;
  assign new_n1413 = ~new_n1410 & ~new_n1412;
  assign new_n1414 = ~py1 & new_n1413;
  assign new_n1415 = ~ph & new_n1414;
  assign new_n1416 = pv2 & new_n1414;
  assign pq6 = new_n1415 | new_n1416;
  assign new_n1418 = ~pa0 & pb0;
  assign new_n1419 = ps & new_n1418;
  assign new_n1420 = ~pa0 & ~pw1;
  assign new_n1421 = ~pb0 & ~pw1;
  assign new_n1422 = ~ps & ~pw1;
  assign new_n1423 = ~new_n1419 & ~new_n1420;
  assign new_n1424 = ~new_n1421 & ~new_n1422;
  assign new_n1425 = new_n1423 & new_n1424;
  assign pr5 = ~py1 & new_n1425;
  assign new_n1427 = ~pp & ~pr;
  assign new_n1428 = pi & new_n1427;
  assign new_n1429 = ~pp & ~px0;
  assign new_n1430 = pr & ~px0;
  assign new_n1431 = ~px0 & ~pi;
  assign new_n1432 = ~new_n1428 & ~new_n1429;
  assign new_n1433 = ~new_n1430 & ~new_n1431;
  assign new_n1434 = new_n1432 & new_n1433;
  assign ps4 = ~py1 & new_n1434;
  assign new_n1436 = pr & ~pm;
  assign new_n1437 = pi & new_n1436;
  assign new_n1438 = ~pc1 & ~pm;
  assign new_n1439 = ~pc1 & ~pr;
  assign new_n1440 = ~pc1 & ~pi;
  assign new_n1441 = ~new_n1437 & ~new_n1438;
  assign new_n1442 = ~new_n1439 & ~new_n1440;
  assign new_n1443 = new_n1441 & new_n1442;
  assign px4 = ~py1 & new_n1443;
  assign new_n1445 = ~pd2 & ~pl0;
  assign new_n1446 = pb & ~new_n1445;
  assign new_n1447 = ~pn0 & new_n1446;
  assign new_n1448 = ~pg2 & new_n1447;
  assign new_n1449 = ~ph2 & new_n1447;
  assign py5 = new_n1448 | new_n1449;
  assign new_n1451 = ~pe3 & ~pf;
  assign new_n1452 = ~pf3 & ph;
  assign new_n1453 = pf & new_n1452;
  assign new_n1454 = ~new_n1451 & ~new_n1453;
  assign new_n1455 = ~py1 & new_n1454;
  assign new_n1456 = ph & new_n1455;
  assign new_n1457 = pe3 & new_n1455;
  assign pz6 = new_n1456 | new_n1457;
  assign new_n1459 = new_n568 & new_n1224;
  assign new_n1460 = new_n1217 & new_n1459;
  assign new_n1461 = new_n527 & ~new_n1460;
  assign new_n1462 = ~pl0 & new_n1461;
  assign new_n1463 = pb2 & ~pn0;
  assign new_n1464 = ~pc2 & new_n1463;
  assign new_n1465 = ~pl0 & new_n1213;
  assign new_n1466 = new_n641 & new_n1464;
  assign new_n1467 = new_n1465 & new_n1466;
  assign px5 = new_n1462 | new_n1467;
  assign new_n1469 = pr & ~pn;
  assign new_n1470 = pi & new_n1469;
  assign new_n1471 = ~pd1 & ~pn;
  assign new_n1472 = ~pr & ~pd1;
  assign new_n1473 = ~pd1 & ~pi;
  assign new_n1474 = ~new_n1470 & ~new_n1471;
  assign new_n1475 = ~new_n1472 & ~new_n1473;
  assign new_n1476 = new_n1474 & new_n1475;
  assign py4 = ~py1 & new_n1476;
  assign new_n1478 = new_n567 & new_n645;
  assign new_n1479 = py3 & new_n1478;
  assign new_n1480 = new_n573 & new_n1479;
  assign new_n1481 = ~py3 & new_n1480;
  assign new_n1482 = ~new_n568 & new_n1480;
  assign new_n1483 = pe4 & new_n573;
  assign new_n1484 = ~new_n568 & new_n1483;
  assign new_n1485 = ~new_n570 & new_n1483;
  assign new_n1486 = ~py3 & new_n1483;
  assign new_n1487 = ~new_n570 & new_n1480;
  assign new_n1488 = ~new_n1481 & ~new_n1482;
  assign new_n1489 = ~new_n1484 & new_n1488;
  assign new_n1490 = ~new_n1485 & ~new_n1486;
  assign new_n1491 = ~new_n1487 & new_n1490;
  assign pz7 = ~new_n1489 | ~new_n1491;
  assign new_n1493 = ~pc3 & ~pf;
  assign new_n1494 = ~pd3 & ph;
  assign new_n1495 = pf & new_n1494;
  assign new_n1496 = ~new_n1493 & ~new_n1495;
  assign new_n1497 = ~py1 & new_n1496;
  assign new_n1498 = ph & new_n1497;
  assign new_n1499 = pc3 & new_n1497;
  assign px6 = new_n1498 | new_n1499;
  assign new_n1501 = py3 & new_n578;
  assign new_n1502 = pz3 & new_n1501;
  assign new_n1503 = new_n573 & new_n1502;
  assign new_n1504 = ~py3 & new_n1503;
  assign new_n1505 = ~new_n567 & new_n1503;
  assign new_n1506 = pd4 & new_n573;
  assign new_n1507 = ~new_n567 & new_n1506;
  assign new_n1508 = ~new_n1210 & new_n1506;
  assign new_n1509 = ~py3 & new_n1506;
  assign new_n1510 = ~new_n1210 & new_n1503;
  assign new_n1511 = ~new_n1504 & ~new_n1505;
  assign new_n1512 = ~new_n1507 & new_n1511;
  assign new_n1513 = ~new_n1508 & ~new_n1509;
  assign new_n1514 = ~new_n1510 & new_n1513;
  assign py7 = ~new_n1512 | ~new_n1514;
  assign new_n1516 = pr & ~po;
  assign new_n1517 = pi & new_n1516;
  assign new_n1518 = ~pe1 & ~po;
  assign new_n1519 = ~pr & ~pe1;
  assign new_n1520 = ~pe1 & ~pi;
  assign new_n1521 = ~new_n1517 & ~new_n1518;
  assign new_n1522 = ~new_n1519 & ~new_n1520;
  assign new_n1523 = new_n1521 & new_n1522;
  assign pz4 = ~py1 & new_n1523;
  assign new_n1525 = py3 & new_n577;
  assign new_n1526 = pz3 & new_n1525;
  assign new_n1527 = new_n573 & new_n1526;
  assign new_n1528 = ~pz3 & new_n1527;
  assign new_n1529 = ~py3 & new_n1527;
  assign new_n1530 = pc4 & new_n573;
  assign new_n1531 = ~py3 & new_n1530;
  assign new_n1532 = ~new_n578 & new_n1530;
  assign new_n1533 = ~pz3 & new_n1530;
  assign new_n1534 = ~new_n578 & new_n1527;
  assign new_n1535 = ~new_n1528 & ~new_n1529;
  assign new_n1536 = ~new_n1531 & new_n1535;
  assign new_n1537 = ~new_n1532 & ~new_n1533;
  assign new_n1538 = ~new_n1534 & new_n1537;
  assign px7 = ~new_n1536 | ~new_n1538;
  assign new_n1540 = ~pd3 & ~pf;
  assign new_n1541 = ~pe3 & ph;
  assign new_n1542 = pf & new_n1541;
  assign new_n1543 = ~new_n1540 & ~new_n1542;
  assign new_n1544 = ~py1 & new_n1543;
  assign new_n1545 = ph & new_n1544;
  assign new_n1546 = pd3 & new_n1544;
  assign py6 = new_n1545 | new_n1546;
  assign new_n1548 = ~pe2 & new_n509;
  assign new_n1549 = ~pn0 & new_n1548;
  assign new_n1550 = ~pa2 & pe2;
  assign new_n1551 = new_n499 & new_n1550;
  assign new_n1552 = ~pn0 & new_n1551;
  assign pz5 = new_n1549 | new_n1552;
endmodule


