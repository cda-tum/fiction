// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    _1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_,
    _259gat_55_, _36gat_6_, _55gat_9_, _75gat_15_, _159gat_40_,
    _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_,
    _153gat_38_, _59gat_10_, _207gat_48_, _261gat_57_, _88gat_20_,
    _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_,
    _116gat_28_, _130gat_31_, _246gat_53_, _89gat_21_, _111gat_27_,
    _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_,
    _143gat_34_, _201gat_47_, _267gat_58_, _101gat_25_, _171gat_42_,
    _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_,
    _87gat_19_, _165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_,
    _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_,
    _195gat_46_, _126gat_30_,
    _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_,
    _850gat_404_, _389gat_132_, _767gat_349_, _874gat_433_, _418gat_168_,
    _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_,
    _879gat_441_, _449gat_176_, _863gat_424_, _446gat_183_, _866gat_426_,
    _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_,
    _864gat_423_  );
  input  _1gat_0_, _85gat_17_, _135gat_32_, _152gat_37_, _210gat_49_,
    _259gat_55_, _36gat_6_, _55gat_9_, _75gat_15_, _159gat_40_,
    _237gat_52_, _138gat_33_, _8gat_1_, _219gat_50_, _26gat_4_, _74gat_14_,
    _153gat_38_, _59gat_10_, _207gat_48_, _261gat_57_, _88gat_20_,
    _183gat_44_, _149gat_36_, _260gat_56_, _13gat_2_, _73gat_13_,
    _116gat_28_, _130gat_31_, _246gat_53_, _89gat_21_, _111gat_27_,
    _189gat_45_, _68gat_11_, _72gat_12_, _268gat_59_, _90gat_22_,
    _143gat_34_, _201gat_47_, _267gat_58_, _101gat_25_, _171gat_42_,
    _29gat_5_, _228gat_51_, _91gat_23_, _146gat_35_, _51gat_8_, _80gat_16_,
    _87gat_19_, _165gat_41_, _255gat_54_, _156gat_39_, _177gat_43_,
    _42gat_7_, _86gat_18_, _17gat_3_, _96gat_24_, _106gat_26_, _121gat_29_,
    _195gat_46_, _126gat_30_;
  output _768gat_334_, _388gat_133_, _420gat_158_, _423gat_155_, _419gat_164_,
    _850gat_404_, _389gat_132_, _767gat_349_, _874gat_433_, _418gat_168_,
    _421gat_162_, _422gat_161_, _878gat_442_, _450gat_173_, _447gat_182_,
    _879gat_441_, _449gat_176_, _863gat_424_, _446gat_183_, _866gat_426_,
    _880gat_440_, _391gat_124_, _448gat_179_, _865gat_422_, _390gat_131_,
    _864gat_423_;
  wire new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n101, new_n102, new_n103, new_n104, new_n105, new_n106, new_n107,
    new_n108, new_n109, new_n110, new_n111, new_n112, new_n114, new_n116,
    new_n118, new_n120, new_n122, new_n123, new_n124, new_n126, new_n127,
    new_n128, new_n129, new_n130, new_n131, new_n132, new_n133, new_n134,
    new_n135, new_n136, new_n137, new_n138, new_n139, new_n140, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n179, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n265,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n337, new_n338, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n356, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n375,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n412,
    new_n413, new_n414;
  assign new_n87 = ~_201gat_47_ & ~_195gat_46_;
  assign new_n88 = _201gat_47_ & _195gat_46_;
  assign new_n89 = ~new_n87 & ~new_n88;
  assign new_n90 = ~_183gat_44_ & ~_189gat_45_;
  assign new_n91 = _183gat_44_ & _189gat_45_;
  assign new_n92 = ~new_n90 & ~new_n91;
  assign new_n93 = new_n89 & new_n92;
  assign new_n94 = ~new_n89 & ~new_n92;
  assign new_n95 = ~new_n93 & ~new_n94;
  assign new_n96 = ~_207gat_48_ & ~new_n95;
  assign new_n97 = _207gat_48_ & new_n95;
  assign new_n98 = ~new_n96 & ~new_n97;
  assign new_n99 = ~_171gat_42_ & ~_177gat_43_;
  assign new_n100 = _171gat_42_ & _177gat_43_;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = ~_159gat_40_ & ~_165gat_41_;
  assign new_n103 = _159gat_40_ & _165gat_41_;
  assign new_n104 = ~new_n102 & ~new_n103;
  assign new_n105 = new_n101 & new_n104;
  assign new_n106 = ~new_n101 & ~new_n104;
  assign new_n107 = ~new_n105 & ~new_n106;
  assign new_n108 = ~_130gat_31_ & ~new_n107;
  assign new_n109 = _130gat_31_ & new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = new_n98 & new_n110;
  assign new_n112 = ~new_n98 & ~new_n110;
  assign _768gat_334_ = ~new_n111 & ~new_n112;
  assign new_n114 = _75gat_15_ & _42gat_7_;
  assign _388gat_133_ = _29gat_5_ & new_n114;
  assign new_n116 = _75gat_15_ & _80gat_16_;
  assign _420gat_158_ = ~_59gat_10_ | ~new_n116;
  assign new_n118 = ~_88gat_20_ & ~_87gat_19_;
  assign _423gat_155_ = _90gat_22_ & ~new_n118;
  assign new_n120 = _36gat_6_ & _42gat_7_;
  assign _390gat_131_ = _29gat_5_ & new_n120;
  assign new_n122 = _26gat_4_ & _17gat_3_;
  assign new_n123 = _13gat_2_ & new_n122;
  assign new_n124 = _1gat_0_ & new_n123;
  assign _419gat_164_ = _390gat_131_ | ~new_n124;
  assign new_n126 = _72gat_12_ & _42gat_7_;
  assign new_n127 = _68gat_11_ & new_n126;
  assign new_n128 = _59gat_10_ & new_n127;
  assign new_n129 = _55gat_9_ & _8gat_1_;
  assign new_n130 = _13gat_2_ & new_n129;
  assign new_n131 = _1gat_0_ & new_n130;
  assign new_n132 = new_n128 & new_n131;
  assign new_n133 = _73gat_13_ & new_n132;
  assign new_n134 = _201gat_47_ & new_n133;
  assign new_n135 = _59gat_10_ & new_n114;
  assign new_n136 = _8gat_1_ & _17gat_3_;
  assign new_n137 = _51gat_8_ & new_n136;
  assign new_n138 = _1gat_0_ & new_n137;
  assign new_n139 = ~new_n135 & new_n138;
  assign new_n140 = _26gat_4_ & _51gat_8_;
  assign _447gat_182_ = _1gat_0_ & new_n140;
  assign new_n142 = _42gat_7_ & _17gat_3_;
  assign new_n143 = ~_42gat_7_ & ~_17gat_3_;
  assign new_n144 = ~new_n142 & ~new_n143;
  assign new_n145 = _59gat_10_ & _447gat_182_;
  assign new_n146 = _156gat_39_ & new_n145;
  assign new_n147 = new_n144 & new_n146;
  assign new_n148 = ~new_n139 & ~new_n147;
  assign new_n149 = _126gat_30_ & ~new_n148;
  assign new_n150 = _59gat_10_ & _156gat_39_;
  assign new_n151 = _17gat_3_ & ~new_n150;
  assign new_n152 = _447gat_182_ & new_n151;
  assign new_n153 = _1gat_0_ & ~new_n152;
  assign new_n154 = _153gat_38_ & ~new_n153;
  assign new_n155 = ~new_n149 & ~new_n154;
  assign new_n156 = _29gat_5_ & new_n116;
  assign new_n157 = _55gat_9_ & new_n156;
  assign new_n158 = _447gat_182_ & new_n157;
  assign new_n159 = ~_268gat_59_ & new_n158;
  assign new_n160 = new_n155 & ~new_n159;
  assign new_n161 = _201gat_47_ & ~new_n160;
  assign new_n162 = _237gat_52_ & new_n161;
  assign new_n163 = ~_201gat_47_ & new_n160;
  assign new_n164 = ~new_n161 & ~new_n163;
  assign new_n165 = _228gat_51_ & new_n164;
  assign new_n166 = ~new_n162 & ~new_n165;
  assign new_n167 = _246gat_53_ & ~new_n160;
  assign new_n168 = _267gat_58_ & _255gat_54_;
  assign new_n169 = ~new_n167 & ~new_n168;
  assign new_n170 = _261gat_57_ & new_n164;
  assign new_n171 = ~_261gat_57_ & ~new_n164;
  assign new_n172 = ~new_n170 & ~new_n171;
  assign new_n173 = _219gat_50_ & new_n172;
  assign new_n174 = _210gat_49_ & _121gat_29_;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176 = ~new_n134 & new_n166;
  assign new_n177 = new_n169 & new_n176;
  assign _850gat_404_ = ~new_n175 | ~new_n177;
  assign new_n179 = _36gat_6_ & _80gat_16_;
  assign _389gat_132_ = _29gat_5_ & new_n179;
  assign new_n181 = ~_121gat_29_ & ~_126gat_30_;
  assign new_n182 = _121gat_29_ & _126gat_30_;
  assign new_n183 = ~new_n181 & ~new_n182;
  assign new_n184 = ~_116gat_28_ & ~_111gat_27_;
  assign new_n185 = _116gat_28_ & _111gat_27_;
  assign new_n186 = ~new_n184 & ~new_n185;
  assign new_n187 = new_n183 & new_n186;
  assign new_n188 = ~new_n183 & ~new_n186;
  assign new_n189 = ~new_n187 & ~new_n188;
  assign new_n190 = ~_135gat_32_ & ~new_n189;
  assign new_n191 = _135gat_32_ & new_n189;
  assign new_n192 = ~new_n190 & ~new_n191;
  assign new_n193 = ~_101gat_25_ & ~_106gat_26_;
  assign new_n194 = _101gat_25_ & _106gat_26_;
  assign new_n195 = ~new_n193 & ~new_n194;
  assign new_n196 = ~_91gat_23_ & ~_96gat_24_;
  assign new_n197 = _91gat_23_ & _96gat_24_;
  assign new_n198 = ~new_n196 & ~new_n197;
  assign new_n199 = new_n195 & new_n198;
  assign new_n200 = ~new_n195 & ~new_n198;
  assign new_n201 = ~new_n199 & ~new_n200;
  assign new_n202 = ~_130gat_31_ & ~new_n201;
  assign new_n203 = _130gat_31_ & new_n201;
  assign new_n204 = ~new_n202 & ~new_n203;
  assign new_n205 = new_n192 & new_n204;
  assign new_n206 = ~new_n192 & ~new_n204;
  assign _767gat_349_ = ~new_n205 & ~new_n206;
  assign new_n208 = _17gat_3_ & new_n156;
  assign new_n209 = _447gat_182_ & new_n208;
  assign new_n210 = ~_268gat_59_ & new_n209;
  assign new_n211 = _55gat_9_ & _447gat_182_;
  assign new_n212 = ~new_n150 & new_n211;
  assign new_n213 = _153gat_38_ & new_n212;
  assign new_n214 = ~new_n210 & ~new_n213;
  assign new_n215 = _106gat_26_ & ~new_n148;
  assign new_n216 = _152gat_37_ & _138gat_33_;
  assign new_n217 = ~new_n215 & ~new_n216;
  assign new_n218 = new_n214 & new_n217;
  assign new_n219 = _177gat_43_ & ~new_n218;
  assign new_n220 = _237gat_52_ & new_n219;
  assign new_n221 = ~_177gat_43_ & new_n218;
  assign new_n222 = ~new_n219 & ~new_n221;
  assign new_n223 = _228gat_51_ & new_n222;
  assign new_n224 = ~new_n220 & ~new_n223;
  assign new_n225 = _177gat_43_ & new_n133;
  assign new_n226 = _246gat_53_ & ~new_n218;
  assign new_n227 = ~new_n225 & ~new_n226;
  assign new_n228 = _111gat_27_ & ~new_n148;
  assign new_n229 = _143gat_34_ & ~new_n153;
  assign new_n230 = ~new_n228 & ~new_n229;
  assign new_n231 = ~new_n159 & new_n230;
  assign new_n232 = _183gat_44_ & ~new_n231;
  assign new_n233 = _121gat_29_ & ~new_n148;
  assign new_n234 = _149gat_36_ & ~new_n153;
  assign new_n235 = ~new_n233 & ~new_n234;
  assign new_n236 = ~new_n159 & new_n235;
  assign new_n237 = ~_195gat_46_ & new_n236;
  assign new_n238 = _116gat_28_ & ~new_n148;
  assign new_n239 = _146gat_35_ & ~new_n153;
  assign new_n240 = ~new_n238 & ~new_n239;
  assign new_n241 = ~new_n159 & new_n240;
  assign new_n242 = ~_189gat_45_ & new_n241;
  assign new_n243 = _261gat_57_ & ~new_n237;
  assign new_n244 = ~new_n163 & new_n243;
  assign new_n245 = ~new_n242 & new_n244;
  assign new_n246 = _195gat_46_ & ~new_n236;
  assign new_n247 = ~new_n242 & new_n246;
  assign new_n248 = new_n161 & ~new_n237;
  assign new_n249 = ~new_n242 & new_n248;
  assign new_n250 = _189gat_45_ & ~new_n241;
  assign new_n251 = ~new_n245 & ~new_n247;
  assign new_n252 = ~new_n249 & new_n251;
  assign new_n253 = ~new_n250 & new_n252;
  assign new_n254 = ~_183gat_44_ & new_n231;
  assign new_n255 = ~new_n253 & ~new_n254;
  assign new_n256 = ~new_n232 & ~new_n255;
  assign new_n257 = new_n222 & ~new_n256;
  assign new_n258 = ~new_n222 & new_n256;
  assign new_n259 = ~new_n257 & ~new_n258;
  assign new_n260 = _219gat_50_ & new_n259;
  assign new_n261 = _210gat_49_ & _101gat_25_;
  assign new_n262 = ~new_n260 & ~new_n261;
  assign new_n263 = new_n224 & new_n227;
  assign _874gat_433_ = ~new_n262 | ~new_n263;
  assign new_n265 = _13gat_2_ & new_n136;
  assign _418gat_168_ = _1gat_0_ & new_n265;
  assign _421gat_162_ = ~_59gat_10_ | ~new_n179;
  assign _422gat_161_ = ~_59gat_10_ | ~new_n120;
  assign new_n269 = _143gat_34_ & new_n212;
  assign new_n270 = ~new_n210 & ~new_n269;
  assign new_n271 = _91gat_23_ & ~new_n148;
  assign new_n272 = _138gat_33_ & _8gat_1_;
  assign new_n273 = ~new_n271 & ~new_n272;
  assign new_n274 = new_n270 & new_n273;
  assign new_n275 = _159gat_40_ & ~new_n274;
  assign new_n276 = _237gat_52_ & new_n275;
  assign new_n277 = ~_159gat_40_ & new_n274;
  assign new_n278 = ~new_n275 & ~new_n277;
  assign new_n279 = _228gat_51_ & new_n278;
  assign new_n280 = ~new_n276 & ~new_n279;
  assign new_n281 = _159gat_40_ & new_n133;
  assign new_n282 = _246gat_53_ & ~new_n274;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = _149gat_36_ & new_n212;
  assign new_n285 = ~new_n210 & ~new_n284;
  assign new_n286 = _101gat_25_ & ~new_n148;
  assign new_n287 = _138gat_33_ & _17gat_3_;
  assign new_n288 = ~new_n286 & ~new_n287;
  assign new_n289 = new_n285 & new_n288;
  assign new_n290 = ~_171gat_42_ & new_n289;
  assign new_n291 = _146gat_35_ & new_n212;
  assign new_n292 = ~new_n210 & ~new_n291;
  assign new_n293 = _96gat_24_ & ~new_n148;
  assign new_n294 = _138gat_33_ & _51gat_8_;
  assign new_n295 = ~new_n293 & ~new_n294;
  assign new_n296 = new_n292 & new_n295;
  assign new_n297 = ~_165gat_41_ & new_n296;
  assign new_n298 = ~new_n256 & ~new_n290;
  assign new_n299 = ~new_n221 & new_n298;
  assign new_n300 = ~new_n297 & new_n299;
  assign new_n301 = _171gat_42_ & ~new_n289;
  assign new_n302 = ~new_n297 & new_n301;
  assign new_n303 = new_n219 & ~new_n290;
  assign new_n304 = ~new_n297 & new_n303;
  assign new_n305 = _165gat_41_ & ~new_n296;
  assign new_n306 = ~new_n300 & ~new_n302;
  assign new_n307 = ~new_n304 & new_n306;
  assign new_n308 = ~new_n305 & new_n307;
  assign new_n309 = new_n278 & ~new_n308;
  assign new_n310 = ~new_n278 & new_n308;
  assign new_n311 = ~new_n309 & ~new_n310;
  assign new_n312 = _219gat_50_ & new_n311;
  assign new_n313 = _210gat_49_ & _268gat_59_;
  assign new_n314 = ~new_n312 & ~new_n313;
  assign new_n315 = new_n280 & new_n283;
  assign _878gat_442_ = ~new_n314 | ~new_n315;
  assign _450gat_173_ = _89gat_21_ & ~new_n118;
  assign new_n318 = _237gat_52_ & new_n305;
  assign new_n319 = ~new_n297 & ~new_n305;
  assign new_n320 = _228gat_51_ & new_n319;
  assign new_n321 = ~new_n318 & ~new_n320;
  assign new_n322 = _165gat_41_ & new_n133;
  assign new_n323 = _246gat_53_ & ~new_n296;
  assign new_n324 = ~new_n322 & ~new_n323;
  assign new_n325 = ~new_n221 & ~new_n256;
  assign new_n326 = ~new_n290 & new_n325;
  assign new_n327 = ~new_n303 & ~new_n326;
  assign new_n328 = ~new_n301 & new_n327;
  assign new_n329 = new_n319 & ~new_n328;
  assign new_n330 = ~new_n319 & new_n328;
  assign new_n331 = ~new_n329 & ~new_n330;
  assign new_n332 = _219gat_50_ & new_n331;
  assign new_n333 = _210gat_49_ & _91gat_23_;
  assign new_n334 = ~new_n332 & ~new_n333;
  assign new_n335 = new_n321 & new_n324;
  assign _879gat_441_ = ~new_n334 | ~new_n335;
  assign new_n337 = _74gat_14_ & _68gat_11_;
  assign new_n338 = _59gat_10_ & new_n337;
  assign _449gat_176_ = new_n131 & new_n338;
  assign new_n340 = _237gat_52_ & new_n232;
  assign new_n341 = ~new_n232 & ~new_n254;
  assign new_n342 = _228gat_51_ & new_n341;
  assign new_n343 = ~new_n340 & ~new_n342;
  assign new_n344 = _183gat_44_ & new_n133;
  assign new_n345 = _246gat_53_ & ~new_n231;
  assign new_n346 = ~new_n344 & ~new_n345;
  assign new_n347 = ~new_n253 & new_n341;
  assign new_n348 = new_n253 & ~new_n341;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = _219gat_50_ & new_n349;
  assign new_n351 = _210gat_49_ & _106gat_26_;
  assign new_n352 = ~new_n350 & ~new_n351;
  assign new_n353 = new_n343 & new_n346;
  assign _863gat_424_ = ~new_n352 | ~new_n353;
  assign _446gat_183_ = ~_390gat_131_ | ~new_n124;
  assign new_n356 = ~new_n277 & ~new_n308;
  assign _866gat_426_ = new_n275 | new_n356;
  assign new_n358 = _237gat_52_ & new_n301;
  assign new_n359 = ~new_n290 & ~new_n301;
  assign new_n360 = _228gat_51_ & new_n359;
  assign new_n361 = ~new_n358 & ~new_n360;
  assign new_n362 = _171gat_42_ & new_n133;
  assign new_n363 = _246gat_53_ & ~new_n289;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = ~new_n219 & ~new_n325;
  assign new_n366 = new_n359 & ~new_n365;
  assign new_n367 = ~new_n359 & new_n365;
  assign new_n368 = ~new_n366 & ~new_n367;
  assign new_n369 = _219gat_50_ & new_n368;
  assign new_n370 = _210gat_49_ & _96gat_24_;
  assign new_n371 = ~new_n369 & ~new_n370;
  assign new_n372 = new_n361 & new_n364;
  assign _880gat_440_ = ~new_n371 | ~new_n372;
  assign _391gat_124_ = _85gat_17_ & _86gat_18_;
  assign new_n375 = _68gat_11_ & _29gat_5_;
  assign _448gat_179_ = new_n131 & new_n375;
  assign new_n377 = _195gat_46_ & new_n133;
  assign new_n378 = _237gat_52_ & new_n246;
  assign new_n379 = ~new_n237 & ~new_n246;
  assign new_n380 = _228gat_51_ & new_n379;
  assign new_n381 = ~new_n378 & ~new_n380;
  assign new_n382 = _246gat_53_ & ~new_n236;
  assign new_n383 = _260gat_56_ & _255gat_54_;
  assign new_n384 = ~new_n382 & ~new_n383;
  assign new_n385 = _261gat_57_ & ~new_n163;
  assign new_n386 = ~new_n161 & ~new_n385;
  assign new_n387 = new_n379 & ~new_n386;
  assign new_n388 = ~new_n379 & new_n386;
  assign new_n389 = ~new_n387 & ~new_n388;
  assign new_n390 = _219gat_50_ & new_n389;
  assign new_n391 = _210gat_49_ & _116gat_28_;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = ~new_n377 & new_n381;
  assign new_n394 = new_n384 & new_n393;
  assign _865gat_422_ = ~new_n392 | ~new_n394;
  assign new_n396 = _189gat_45_ & new_n133;
  assign new_n397 = _237gat_52_ & new_n250;
  assign new_n398 = ~new_n242 & ~new_n250;
  assign new_n399 = _228gat_51_ & new_n398;
  assign new_n400 = ~new_n397 & ~new_n399;
  assign new_n401 = _246gat_53_ & ~new_n241;
  assign new_n402 = _259gat_55_ & _255gat_54_;
  assign new_n403 = ~new_n401 & ~new_n402;
  assign new_n404 = ~new_n237 & new_n385;
  assign new_n405 = ~new_n248 & ~new_n404;
  assign new_n406 = ~new_n246 & new_n405;
  assign new_n407 = new_n398 & ~new_n406;
  assign new_n408 = ~new_n398 & new_n406;
  assign new_n409 = ~new_n407 & ~new_n408;
  assign new_n410 = _219gat_50_ & new_n409;
  assign new_n411 = _210gat_49_ & _111gat_27_;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign new_n413 = ~new_n396 & new_n400;
  assign new_n414 = new_n403 & new_n413;
  assign _864gat_423_ = ~new_n412 | ~new_n414;
endmodule


