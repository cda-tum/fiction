// Benchmark "top" written by ABC on Mon Nov 27 17:03:58 2023

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi084, pi085, pi086, pi087, pi088, pi089, pi090,
    pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100,
    pi106, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117,
    pi118, pi119, pi120, pi122, pi123, pi124, pi125, pi126, pi127, pi129,
    pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140,
    pi141, pi142, pi143, pi144, pi145, pi146,
    po015, po016, po017, po018, po019, po020, po021, po022, po023, po024,
    po025, po026, po027, po028, po029, po030, po031, po032, po033, po034,
    po035, po036, po037, po038, po039, po040, po041, po042, po043, po044,
    po045, po046, po047, po048, po049, po050, po051, po052, po053, po054,
    po055, po056, po057, po058, po059, po060, po061, po062, po063, po064,
    po065, po066, po067, po068, po069, po070, po071, po072, po073, po074,
    po075, po076, po077, po078, po079, po080, po081, po082, po083, po084,
    po085, po086, po087, po088, po089, po090, po091, po092, po093, po094,
    po095, po096, po097, po098, po099, po100, po101, po102, po103, po104,
    po105, po106, po107, po108, po109, po110, po111, po112, po113, po114,
    po115, po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi106, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi122, pi123, pi124, pi125, pi126, pi127,
    pi129, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po015, po016, po017, po018, po019, po020, po021, po022, po023, po024,
    po025, po026, po027, po028, po029, po030, po031, po032, po033, po034,
    po035, po036, po037, po038, po039, po040, po041, po042, po043, po044,
    po045, po046, po047, po048, po049, po050, po051, po052, po053, po054,
    po055, po056, po057, po058, po059, po060, po061, po062, po063, po064,
    po065, po066, po067, po068, po069, po070, po071, po072, po073, po074,
    po075, po076, po077, po078, po079, po080, po081, po082, po083, po084,
    po085, po086, po087, po088, po089, po090, po091, po092, po093, po094,
    po095, po096, po097, po098, po099, po100, po101, po102, po103, po104,
    po105, po106, po107, po108, po109, po110, po111, po112, po113, po114,
    po115, po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141;
  wire new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337, new_n338, new_n339, new_n340, new_n341, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n369, new_n370, new_n371, new_n372,
    new_n374, new_n375, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n392, new_n393, new_n394, new_n395, new_n397, new_n398,
    new_n399, new_n401, new_n402, new_n404, new_n405, new_n406, new_n407,
    new_n409, new_n410, new_n411, new_n412, new_n414, new_n415, new_n416,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n426, new_n427, new_n428, new_n429, new_n431, new_n432, new_n433,
    new_n434, new_n436, new_n437, new_n438, new_n439, new_n441, new_n442,
    new_n444, new_n445, new_n446, new_n448, new_n449, new_n450, new_n452,
    new_n453, new_n454, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n462, new_n463, new_n464, new_n465, new_n467, new_n468, new_n470,
    new_n471, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n805, new_n806, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n891, new_n892, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n918, new_n919, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1052, new_n1053,
    new_n1054, new_n1057, new_n1058, new_n1060, new_n1065, new_n1066;
  assign new_n264 = ~pi003 & ~pi129;
  assign new_n265 = pi000 & ~pi054;
  assign new_n266 = ~pi008 & ~pi021;
  assign new_n267 = ~pi007 & ~pi013;
  assign new_n268 = ~pi014 & new_n267;
  assign new_n269 = ~pi005 & ~pi006;
  assign new_n270 = ~pi012 & new_n269;
  assign new_n271 = new_n268 & new_n270;
  assign new_n272 = new_n266 & new_n271;
  assign new_n273 = ~pi009 & ~pi011;
  assign new_n274 = ~pi004 & ~pi019;
  assign new_n275 = ~pi018 & new_n274;
  assign new_n276 = ~pi016 & new_n275;
  assign new_n277 = ~pi017 & ~pi022;
  assign new_n278 = new_n273 & new_n277;
  assign new_n279 = new_n276 & new_n278;
  assign new_n280 = new_n272 & new_n279;
  assign new_n281 = pi054 & ~new_n280;
  assign new_n282 = pi000 & ~pi010;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = ~pi005 & ~pi022;
  assign new_n285 = new_n273 & new_n284;
  assign new_n286 = ~new_n273 & ~new_n284;
  assign new_n287 = ~pi056 & ~new_n285;
  assign new_n288 = ~new_n286 & new_n287;
  assign new_n289 = pi007 & pi013;
  assign new_n290 = new_n270 & ~new_n289;
  assign new_n291 = pi008 & ~pi021;
  assign new_n292 = pi014 & new_n267;
  assign new_n293 = ~pi008 & pi021;
  assign new_n294 = ~pi014 & ~new_n267;
  assign new_n295 = ~new_n291 & ~new_n293;
  assign new_n296 = ~new_n292 & new_n295;
  assign new_n297 = ~new_n294 & new_n296;
  assign new_n298 = ~new_n266 & ~new_n268;
  assign new_n299 = ~pi010 & new_n290;
  assign new_n300 = ~new_n298 & new_n299;
  assign new_n301 = new_n279 & ~new_n297;
  assign new_n302 = new_n300 & new_n301;
  assign new_n303 = ~new_n288 & ~new_n302;
  assign new_n304 = ~new_n283 & new_n303;
  assign new_n305 = new_n264 & ~new_n265;
  assign po015 = new_n304 | ~new_n305;
  assign new_n307 = ~pi009 & ~pi014;
  assign new_n308 = ~new_n271 & ~new_n307;
  assign new_n309 = ~pi010 & ~pi022;
  assign new_n310 = new_n264 & new_n309;
  assign new_n311 = ~pi017 & pi054;
  assign new_n312 = new_n276 & new_n311;
  assign new_n313 = ~pi011 & new_n310;
  assign new_n314 = new_n312 & new_n313;
  assign new_n315 = new_n266 & new_n314;
  assign new_n316 = ~new_n267 & new_n290;
  assign new_n317 = pi005 & pi006;
  assign new_n318 = pi012 & ~new_n269;
  assign new_n319 = new_n267 & ~new_n317;
  assign new_n320 = ~new_n270 & new_n319;
  assign new_n321 = ~new_n318 & new_n320;
  assign new_n322 = ~pi009 & ~new_n316;
  assign new_n323 = ~new_n321 & new_n322;
  assign new_n324 = ~new_n308 & new_n315;
  assign new_n325 = ~new_n323 & new_n324;
  assign new_n326 = ~pi009 & new_n271;
  assign new_n327 = new_n315 & new_n326;
  assign new_n328 = new_n311 & ~new_n327;
  assign new_n329 = ~pi001 & new_n264;
  assign new_n330 = ~new_n328 & new_n329;
  assign po016 = ~new_n325 & ~new_n330;
  assign new_n332 = ~pi045 & ~pi048;
  assign new_n333 = ~pi024 & new_n332;
  assign new_n334 = ~pi002 & ~pi015;
  assign new_n335 = ~pi020 & new_n334;
  assign new_n336 = ~pi049 & new_n335;
  assign new_n337 = new_n333 & new_n336;
  assign new_n338 = pi082 & ~new_n337;
  assign new_n339 = ~pi038 & ~pi050;
  assign new_n340 = ~pi046 & new_n339;
  assign new_n341 = ~pi041 & ~pi043;
  assign new_n342 = ~pi047 & new_n341;
  assign new_n343 = new_n340 & new_n342;
  assign new_n344 = pi082 & ~new_n343;
  assign new_n345 = ~new_n338 & ~new_n344;
  assign new_n346 = ~pi042 & ~pi044;
  assign new_n347 = ~pi040 & new_n346;
  assign new_n348 = pi082 & ~new_n347;
  assign new_n349 = pi122 & pi127;
  assign new_n350 = ~new_n338 & new_n349;
  assign new_n351 = ~new_n344 & new_n350;
  assign new_n352 = ~new_n348 & ~new_n351;
  assign new_n353 = pi082 & ~new_n339;
  assign new_n354 = new_n352 & ~new_n353;
  assign new_n355 = new_n345 & new_n354;
  assign new_n356 = ~pi129 & new_n355;
  assign new_n357 = ~pi065 & new_n356;
  assign po069 = pi129 | new_n355;
  assign new_n359 = new_n343 & new_n347;
  assign new_n360 = pi082 & new_n359;
  assign new_n361 = new_n333 & new_n360;
  assign new_n362 = ~pi049 & new_n361;
  assign new_n363 = ~new_n335 & new_n362;
  assign new_n364 = ~pi015 & new_n363;
  assign new_n365 = ~pi020 & new_n364;
  assign new_n366 = pi002 & ~new_n365;
  assign new_n367 = ~po069 & new_n366;
  assign po017 = new_n357 | new_n367;
  assign new_n369 = new_n280 & new_n309;
  assign new_n370 = ~pi061 & ~pi118;
  assign new_n371 = ~pi129 & new_n370;
  assign new_n372 = ~new_n369 & new_n371;
  assign po129 = pi123 | pi129;
  assign new_n374 = pi000 & ~pi113;
  assign new_n375 = ~po129 & new_n374;
  assign po018 = new_n372 | new_n375;
  assign new_n377 = ~pi054 & new_n264;
  assign new_n378 = pi004 & new_n377;
  assign new_n379 = new_n272 & new_n312;
  assign new_n380 = pi054 & new_n264;
  assign new_n381 = new_n273 & new_n380;
  assign new_n382 = new_n379 & new_n381;
  assign new_n383 = pi010 & ~pi022;
  assign new_n384 = new_n382 & new_n383;
  assign po019 = new_n378 | new_n384;
  assign new_n386 = pi005 & new_n377;
  assign new_n387 = ~pi029 & new_n327;
  assign new_n388 = ~pi025 & ~pi059;
  assign new_n389 = pi028 & new_n388;
  assign new_n390 = new_n387 & new_n389;
  assign po020 = new_n386 | new_n390;
  assign new_n392 = pi006 & new_n377;
  assign new_n393 = ~pi028 & new_n387;
  assign new_n394 = pi025 & ~pi059;
  assign new_n395 = new_n393 & new_n394;
  assign po021 = new_n392 | new_n395;
  assign new_n397 = new_n314 & new_n326;
  assign new_n398 = new_n291 & new_n397;
  assign new_n399 = pi007 & new_n377;
  assign po022 = new_n398 | new_n399;
  assign new_n401 = pi008 & new_n377;
  assign new_n402 = new_n293 & new_n397;
  assign po023 = new_n401 | new_n402;
  assign new_n404 = pi009 & new_n377;
  assign new_n405 = ~pi009 & pi011;
  assign new_n406 = new_n310 & new_n405;
  assign new_n407 = new_n379 & new_n406;
  assign po024 = new_n404 | new_n407;
  assign new_n409 = pi010 & new_n377;
  assign new_n410 = new_n270 & new_n315;
  assign new_n411 = ~pi009 & new_n292;
  assign new_n412 = new_n410 & new_n411;
  assign po025 = new_n409 | new_n412;
  assign new_n414 = pi011 & new_n377;
  assign new_n415 = ~pi010 & pi022;
  assign new_n416 = new_n382 & new_n415;
  assign po026 = new_n414 | new_n416;
  assign new_n418 = pi012 & new_n377;
  assign new_n419 = new_n309 & new_n381;
  assign new_n420 = new_n272 & new_n419;
  assign new_n421 = ~pi017 & new_n420;
  assign new_n422 = ~pi016 & new_n421;
  assign new_n423 = pi018 & new_n274;
  assign new_n424 = new_n422 & new_n423;
  assign po027 = new_n418 | new_n424;
  assign new_n426 = ~pi028 & pi029;
  assign new_n427 = new_n388 & new_n426;
  assign new_n428 = new_n327 & new_n427;
  assign new_n429 = pi013 & new_n377;
  assign po028 = new_n428 | new_n429;
  assign new_n431 = pi014 & new_n377;
  assign new_n432 = ~pi007 & pi013;
  assign new_n433 = new_n307 & new_n432;
  assign new_n434 = new_n410 & new_n433;
  assign po029 = new_n431 | new_n434;
  assign new_n436 = ~pi070 & new_n356;
  assign new_n437 = pi015 & ~new_n362;
  assign new_n438 = ~new_n364 & ~new_n437;
  assign new_n439 = ~po069 & ~new_n438;
  assign po030 = new_n436 | new_n439;
  assign new_n441 = pi016 & new_n377;
  assign new_n442 = pi006 & new_n325;
  assign po031 = new_n441 | new_n442;
  assign new_n444 = pi017 & new_n377;
  assign new_n445 = ~pi025 & pi059;
  assign new_n446 = new_n393 & new_n445;
  assign po032 = new_n444 | new_n446;
  assign new_n448 = pi018 & new_n377;
  assign new_n449 = pi016 & new_n275;
  assign new_n450 = new_n421 & new_n449;
  assign po033 = new_n448 | new_n450;
  assign new_n452 = pi019 & new_n377;
  assign new_n453 = pi017 & new_n276;
  assign new_n454 = new_n420 & new_n453;
  assign po034 = new_n452 | new_n454;
  assign new_n456 = pi071 & new_n355;
  assign new_n457 = ~pi020 & ~new_n355;
  assign new_n458 = ~new_n364 & ~new_n457;
  assign new_n459 = ~new_n365 & ~new_n458;
  assign new_n460 = ~pi129 & ~new_n456;
  assign po035 = ~new_n459 & new_n460;
  assign new_n462 = pi021 & new_n377;
  assign new_n463 = ~pi004 & ~pi018;
  assign new_n464 = pi019 & new_n463;
  assign new_n465 = new_n422 & new_n464;
  assign po036 = new_n462 | new_n465;
  assign new_n467 = pi022 & new_n377;
  assign new_n468 = pi005 & new_n325;
  assign po037 = new_n467 | new_n468;
  assign new_n470 = ~pi023 & pi055;
  assign new_n471 = pi061 & ~pi129;
  assign po038 = ~new_n470 & new_n471;
  assign new_n473 = new_n332 & new_n359;
  assign new_n474 = pi082 & ~new_n473;
  assign new_n475 = ~new_n350 & ~new_n474;
  assign new_n476 = ~pi024 & ~new_n475;
  assign new_n477 = pi024 & pi082;
  assign new_n478 = new_n475 & new_n477;
  assign new_n479 = new_n336 & new_n473;
  assign new_n480 = pi082 & ~new_n479;
  assign new_n481 = pi063 & ~new_n349;
  assign new_n482 = ~new_n480 & new_n481;
  assign new_n483 = ~pi129 & ~new_n476;
  assign new_n484 = ~new_n478 & ~new_n482;
  assign po039 = new_n483 & new_n484;
  assign new_n486 = pi085 & pi116;
  assign new_n487 = ~pi096 & ~pi110;
  assign new_n488 = ~pi085 & new_n487;
  assign new_n489 = ~new_n486 & ~new_n488;
  assign new_n490 = pi100 & ~new_n489;
  assign new_n491 = ~pi026 & ~pi027;
  assign new_n492 = ~pi053 & new_n491;
  assign new_n493 = ~pi053 & ~pi085;
  assign new_n494 = pi026 & pi027;
  assign new_n495 = new_n493 & ~new_n494;
  assign new_n496 = ~pi025 & ~pi116;
  assign new_n497 = new_n495 & ~new_n496;
  assign new_n498 = ~pi039 & ~pi052;
  assign new_n499 = ~pi051 & pi116;
  assign new_n500 = new_n498 & new_n499;
  assign new_n501 = pi026 & ~new_n500;
  assign new_n502 = pi027 & ~new_n500;
  assign new_n503 = ~pi026 & ~new_n502;
  assign new_n504 = pi116 & ~new_n494;
  assign new_n505 = ~new_n503 & new_n504;
  assign new_n506 = ~new_n501 & new_n505;
  assign new_n507 = new_n497 & ~new_n506;
  assign new_n508 = ~new_n492 & ~new_n507;
  assign new_n509 = ~pi095 & ~pi100;
  assign new_n510 = ~pi097 & new_n509;
  assign new_n511 = ~pi110 & ~new_n510;
  assign new_n512 = ~pi085 & new_n511;
  assign new_n513 = pi025 & ~new_n512;
  assign new_n514 = new_n491 & ~new_n513;
  assign new_n515 = ~new_n486 & ~new_n514;
  assign new_n516 = ~new_n490 & ~new_n515;
  assign new_n517 = ~new_n508 & new_n516;
  assign new_n518 = ~pi058 & new_n264;
  assign new_n519 = ~pi085 & new_n491;
  assign new_n520 = pi025 & ~pi116;
  assign new_n521 = new_n519 & new_n520;
  assign new_n522 = new_n508 & ~new_n521;
  assign new_n523 = ~new_n517 & new_n518;
  assign new_n524 = ~new_n522 & new_n523;
  assign new_n525 = ~pi058 & new_n495;
  assign new_n526 = ~new_n495 & ~new_n519;
  assign new_n527 = ~pi058 & ~new_n526;
  assign new_n528 = ~new_n492 & ~new_n527;
  assign new_n529 = new_n264 & ~new_n528;
  assign new_n530 = pi058 & ~new_n519;
  assign new_n531 = new_n529 & ~new_n530;
  assign new_n532 = ~new_n525 & new_n531;
  assign new_n533 = pi058 & pi116;
  assign new_n534 = new_n497 & ~new_n533;
  assign new_n535 = new_n532 & new_n534;
  assign po040 = new_n524 | new_n535;
  assign new_n537 = ~pi053 & ~pi058;
  assign new_n538 = new_n529 & new_n537;
  assign new_n539 = new_n490 & new_n491;
  assign new_n540 = ~new_n501 & ~new_n539;
  assign po041 = new_n538 & ~new_n540;
  assign new_n542 = ~pi100 & new_n486;
  assign new_n543 = ~pi027 & pi095;
  assign new_n544 = ~pi100 & new_n543;
  assign new_n545 = new_n487 & new_n544;
  assign new_n546 = ~new_n502 & ~new_n545;
  assign new_n547 = ~pi026 & ~pi085;
  assign new_n548 = ~new_n546 & new_n547;
  assign new_n549 = ~new_n542 & ~new_n548;
  assign po042 = new_n538 & ~new_n549;
  assign new_n551 = pi028 & ~pi116;
  assign new_n552 = ~new_n542 & ~new_n551;
  assign new_n553 = new_n532 & ~new_n552;
  assign new_n554 = ~new_n493 & ~new_n553;
  assign new_n555 = ~pi028 & ~new_n511;
  assign new_n556 = new_n511 & new_n546;
  assign new_n557 = new_n491 & ~new_n555;
  assign new_n558 = ~new_n556 & new_n557;
  assign new_n559 = ~new_n506 & ~new_n558;
  assign new_n560 = new_n518 & ~new_n559;
  assign new_n561 = ~new_n491 & ~new_n494;
  assign new_n562 = new_n518 & new_n561;
  assign new_n563 = ~new_n532 & ~new_n562;
  assign new_n564 = new_n551 & ~new_n563;
  assign new_n565 = new_n493 & ~new_n560;
  assign new_n566 = ~new_n564 & new_n565;
  assign po043 = ~new_n554 & ~new_n566;
  assign new_n568 = new_n264 & new_n519;
  assign new_n569 = new_n537 & new_n568;
  assign new_n570 = ~new_n511 & new_n569;
  assign new_n571 = ~pi116 & ~new_n569;
  assign new_n572 = new_n531 & new_n571;
  assign new_n573 = ~new_n570 & ~new_n572;
  assign new_n574 = pi029 & ~new_n573;
  assign new_n575 = ~pi053 & pi097;
  assign new_n576 = ~pi058 & new_n487;
  assign new_n577 = new_n509 & new_n576;
  assign new_n578 = ~new_n533 & ~new_n577;
  assign new_n579 = new_n568 & new_n575;
  assign new_n580 = ~new_n578 & new_n579;
  assign po044 = new_n574 | new_n580;
  assign new_n582 = ~pi106 & ~pi129;
  assign new_n583 = pi109 & new_n582;
  assign new_n584 = pi060 & new_n583;
  assign new_n585 = pi106 & ~pi129;
  assign new_n586 = pi088 & new_n585;
  assign new_n587 = ~pi109 & new_n582;
  assign new_n588 = pi030 & new_n587;
  assign new_n589 = ~new_n584 & ~new_n586;
  assign po045 = new_n588 | ~new_n589;
  assign new_n591 = pi031 & new_n587;
  assign new_n592 = pi089 & new_n585;
  assign new_n593 = pi030 & new_n583;
  assign new_n594 = ~new_n591 & ~new_n592;
  assign po046 = new_n593 | ~new_n594;
  assign new_n596 = pi032 & new_n587;
  assign new_n597 = pi099 & new_n585;
  assign new_n598 = pi031 & new_n583;
  assign new_n599 = ~new_n596 & ~new_n597;
  assign po047 = new_n598 | ~new_n599;
  assign new_n601 = pi033 & new_n587;
  assign new_n602 = pi090 & new_n585;
  assign new_n603 = pi032 & new_n583;
  assign new_n604 = ~new_n601 & ~new_n602;
  assign po048 = new_n603 | ~new_n604;
  assign new_n606 = pi034 & new_n587;
  assign new_n607 = pi091 & new_n585;
  assign new_n608 = pi033 & new_n583;
  assign new_n609 = ~new_n606 & ~new_n607;
  assign po049 = new_n608 | ~new_n609;
  assign new_n611 = pi035 & new_n587;
  assign new_n612 = pi092 & new_n585;
  assign new_n613 = pi034 & new_n583;
  assign new_n614 = ~new_n611 & ~new_n612;
  assign po050 = new_n613 | ~new_n614;
  assign new_n616 = pi036 & new_n587;
  assign new_n617 = pi098 & new_n585;
  assign new_n618 = pi035 & new_n583;
  assign new_n619 = ~new_n616 & ~new_n617;
  assign po051 = new_n618 | ~new_n619;
  assign new_n621 = pi037 & new_n587;
  assign new_n622 = pi093 & new_n585;
  assign new_n623 = pi036 & new_n583;
  assign new_n624 = ~new_n621 & ~new_n622;
  assign po052 = new_n623 | ~new_n624;
  assign new_n626 = ~pi038 & ~new_n352;
  assign new_n627 = pi038 & ~new_n345;
  assign new_n628 = pi074 & new_n345;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = new_n352 & ~new_n629;
  assign new_n631 = ~pi129 & ~new_n626;
  assign po053 = ~new_n630 & new_n631;
  assign new_n633 = ~pi051 & pi109;
  assign new_n634 = ~pi052 & new_n633;
  assign new_n635 = pi039 & ~new_n634;
  assign new_n636 = new_n498 & new_n633;
  assign new_n637 = ~pi106 & ~new_n636;
  assign new_n638 = ~new_n635 & new_n637;
  assign po054 = ~pi129 & ~new_n638;
  assign new_n640 = ~new_n338 & ~new_n349;
  assign new_n641 = pi082 & ~new_n346;
  assign new_n642 = pi073 & ~new_n641;
  assign new_n643 = ~new_n344 & new_n642;
  assign new_n644 = new_n640 & new_n643;
  assign new_n645 = ~pi040 & ~new_n352;
  assign new_n646 = pi040 & pi082;
  assign new_n647 = new_n346 & new_n646;
  assign new_n648 = ~pi129 & ~new_n647;
  assign new_n649 = ~new_n644 & new_n648;
  assign po055 = ~new_n645 & new_n649;
  assign new_n651 = new_n340 & new_n347;
  assign new_n652 = ~pi041 & new_n651;
  assign new_n653 = pi041 & ~new_n651;
  assign new_n654 = pi082 & ~new_n652;
  assign new_n655 = ~new_n653 & new_n654;
  assign new_n656 = pi076 & new_n355;
  assign new_n657 = ~pi041 & new_n351;
  assign new_n658 = ~pi129 & ~new_n655;
  assign new_n659 = ~new_n657 & new_n658;
  assign po056 = ~new_n656 & new_n659;
  assign new_n661 = pi042 & pi044;
  assign new_n662 = new_n641 & ~new_n661;
  assign new_n663 = ~pi082 & ~new_n349;
  assign new_n664 = pi042 & ~new_n663;
  assign new_n665 = ~pi072 & ~new_n349;
  assign new_n666 = ~new_n646 & ~new_n665;
  assign new_n667 = ~new_n664 & new_n666;
  assign new_n668 = new_n345 & new_n667;
  assign new_n669 = ~pi129 & ~new_n662;
  assign po057 = ~new_n668 & new_n669;
  assign new_n671 = pi077 & new_n355;
  assign new_n672 = pi043 & ~new_n652;
  assign new_n673 = ~pi043 & new_n652;
  assign new_n674 = pi082 & ~new_n673;
  assign new_n675 = ~new_n672 & new_n674;
  assign new_n676 = ~pi043 & new_n351;
  assign new_n677 = ~pi129 & ~new_n675;
  assign new_n678 = ~new_n676 & new_n677;
  assign po058 = ~new_n671 & new_n678;
  assign new_n680 = pi044 & new_n480;
  assign new_n681 = ~pi044 & new_n351;
  assign new_n682 = pi067 & new_n640;
  assign new_n683 = ~new_n681 & ~new_n682;
  assign new_n684 = ~new_n480 & ~new_n683;
  assign new_n685 = ~pi129 & ~new_n680;
  assign po059 = ~new_n684 & new_n685;
  assign new_n687 = pi068 & new_n640;
  assign new_n688 = ~pi048 & new_n360;
  assign new_n689 = pi045 & ~new_n688;
  assign new_n690 = ~new_n475 & ~new_n689;
  assign new_n691 = ~pi129 & ~new_n687;
  assign po060 = ~new_n690 & new_n691;
  assign new_n693 = ~pi046 & ~new_n354;
  assign new_n694 = pi046 & ~new_n345;
  assign new_n695 = pi075 & new_n345;
  assign new_n696 = ~new_n694 & ~new_n695;
  assign new_n697 = new_n354 & ~new_n696;
  assign new_n698 = ~pi129 & ~new_n693;
  assign po061 = ~new_n697 & new_n698;
  assign new_n700 = ~pi047 & new_n350;
  assign new_n701 = pi064 & new_n640;
  assign new_n702 = pi082 & ~new_n359;
  assign new_n703 = ~new_n701 & ~new_n702;
  assign new_n704 = pi047 & new_n674;
  assign new_n705 = ~new_n703 & ~new_n704;
  assign new_n706 = ~pi129 & ~new_n700;
  assign po062 = ~new_n705 & new_n706;
  assign new_n708 = ~new_n337 & new_n688;
  assign new_n709 = ~pi062 & new_n355;
  assign new_n710 = pi048 & ~new_n360;
  assign new_n711 = ~new_n640 & new_n710;
  assign new_n712 = ~new_n708 & ~new_n711;
  assign new_n713 = ~new_n709 & new_n712;
  assign po063 = ~pi129 & ~new_n713;
  assign new_n715 = ~pi069 & new_n355;
  assign new_n716 = pi049 & ~new_n663;
  assign new_n717 = ~new_n361 & new_n716;
  assign new_n718 = ~new_n363 & ~new_n717;
  assign new_n719 = ~new_n715 & new_n718;
  assign po064 = ~pi129 & ~new_n719;
  assign new_n721 = ~pi050 & ~new_n352;
  assign new_n722 = pi066 & new_n355;
  assign new_n723 = ~pi038 & new_n352;
  assign new_n724 = pi050 & ~new_n723;
  assign new_n725 = new_n353 & ~new_n724;
  assign new_n726 = ~pi129 & ~new_n721;
  assign new_n727 = ~new_n722 & new_n726;
  assign po065 = ~new_n725 & new_n727;
  assign new_n729 = pi051 & ~pi109;
  assign new_n730 = ~pi106 & ~new_n633;
  assign new_n731 = ~new_n729 & new_n730;
  assign po066 = ~pi129 & ~new_n731;
  assign new_n733 = pi052 & ~new_n633;
  assign new_n734 = ~pi106 & ~new_n634;
  assign new_n735 = ~new_n733 & new_n734;
  assign po067 = ~pi129 & ~new_n735;
  assign new_n737 = pi053 & new_n572;
  assign po068 = new_n580 | new_n737;
  assign new_n739 = pi114 & ~pi122;
  assign po070 = ~po129 & new_n739;
  assign new_n741 = pi026 & pi116;
  assign new_n742 = ~pi037 & ~pi058;
  assign new_n743 = ~new_n741 & new_n742;
  assign new_n744 = pi058 & ~pi116;
  assign new_n745 = ~new_n741 & ~new_n744;
  assign new_n746 = ~pi094 & ~new_n745;
  assign new_n747 = ~new_n743 & ~new_n746;
  assign po071 = new_n531 & new_n747;
  assign new_n749 = pi057 & new_n538;
  assign new_n750 = ~pi057 & ~new_n533;
  assign new_n751 = ~pi060 & new_n533;
  assign new_n752 = ~new_n750 & ~new_n751;
  assign new_n753 = new_n532 & new_n752;
  assign po072 = new_n749 | new_n753;
  assign new_n755 = new_n491 & new_n744;
  assign new_n756 = ~pi058 & new_n500;
  assign new_n757 = new_n561 & new_n756;
  assign new_n758 = ~new_n755 & ~new_n757;
  assign new_n759 = new_n264 & new_n493;
  assign po073 = ~new_n758 & new_n759;
  assign new_n761 = pi059 & new_n572;
  assign new_n762 = ~pi096 & new_n511;
  assign new_n763 = new_n492 & new_n518;
  assign new_n764 = ~pi059 & ~new_n511;
  assign new_n765 = ~new_n762 & new_n763;
  assign new_n766 = ~new_n764 & new_n765;
  assign new_n767 = new_n563 & new_n766;
  assign po074 = new_n761 | new_n767;
  assign new_n769 = ~pi117 & ~pi122;
  assign new_n770 = pi060 & ~new_n769;
  assign new_n771 = pi123 & new_n769;
  assign po075 = new_n770 | new_n771;
  assign new_n773 = ~pi114 & ~pi122;
  assign new_n774 = pi123 & ~pi129;
  assign po076 = new_n773 & new_n774;
  assign new_n776 = pi136 & ~pi138;
  assign new_n777 = ~pi137 & new_n776;
  assign new_n778 = pi132 & pi133;
  assign new_n779 = ~pi129 & pi131;
  assign new_n780 = new_n778 & new_n779;
  assign new_n781 = new_n777 & new_n780;
  assign new_n782 = ~pi140 & new_n781;
  assign new_n783 = ~pi129 & ~new_n781;
  assign new_n784 = pi062 & new_n783;
  assign po077 = ~new_n782 & ~new_n784;
  assign new_n786 = ~pi142 & new_n781;
  assign new_n787 = pi063 & new_n783;
  assign po078 = ~new_n786 & ~new_n787;
  assign new_n789 = ~pi139 & new_n781;
  assign new_n790 = pi064 & new_n783;
  assign po079 = ~new_n789 & ~new_n790;
  assign new_n792 = ~pi146 & new_n781;
  assign new_n793 = pi065 & new_n783;
  assign po080 = ~new_n792 & ~new_n793;
  assign new_n795 = ~pi136 & ~pi138;
  assign new_n796 = ~pi137 & new_n795;
  assign new_n797 = new_n780 & new_n796;
  assign new_n798 = ~pi143 & new_n797;
  assign new_n799 = ~pi129 & ~new_n797;
  assign new_n800 = pi066 & new_n799;
  assign po081 = ~new_n798 & ~new_n800;
  assign new_n802 = ~pi139 & new_n797;
  assign new_n803 = pi067 & new_n799;
  assign po082 = ~new_n802 & ~new_n803;
  assign new_n805 = ~pi141 & new_n781;
  assign new_n806 = pi068 & new_n783;
  assign po083 = ~new_n805 & ~new_n806;
  assign new_n808 = ~pi143 & new_n781;
  assign new_n809 = pi069 & new_n783;
  assign po084 = ~new_n808 & ~new_n809;
  assign new_n811 = ~pi144 & new_n781;
  assign new_n812 = pi070 & new_n783;
  assign po085 = ~new_n811 & ~new_n812;
  assign new_n814 = ~pi145 & new_n781;
  assign new_n815 = pi071 & new_n783;
  assign po086 = ~new_n814 & ~new_n815;
  assign new_n817 = ~pi140 & new_n797;
  assign new_n818 = pi072 & new_n799;
  assign po087 = ~new_n817 & ~new_n818;
  assign new_n820 = ~pi141 & new_n797;
  assign new_n821 = pi073 & new_n799;
  assign po088 = ~new_n820 & ~new_n821;
  assign new_n823 = ~pi142 & new_n797;
  assign new_n824 = pi074 & new_n799;
  assign po089 = ~new_n823 & ~new_n824;
  assign new_n826 = ~pi144 & new_n797;
  assign new_n827 = pi075 & new_n799;
  assign po090 = ~new_n826 & ~new_n827;
  assign new_n829 = ~pi145 & new_n797;
  assign new_n830 = pi076 & new_n799;
  assign po091 = ~new_n829 & ~new_n830;
  assign new_n832 = ~pi146 & new_n797;
  assign new_n833 = pi077 & new_n799;
  assign po092 = ~new_n832 & ~new_n833;
  assign new_n835 = ~pi136 & pi137;
  assign new_n836 = ~pi138 & new_n835;
  assign new_n837 = new_n780 & new_n836;
  assign new_n838 = pi142 & new_n837;
  assign new_n839 = ~pi129 & ~new_n837;
  assign new_n840 = pi078 & new_n839;
  assign po093 = new_n838 | new_n840;
  assign new_n842 = pi143 & new_n837;
  assign new_n843 = pi079 & new_n839;
  assign po094 = new_n842 | new_n843;
  assign new_n845 = pi144 & new_n837;
  assign new_n846 = pi080 & new_n839;
  assign po095 = new_n845 | new_n846;
  assign new_n848 = pi145 & new_n837;
  assign new_n849 = pi081 & new_n839;
  assign po096 = new_n848 | new_n849;
  assign new_n851 = pi146 & new_n837;
  assign new_n852 = pi082 & new_n839;
  assign po097 = new_n851 | new_n852;
  assign new_n854 = pi072 & new_n796;
  assign new_n855 = pi087 & new_n795;
  assign new_n856 = pi031 & new_n776;
  assign new_n857 = ~pi136 & pi138;
  assign new_n858 = ~pi115 & new_n857;
  assign new_n859 = pi137 & ~new_n855;
  assign new_n860 = ~new_n856 & ~new_n858;
  assign new_n861 = new_n859 & new_n860;
  assign new_n862 = pi136 & pi138;
  assign new_n863 = ~pi089 & new_n862;
  assign new_n864 = ~pi137 & new_n857;
  assign new_n865 = ~pi119 & new_n864;
  assign new_n866 = pi062 & new_n777;
  assign new_n867 = ~new_n854 & ~new_n863;
  assign new_n868 = ~new_n865 & ~new_n866;
  assign new_n869 = new_n867 & new_n868;
  assign po098 = ~new_n861 & new_n869;
  assign new_n871 = pi141 & new_n837;
  assign new_n872 = pi084 & new_n839;
  assign po099 = new_n871 | new_n872;
  assign new_n874 = new_n489 & new_n763;
  assign po100 = ~new_n570 & new_n874;
  assign new_n876 = pi139 & new_n837;
  assign new_n877 = pi086 & new_n839;
  assign po101 = new_n876 | new_n877;
  assign new_n879 = pi140 & new_n837;
  assign new_n880 = pi087 & new_n839;
  assign po102 = new_n879 | new_n880;
  assign new_n882 = pi137 & new_n776;
  assign new_n883 = new_n780 & new_n882;
  assign new_n884 = pi139 & new_n883;
  assign new_n885 = ~pi129 & ~new_n883;
  assign new_n886 = pi088 & new_n885;
  assign po103 = new_n884 | new_n886;
  assign new_n888 = pi140 & new_n883;
  assign new_n889 = pi089 & new_n885;
  assign po104 = new_n888 | new_n889;
  assign new_n891 = pi142 & new_n883;
  assign new_n892 = pi090 & new_n885;
  assign po105 = new_n891 | new_n892;
  assign new_n894 = pi143 & new_n883;
  assign new_n895 = pi091 & new_n885;
  assign po106 = new_n894 | new_n895;
  assign new_n897 = pi144 & new_n883;
  assign new_n898 = pi092 & new_n885;
  assign po107 = new_n897 | new_n898;
  assign new_n900 = pi146 & new_n883;
  assign new_n901 = pi093 & new_n885;
  assign po108 = new_n900 | new_n901;
  assign new_n903 = pi082 & new_n864;
  assign new_n904 = new_n780 & new_n903;
  assign new_n905 = pi142 & new_n904;
  assign new_n906 = ~pi129 & ~new_n904;
  assign new_n907 = pi094 & new_n906;
  assign po109 = new_n905 | new_n907;
  assign new_n909 = pi143 & new_n904;
  assign new_n910 = ~pi003 & ~pi110;
  assign new_n911 = ~new_n780 & ~new_n910;
  assign new_n912 = new_n906 & ~new_n911;
  assign new_n913 = pi095 & new_n912;
  assign po110 = new_n909 | new_n913;
  assign new_n915 = pi146 & new_n904;
  assign new_n916 = pi096 & new_n912;
  assign po111 = new_n915 | new_n916;
  assign new_n918 = pi145 & new_n904;
  assign new_n919 = pi097 & new_n912;
  assign po112 = new_n918 | new_n919;
  assign new_n921 = pi145 & new_n883;
  assign new_n922 = pi098 & new_n885;
  assign po113 = new_n921 | new_n922;
  assign new_n924 = pi141 & new_n883;
  assign new_n925 = pi099 & new_n885;
  assign po114 = new_n924 | new_n925;
  assign new_n927 = pi144 & new_n904;
  assign new_n928 = pi100 & new_n912;
  assign po115 = new_n927 | new_n928;
  assign new_n930 = pi077 & new_n796;
  assign new_n931 = pi096 & new_n857;
  assign new_n932 = pi037 & new_n776;
  assign new_n933 = pi137 & ~new_n932;
  assign new_n934 = pi065 & new_n777;
  assign new_n935 = ~new_n933 & ~new_n934;
  assign new_n936 = pi082 & new_n795;
  assign new_n937 = ~new_n931 & ~new_n936;
  assign new_n938 = ~new_n935 & new_n937;
  assign new_n939 = ~pi093 & new_n862;
  assign new_n940 = ~pi124 & new_n864;
  assign new_n941 = ~new_n930 & ~new_n939;
  assign new_n942 = ~new_n940 & new_n941;
  assign po116 = ~new_n938 & new_n942;
  assign new_n944 = ~pi069 & new_n777;
  assign new_n945 = pi034 & new_n882;
  assign new_n946 = ~pi066 & new_n796;
  assign new_n947 = ~pi137 & new_n862;
  assign new_n948 = pi091 & new_n947;
  assign new_n949 = ~pi079 & ~pi138;
  assign new_n950 = ~pi095 & pi138;
  assign new_n951 = new_n835 & ~new_n949;
  assign new_n952 = ~new_n950 & new_n951;
  assign new_n953 = ~new_n944 & ~new_n945;
  assign new_n954 = ~new_n946 & ~new_n948;
  assign new_n955 = ~new_n952 & new_n954;
  assign po117 = ~new_n953 | ~new_n955;
  assign new_n957 = pi033 & new_n882;
  assign new_n958 = ~pi063 & new_n777;
  assign new_n959 = ~pi074 & new_n796;
  assign new_n960 = pi090 & new_n947;
  assign new_n961 = ~pi078 & ~pi138;
  assign new_n962 = ~pi094 & pi138;
  assign new_n963 = new_n835 & ~new_n961;
  assign new_n964 = ~new_n962 & new_n963;
  assign new_n965 = ~new_n957 & ~new_n958;
  assign new_n966 = ~new_n959 & ~new_n960;
  assign new_n967 = ~new_n964 & new_n966;
  assign po118 = ~new_n965 | ~new_n967;
  assign new_n969 = ~pi073 & new_n796;
  assign new_n970 = ~pi112 & new_n857;
  assign new_n971 = pi084 & new_n795;
  assign new_n972 = ~new_n970 & ~new_n971;
  assign new_n973 = pi137 & ~new_n972;
  assign new_n974 = ~pi068 & new_n777;
  assign new_n975 = pi099 & new_n947;
  assign new_n976 = pi032 & new_n882;
  assign new_n977 = ~new_n969 & ~new_n974;
  assign new_n978 = ~new_n975 & ~new_n976;
  assign new_n979 = new_n977 & new_n978;
  assign po119 = new_n973 | ~new_n979;
  assign new_n981 = pi075 & new_n796;
  assign new_n982 = pi080 & new_n795;
  assign new_n983 = pi035 & new_n776;
  assign new_n984 = pi100 & new_n857;
  assign new_n985 = pi137 & ~new_n982;
  assign new_n986 = ~new_n983 & ~new_n984;
  assign new_n987 = new_n985 & new_n986;
  assign new_n988 = ~pi092 & new_n862;
  assign new_n989 = ~pi125 & new_n864;
  assign new_n990 = pi070 & new_n777;
  assign new_n991 = ~new_n981 & ~new_n988;
  assign new_n992 = ~new_n989 & ~new_n990;
  assign new_n993 = new_n991 & new_n992;
  assign po120 = ~new_n987 & new_n993;
  assign new_n995 = new_n511 & new_n569;
  assign new_n996 = pi116 & new_n264;
  assign new_n997 = pi085 & new_n996;
  assign po121 = new_n995 | new_n997;
  assign new_n999 = pi076 & new_n796;
  assign new_n1000 = pi081 & new_n795;
  assign new_n1001 = ~pi098 & new_n862;
  assign new_n1002 = ~pi137 & ~new_n1001;
  assign new_n1003 = pi097 & new_n857;
  assign new_n1004 = pi036 & new_n776;
  assign new_n1005 = ~new_n1000 & ~new_n1003;
  assign new_n1006 = ~new_n1004 & new_n1005;
  assign new_n1007 = ~new_n1002 & new_n1006;
  assign new_n1008 = ~pi023 & new_n864;
  assign new_n1009 = pi071 & new_n777;
  assign new_n1010 = ~new_n999 & ~new_n1008;
  assign new_n1011 = ~new_n1009 & new_n1010;
  assign po122 = ~new_n1007 & new_n1011;
  assign new_n1013 = pi067 & new_n796;
  assign new_n1014 = pi086 & new_n795;
  assign new_n1015 = pi030 & new_n776;
  assign new_n1016 = pi111 & new_n857;
  assign new_n1017 = pi137 & ~new_n1014;
  assign new_n1018 = ~new_n1015 & ~new_n1016;
  assign new_n1019 = new_n1017 & new_n1018;
  assign new_n1020 = ~pi088 & new_n862;
  assign new_n1021 = ~pi120 & new_n864;
  assign new_n1022 = pi064 & new_n777;
  assign new_n1023 = ~new_n1013 & ~new_n1020;
  assign new_n1024 = ~new_n1021 & ~new_n1022;
  assign new_n1025 = new_n1023 & new_n1024;
  assign po123 = ~new_n1019 & new_n1025;
  assign po124 = new_n264 & new_n505;
  assign new_n1028 = pi053 & pi058;
  assign new_n1029 = ~new_n537 & ~new_n575;
  assign new_n1030 = ~new_n1028 & new_n1029;
  assign po125 = new_n996 & new_n1030;
  assign new_n1032 = pi139 & new_n904;
  assign new_n1033 = new_n780 & ~new_n903;
  assign new_n1034 = pi111 & new_n1033;
  assign po126 = new_n1032 | new_n1034;
  assign new_n1036 = pi141 & new_n904;
  assign new_n1037 = ~pi112 & new_n1033;
  assign po127 = new_n1036 | new_n1037;
  assign new_n1039 = ~pi054 & pi113;
  assign new_n1040 = ~pi011 & ~pi022;
  assign new_n1041 = pi054 & new_n1040;
  assign new_n1042 = new_n264 & ~new_n1039;
  assign po128 = ~new_n1041 & new_n1042;
  assign new_n1044 = pi140 & new_n904;
  assign new_n1045 = ~pi115 & new_n1033;
  assign po130 = new_n1044 | new_n1045;
  assign new_n1047 = ~pi004 & ~pi007;
  assign new_n1048 = ~pi009 & ~pi012;
  assign new_n1049 = new_n1047 & new_n1048;
  assign po131 = new_n380 & ~new_n1049;
  assign po132 = ~pi122 | pi129;
  assign new_n1052 = ~pi054 & ~pi118;
  assign new_n1053 = pi054 & ~new_n427;
  assign new_n1054 = ~pi129 & ~new_n1052;
  assign po133 = ~new_n1053 & new_n1054;
  assign po134 = ~pi129 & ~new_n509;
  assign new_n1057 = ~pi120 & new_n910;
  assign new_n1058 = ~pi111 & ~pi129;
  assign po135 = ~new_n1057 & new_n1058;
  assign new_n1060 = pi081 & pi120;
  assign po136 = ~pi129 & new_n1060;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi057 & ~pi129;
  assign new_n1065 = ~pi096 & pi125;
  assign new_n1066 = ~pi003 & ~new_n1065;
  assign po140 = ~pi129 & ~new_n1066;
  assign po141 = ~pi126 & new_n778;
endmodule


