// Benchmark "b17" written by ABC on Wed Sep  5 10:17:20 2018

module b17 ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P3_DATAO_REG_31_, P3_DATAO_REG_30_, P3_DATAO_REG_29_, P3_DATAO_REG_28_,
    P3_DATAO_REG_27_, P3_DATAO_REG_26_, P3_DATAO_REG_25_, P3_DATAO_REG_24_,
    P3_DATAO_REG_23_, P3_DATAO_REG_22_, P3_DATAO_REG_21_, P3_DATAO_REG_20_,
    P3_DATAO_REG_19_, P3_DATAO_REG_18_, P3_DATAO_REG_17_, P3_DATAO_REG_16_,
    P3_DATAO_REG_15_, P3_DATAO_REG_14_, P3_DATAO_REG_13_, P3_DATAO_REG_12_,
    P3_DATAO_REG_11_, P3_DATAO_REG_10_, P3_DATAO_REG_9_, P3_DATAO_REG_8_,
    P3_DATAO_REG_7_, P3_DATAO_REG_6_, P3_DATAO_REG_5_, P3_DATAO_REG_4_,
    P3_DATAO_REG_3_, P3_DATAO_REG_2_, P3_DATAO_REG_1_, P3_DATAO_REG_0_,
    P1_ADDRESS_REG_29_, P1_ADDRESS_REG_28_, P1_ADDRESS_REG_27_,
    P1_ADDRESS_REG_26_, P1_ADDRESS_REG_25_, P1_ADDRESS_REG_24_,
    P1_ADDRESS_REG_23_, P1_ADDRESS_REG_22_, P1_ADDRESS_REG_21_,
    P1_ADDRESS_REG_20_, P1_ADDRESS_REG_19_, P1_ADDRESS_REG_18_,
    P1_ADDRESS_REG_17_, P1_ADDRESS_REG_16_, P1_ADDRESS_REG_15_,
    P1_ADDRESS_REG_14_, P1_ADDRESS_REG_13_, P1_ADDRESS_REG_12_,
    P1_ADDRESS_REG_11_, P1_ADDRESS_REG_10_, P1_ADDRESS_REG_9_,
    P1_ADDRESS_REG_8_, P1_ADDRESS_REG_7_, P1_ADDRESS_REG_6_,
    P1_ADDRESS_REG_5_, P1_ADDRESS_REG_4_, P1_ADDRESS_REG_3_,
    P1_ADDRESS_REG_2_, P1_ADDRESS_REG_1_, P1_ADDRESS_REG_0_, U355, U356,
    U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369,
    U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352,
    U353, U354, U365, U376, P3_W_R_N_REG, P3_D_C_N_REG, P3_M_IO_N_REG,
    P1_ADS_N_REG, P3_ADS_N_REG  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2;
  output P3_DATAO_REG_31_, P3_DATAO_REG_30_, P3_DATAO_REG_29_,
    P3_DATAO_REG_28_, P3_DATAO_REG_27_, P3_DATAO_REG_26_, P3_DATAO_REG_25_,
    P3_DATAO_REG_24_, P3_DATAO_REG_23_, P3_DATAO_REG_22_, P3_DATAO_REG_21_,
    P3_DATAO_REG_20_, P3_DATAO_REG_19_, P3_DATAO_REG_18_, P3_DATAO_REG_17_,
    P3_DATAO_REG_16_, P3_DATAO_REG_15_, P3_DATAO_REG_14_, P3_DATAO_REG_13_,
    P3_DATAO_REG_12_, P3_DATAO_REG_11_, P3_DATAO_REG_10_, P3_DATAO_REG_9_,
    P3_DATAO_REG_8_, P3_DATAO_REG_7_, P3_DATAO_REG_6_, P3_DATAO_REG_5_,
    P3_DATAO_REG_4_, P3_DATAO_REG_3_, P3_DATAO_REG_2_, P3_DATAO_REG_1_,
    P3_DATAO_REG_0_, P1_ADDRESS_REG_29_, P1_ADDRESS_REG_28_,
    P1_ADDRESS_REG_27_, P1_ADDRESS_REG_26_, P1_ADDRESS_REG_25_,
    P1_ADDRESS_REG_24_, P1_ADDRESS_REG_23_, P1_ADDRESS_REG_22_,
    P1_ADDRESS_REG_21_, P1_ADDRESS_REG_20_, P1_ADDRESS_REG_19_,
    P1_ADDRESS_REG_18_, P1_ADDRESS_REG_17_, P1_ADDRESS_REG_16_,
    P1_ADDRESS_REG_15_, P1_ADDRESS_REG_14_, P1_ADDRESS_REG_13_,
    P1_ADDRESS_REG_12_, P1_ADDRESS_REG_11_, P1_ADDRESS_REG_10_,
    P1_ADDRESS_REG_9_, P1_ADDRESS_REG_8_, P1_ADDRESS_REG_7_,
    P1_ADDRESS_REG_6_, P1_ADDRESS_REG_5_, P1_ADDRESS_REG_4_,
    P1_ADDRESS_REG_3_, P1_ADDRESS_REG_2_, P1_ADDRESS_REG_1_,
    P1_ADDRESS_REG_0_, U355, U356, U357, U358, U359, U360, U361, U362,
    U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, U375,
    U347, U348, U349, U350, U351, U352, U353, U354, U365, U376,
    P3_W_R_N_REG, P3_D_C_N_REG, P3_M_IO_N_REG, P1_ADS_N_REG, P3_ADS_N_REG;
  reg BUF1_REG_0_, BUF1_REG_1_, BUF1_REG_2_, BUF1_REG_3_, BUF1_REG_4_,
    BUF1_REG_5_, BUF1_REG_6_, BUF1_REG_7_, BUF1_REG_8_, BUF1_REG_9_,
    BUF1_REG_10_, BUF1_REG_11_, BUF1_REG_12_, BUF1_REG_13_, BUF1_REG_14_,
    BUF1_REG_15_, BUF1_REG_16_, BUF1_REG_17_, BUF1_REG_18_, BUF1_REG_19_,
    BUF1_REG_20_, BUF1_REG_21_, BUF1_REG_22_, BUF1_REG_23_, BUF1_REG_24_,
    BUF1_REG_25_, BUF1_REG_26_, BUF1_REG_27_, BUF1_REG_28_, BUF1_REG_29_,
    BUF1_REG_30_, BUF1_REG_31_, BUF2_REG_0_, BUF2_REG_1_, BUF2_REG_2_,
    BUF2_REG_3_, BUF2_REG_4_, BUF2_REG_5_, BUF2_REG_6_, BUF2_REG_7_,
    BUF2_REG_8_, BUF2_REG_9_, BUF2_REG_10_, BUF2_REG_11_, BUF2_REG_12_,
    BUF2_REG_13_, BUF2_REG_14_, BUF2_REG_15_, BUF2_REG_16_, BUF2_REG_17_,
    BUF2_REG_18_, BUF2_REG_19_, BUF2_REG_20_, BUF2_REG_21_, BUF2_REG_22_,
    BUF2_REG_23_, BUF2_REG_24_, BUF2_REG_25_, BUF2_REG_26_, BUF2_REG_27_,
    BUF2_REG_28_, BUF2_REG_29_, BUF2_REG_30_, BUF2_REG_31_, READY12_REG,
    READY21_REG, READY22_REG, READY11_REG, P3_BE_N_REG_3_, P3_BE_N_REG_2_,
    P3_BE_N_REG_1_, P3_BE_N_REG_0_, P3_ADDRESS_REG_29_, P3_ADDRESS_REG_28_,
    P3_ADDRESS_REG_27_, P3_ADDRESS_REG_26_, P3_ADDRESS_REG_25_,
    P3_ADDRESS_REG_24_, P3_ADDRESS_REG_23_, P3_ADDRESS_REG_22_,
    P3_ADDRESS_REG_21_, P3_ADDRESS_REG_20_, P3_ADDRESS_REG_19_,
    P3_ADDRESS_REG_18_, P3_ADDRESS_REG_17_, P3_ADDRESS_REG_16_,
    P3_ADDRESS_REG_15_, P3_ADDRESS_REG_14_, P3_ADDRESS_REG_13_,
    P3_ADDRESS_REG_12_, P3_ADDRESS_REG_11_, P3_ADDRESS_REG_10_,
    P3_ADDRESS_REG_9_, P3_ADDRESS_REG_8_, P3_ADDRESS_REG_7_,
    P3_ADDRESS_REG_6_, P3_ADDRESS_REG_5_, P3_ADDRESS_REG_4_,
    P3_ADDRESS_REG_3_, P3_ADDRESS_REG_2_, P3_ADDRESS_REG_1_,
    P3_ADDRESS_REG_0_, P3_STATE_REG_2_, P3_STATE_REG_1_, P3_STATE_REG_0_,
    P3_DATAWIDTH_REG_0_, P3_DATAWIDTH_REG_1_, P3_DATAWIDTH_REG_2_,
    P3_DATAWIDTH_REG_3_, P3_DATAWIDTH_REG_4_, P3_DATAWIDTH_REG_5_,
    P3_DATAWIDTH_REG_6_, P3_DATAWIDTH_REG_7_, P3_DATAWIDTH_REG_8_,
    P3_DATAWIDTH_REG_9_, P3_DATAWIDTH_REG_10_, P3_DATAWIDTH_REG_11_,
    P3_DATAWIDTH_REG_12_, P3_DATAWIDTH_REG_13_, P3_DATAWIDTH_REG_14_,
    P3_DATAWIDTH_REG_15_, P3_DATAWIDTH_REG_16_, P3_DATAWIDTH_REG_17_,
    P3_DATAWIDTH_REG_18_, P3_DATAWIDTH_REG_19_, P3_DATAWIDTH_REG_20_,
    P3_DATAWIDTH_REG_21_, P3_DATAWIDTH_REG_22_, P3_DATAWIDTH_REG_23_,
    P3_DATAWIDTH_REG_24_, P3_DATAWIDTH_REG_25_, P3_DATAWIDTH_REG_26_,
    P3_DATAWIDTH_REG_27_, P3_DATAWIDTH_REG_28_, P3_DATAWIDTH_REG_29_,
    P3_DATAWIDTH_REG_30_, P3_DATAWIDTH_REG_31_, P3_STATE2_REG_3_,
    P3_STATE2_REG_2_, P3_STATE2_REG_1_, P3_STATE2_REG_0_,
    P3_INSTQUEUE_REG_15__7_, P3_INSTQUEUE_REG_15__6_,
    P3_INSTQUEUE_REG_15__5_, P3_INSTQUEUE_REG_15__4_,
    P3_INSTQUEUE_REG_15__3_, P3_INSTQUEUE_REG_15__2_,
    P3_INSTQUEUE_REG_15__1_, P3_INSTQUEUE_REG_15__0_,
    P3_INSTQUEUE_REG_14__7_, P3_INSTQUEUE_REG_14__6_,
    P3_INSTQUEUE_REG_14__5_, P3_INSTQUEUE_REG_14__4_,
    P3_INSTQUEUE_REG_14__3_, P3_INSTQUEUE_REG_14__2_,
    P3_INSTQUEUE_REG_14__1_, P3_INSTQUEUE_REG_14__0_,
    P3_INSTQUEUE_REG_13__7_, P3_INSTQUEUE_REG_13__6_,
    P3_INSTQUEUE_REG_13__5_, P3_INSTQUEUE_REG_13__4_,
    P3_INSTQUEUE_REG_13__3_, P3_INSTQUEUE_REG_13__2_,
    P3_INSTQUEUE_REG_13__1_, P3_INSTQUEUE_REG_13__0_,
    P3_INSTQUEUE_REG_12__7_, P3_INSTQUEUE_REG_12__6_,
    P3_INSTQUEUE_REG_12__5_, P3_INSTQUEUE_REG_12__4_,
    P3_INSTQUEUE_REG_12__3_, P3_INSTQUEUE_REG_12__2_,
    P3_INSTQUEUE_REG_12__1_, P3_INSTQUEUE_REG_12__0_,
    P3_INSTQUEUE_REG_11__7_, P3_INSTQUEUE_REG_11__6_,
    P3_INSTQUEUE_REG_11__5_, P3_INSTQUEUE_REG_11__4_,
    P3_INSTQUEUE_REG_11__3_, P3_INSTQUEUE_REG_11__2_,
    P3_INSTQUEUE_REG_11__1_, P3_INSTQUEUE_REG_11__0_,
    P3_INSTQUEUE_REG_10__7_, P3_INSTQUEUE_REG_10__6_,
    P3_INSTQUEUE_REG_10__5_, P3_INSTQUEUE_REG_10__4_,
    P3_INSTQUEUE_REG_10__3_, P3_INSTQUEUE_REG_10__2_,
    P3_INSTQUEUE_REG_10__1_, P3_INSTQUEUE_REG_10__0_,
    P3_INSTQUEUE_REG_9__7_, P3_INSTQUEUE_REG_9__6_, P3_INSTQUEUE_REG_9__5_,
    P3_INSTQUEUE_REG_9__4_, P3_INSTQUEUE_REG_9__3_, P3_INSTQUEUE_REG_9__2_,
    P3_INSTQUEUE_REG_9__1_, P3_INSTQUEUE_REG_9__0_, P3_INSTQUEUE_REG_8__7_,
    P3_INSTQUEUE_REG_8__6_, P3_INSTQUEUE_REG_8__5_, P3_INSTQUEUE_REG_8__4_,
    P3_INSTQUEUE_REG_8__3_, P3_INSTQUEUE_REG_8__2_, P3_INSTQUEUE_REG_8__1_,
    P3_INSTQUEUE_REG_8__0_, P3_INSTQUEUE_REG_7__7_, P3_INSTQUEUE_REG_7__6_,
    P3_INSTQUEUE_REG_7__5_, P3_INSTQUEUE_REG_7__4_, P3_INSTQUEUE_REG_7__3_,
    P3_INSTQUEUE_REG_7__2_, P3_INSTQUEUE_REG_7__1_, P3_INSTQUEUE_REG_7__0_,
    P3_INSTQUEUE_REG_6__7_, P3_INSTQUEUE_REG_6__6_, P3_INSTQUEUE_REG_6__5_,
    P3_INSTQUEUE_REG_6__4_, P3_INSTQUEUE_REG_6__3_, P3_INSTQUEUE_REG_6__2_,
    P3_INSTQUEUE_REG_6__1_, P3_INSTQUEUE_REG_6__0_, P3_INSTQUEUE_REG_5__7_,
    P3_INSTQUEUE_REG_5__6_, P3_INSTQUEUE_REG_5__5_, P3_INSTQUEUE_REG_5__4_,
    P3_INSTQUEUE_REG_5__3_, P3_INSTQUEUE_REG_5__2_, P3_INSTQUEUE_REG_5__1_,
    P3_INSTQUEUE_REG_5__0_, P3_INSTQUEUE_REG_4__7_, P3_INSTQUEUE_REG_4__6_,
    P3_INSTQUEUE_REG_4__5_, P3_INSTQUEUE_REG_4__4_, P3_INSTQUEUE_REG_4__3_,
    P3_INSTQUEUE_REG_4__2_, P3_INSTQUEUE_REG_4__1_, P3_INSTQUEUE_REG_4__0_,
    P3_INSTQUEUE_REG_3__7_, P3_INSTQUEUE_REG_3__6_, P3_INSTQUEUE_REG_3__5_,
    P3_INSTQUEUE_REG_3__4_, P3_INSTQUEUE_REG_3__3_, P3_INSTQUEUE_REG_3__2_,
    P3_INSTQUEUE_REG_3__1_, P3_INSTQUEUE_REG_3__0_, P3_INSTQUEUE_REG_2__7_,
    P3_INSTQUEUE_REG_2__6_, P3_INSTQUEUE_REG_2__5_, P3_INSTQUEUE_REG_2__4_,
    P3_INSTQUEUE_REG_2__3_, P3_INSTQUEUE_REG_2__2_, P3_INSTQUEUE_REG_2__1_,
    P3_INSTQUEUE_REG_2__0_, P3_INSTQUEUE_REG_1__7_, P3_INSTQUEUE_REG_1__6_,
    P3_INSTQUEUE_REG_1__5_, P3_INSTQUEUE_REG_1__4_, P3_INSTQUEUE_REG_1__3_,
    P3_INSTQUEUE_REG_1__2_, P3_INSTQUEUE_REG_1__1_, P3_INSTQUEUE_REG_1__0_,
    P3_INSTQUEUE_REG_0__7_, P3_INSTQUEUE_REG_0__6_, P3_INSTQUEUE_REG_0__5_,
    P3_INSTQUEUE_REG_0__4_, P3_INSTQUEUE_REG_0__3_, P3_INSTQUEUE_REG_0__2_,
    P3_INSTQUEUE_REG_0__1_, P3_INSTQUEUE_REG_0__0_,
    P3_INSTQUEUERD_ADDR_REG_4_, P3_INSTQUEUERD_ADDR_REG_3_,
    P3_INSTQUEUERD_ADDR_REG_2_, P3_INSTQUEUERD_ADDR_REG_1_,
    P3_INSTQUEUERD_ADDR_REG_0_, P3_INSTQUEUEWR_ADDR_REG_4_,
    P3_INSTQUEUEWR_ADDR_REG_3_, P3_INSTQUEUEWR_ADDR_REG_2_,
    P3_INSTQUEUEWR_ADDR_REG_1_, P3_INSTQUEUEWR_ADDR_REG_0_,
    P3_INSTADDRPOINTER_REG_0_, P3_INSTADDRPOINTER_REG_1_,
    P3_INSTADDRPOINTER_REG_2_, P3_INSTADDRPOINTER_REG_3_,
    P3_INSTADDRPOINTER_REG_4_, P3_INSTADDRPOINTER_REG_5_,
    P3_INSTADDRPOINTER_REG_6_, P3_INSTADDRPOINTER_REG_7_,
    P3_INSTADDRPOINTER_REG_8_, P3_INSTADDRPOINTER_REG_9_,
    P3_INSTADDRPOINTER_REG_10_, P3_INSTADDRPOINTER_REG_11_,
    P3_INSTADDRPOINTER_REG_12_, P3_INSTADDRPOINTER_REG_13_,
    P3_INSTADDRPOINTER_REG_14_, P3_INSTADDRPOINTER_REG_15_,
    P3_INSTADDRPOINTER_REG_16_, P3_INSTADDRPOINTER_REG_17_,
    P3_INSTADDRPOINTER_REG_18_, P3_INSTADDRPOINTER_REG_19_,
    P3_INSTADDRPOINTER_REG_20_, P3_INSTADDRPOINTER_REG_21_,
    P3_INSTADDRPOINTER_REG_22_, P3_INSTADDRPOINTER_REG_23_,
    P3_INSTADDRPOINTER_REG_24_, P3_INSTADDRPOINTER_REG_25_,
    P3_INSTADDRPOINTER_REG_26_, P3_INSTADDRPOINTER_REG_27_,
    P3_INSTADDRPOINTER_REG_28_, P3_INSTADDRPOINTER_REG_29_,
    P3_INSTADDRPOINTER_REG_30_, P3_INSTADDRPOINTER_REG_31_,
    P3_PHYADDRPOINTER_REG_0_, P3_PHYADDRPOINTER_REG_1_,
    P3_PHYADDRPOINTER_REG_2_, P3_PHYADDRPOINTER_REG_3_,
    P3_PHYADDRPOINTER_REG_4_, P3_PHYADDRPOINTER_REG_5_,
    P3_PHYADDRPOINTER_REG_6_, P3_PHYADDRPOINTER_REG_7_,
    P3_PHYADDRPOINTER_REG_8_, P3_PHYADDRPOINTER_REG_9_,
    P3_PHYADDRPOINTER_REG_10_, P3_PHYADDRPOINTER_REG_11_,
    P3_PHYADDRPOINTER_REG_12_, P3_PHYADDRPOINTER_REG_13_,
    P3_PHYADDRPOINTER_REG_14_, P3_PHYADDRPOINTER_REG_15_,
    P3_PHYADDRPOINTER_REG_16_, P3_PHYADDRPOINTER_REG_17_,
    P3_PHYADDRPOINTER_REG_18_, P3_PHYADDRPOINTER_REG_19_,
    P3_PHYADDRPOINTER_REG_20_, P3_PHYADDRPOINTER_REG_21_,
    P3_PHYADDRPOINTER_REG_22_, P3_PHYADDRPOINTER_REG_23_,
    P3_PHYADDRPOINTER_REG_24_, P3_PHYADDRPOINTER_REG_25_,
    P3_PHYADDRPOINTER_REG_26_, P3_PHYADDRPOINTER_REG_27_,
    P3_PHYADDRPOINTER_REG_28_, P3_PHYADDRPOINTER_REG_29_,
    P3_PHYADDRPOINTER_REG_30_, P3_PHYADDRPOINTER_REG_31_, P3_LWORD_REG_15_,
    P3_LWORD_REG_14_, P3_LWORD_REG_13_, P3_LWORD_REG_12_, P3_LWORD_REG_11_,
    P3_LWORD_REG_10_, P3_LWORD_REG_9_, P3_LWORD_REG_8_, P3_LWORD_REG_7_,
    P3_LWORD_REG_6_, P3_LWORD_REG_5_, P3_LWORD_REG_4_, P3_LWORD_REG_3_,
    P3_LWORD_REG_2_, P3_LWORD_REG_1_, P3_LWORD_REG_0_, P3_UWORD_REG_14_,
    P3_UWORD_REG_13_, P3_UWORD_REG_12_, P3_UWORD_REG_11_, P3_UWORD_REG_10_,
    P3_UWORD_REG_9_, P3_UWORD_REG_8_, P3_UWORD_REG_7_, P3_UWORD_REG_6_,
    P3_UWORD_REG_5_, P3_UWORD_REG_4_, P3_UWORD_REG_3_, P3_UWORD_REG_2_,
    P3_UWORD_REG_1_, P3_UWORD_REG_0_, P3_DATAO_REG_0_, P3_DATAO_REG_1_,
    P3_DATAO_REG_2_, P3_DATAO_REG_3_, P3_DATAO_REG_4_, P3_DATAO_REG_5_,
    P3_DATAO_REG_6_, P3_DATAO_REG_7_, P3_DATAO_REG_8_, P3_DATAO_REG_9_,
    P3_DATAO_REG_10_, P3_DATAO_REG_11_, P3_DATAO_REG_12_, P3_DATAO_REG_13_,
    P3_DATAO_REG_14_, P3_DATAO_REG_15_, P3_DATAO_REG_16_, P3_DATAO_REG_17_,
    P3_DATAO_REG_18_, P3_DATAO_REG_19_, P3_DATAO_REG_20_, P3_DATAO_REG_21_,
    P3_DATAO_REG_22_, P3_DATAO_REG_23_, P3_DATAO_REG_24_, P3_DATAO_REG_25_,
    P3_DATAO_REG_26_, P3_DATAO_REG_27_, P3_DATAO_REG_28_, P3_DATAO_REG_29_,
    P3_DATAO_REG_30_, P3_DATAO_REG_31_, P3_EAX_REG_0_, P3_EAX_REG_1_,
    P3_EAX_REG_2_, P3_EAX_REG_3_, P3_EAX_REG_4_, P3_EAX_REG_5_,
    P3_EAX_REG_6_, P3_EAX_REG_7_, P3_EAX_REG_8_, P3_EAX_REG_9_,
    P3_EAX_REG_10_, P3_EAX_REG_11_, P3_EAX_REG_12_, P3_EAX_REG_13_,
    P3_EAX_REG_14_, P3_EAX_REG_15_, P3_EAX_REG_16_, P3_EAX_REG_17_,
    P3_EAX_REG_18_, P3_EAX_REG_19_, P3_EAX_REG_20_, P3_EAX_REG_21_,
    P3_EAX_REG_22_, P3_EAX_REG_23_, P3_EAX_REG_24_, P3_EAX_REG_25_,
    P3_EAX_REG_26_, P3_EAX_REG_27_, P3_EAX_REG_28_, P3_EAX_REG_29_,
    P3_EAX_REG_30_, P3_EAX_REG_31_, P3_EBX_REG_0_, P3_EBX_REG_1_,
    P3_EBX_REG_2_, P3_EBX_REG_3_, P3_EBX_REG_4_, P3_EBX_REG_5_,
    P3_EBX_REG_6_, P3_EBX_REG_7_, P3_EBX_REG_8_, P3_EBX_REG_9_,
    P3_EBX_REG_10_, P3_EBX_REG_11_, P3_EBX_REG_12_, P3_EBX_REG_13_,
    P3_EBX_REG_14_, P3_EBX_REG_15_, P3_EBX_REG_16_, P3_EBX_REG_17_,
    P3_EBX_REG_18_, P3_EBX_REG_19_, P3_EBX_REG_20_, P3_EBX_REG_21_,
    P3_EBX_REG_22_, P3_EBX_REG_23_, P3_EBX_REG_24_, P3_EBX_REG_25_,
    P3_EBX_REG_26_, P3_EBX_REG_27_, P3_EBX_REG_28_, P3_EBX_REG_29_,
    P3_EBX_REG_30_, P3_EBX_REG_31_, P3_REIP_REG_0_, P3_REIP_REG_1_,
    P3_REIP_REG_2_, P3_REIP_REG_3_, P3_REIP_REG_4_, P3_REIP_REG_5_,
    P3_REIP_REG_6_, P3_REIP_REG_7_, P3_REIP_REG_8_, P3_REIP_REG_9_,
    P3_REIP_REG_10_, P3_REIP_REG_11_, P3_REIP_REG_12_, P3_REIP_REG_13_,
    P3_REIP_REG_14_, P3_REIP_REG_15_, P3_REIP_REG_16_, P3_REIP_REG_17_,
    P3_REIP_REG_18_, P3_REIP_REG_19_, P3_REIP_REG_20_, P3_REIP_REG_21_,
    P3_REIP_REG_22_, P3_REIP_REG_23_, P3_REIP_REG_24_, P3_REIP_REG_25_,
    P3_REIP_REG_26_, P3_REIP_REG_27_, P3_REIP_REG_28_, P3_REIP_REG_29_,
    P3_REIP_REG_30_, P3_REIP_REG_31_, P3_BYTEENABLE_REG_3_,
    P3_BYTEENABLE_REG_2_, P3_BYTEENABLE_REG_1_, P3_BYTEENABLE_REG_0_,
    P3_W_R_N_REG, P3_FLUSH_REG, P3_MORE_REG, P3_STATEBS16_REG,
    P3_REQUESTPENDING_REG, P3_D_C_N_REG, P3_M_IO_N_REG, P3_CODEFETCH_REG,
    P3_ADS_N_REG, P3_READREQUEST_REG, P3_MEMORYFETCH_REG, P2_BE_N_REG_3_,
    P2_BE_N_REG_2_, P2_BE_N_REG_1_, P2_BE_N_REG_0_, P2_ADDRESS_REG_29_,
    P2_ADDRESS_REG_28_, P2_ADDRESS_REG_27_, P2_ADDRESS_REG_26_,
    P2_ADDRESS_REG_25_, P2_ADDRESS_REG_24_, P2_ADDRESS_REG_23_,
    P2_ADDRESS_REG_22_, P2_ADDRESS_REG_21_, P2_ADDRESS_REG_20_,
    P2_ADDRESS_REG_19_, P2_ADDRESS_REG_18_, P2_ADDRESS_REG_17_,
    P2_ADDRESS_REG_16_, P2_ADDRESS_REG_15_, P2_ADDRESS_REG_14_,
    P2_ADDRESS_REG_13_, P2_ADDRESS_REG_12_, P2_ADDRESS_REG_11_,
    P2_ADDRESS_REG_10_, P2_ADDRESS_REG_9_, P2_ADDRESS_REG_8_,
    P2_ADDRESS_REG_7_, P2_ADDRESS_REG_6_, P2_ADDRESS_REG_5_,
    P2_ADDRESS_REG_4_, P2_ADDRESS_REG_3_, P2_ADDRESS_REG_2_,
    P2_ADDRESS_REG_1_, P2_ADDRESS_REG_0_, P2_STATE_REG_2_, P2_STATE_REG_1_,
    P2_STATE_REG_0_, P2_DATAWIDTH_REG_0_, P2_DATAWIDTH_REG_1_,
    P2_DATAWIDTH_REG_2_, P2_DATAWIDTH_REG_3_, P2_DATAWIDTH_REG_4_,
    P2_DATAWIDTH_REG_5_, P2_DATAWIDTH_REG_6_, P2_DATAWIDTH_REG_7_,
    P2_DATAWIDTH_REG_8_, P2_DATAWIDTH_REG_9_, P2_DATAWIDTH_REG_10_,
    P2_DATAWIDTH_REG_11_, P2_DATAWIDTH_REG_12_, P2_DATAWIDTH_REG_13_,
    P2_DATAWIDTH_REG_14_, P2_DATAWIDTH_REG_15_, P2_DATAWIDTH_REG_16_,
    P2_DATAWIDTH_REG_17_, P2_DATAWIDTH_REG_18_, P2_DATAWIDTH_REG_19_,
    P2_DATAWIDTH_REG_20_, P2_DATAWIDTH_REG_21_, P2_DATAWIDTH_REG_22_,
    P2_DATAWIDTH_REG_23_, P2_DATAWIDTH_REG_24_, P2_DATAWIDTH_REG_25_,
    P2_DATAWIDTH_REG_26_, P2_DATAWIDTH_REG_27_, P2_DATAWIDTH_REG_28_,
    P2_DATAWIDTH_REG_29_, P2_DATAWIDTH_REG_30_, P2_DATAWIDTH_REG_31_,
    P2_STATE2_REG_3_, P2_STATE2_REG_2_, P2_STATE2_REG_1_, P2_STATE2_REG_0_,
    P2_INSTQUEUE_REG_15__7_, P2_INSTQUEUE_REG_15__6_,
    P2_INSTQUEUE_REG_15__5_, P2_INSTQUEUE_REG_15__4_,
    P2_INSTQUEUE_REG_15__3_, P2_INSTQUEUE_REG_15__2_,
    P2_INSTQUEUE_REG_15__1_, P2_INSTQUEUE_REG_15__0_,
    P2_INSTQUEUE_REG_14__7_, P2_INSTQUEUE_REG_14__6_,
    P2_INSTQUEUE_REG_14__5_, P2_INSTQUEUE_REG_14__4_,
    P2_INSTQUEUE_REG_14__3_, P2_INSTQUEUE_REG_14__2_,
    P2_INSTQUEUE_REG_14__1_, P2_INSTQUEUE_REG_14__0_,
    P2_INSTQUEUE_REG_13__7_, P2_INSTQUEUE_REG_13__6_,
    P2_INSTQUEUE_REG_13__5_, P2_INSTQUEUE_REG_13__4_,
    P2_INSTQUEUE_REG_13__3_, P2_INSTQUEUE_REG_13__2_,
    P2_INSTQUEUE_REG_13__1_, P2_INSTQUEUE_REG_13__0_,
    P2_INSTQUEUE_REG_12__7_, P2_INSTQUEUE_REG_12__6_,
    P2_INSTQUEUE_REG_12__5_, P2_INSTQUEUE_REG_12__4_,
    P2_INSTQUEUE_REG_12__3_, P2_INSTQUEUE_REG_12__2_,
    P2_INSTQUEUE_REG_12__1_, P2_INSTQUEUE_REG_12__0_,
    P2_INSTQUEUE_REG_11__7_, P2_INSTQUEUE_REG_11__6_,
    P2_INSTQUEUE_REG_11__5_, P2_INSTQUEUE_REG_11__4_,
    P2_INSTQUEUE_REG_11__3_, P2_INSTQUEUE_REG_11__2_,
    P2_INSTQUEUE_REG_11__1_, P2_INSTQUEUE_REG_11__0_,
    P2_INSTQUEUE_REG_10__7_, P2_INSTQUEUE_REG_10__6_,
    P2_INSTQUEUE_REG_10__5_, P2_INSTQUEUE_REG_10__4_,
    P2_INSTQUEUE_REG_10__3_, P2_INSTQUEUE_REG_10__2_,
    P2_INSTQUEUE_REG_10__1_, P2_INSTQUEUE_REG_10__0_,
    P2_INSTQUEUE_REG_9__7_, P2_INSTQUEUE_REG_9__6_, P2_INSTQUEUE_REG_9__5_,
    P2_INSTQUEUE_REG_9__4_, P2_INSTQUEUE_REG_9__3_, P2_INSTQUEUE_REG_9__2_,
    P2_INSTQUEUE_REG_9__1_, P2_INSTQUEUE_REG_9__0_, P2_INSTQUEUE_REG_8__7_,
    P2_INSTQUEUE_REG_8__6_, P2_INSTQUEUE_REG_8__5_, P2_INSTQUEUE_REG_8__4_,
    P2_INSTQUEUE_REG_8__3_, P2_INSTQUEUE_REG_8__2_, P2_INSTQUEUE_REG_8__1_,
    P2_INSTQUEUE_REG_8__0_, P2_INSTQUEUE_REG_7__7_, P2_INSTQUEUE_REG_7__6_,
    P2_INSTQUEUE_REG_7__5_, P2_INSTQUEUE_REG_7__4_, P2_INSTQUEUE_REG_7__3_,
    P2_INSTQUEUE_REG_7__2_, P2_INSTQUEUE_REG_7__1_, P2_INSTQUEUE_REG_7__0_,
    P2_INSTQUEUE_REG_6__7_, P2_INSTQUEUE_REG_6__6_, P2_INSTQUEUE_REG_6__5_,
    P2_INSTQUEUE_REG_6__4_, P2_INSTQUEUE_REG_6__3_, P2_INSTQUEUE_REG_6__2_,
    P2_INSTQUEUE_REG_6__1_, P2_INSTQUEUE_REG_6__0_, P2_INSTQUEUE_REG_5__7_,
    P2_INSTQUEUE_REG_5__6_, P2_INSTQUEUE_REG_5__5_, P2_INSTQUEUE_REG_5__4_,
    P2_INSTQUEUE_REG_5__3_, P2_INSTQUEUE_REG_5__2_, P2_INSTQUEUE_REG_5__1_,
    P2_INSTQUEUE_REG_5__0_, P2_INSTQUEUE_REG_4__7_, P2_INSTQUEUE_REG_4__6_,
    P2_INSTQUEUE_REG_4__5_, P2_INSTQUEUE_REG_4__4_, P2_INSTQUEUE_REG_4__3_,
    P2_INSTQUEUE_REG_4__2_, P2_INSTQUEUE_REG_4__1_, P2_INSTQUEUE_REG_4__0_,
    P2_INSTQUEUE_REG_3__7_, P2_INSTQUEUE_REG_3__6_, P2_INSTQUEUE_REG_3__5_,
    P2_INSTQUEUE_REG_3__4_, P2_INSTQUEUE_REG_3__3_, P2_INSTQUEUE_REG_3__2_,
    P2_INSTQUEUE_REG_3__1_, P2_INSTQUEUE_REG_3__0_, P2_INSTQUEUE_REG_2__7_,
    P2_INSTQUEUE_REG_2__6_, P2_INSTQUEUE_REG_2__5_, P2_INSTQUEUE_REG_2__4_,
    P2_INSTQUEUE_REG_2__3_, P2_INSTQUEUE_REG_2__2_, P2_INSTQUEUE_REG_2__1_,
    P2_INSTQUEUE_REG_2__0_, P2_INSTQUEUE_REG_1__7_, P2_INSTQUEUE_REG_1__6_,
    P2_INSTQUEUE_REG_1__5_, P2_INSTQUEUE_REG_1__4_, P2_INSTQUEUE_REG_1__3_,
    P2_INSTQUEUE_REG_1__2_, P2_INSTQUEUE_REG_1__1_, P2_INSTQUEUE_REG_1__0_,
    P2_INSTQUEUE_REG_0__7_, P2_INSTQUEUE_REG_0__6_, P2_INSTQUEUE_REG_0__5_,
    P2_INSTQUEUE_REG_0__4_, P2_INSTQUEUE_REG_0__3_, P2_INSTQUEUE_REG_0__2_,
    P2_INSTQUEUE_REG_0__1_, P2_INSTQUEUE_REG_0__0_,
    P2_INSTQUEUERD_ADDR_REG_4_, P2_INSTQUEUERD_ADDR_REG_3_,
    P2_INSTQUEUERD_ADDR_REG_2_, P2_INSTQUEUERD_ADDR_REG_1_,
    P2_INSTQUEUERD_ADDR_REG_0_, P2_INSTQUEUEWR_ADDR_REG_4_,
    P2_INSTQUEUEWR_ADDR_REG_3_, P2_INSTQUEUEWR_ADDR_REG_2_,
    P2_INSTQUEUEWR_ADDR_REG_1_, P2_INSTQUEUEWR_ADDR_REG_0_,
    P2_INSTADDRPOINTER_REG_0_, P2_INSTADDRPOINTER_REG_1_,
    P2_INSTADDRPOINTER_REG_2_, P2_INSTADDRPOINTER_REG_3_,
    P2_INSTADDRPOINTER_REG_4_, P2_INSTADDRPOINTER_REG_5_,
    P2_INSTADDRPOINTER_REG_6_, P2_INSTADDRPOINTER_REG_7_,
    P2_INSTADDRPOINTER_REG_8_, P2_INSTADDRPOINTER_REG_9_,
    P2_INSTADDRPOINTER_REG_10_, P2_INSTADDRPOINTER_REG_11_,
    P2_INSTADDRPOINTER_REG_12_, P2_INSTADDRPOINTER_REG_13_,
    P2_INSTADDRPOINTER_REG_14_, P2_INSTADDRPOINTER_REG_15_,
    P2_INSTADDRPOINTER_REG_16_, P2_INSTADDRPOINTER_REG_17_,
    P2_INSTADDRPOINTER_REG_18_, P2_INSTADDRPOINTER_REG_19_,
    P2_INSTADDRPOINTER_REG_20_, P2_INSTADDRPOINTER_REG_21_,
    P2_INSTADDRPOINTER_REG_22_, P2_INSTADDRPOINTER_REG_23_,
    P2_INSTADDRPOINTER_REG_24_, P2_INSTADDRPOINTER_REG_25_,
    P2_INSTADDRPOINTER_REG_26_, P2_INSTADDRPOINTER_REG_27_,
    P2_INSTADDRPOINTER_REG_28_, P2_INSTADDRPOINTER_REG_29_,
    P2_INSTADDRPOINTER_REG_30_, P2_INSTADDRPOINTER_REG_31_,
    P2_PHYADDRPOINTER_REG_0_, P2_PHYADDRPOINTER_REG_1_,
    P2_PHYADDRPOINTER_REG_2_, P2_PHYADDRPOINTER_REG_3_,
    P2_PHYADDRPOINTER_REG_4_, P2_PHYADDRPOINTER_REG_5_,
    P2_PHYADDRPOINTER_REG_6_, P2_PHYADDRPOINTER_REG_7_,
    P2_PHYADDRPOINTER_REG_8_, P2_PHYADDRPOINTER_REG_9_,
    P2_PHYADDRPOINTER_REG_10_, P2_PHYADDRPOINTER_REG_11_,
    P2_PHYADDRPOINTER_REG_12_, P2_PHYADDRPOINTER_REG_13_,
    P2_PHYADDRPOINTER_REG_14_, P2_PHYADDRPOINTER_REG_15_,
    P2_PHYADDRPOINTER_REG_16_, P2_PHYADDRPOINTER_REG_17_,
    P2_PHYADDRPOINTER_REG_18_, P2_PHYADDRPOINTER_REG_19_,
    P2_PHYADDRPOINTER_REG_20_, P2_PHYADDRPOINTER_REG_21_,
    P2_PHYADDRPOINTER_REG_22_, P2_PHYADDRPOINTER_REG_23_,
    P2_PHYADDRPOINTER_REG_24_, P2_PHYADDRPOINTER_REG_25_,
    P2_PHYADDRPOINTER_REG_26_, P2_PHYADDRPOINTER_REG_27_,
    P2_PHYADDRPOINTER_REG_28_, P2_PHYADDRPOINTER_REG_29_,
    P2_PHYADDRPOINTER_REG_30_, P2_PHYADDRPOINTER_REG_31_, P2_LWORD_REG_15_,
    P2_LWORD_REG_14_, P2_LWORD_REG_13_, P2_LWORD_REG_12_, P2_LWORD_REG_11_,
    P2_LWORD_REG_10_, P2_LWORD_REG_9_, P2_LWORD_REG_8_, P2_LWORD_REG_7_,
    P2_LWORD_REG_6_, P2_LWORD_REG_5_, P2_LWORD_REG_4_, P2_LWORD_REG_3_,
    P2_LWORD_REG_2_, P2_LWORD_REG_1_, P2_LWORD_REG_0_, P2_UWORD_REG_14_,
    P2_UWORD_REG_13_, P2_UWORD_REG_12_, P2_UWORD_REG_11_, P2_UWORD_REG_10_,
    P2_UWORD_REG_9_, P2_UWORD_REG_8_, P2_UWORD_REG_7_, P2_UWORD_REG_6_,
    P2_UWORD_REG_5_, P2_UWORD_REG_4_, P2_UWORD_REG_3_, P2_UWORD_REG_2_,
    P2_UWORD_REG_1_, P2_UWORD_REG_0_, P2_DATAO_REG_0_, P2_DATAO_REG_1_,
    P2_DATAO_REG_2_, P2_DATAO_REG_3_, P2_DATAO_REG_4_, P2_DATAO_REG_5_,
    P2_DATAO_REG_6_, P2_DATAO_REG_7_, P2_DATAO_REG_8_, P2_DATAO_REG_9_,
    P2_DATAO_REG_10_, P2_DATAO_REG_11_, P2_DATAO_REG_12_, P2_DATAO_REG_13_,
    P2_DATAO_REG_14_, P2_DATAO_REG_15_, P2_DATAO_REG_16_, P2_DATAO_REG_17_,
    P2_DATAO_REG_18_, P2_DATAO_REG_19_, P2_DATAO_REG_20_, P2_DATAO_REG_21_,
    P2_DATAO_REG_22_, P2_DATAO_REG_23_, P2_DATAO_REG_24_, P2_DATAO_REG_25_,
    P2_DATAO_REG_26_, P2_DATAO_REG_27_, P2_DATAO_REG_28_, P2_DATAO_REG_29_,
    P2_DATAO_REG_30_, P2_DATAO_REG_31_, P2_EAX_REG_0_, P2_EAX_REG_1_,
    P2_EAX_REG_2_, P2_EAX_REG_3_, P2_EAX_REG_4_, P2_EAX_REG_5_,
    P2_EAX_REG_6_, P2_EAX_REG_7_, P2_EAX_REG_8_, P2_EAX_REG_9_,
    P2_EAX_REG_10_, P2_EAX_REG_11_, P2_EAX_REG_12_, P2_EAX_REG_13_,
    P2_EAX_REG_14_, P2_EAX_REG_15_, P2_EAX_REG_16_, P2_EAX_REG_17_,
    P2_EAX_REG_18_, P2_EAX_REG_19_, P2_EAX_REG_20_, P2_EAX_REG_21_,
    P2_EAX_REG_22_, P2_EAX_REG_23_, P2_EAX_REG_24_, P2_EAX_REG_25_,
    P2_EAX_REG_26_, P2_EAX_REG_27_, P2_EAX_REG_28_, P2_EAX_REG_29_,
    P2_EAX_REG_30_, P2_EAX_REG_31_, P2_EBX_REG_0_, P2_EBX_REG_1_,
    P2_EBX_REG_2_, P2_EBX_REG_3_, P2_EBX_REG_4_, P2_EBX_REG_5_,
    P2_EBX_REG_6_, P2_EBX_REG_7_, P2_EBX_REG_8_, P2_EBX_REG_9_,
    P2_EBX_REG_10_, P2_EBX_REG_11_, P2_EBX_REG_12_, P2_EBX_REG_13_,
    P2_EBX_REG_14_, P2_EBX_REG_15_, P2_EBX_REG_16_, P2_EBX_REG_17_,
    P2_EBX_REG_18_, P2_EBX_REG_19_, P2_EBX_REG_20_, P2_EBX_REG_21_,
    P2_EBX_REG_22_, P2_EBX_REG_23_, P2_EBX_REG_24_, P2_EBX_REG_25_,
    P2_EBX_REG_26_, P2_EBX_REG_27_, P2_EBX_REG_28_, P2_EBX_REG_29_,
    P2_EBX_REG_30_, P2_EBX_REG_31_, P2_REIP_REG_0_, P2_REIP_REG_1_,
    P2_REIP_REG_2_, P2_REIP_REG_3_, P2_REIP_REG_4_, P2_REIP_REG_5_,
    P2_REIP_REG_6_, P2_REIP_REG_7_, P2_REIP_REG_8_, P2_REIP_REG_9_,
    P2_REIP_REG_10_, P2_REIP_REG_11_, P2_REIP_REG_12_, P2_REIP_REG_13_,
    P2_REIP_REG_14_, P2_REIP_REG_15_, P2_REIP_REG_16_, P2_REIP_REG_17_,
    P2_REIP_REG_18_, P2_REIP_REG_19_, P2_REIP_REG_20_, P2_REIP_REG_21_,
    P2_REIP_REG_22_, P2_REIP_REG_23_, P2_REIP_REG_24_, P2_REIP_REG_25_,
    P2_REIP_REG_26_, P2_REIP_REG_27_, P2_REIP_REG_28_, P2_REIP_REG_29_,
    P2_REIP_REG_30_, P2_REIP_REG_31_, P2_BYTEENABLE_REG_3_,
    P2_BYTEENABLE_REG_2_, P2_BYTEENABLE_REG_1_, P2_BYTEENABLE_REG_0_,
    P2_W_R_N_REG, P2_FLUSH_REG, P2_MORE_REG, P2_STATEBS16_REG,
    P2_REQUESTPENDING_REG, P2_D_C_N_REG, P2_M_IO_N_REG, P2_CODEFETCH_REG,
    P2_ADS_N_REG, P2_READREQUEST_REG, P2_MEMORYFETCH_REG, P1_BE_N_REG_3_,
    P1_BE_N_REG_2_, P1_BE_N_REG_1_, P1_BE_N_REG_0_, P1_ADDRESS_REG_29_,
    P1_ADDRESS_REG_28_, P1_ADDRESS_REG_27_, P1_ADDRESS_REG_26_,
    P1_ADDRESS_REG_25_, P1_ADDRESS_REG_24_, P1_ADDRESS_REG_23_,
    P1_ADDRESS_REG_22_, P1_ADDRESS_REG_21_, P1_ADDRESS_REG_20_,
    P1_ADDRESS_REG_19_, P1_ADDRESS_REG_18_, P1_ADDRESS_REG_17_,
    P1_ADDRESS_REG_16_, P1_ADDRESS_REG_15_, P1_ADDRESS_REG_14_,
    P1_ADDRESS_REG_13_, P1_ADDRESS_REG_12_, P1_ADDRESS_REG_11_,
    P1_ADDRESS_REG_10_, P1_ADDRESS_REG_9_, P1_ADDRESS_REG_8_,
    P1_ADDRESS_REG_7_, P1_ADDRESS_REG_6_, P1_ADDRESS_REG_5_,
    P1_ADDRESS_REG_4_, P1_ADDRESS_REG_3_, P1_ADDRESS_REG_2_,
    P1_ADDRESS_REG_1_, P1_ADDRESS_REG_0_, P1_STATE_REG_2_, P1_STATE_REG_1_,
    P1_STATE_REG_0_, P1_DATAWIDTH_REG_0_, P1_DATAWIDTH_REG_1_,
    P1_DATAWIDTH_REG_2_, P1_DATAWIDTH_REG_3_, P1_DATAWIDTH_REG_4_,
    P1_DATAWIDTH_REG_5_, P1_DATAWIDTH_REG_6_, P1_DATAWIDTH_REG_7_,
    P1_DATAWIDTH_REG_8_, P1_DATAWIDTH_REG_9_, P1_DATAWIDTH_REG_10_,
    P1_DATAWIDTH_REG_11_, P1_DATAWIDTH_REG_12_, P1_DATAWIDTH_REG_13_,
    P1_DATAWIDTH_REG_14_, P1_DATAWIDTH_REG_15_, P1_DATAWIDTH_REG_16_,
    P1_DATAWIDTH_REG_17_, P1_DATAWIDTH_REG_18_, P1_DATAWIDTH_REG_19_,
    P1_DATAWIDTH_REG_20_, P1_DATAWIDTH_REG_21_, P1_DATAWIDTH_REG_22_,
    P1_DATAWIDTH_REG_23_, P1_DATAWIDTH_REG_24_, P1_DATAWIDTH_REG_25_,
    P1_DATAWIDTH_REG_26_, P1_DATAWIDTH_REG_27_, P1_DATAWIDTH_REG_28_,
    P1_DATAWIDTH_REG_29_, P1_DATAWIDTH_REG_30_, P1_DATAWIDTH_REG_31_,
    P1_STATE2_REG_3_, P1_STATE2_REG_2_, P1_STATE2_REG_1_, P1_STATE2_REG_0_,
    P1_INSTQUEUE_REG_15__7_, P1_INSTQUEUE_REG_15__6_,
    P1_INSTQUEUE_REG_15__5_, P1_INSTQUEUE_REG_15__4_,
    P1_INSTQUEUE_REG_15__3_, P1_INSTQUEUE_REG_15__2_,
    P1_INSTQUEUE_REG_15__1_, P1_INSTQUEUE_REG_15__0_,
    P1_INSTQUEUE_REG_14__7_, P1_INSTQUEUE_REG_14__6_,
    P1_INSTQUEUE_REG_14__5_, P1_INSTQUEUE_REG_14__4_,
    P1_INSTQUEUE_REG_14__3_, P1_INSTQUEUE_REG_14__2_,
    P1_INSTQUEUE_REG_14__1_, P1_INSTQUEUE_REG_14__0_,
    P1_INSTQUEUE_REG_13__7_, P1_INSTQUEUE_REG_13__6_,
    P1_INSTQUEUE_REG_13__5_, P1_INSTQUEUE_REG_13__4_,
    P1_INSTQUEUE_REG_13__3_, P1_INSTQUEUE_REG_13__2_,
    P1_INSTQUEUE_REG_13__1_, P1_INSTQUEUE_REG_13__0_,
    P1_INSTQUEUE_REG_12__7_, P1_INSTQUEUE_REG_12__6_,
    P1_INSTQUEUE_REG_12__5_, P1_INSTQUEUE_REG_12__4_,
    P1_INSTQUEUE_REG_12__3_, P1_INSTQUEUE_REG_12__2_,
    P1_INSTQUEUE_REG_12__1_, P1_INSTQUEUE_REG_12__0_,
    P1_INSTQUEUE_REG_11__7_, P1_INSTQUEUE_REG_11__6_,
    P1_INSTQUEUE_REG_11__5_, P1_INSTQUEUE_REG_11__4_,
    P1_INSTQUEUE_REG_11__3_, P1_INSTQUEUE_REG_11__2_,
    P1_INSTQUEUE_REG_11__1_, P1_INSTQUEUE_REG_11__0_,
    P1_INSTQUEUE_REG_10__7_, P1_INSTQUEUE_REG_10__6_,
    P1_INSTQUEUE_REG_10__5_, P1_INSTQUEUE_REG_10__4_,
    P1_INSTQUEUE_REG_10__3_, P1_INSTQUEUE_REG_10__2_,
    P1_INSTQUEUE_REG_10__1_, P1_INSTQUEUE_REG_10__0_,
    P1_INSTQUEUE_REG_9__7_, P1_INSTQUEUE_REG_9__6_, P1_INSTQUEUE_REG_9__5_,
    P1_INSTQUEUE_REG_9__4_, P1_INSTQUEUE_REG_9__3_, P1_INSTQUEUE_REG_9__2_,
    P1_INSTQUEUE_REG_9__1_, P1_INSTQUEUE_REG_9__0_, P1_INSTQUEUE_REG_8__7_,
    P1_INSTQUEUE_REG_8__6_, P1_INSTQUEUE_REG_8__5_, P1_INSTQUEUE_REG_8__4_,
    P1_INSTQUEUE_REG_8__3_, P1_INSTQUEUE_REG_8__2_, P1_INSTQUEUE_REG_8__1_,
    P1_INSTQUEUE_REG_8__0_, P1_INSTQUEUE_REG_7__7_, P1_INSTQUEUE_REG_7__6_,
    P1_INSTQUEUE_REG_7__5_, P1_INSTQUEUE_REG_7__4_, P1_INSTQUEUE_REG_7__3_,
    P1_INSTQUEUE_REG_7__2_, P1_INSTQUEUE_REG_7__1_, P1_INSTQUEUE_REG_7__0_,
    P1_INSTQUEUE_REG_6__7_, P1_INSTQUEUE_REG_6__6_, P1_INSTQUEUE_REG_6__5_,
    P1_INSTQUEUE_REG_6__4_, P1_INSTQUEUE_REG_6__3_, P1_INSTQUEUE_REG_6__2_,
    P1_INSTQUEUE_REG_6__1_, P1_INSTQUEUE_REG_6__0_, P1_INSTQUEUE_REG_5__7_,
    P1_INSTQUEUE_REG_5__6_, P1_INSTQUEUE_REG_5__5_, P1_INSTQUEUE_REG_5__4_,
    P1_INSTQUEUE_REG_5__3_, P1_INSTQUEUE_REG_5__2_, P1_INSTQUEUE_REG_5__1_,
    P1_INSTQUEUE_REG_5__0_, P1_INSTQUEUE_REG_4__7_, P1_INSTQUEUE_REG_4__6_,
    P1_INSTQUEUE_REG_4__5_, P1_INSTQUEUE_REG_4__4_, P1_INSTQUEUE_REG_4__3_,
    P1_INSTQUEUE_REG_4__2_, P1_INSTQUEUE_REG_4__1_, P1_INSTQUEUE_REG_4__0_,
    P1_INSTQUEUE_REG_3__7_, P1_INSTQUEUE_REG_3__6_, P1_INSTQUEUE_REG_3__5_,
    P1_INSTQUEUE_REG_3__4_, P1_INSTQUEUE_REG_3__3_, P1_INSTQUEUE_REG_3__2_,
    P1_INSTQUEUE_REG_3__1_, P1_INSTQUEUE_REG_3__0_, P1_INSTQUEUE_REG_2__7_,
    P1_INSTQUEUE_REG_2__6_, P1_INSTQUEUE_REG_2__5_, P1_INSTQUEUE_REG_2__4_,
    P1_INSTQUEUE_REG_2__3_, P1_INSTQUEUE_REG_2__2_, P1_INSTQUEUE_REG_2__1_,
    P1_INSTQUEUE_REG_2__0_, P1_INSTQUEUE_REG_1__7_, P1_INSTQUEUE_REG_1__6_,
    P1_INSTQUEUE_REG_1__5_, P1_INSTQUEUE_REG_1__4_, P1_INSTQUEUE_REG_1__3_,
    P1_INSTQUEUE_REG_1__2_, P1_INSTQUEUE_REG_1__1_, P1_INSTQUEUE_REG_1__0_,
    P1_INSTQUEUE_REG_0__7_, P1_INSTQUEUE_REG_0__6_, P1_INSTQUEUE_REG_0__5_,
    P1_INSTQUEUE_REG_0__4_, P1_INSTQUEUE_REG_0__3_, P1_INSTQUEUE_REG_0__2_,
    P1_INSTQUEUE_REG_0__1_, P1_INSTQUEUE_REG_0__0_,
    P1_INSTQUEUERD_ADDR_REG_4_, P1_INSTQUEUERD_ADDR_REG_3_,
    P1_INSTQUEUERD_ADDR_REG_2_, P1_INSTQUEUERD_ADDR_REG_1_,
    P1_INSTQUEUERD_ADDR_REG_0_, P1_INSTQUEUEWR_ADDR_REG_4_,
    P1_INSTQUEUEWR_ADDR_REG_3_, P1_INSTQUEUEWR_ADDR_REG_2_,
    P1_INSTQUEUEWR_ADDR_REG_1_, P1_INSTQUEUEWR_ADDR_REG_0_,
    P1_INSTADDRPOINTER_REG_0_, P1_INSTADDRPOINTER_REG_1_,
    P1_INSTADDRPOINTER_REG_2_, P1_INSTADDRPOINTER_REG_3_,
    P1_INSTADDRPOINTER_REG_4_, P1_INSTADDRPOINTER_REG_5_,
    P1_INSTADDRPOINTER_REG_6_, P1_INSTADDRPOINTER_REG_7_,
    P1_INSTADDRPOINTER_REG_8_, P1_INSTADDRPOINTER_REG_9_,
    P1_INSTADDRPOINTER_REG_10_, P1_INSTADDRPOINTER_REG_11_,
    P1_INSTADDRPOINTER_REG_12_, P1_INSTADDRPOINTER_REG_13_,
    P1_INSTADDRPOINTER_REG_14_, P1_INSTADDRPOINTER_REG_15_,
    P1_INSTADDRPOINTER_REG_16_, P1_INSTADDRPOINTER_REG_17_,
    P1_INSTADDRPOINTER_REG_18_, P1_INSTADDRPOINTER_REG_19_,
    P1_INSTADDRPOINTER_REG_20_, P1_INSTADDRPOINTER_REG_21_,
    P1_INSTADDRPOINTER_REG_22_, P1_INSTADDRPOINTER_REG_23_,
    P1_INSTADDRPOINTER_REG_24_, P1_INSTADDRPOINTER_REG_25_,
    P1_INSTADDRPOINTER_REG_26_, P1_INSTADDRPOINTER_REG_27_,
    P1_INSTADDRPOINTER_REG_28_, P1_INSTADDRPOINTER_REG_29_,
    P1_INSTADDRPOINTER_REG_30_, P1_INSTADDRPOINTER_REG_31_,
    P1_PHYADDRPOINTER_REG_0_, P1_PHYADDRPOINTER_REG_1_,
    P1_PHYADDRPOINTER_REG_2_, P1_PHYADDRPOINTER_REG_3_,
    P1_PHYADDRPOINTER_REG_4_, P1_PHYADDRPOINTER_REG_5_,
    P1_PHYADDRPOINTER_REG_6_, P1_PHYADDRPOINTER_REG_7_,
    P1_PHYADDRPOINTER_REG_8_, P1_PHYADDRPOINTER_REG_9_,
    P1_PHYADDRPOINTER_REG_10_, P1_PHYADDRPOINTER_REG_11_,
    P1_PHYADDRPOINTER_REG_12_, P1_PHYADDRPOINTER_REG_13_,
    P1_PHYADDRPOINTER_REG_14_, P1_PHYADDRPOINTER_REG_15_,
    P1_PHYADDRPOINTER_REG_16_, P1_PHYADDRPOINTER_REG_17_,
    P1_PHYADDRPOINTER_REG_18_, P1_PHYADDRPOINTER_REG_19_,
    P1_PHYADDRPOINTER_REG_20_, P1_PHYADDRPOINTER_REG_21_,
    P1_PHYADDRPOINTER_REG_22_, P1_PHYADDRPOINTER_REG_23_,
    P1_PHYADDRPOINTER_REG_24_, P1_PHYADDRPOINTER_REG_25_,
    P1_PHYADDRPOINTER_REG_26_, P1_PHYADDRPOINTER_REG_27_,
    P1_PHYADDRPOINTER_REG_28_, P1_PHYADDRPOINTER_REG_29_,
    P1_PHYADDRPOINTER_REG_30_, P1_PHYADDRPOINTER_REG_31_, P1_LWORD_REG_15_,
    P1_LWORD_REG_14_, P1_LWORD_REG_13_, P1_LWORD_REG_12_, P1_LWORD_REG_11_,
    P1_LWORD_REG_10_, P1_LWORD_REG_9_, P1_LWORD_REG_8_, P1_LWORD_REG_7_,
    P1_LWORD_REG_6_, P1_LWORD_REG_5_, P1_LWORD_REG_4_, P1_LWORD_REG_3_,
    P1_LWORD_REG_2_, P1_LWORD_REG_1_, P1_LWORD_REG_0_, P1_UWORD_REG_14_,
    P1_UWORD_REG_13_, P1_UWORD_REG_12_, P1_UWORD_REG_11_, P1_UWORD_REG_10_,
    P1_UWORD_REG_9_, P1_UWORD_REG_8_, P1_UWORD_REG_7_, P1_UWORD_REG_6_,
    P1_UWORD_REG_5_, P1_UWORD_REG_4_, P1_UWORD_REG_3_, P1_UWORD_REG_2_,
    P1_UWORD_REG_1_, P1_UWORD_REG_0_, P1_DATAO_REG_0_, P1_DATAO_REG_1_,
    P1_DATAO_REG_2_, P1_DATAO_REG_3_, P1_DATAO_REG_4_, P1_DATAO_REG_5_,
    P1_DATAO_REG_6_, P1_DATAO_REG_7_, P1_DATAO_REG_8_, P1_DATAO_REG_9_,
    P1_DATAO_REG_10_, P1_DATAO_REG_11_, P1_DATAO_REG_12_, P1_DATAO_REG_13_,
    P1_DATAO_REG_14_, P1_DATAO_REG_15_, P1_DATAO_REG_16_, P1_DATAO_REG_17_,
    P1_DATAO_REG_18_, P1_DATAO_REG_19_, P1_DATAO_REG_20_, P1_DATAO_REG_21_,
    P1_DATAO_REG_22_, P1_DATAO_REG_23_, P1_DATAO_REG_24_, P1_DATAO_REG_25_,
    P1_DATAO_REG_26_, P1_DATAO_REG_27_, P1_DATAO_REG_28_, P1_DATAO_REG_29_,
    P1_DATAO_REG_30_, P1_DATAO_REG_31_, P1_EAX_REG_0_, P1_EAX_REG_1_,
    P1_EAX_REG_2_, P1_EAX_REG_3_, P1_EAX_REG_4_, P1_EAX_REG_5_,
    P1_EAX_REG_6_, P1_EAX_REG_7_, P1_EAX_REG_8_, P1_EAX_REG_9_,
    P1_EAX_REG_10_, P1_EAX_REG_11_, P1_EAX_REG_12_, P1_EAX_REG_13_,
    P1_EAX_REG_14_, P1_EAX_REG_15_, P1_EAX_REG_16_, P1_EAX_REG_17_,
    P1_EAX_REG_18_, P1_EAX_REG_19_, P1_EAX_REG_20_, P1_EAX_REG_21_,
    P1_EAX_REG_22_, P1_EAX_REG_23_, P1_EAX_REG_24_, P1_EAX_REG_25_,
    P1_EAX_REG_26_, P1_EAX_REG_27_, P1_EAX_REG_28_, P1_EAX_REG_29_,
    P1_EAX_REG_30_, P1_EAX_REG_31_, P1_EBX_REG_0_, P1_EBX_REG_1_,
    P1_EBX_REG_2_, P1_EBX_REG_3_, P1_EBX_REG_4_, P1_EBX_REG_5_,
    P1_EBX_REG_6_, P1_EBX_REG_7_, P1_EBX_REG_8_, P1_EBX_REG_9_,
    P1_EBX_REG_10_, P1_EBX_REG_11_, P1_EBX_REG_12_, P1_EBX_REG_13_,
    P1_EBX_REG_14_, P1_EBX_REG_15_, P1_EBX_REG_16_, P1_EBX_REG_17_,
    P1_EBX_REG_18_, P1_EBX_REG_19_, P1_EBX_REG_20_, P1_EBX_REG_21_,
    P1_EBX_REG_22_, P1_EBX_REG_23_, P1_EBX_REG_24_, P1_EBX_REG_25_,
    P1_EBX_REG_26_, P1_EBX_REG_27_, P1_EBX_REG_28_, P1_EBX_REG_29_,
    P1_EBX_REG_30_, P1_EBX_REG_31_, P1_REIP_REG_0_, P1_REIP_REG_1_,
    P1_REIP_REG_2_, P1_REIP_REG_3_, P1_REIP_REG_4_, P1_REIP_REG_5_,
    P1_REIP_REG_6_, P1_REIP_REG_7_, P1_REIP_REG_8_, P1_REIP_REG_9_,
    P1_REIP_REG_10_, P1_REIP_REG_11_, P1_REIP_REG_12_, P1_REIP_REG_13_,
    P1_REIP_REG_14_, P1_REIP_REG_15_, P1_REIP_REG_16_, P1_REIP_REG_17_,
    P1_REIP_REG_18_, P1_REIP_REG_19_, P1_REIP_REG_20_, P1_REIP_REG_21_,
    P1_REIP_REG_22_, P1_REIP_REG_23_, P1_REIP_REG_24_, P1_REIP_REG_25_,
    P1_REIP_REG_26_, P1_REIP_REG_27_, P1_REIP_REG_28_, P1_REIP_REG_29_,
    P1_REIP_REG_30_, P1_REIP_REG_31_, P1_BYTEENABLE_REG_3_,
    P1_BYTEENABLE_REG_2_, P1_BYTEENABLE_REG_1_, P1_BYTEENABLE_REG_0_,
    P1_W_R_N_REG, P1_FLUSH_REG, P1_MORE_REG, P1_STATEBS16_REG,
    P1_REQUESTPENDING_REG, P1_D_C_N_REG, P1_M_IO_N_REG, P1_CODEFETCH_REG,
    P1_ADS_N_REG, P1_READREQUEST_REG, P1_MEMORYFETCH_REG;
  wire n4380, n4381, n4382, n4383, n4384_1, n4385, n4386, n4388, n4389_1,
    n4391, n4392, n4394_1, n4395, n4397, n4398, n4400, n4401, n4403,
    n4404_1, n4406, n4407, n4409_1, n4410, n4412, n4413, n4415, n4416,
    n4418, n4419_1, n4421, n4422, n4424_1, n4425, n4427, n4428, n4430,
    n4431, n4433, n4434_1, n4436, n4437, n4439_1, n4440, n4442, n4443,
    n4445, n4446, n4448, n4449_1, n4451, n4452, n4454_1, n4455, n4457,
    n4458, n4460, n4461, n4463, n4464_1, n4466, n4467, n4469_1, n4470,
    n4472, n4473, n4475, n4476, n4477, n4478, n4479_1, n4480, n4481, n4482,
    n4483, n4484_1, n4485, n4486, n4487, n4488, n4489_1, n4490, n4491,
    n4492, n4493, n4494_1, n4495, n4496, n4497, n4498, n4499_1, n4500,
    n4501, n4502, n4503, n4504_1, n4505, n4506, n4507, n4508, n4509_1,
    n4510, n4512, n4513, n4514_1, n4515, n4516, n4517, n4518, n4519_1,
    n4520, n4521, n4522, n4523, n4524_1, n4525, n4526, n4527, n4528,
    n4529_1, n4530, n4531, n4532, n4533, n4534_1, n4535, n4536, n4537,
    n4538, n4539_1, n4540, n4541, n4542, n4543, n4544_1, n4545, n4546,
    n4547, n4548, n4549_1, n4550, n4551, n4552, n4553, n4554_1, n4556,
    n4557, n4558, n4559_1, n4561, n4562, n4563, n4564_1, n4566, n4567,
    n4568, n4569_1, n4571, n4572, n4573, n4574_1, n4576, n4577, n4578,
    n4579_1, n4581, n4582, n4583, n4584_1, n4586, n4587, n4588, n4589_1,
    n4591, n4592, n4593, n4594_1, n4596, n4597, n4598, n4599_1, n4601,
    n4602, n4603, n4604_1, n4606, n4607, n4608, n4609_1, n4611, n4612,
    n4613, n4614_1, n4616, n4617, n4618, n4619_1, n4621, n4622, n4623,
    n4624_1, n4626, n4627, n4628, n4629_1, n4631, n4632, n4633, n4634_1,
    n4636, n4637, n4638, n4639_1, n4641, n4642, n4643, n4644_1, n4646,
    n4647, n4648, n4649_1, n4651, n4652, n4653, n4654_1, n4656, n4657,
    n4658, n4659_1, n4661, n4662, n4663, n4664_1, n4666, n4667, n4668,
    n4669_1, n4671, n4672, n4673, n4674_1, n4676, n4677, n4678, n4679_1,
    n4681, n4682, n4683, n4684_1, n4686, n4687, n4688, n4689_1, n4691,
    n4692, n4693, n4694_1, n4696, n4697, n4698, n4699_1, n4701, n4702,
    n4703, n4704_1, n4706, n4707, n4708, n4709_1, n4712, n4713, n4715,
    n4716, n4718, n4719_1, n4721, n4722, n4724_1, n4725, n4727, n4728,
    n4730, n4731, n4733, n4734_1, n4736, n4737, n4739_1, n4740, n4742,
    n4743, n4745, n4746, n4748, n4749_1, n4751, n4752, n4754_1, n4755,
    n4757, n4758, n4760, n4761, n4763, n4764_1, n4766, n4767, n4769_1,
    n4770, n4772, n4773, n4775, n4776, n4778, n4779_1, n4781, n4782,
    n4784_1, n4785, n4787, n4788, n4790, n4791, n4793, n4794_1, n4796,
    n4797, n4799_1, n4800, n4802, n4803, n4805, n4806, n4809_1, n4810,
    n4811, n4812, n4813, n4814_1, n4815, n4817, n4818, n4819_1, n4821,
    n4822, n4824_1, n4825, n4827, n4828, n4830, n4831, n4832, n4833,
    n4834_1, n4835, n4837, n4838, n4839_1, n4840, n4842, n4843, n4844_1,
    n4845, n4847, n4848, n4849_1, n4850, n4852, n4853, n4854_1, n4855,
    n4857, n4858, n4859_1, n4860, n4862, n4863, n4864_1, n4865, n4867,
    n4868, n4869_1, n4870, n4872, n4873, n4874_1, n4875, n4877, n4878,
    n4879_1, n4880, n4882, n4883, n4884_1, n4885, n4887, n4888, n4889_1,
    n4890, n4892, n4893, n4894_1, n4895, n4897, n4898, n4899_1, n4900,
    n4902, n4903, n4904_1, n4905, n4907, n4908, n4909_1, n4910, n4912,
    n4913, n4914_1, n4915, n4917, n4918, n4919_1, n4920, n4922, n4923,
    n4924_1, n4925, n4927, n4928, n4929_1, n4930, n4932, n4933, n4934_1,
    n4935, n4937, n4938, n4939_1, n4940, n4942, n4943, n4944_1, n4945,
    n4947, n4948, n4949_1, n4950, n4952, n4953, n4954_1, n4955, n4957,
    n4958, n4959_1, n4960, n4962, n4963, n4964_1, n4965, n4967, n4968,
    n4969_1, n4970, n4972, n4973, n4974_1, n4975, n4977, n4978, n4979_1,
    n4980, n4982, n4983, n4984_1, n4985, n4986, n4987, n4988, n4989_1,
    n4990, n4991, n4992, n4993, n4994_1, n4995, n4996, n4997, n4998,
    n4999_1, n5000, n5001, n5002, n5003, n5004_1, n5005, n5007, n5008,
    n5009_1, n5010, n5011, n5012, n5013, n5014_1, n5015, n5016, n5017,
    n5018, n5019_1, n5021, n5022, n5023, n5024_1, n5025, n5026, n5027,
    n5028, n5029_1, n5031, n5032, n5033, n5034_1, n5035, n5036, n5038,
    n5039_1, n5071, n5072, n5073, n5074_1, n5075, n5076, n5077, n5078,
    n5079_1, n5080, n5081, n5082, n5083, n5084_1, n5085, n5086, n5087,
    n5088_1, n5089, n5090, n5091, n5092_1, n5093, n5094, n5095, n5096_1,
    n5097, n5098, n5099, n5100_1, n5101, n5102, n5103, n5104_1, n5105,
    n5106, n5107, n5108_1, n5109, n5110, n5111, n5112_1, n5113, n5114,
    n5115, n5116_1, n5117, n5118, n5119, n5120_1, n5121, n5122, n5123,
    n5124_1, n5125, n5126, n5127, n5128_1, n5129, n5130, n5131, n5132_1,
    n5133, n5134, n5135, n5136_1, n5137, n5138, n5139, n5140_1, n5141,
    n5142, n5143, n5144_1, n5145, n5146, n5147, n5148_1, n5149, n5150,
    n5151, n5152_1, n5153, n5154, n5155, n5156_1, n5157, n5158, n5159,
    n5160_1, n5161, n5162, n5163, n5164_1, n5165, n5166, n5167, n5168_1,
    n5169, n5170, n5171, n5172_1, n5173, n5174, n5175, n5176_1, n5177,
    n5178, n5179, n5180_1, n5181, n5182, n5183, n5184_1, n5185, n5186,
    n5187, n5188_1, n5189, n5190, n5191, n5192_1, n5193, n5194, n5195,
    n5196_1, n5197, n5198, n5199, n5200_1, n5201, n5202, n5203, n5204_1,
    n5205, n5206, n5207, n5208, n5209_1, n5210, n5211, n5212, n5213,
    n5214_1, n5215, n5216, n5217, n5218, n5219_1, n5220, n5221, n5222,
    n5223, n5224_1, n5225, n5226, n5227, n5228, n5229_1, n5230, n5231,
    n5232, n5233, n5234_1, n5235, n5236, n5237, n5238, n5239_1, n5240,
    n5241, n5242, n5243, n5244_1, n5245, n5246, n5247, n5248, n5249_1,
    n5250, n5251, n5252, n5253, n5254_1, n5255, n5256, n5257, n5258,
    n5259_1, n5260, n5261, n5262, n5263, n5264_1, n5265, n5266, n5267,
    n5268, n5269_1, n5270, n5271, n5272, n5273, n5274_1, n5275, n5276,
    n5277, n5278, n5279_1, n5280, n5281, n5282, n5283, n5284_1, n5285,
    n5286, n5287, n5288, n5289_1, n5290, n5291, n5292, n5293, n5294_1,
    n5295, n5296, n5297, n5298, n5299_1, n5300, n5301, n5302, n5303,
    n5304_1, n5305, n5306, n5307, n5308, n5309_1, n5310, n5311, n5312,
    n5313, n5314_1, n5315, n5316, n5317, n5318, n5319_1, n5320, n5321,
    n5322, n5323, n5324_1, n5325, n5326, n5327, n5328, n5329_1, n5330,
    n5331, n5332, n5333, n5334_1, n5335, n5336, n5337, n5338, n5339_1,
    n5340, n5341, n5342, n5343, n5344_1, n5345, n5346, n5347, n5348,
    n5349_1, n5350, n5351, n5352, n5353, n5354_1, n5355, n5356, n5357,
    n5358, n5359_1, n5360, n5361, n5362, n5363, n5364_1, n5365, n5366,
    n5367, n5368, n5369_1, n5370, n5371, n5372, n5373, n5374_1, n5375,
    n5376, n5377, n5378, n5379_1, n5380, n5381, n5382, n5383, n5384_1,
    n5385, n5386, n5387, n5388, n5389_1, n5390, n5391, n5392, n5393,
    n5394_1, n5395, n5396, n5397, n5398, n5399_1, n5400, n5401, n5402,
    n5403, n5404_1, n5405, n5406, n5407, n5408, n5409_1, n5410, n5411,
    n5412, n5413, n5414_1, n5415, n5416, n5417, n5418, n5419_1, n5420,
    n5421, n5422, n5423, n5424_1, n5425, n5426, n5427, n5428, n5429_1,
    n5430, n5431, n5432, n5433, n5434_1, n5435, n5436, n5437, n5438,
    n5439_1, n5440, n5441, n5442, n5443, n5444_1, n5445, n5446, n5447,
    n5448, n5449_1, n5450, n5451, n5452, n5453, n5454_1, n5455, n5456,
    n5457, n5458, n5459_1, n5460, n5461, n5462, n5463, n5464_1, n5465,
    n5466, n5467, n5468, n5469_1, n5470, n5471, n5472, n5473, n5474_1,
    n5475, n5476, n5477, n5478, n5479_1, n5480, n5481, n5482, n5483,
    n5484_1, n5485, n5486, n5487, n5488, n5489_1, n5490, n5491, n5492,
    n5493, n5494_1, n5495, n5496, n5497, n5498, n5499_1, n5500, n5501,
    n5502, n5503, n5504_1, n5505, n5506, n5507, n5508, n5509_1, n5510,
    n5511, n5512, n5513, n5514_1, n5515, n5516, n5517, n5518, n5519_1,
    n5520, n5521, n5522, n5523, n5524_1, n5525, n5526, n5527, n5528,
    n5529_1, n5530, n5531, n5532, n5533, n5534_1, n5535, n5536, n5537,
    n5538, n5539_1, n5540, n5541, n5542, n5543, n5544_1, n5545, n5546,
    n5547, n5548, n5549_1, n5550, n5551, n5552, n5553, n5554_1, n5555,
    n5556, n5557, n5558, n5559_1, n5560, n5561, n5562, n5563, n5564_1,
    n5565, n5566, n5567, n5568, n5569_1, n5570, n5571, n5572, n5573,
    n5574_1, n5575, n5576, n5577, n5578, n5579_1, n5580, n5581, n5582,
    n5583, n5584_1, n5585, n5586, n5587, n5588, n5589_1, n5590, n5591,
    n5592, n5593, n5594_1, n5595, n5596, n5597, n5598, n5599_1, n5600,
    n5601, n5602, n5603, n5604_1, n5605, n5606, n5607, n5608, n5609_1,
    n5610, n5611, n5612, n5613, n5614_1, n5615, n5616, n5617, n5618,
    n5619_1, n5620, n5621, n5622, n5623, n5624_1, n5625, n5626, n5627,
    n5628, n5629_1, n5630, n5631, n5632, n5633, n5634_1, n5635, n5636,
    n5637, n5638, n5639_1, n5640, n5641, n5642, n5643, n5644_1, n5645,
    n5646, n5647, n5648, n5649_1, n5650, n5651, n5652, n5653, n5654_1,
    n5655, n5656, n5657, n5658, n5659_1, n5660, n5661, n5662, n5663,
    n5664_1, n5665, n5666, n5667, n5668, n5669_1, n5670, n5671, n5672,
    n5673, n5674_1, n5675, n5676, n5677, n5678, n5679_1, n5680, n5681,
    n5682, n5683, n5684_1, n5685, n5686, n5687, n5688, n5689_1, n5690,
    n5691, n5692, n5693, n5694_1, n5695, n5696, n5697, n5698, n5699_1,
    n5700, n5701, n5702, n5704_1, n5705, n5706, n5707, n5708, n5709_1,
    n5710, n5711, n5713, n5714_1, n5715, n5716, n5717, n5718, n5719_1,
    n5720, n5721, n5722, n5723, n5724_1, n5725, n5726, n5728, n5729_1,
    n5730, n5731, n5732, n5733, n5734_1, n5735, n5736, n5737, n5738,
    n5739_1, n5740, n5741, n5742, n5743, n5744_1, n5745, n5746, n5747,
    n5748, n5749_1, n5750, n5751, n5752, n5753, n5754_1, n5755, n5756,
    n5757, n5758, n5759_1, n5760, n5761, n5762, n5763, n5764_1, n5765,
    n5766, n5767, n5769_1, n5770, n5771, n5772, n5773, n5774_1, n5775,
    n5776, n5777, n5778, n5779_1, n5780, n5781, n5782, n5783, n5784_1,
    n5785, n5786, n5787, n5788, n5789_1, n5790, n5791, n5792, n5793,
    n5794_1, n5795, n5796, n5797, n5798, n5799_1, n5800, n5801, n5802,
    n5803, n5804_1, n5805, n5806, n5807, n5808, n5809_1, n5810, n5811,
    n5812, n5813, n5814_1, n5815, n5816, n5817, n5818, n5819_1, n5820,
    n5821, n5822, n5823, n5824_1, n5825, n5826, n5827, n5828, n5829_1,
    n5830, n5831, n5832, n5833, n5834_1, n5835, n5836, n5837, n5838,
    n5839_1, n5840, n5841, n5842, n5843, n5844_1, n5846, n5847, n5848,
    n5849_1, n5850, n5851, n5852, n5853, n5854_1, n5855, n5856, n5857,
    n5859_1, n5860, n5861, n5862, n5863, n5864_1, n5865, n5866, n5867,
    n5868, n5869_1, n5870, n5872, n5873, n5874_1, n5875, n5876, n5877,
    n5878, n5879_1, n5880, n5881, n5882, n5883, n5885, n5886, n5887, n5888,
    n5889_1, n5890, n5891, n5892, n5893, n5894_1, n5895, n5896, n5898,
    n5899_1, n5900, n5901, n5902, n5903, n5904_1, n5905, n5906, n5907,
    n5908, n5909_1, n5911, n5912, n5913, n5914_1, n5915, n5916, n5917,
    n5918, n5919_1, n5920, n5921, n5922, n5924_1, n5925, n5926, n5927,
    n5928, n5929_1, n5930, n5931, n5932, n5933, n5934_1, n5935, n5937,
    n5938, n5939_1, n5940, n5941, n5942, n5943, n5944_1, n5945, n5946,
    n5947, n5948, n5949_1, n5950, n5951, n5952, n5953, n5954_1, n5955,
    n5956, n5957, n5958, n5959_1, n5960, n5961, n5963, n5964_1, n5965,
    n5966, n5967, n5968, n5969_1, n5970, n5972, n5973, n5974_1, n5975,
    n5976, n5977, n5978, n5979_1, n5981, n5982, n5983, n5984_1, n5985,
    n5986, n5987, n5988, n5990, n5991, n5992, n5993, n5994_1, n5995, n5996,
    n5997, n5999_1, n6000, n6001, n6002, n6003, n6004_1, n6005, n6006,
    n6008, n6009_1, n6010, n6011, n6012, n6013, n6014_1, n6015, n6017,
    n6018, n6019_1, n6020, n6021, n6022, n6023, n6024_1, n6026, n6027,
    n6028, n6029_1, n6030, n6031, n6032, n6033, n6034_1, n6035, n6036,
    n6037, n6038, n6039_1, n6040, n6041, n6042, n6043, n6044_1, n6045,
    n6046, n6047, n6048, n6049_1, n6051, n6052, n6053, n6054_1, n6055,
    n6056, n6057, n6058, n6060, n6061, n6062, n6063, n6064_1, n6065, n6066,
    n6067, n6069_1, n6070, n6071, n6072, n6073, n6074_1, n6075, n6076,
    n6078, n6079_1, n6080, n6081, n6082, n6083, n6084_1, n6085, n6087,
    n6088, n6089_1, n6090, n6091, n6092, n6093, n6094_1, n6096, n6097,
    n6098, n6099_1, n6100, n6101, n6102, n6103, n6105, n6106, n6107, n6108,
    n6109_1, n6110, n6111, n6112, n6114_1, n6115, n6116, n6117, n6118,
    n6119_1, n6120, n6121, n6122, n6123, n6124_1, n6125, n6126, n6127,
    n6128, n6129_1, n6130, n6131, n6132, n6133, n6134_1, n6135, n6136,
    n6137, n6139_1, n6140, n6141, n6142, n6143, n6144_1, n6145, n6146,
    n6148, n6149_1, n6150, n6151, n6152, n6153, n6154_1, n6155, n6157,
    n6158, n6159_1, n6160, n6161, n6162, n6163, n6164_1, n6166, n6167,
    n6168, n6169_1, n6170, n6171, n6172, n6173, n6175, n6176, n6177, n6178,
    n6179_1, n6180, n6181, n6182, n6184_1, n6185, n6186, n6187, n6188,
    n6189_1, n6190, n6191, n6193, n6194_1, n6195, n6196, n6197, n6198,
    n6199_1, n6200, n6202, n6203, n6204_1, n6205, n6206, n6207, n6208,
    n6209_1, n6210, n6211, n6212, n6213, n6214_1, n6215, n6216, n6217,
    n6218, n6219_1, n6220, n6221, n6222, n6223, n6224_1, n6225, n6226,
    n6228, n6229_1, n6230, n6231, n6232, n6233, n6234_1, n6235, n6237,
    n6238, n6239_1, n6240, n6241, n6242, n6243, n6244_1, n6246, n6247,
    n6248, n6249_1, n6250, n6251, n6252, n6253, n6255, n6256, n6257, n6258,
    n6259_1, n6260, n6261, n6262, n6264_1, n6265, n6266, n6267, n6268,
    n6269_1, n6270, n6271, n6273, n6274_1, n6275, n6276, n6277, n6278,
    n6279_1, n6280, n6282, n6283, n6284_1, n6285, n6286, n6287, n6288,
    n6289_1, n6291, n6292, n6293, n6294_1, n6295, n6296, n6297, n6298,
    n6299_1, n6300, n6301, n6302, n6303, n6304_1, n6305, n6306, n6307,
    n6308, n6309_1, n6310, n6311, n6312, n6313, n6315, n6316, n6317, n6318,
    n6319_1, n6320, n6321, n6322, n6324_1, n6325, n6326, n6327, n6328,
    n6329_1, n6330, n6331, n6333, n6334_1, n6335, n6336, n6337, n6338,
    n6339_1, n6340, n6342, n6343, n6344_1, n6345, n6346, n6347, n6348,
    n6349_1, n6351, n6352, n6353, n6354_1, n6355, n6356, n6357, n6358,
    n6360, n6361, n6362, n6363, n6364_1, n6365, n6366, n6367, n6369_1,
    n6370, n6371, n6372, n6373, n6374_1, n6375, n6376, n6378, n6379_1,
    n6380, n6381, n6382, n6383, n6384_1, n6385, n6386, n6387, n6388,
    n6389_1, n6390, n6391, n6392, n6393, n6394_1, n6395, n6396, n6397,
    n6398, n6399_1, n6401, n6402, n6403, n6404_1, n6405, n6406, n6407,
    n6408, n6410, n6411, n6412, n6413, n6414_1, n6415, n6416, n6417,
    n6419_1, n6420, n6421, n6422, n6423, n6424_1, n6425, n6426, n6428,
    n6429_1, n6430, n6431, n6432, n6433, n6434_1, n6435, n6437, n6438,
    n6439_1, n6440, n6441, n6442, n6443, n6444_1, n6446, n6447, n6448,
    n6449_1, n6450, n6451, n6452, n6453, n6455, n6456, n6457, n6458,
    n6459_1, n6460, n6461, n6462, n6464_1, n6465, n6466, n6467, n6468,
    n6469_1, n6470, n6471, n6472, n6473, n6474_1, n6475, n6476, n6477,
    n6478, n6479_1, n6480, n6481, n6482, n6483, n6484_1, n6486, n6487,
    n6488, n6489_1, n6490, n6491, n6492, n6493, n6495, n6496, n6497, n6498,
    n6499_1, n6500, n6501, n6502, n6504_1, n6505, n6506, n6507, n6508,
    n6509_1, n6510, n6511, n6513, n6514_1, n6515, n6516, n6517, n6518,
    n6519_1, n6520, n6522, n6523, n6524_1, n6525, n6526, n6527, n6528,
    n6529_1, n6531, n6532, n6533, n6534_1, n6535, n6536, n6537, n6538,
    n6540, n6541, n6542, n6543, n6544_1, n6545, n6546, n6547, n6549_1,
    n6550, n6551, n6552, n6553, n6554_1, n6555, n6556, n6557, n6558,
    n6559_1, n6560, n6561, n6562, n6563, n6564_1, n6565, n6566, n6567,
    n6568, n6570, n6571, n6572, n6573, n6574_1, n6575, n6576, n6577,
    n6579_1, n6580, n6581, n6582, n6583, n6584_1, n6585, n6586, n6588,
    n6589_1, n6590, n6591, n6592, n6593, n6594_1, n6595, n6597, n6598,
    n6599_1, n6600, n6601, n6602, n6603, n6604_1, n6606, n6607, n6608,
    n6609_1, n6610, n6611, n6612, n6613, n6615, n6616, n6617, n6618,
    n6619_1, n6620, n6621, n6622, n6624_1, n6625, n6626, n6627, n6628,
    n6629_1, n6630, n6631, n6633, n6634_1, n6635, n6636, n6637, n6638,
    n6639_1, n6640, n6641, n6642, n6643, n6644_1, n6645, n6646, n6647,
    n6648, n6649_1, n6650, n6651, n6652, n6653, n6654_1, n6655, n6657,
    n6658, n6659_1, n6660, n6661, n6662, n6663, n6664_1, n6666, n6667,
    n6668, n6669_1, n6670, n6671, n6672, n6673, n6675, n6676, n6677, n6678,
    n6679_1, n6680, n6681, n6682, n6684_1, n6685, n6686, n6687, n6688,
    n6689_1, n6690, n6691, n6693, n6694_1, n6695, n6696, n6697, n6698,
    n6699_1, n6700, n6702, n6703, n6704_1, n6705, n6706, n6707, n6708,
    n6709_1, n6711, n6712, n6713, n6714_1, n6715, n6716, n6717, n6718,
    n6720, n6721, n6722, n6723, n6724_1, n6725, n6726, n6727, n6728,
    n6729_1, n6730, n6731, n6732, n6733, n6734_1, n6735, n6736, n6737,
    n6738, n6739_1, n6740, n6741, n6742, n6744_1, n6745, n6746, n6747,
    n6748, n6749_1, n6750, n6751, n6753, n6754_1, n6755, n6756, n6757,
    n6758, n6759_1, n6760, n6762, n6763, n6764_1, n6765, n6766, n6767,
    n6768, n6769_1, n6771, n6772, n6773, n6774_1, n6775, n6776, n6777,
    n6778, n6780, n6781, n6782, n6783, n6784_1, n6785, n6786, n6787,
    n6789_1, n6790, n6791, n6792, n6793, n6794_1, n6795, n6796, n6798,
    n6799_1, n6800, n6801, n6802, n6803, n6804_1, n6805, n6807, n6808,
    n6809_1, n6810, n6811, n6812, n6813, n6814_1, n6815, n6816, n6817,
    n6818, n6819_1, n6820, n6821, n6822, n6823, n6824_1, n6825, n6826,
    n6827, n6829_1, n6830, n6831, n6832, n6833, n6834_1, n6835, n6836,
    n6838, n6839_1, n6840, n6841, n6842, n6843, n6844_1, n6845, n6847,
    n6848, n6849_1, n6850, n6851, n6852, n6853, n6854_1, n6856, n6857,
    n6858, n6859_1, n6860, n6861, n6862, n6863, n6865, n6866, n6867, n6868,
    n6869_1, n6870, n6871, n6872, n6874_1, n6875, n6876, n6877, n6878,
    n6879_1, n6880, n6881, n6883, n6884_1, n6885, n6886, n6887, n6888,
    n6889_1, n6890, n6892, n6893, n6894_1, n6895, n6896, n6897, n6898,
    n6899_1, n6900, n6901, n6902, n6903, n6904_1, n6905, n6906, n6907,
    n6908, n6909_1, n6910, n6911, n6912, n6913, n6914_1, n6915, n6917,
    n6918, n6919_1, n6920, n6921, n6922, n6923, n6924_1, n6926, n6927,
    n6928, n6929_1, n6930, n6931, n6932, n6933, n6935, n6936, n6937, n6938,
    n6939_1, n6940, n6941, n6942, n6944_1, n6945, n6946, n6947, n6948,
    n6949_1, n6950, n6951, n6953, n6954_1, n6955, n6956, n6957, n6958,
    n6959_1, n6960, n6962, n6963, n6964_1, n6965, n6966, n6967, n6968,
    n6969_1, n6971, n6972, n6973, n6974_1, n6975, n6976, n6977, n6978,
    n6980, n6981, n6982, n6983, n6984_1, n6985, n6986, n6987, n6988,
    n6989_1, n6990, n6991, n6992, n6993, n6994_1, n6995, n6996, n6997,
    n6998, n6999_1, n7001, n7002, n7003, n7004_1, n7005, n7006, n7007,
    n7008, n7010, n7011, n7012, n7013, n7014_1, n7015, n7016, n7017,
    n7019_1, n7020, n7021, n7022, n7023, n7024_1, n7025, n7026, n7028,
    n7029_1, n7030, n7031, n7032, n7033, n7034_1, n7035, n7037, n7038,
    n7039_1, n7040, n7041, n7042, n7043, n7044_1, n7046, n7047, n7048,
    n7049_1, n7050, n7051, n7052, n7053, n7055, n7056, n7057, n7058,
    n7059_1, n7060, n7061, n7062, n7064_1, n7065, n7066, n7067, n7068,
    n7069_1, n7070, n7071, n7072, n7073, n7074_1, n7075, n7076, n7077,
    n7078, n7079_1, n7080, n7081, n7082, n7083, n7085, n7086, n7087, n7088,
    n7089_1, n7090, n7091, n7092, n7094_1, n7095, n7096, n7097, n7098,
    n7099_1, n7100, n7101, n7103, n7104_1, n7105, n7106, n7107, n7108,
    n7109_1, n7110, n7112, n7113, n7114_1, n7115, n7116, n7117, n7118,
    n7119_1, n7121, n7122, n7123, n7124_1, n7125, n7126, n7127, n7128,
    n7130, n7131, n7132, n7133, n7134_1, n7135, n7136, n7137, n7139_1,
    n7140, n7141, n7142, n7143, n7144_1, n7145, n7146, n7148, n7149_1,
    n7150, n7151, n7152, n7153, n7154_1, n7155, n7156, n7157, n7158,
    n7159_1, n7160, n7161, n7162, n7163, n7164_1, n7165, n7166, n7168,
    n7169_1, n7170, n7171, n7172, n7173, n7174_1, n7175, n7177, n7178,
    n7179_1, n7180, n7181, n7182, n7183, n7184_1, n7186, n7187, n7188,
    n7189_1, n7190, n7191, n7192, n7193, n7195, n7196, n7197, n7198,
    n7199_1, n7200, n7201, n7202, n7204_1, n7205, n7206, n7207, n7208,
    n7209_1, n7210, n7211, n7213, n7214_1, n7215, n7216, n7217, n7218,
    n7219_1, n7220, n7222, n7223, n7224_1, n7225, n7226, n7227, n7228,
    n7229_1, n7231, n7232, n7233, n7234_1, n7235, n7236, n7237, n7238,
    n7239_1, n7240, n7242, n7243, n7244_1, n7245, n7246, n7247, n7249_1,
    n7250, n7251, n7252, n7253, n7254_1, n7255, n7256, n7258, n7259_1,
    n7260, n7261, n7262, n7263, n7264_1, n7266, n7267, n7268_1, n7269,
    n7270, n7271, n7272, n7274, n7275, n7276, n7277, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7320, n7321, n7322, n7323, n7324,
    n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
    n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
    n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
    n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7859,
    n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
    n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
    n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
    n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
    n8464, n8465, n8466, n8467, n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
    n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
    n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
    n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
    n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
    n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
    n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9431, n9432, n9433, n9434, n9435, n9436,
    n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
    n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
    n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
    n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
    n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
    n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9988, n9989, n9990, n9991, n9992, n9993,
    n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10072, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
    n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
    n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
    n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
    n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
    n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
    n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10358, n10359,
    n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
    n10369, n10370, n10371, n10372, n10373, n10374, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
    n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
    n10416, n10417, n10418, n10419, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
    n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
    n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
    n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
    n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
    n10943, n10944, n10945, n10946, n10947, n10948, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
    n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11053, n11054, n11055, n11056,
    n11058, n11059, n11060, n11061, n11063, n11064, n11065, n11066, n11068,
    n11069, n11070, n11071, n11073, n11074, n11075, n11076, n11078, n11079,
    n11080, n11081, n11083, n11084, n11085, n11086, n11088, n11089, n11090,
    n11091, n11093, n11094, n11095, n11096, n11098, n11099, n11100, n11101,
    n11103, n11104, n11105, n11106, n11108, n11109, n11110, n11111, n11113,
    n11114, n11115, n11116, n11118, n11119, n11120, n11121, n11123, n11124,
    n11125, n11126, n11128, n11129, n11130, n11132, n11133, n11134, n11136,
    n11137, n11138, n11140, n11141, n11142, n11144, n11145, n11146, n11148,
    n11149, n11150, n11152, n11153, n11154, n11156, n11157, n11158, n11160,
    n11161, n11162, n11164, n11165, n11166, n11168, n11169, n11170, n11172,
    n11173, n11174, n11176, n11177, n11178, n11180, n11181, n11182, n11184,
    n11185, n11186, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11199, n11200, n11201, n11202, n11204, n11205,
    n11206, n11207, n11209, n11210, n11211, n11212, n11214, n11215, n11216,
    n11217, n11219, n11220, n11221, n11222, n11224, n11225, n11226, n11227,
    n11229, n11230, n11231, n11232, n11234, n11235, n11236, n11237, n11239,
    n11240, n11241, n11242, n11244, n11245, n11246, n11247, n11249, n11250,
    n11251, n11252, n11254, n11255, n11256, n11257, n11259, n11260, n11261,
    n11262, n11264, n11265, n11266, n11267, n11269, n11270, n11271, n11272,
    n11274, n11275, n11276, n11277, n11278, n11280, n11281, n11282, n11283,
    n11285, n11286, n11287, n11288, n11290, n11291, n11292, n11293, n11295,
    n11296, n11297, n11298, n11300, n11301, n11302, n11303, n11305, n11306,
    n11307, n11308, n11310, n11311, n11312, n11313, n11315, n11316, n11317,
    n11318, n11320, n11321, n11322, n11323, n11325, n11326, n11327, n11328,
    n11330, n11331, n11332, n11333, n11335, n11336, n11337, n11338, n11340,
    n11341, n11342, n11343, n11345, n11346, n11347, n11348, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
    n11382, n11383, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
    n11392, n11393, n11394, n11395, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11408, n11409, n11410, n11411,
    n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
    n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
    n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
    n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
    n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
    n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
    n11542, n11543, n11544, n11545, n11546, n11547, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759, n11761, n11762, n11763,
    n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
    n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
    n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
    n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
    n11800, n11801, n11802, n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
    n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
    n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
    n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
    n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
    n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12053, n12054, n12055, n12056, n12057,
    n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
    n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
    n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
    n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
    n12094, n12095, n12096, n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
    n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
    n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
    n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12386, n12387,
    n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
    n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
    n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
    n12433, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
    n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530, n12532, n12533, n12534,
    n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
    n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
    n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
    n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
    n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12598, n12599, n12600,
    n12601, n12602, n12603, n12604, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12625, n12626, n12627, n12628, n12629, n12630,
    n12631, n12632, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
    n12661, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12710, n12711,
    n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12796, n12797, n12798, n12799, n12800, n12801,
    n12802, n12803, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
    n12832, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12881, n12882,
    n12883, n12884, n12885, n12886, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12954, n12955, n12956, n12957,
    n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
    n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
    n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
    n13162, n13163, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
    n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
    n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
    n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
    n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
    n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
    n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
    n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
    n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
    n13667, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
    n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
    n13714, n13715, n13716, n13717, n13718, n13719, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
    n13770, n13771, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
    n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
    n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13812, n13813, n13814, n13815, n13816,
    n13817, n13818, n13819, n13821, n13822, n13823, n13825, n13826, n13827,
    n13829, n13830, n13832, n13833, n13834, n13836, n13837, n13839, n13840,
    n13841, n13842, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13860,
    n13861, n13862, n13864, n13865, n13867, n13868, n13869, n13871, n13873,
    n13874, n13875, n13876, n13877, n13879, n13880, n13881, n13883, n13884,
    n13885, n13887, n13888, n13890, n13891, n13893, n13894, n13896, n13897,
    n13898, n13899, n13900, n13901, n13903, n13904, n13905, n13906, n13908,
    n13909, n13910, n13911, n13913, n13914, n13915, n13916, n13918, n13919,
    n13920, n13921, n13923, n13924, n13925, n13926, n13928, n13929, n13930,
    n13931, n13933, n13934, n13935, n13936, n13938, n13939, n13940, n13941,
    n13943, n13944, n13945, n13946, n13948, n13949, n13950, n13951, n13953,
    n13954, n13955, n13956, n13958, n13959, n13960, n13961, n13963, n13964,
    n13965, n13966, n13968, n13969, n13970, n13971, n13973, n13974, n13975,
    n13976, n13978, n13979, n13980, n13981, n13983, n13984, n13985, n13986,
    n13988, n13989, n13990, n13991, n13993, n13994, n13995, n13996, n13998,
    n13999, n14000, n14001, n14003, n14004, n14005, n14006, n14008, n14009,
    n14010, n14011, n14013, n14014, n14015, n14016, n14018, n14019, n14020,
    n14021, n14023, n14024, n14025, n14026, n14028, n14029, n14030, n14031,
    n14033, n14034, n14035, n14036, n14038, n14039, n14040, n14041, n14043,
    n14044, n14045, n14046, n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
    n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
    n14082, n14083, n14084, n14085, n14086, n14087, n14089, n14090, n14091,
    n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14101,
    n14102, n14103, n14104, n14105, n14106, n14108, n14109, n14141, n14142,
    n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
    n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
    n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
    n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
    n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
    n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
    n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
    n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
    n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
    n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
    n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
    n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
    n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
    n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
    n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
    n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
    n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
    n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
    n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
    n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
    n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
    n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
    n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
    n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
    n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
    n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
    n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
    n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
    n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
    n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
    n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
    n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
    n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
    n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
    n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
    n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
    n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
    n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
    n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
    n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
    n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
    n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
    n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
    n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
    n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
    n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
    n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
    n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
    n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
    n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
    n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
    n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
    n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
    n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
    n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
    n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
    n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
    n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
    n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
    n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
    n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
    n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
    n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
    n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
    n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
    n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
    n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
    n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
    n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
    n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
    n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
    n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
    n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
    n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
    n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
    n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
    n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
    n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
    n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
    n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
    n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
    n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
    n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
    n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
    n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
    n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
    n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
    n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
    n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
    n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
    n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
    n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
    n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
    n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
    n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
    n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
    n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
    n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
    n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15446, n15447, n15448, n15449, n15450,
    n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
    n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
    n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
    n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
    n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
    n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
    n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
    n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
    n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
    n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
    n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
    n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
    n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
    n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
    n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
    n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
    n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15637, n15638, n15639, n15640, n15641, n15642,
    n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
    n15652, n15653, n15654, n15655, n15656, n15657, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
    n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15703, n15704, n15705, n15706, n15707, n15708,
    n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
    n15718, n15719, n15720, n15721, n15722, n15723, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
    n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
    n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15769, n15770, n15771, n15772, n15773, n15774,
    n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
    n15793, n15794, n15795, n15796, n15797, n15798, n15800, n15801, n15802,
    n15803, n15804, n15805, n15806, n15807, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15818, n15819, n15820, n15821, n15822,
    n15823, n15824, n15825, n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
    n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15863,
    n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
    n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15896, n15897, n15898, n15899, n15900,
    n15901, n15902, n15903, n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
    n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15941,
    n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15950, n15951,
    n15952, n15953, n15954, n15955, n15956, n15957, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
    n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16028, n16029,
    n16030, n16031, n16032, n16033, n16034, n16035, n16037, n16038, n16039,
    n16040, n16041, n16042, n16043, n16044, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16055, n16056, n16057, n16058, n16059,
    n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
    n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
    n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
    n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16097,
    n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16113, n16115, n16116, n16117,
    n16118, n16119, n16120, n16121, n16122, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16133, n16134, n16135, n16136, n16137,
    n16138, n16139, n16140, n16142, n16143, n16144, n16145, n16146, n16147,
    n16148, n16149, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
    n16196, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
    n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16216,
    n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232, n16234, n16235, n16236,
    n16237, n16238, n16239, n16240, n16241, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16282, n16283, n16284,
    n16285, n16286, n16287, n16288, n16289, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16309, n16310, n16311, n16312, n16313, n16314,
    n16315, n16316, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
    n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
    n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
    n16363, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16419, n16420, n16421, n16422, n16423,
    n16424, n16425, n16426, n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457, n16459, n16460, n16461,
    n16462, n16463, n16464, n16465, n16466, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
    n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16522,
    n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
    n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
    n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16587, n16588, n16589, n16590,
    n16591, n16592, n16593, n16594, n16596, n16597, n16598, n16599, n16600,
    n16601, n16602, n16603, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
    n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
    n16639, n16640, n16641, n16642, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
    n16669, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
    n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16736, n16737,
    n16738, n16739, n16740, n16741, n16742, n16743, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
    n16788, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
    n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841, n16843, n16844, n16845,
    n16846, n16847, n16848, n16849, n16850, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
    n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
    n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
    n16924, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
    n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
    n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17019, n17020, n17021, n17022,
    n17023, n17024, n17025, n17026, n17028, n17029, n17030, n17031, n17032,
    n17033, n17034, n17035, n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
    n17053, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
    n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17138, n17139, n17140, n17141,
    n17142, n17143, n17144, n17145, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17185, n17186, n17187, n17188, n17189, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17199, n17200, n17201, n17202,
    n17203, n17204, n17205, n17206, n17208, n17209, n17210, n17211, n17212,
    n17213, n17214, n17216, n17217, n17218, n17219, n17221, n17222, n17223,
    n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
    n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
    n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
    n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
    n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
    n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
    n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
    n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
    n17296, n17297, n17298, n17300, n17301, n17302, n17303, n17304, n17305,
    n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
    n17315, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
    n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
    n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
    n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
    n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
    n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
    n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
    n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485, n17487, n17488, n17489,
    n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
    n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
    n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
    n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
    n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
    n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
    n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
    n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
    n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
    n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
    n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
    n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
    n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
    n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
    n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
    n17671, n17672, n17673, n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17766, n17767, n17768, n17769, n17770, n17771,
    n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
    n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
    n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
    n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
    n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
    n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
    n17880, n17881, n17882, n17883, n17884, n17885, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
    n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
    n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
    n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
    n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
    n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
    n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
    n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
    n17998, n17999, n18000, n18001, n18003, n18004, n18005, n18006, n18007,
    n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
    n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
    n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
    n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
    n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
    n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
    n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
    n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
    n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
    n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
    n18116, n18117, n18118, n18119, n18120, n18121, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18249, n18250, n18251, n18252,
    n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
    n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
    n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
    n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
    n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
    n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
    n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
    n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
    n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
    n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18492, n18493, n18494, n18495, n18496, n18497,
    n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
    n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
    n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
    n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
    n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
    n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
    n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
    n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
    n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18887, n18888,
    n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
    n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
    n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
    n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
    n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
    n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
    n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
    n18979, n18980, n18981, n18982, n18983, n18984, n18986, n18987, n18988,
    n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
    n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
    n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
    n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
    n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
    n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
    n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
    n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
    n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
    n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
    n19079, n19080, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
    n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
    n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
    n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
    n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349, n19351, n19352, n19353,
    n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
    n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
    n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
    n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
    n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
    n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
    n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
    n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
    n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
    n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
    n19481, n19482, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
    n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
    n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
    n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
    n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
    n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
    n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
    n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
    n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
    n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
    n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
    n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
    n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
    n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
    n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
    n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
    n19810, n19811, n19812, n19813, n19814, n19815, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
    n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
    n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
    n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19880, n19881, n19882, n19883,
    n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
    n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
    n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
    n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20157,
    n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
    n20176, n20177, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20190, n20191, n20192, n20193, n20194, n20195,
    n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20204, n20205,
    n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
    n20244, n20245, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
    n20254, n20255, n20256, n20257, n20258, n20259, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
    n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20331,
    n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20345, n20346, n20347, n20348, n20349, n20350,
    n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
    n20370, n20371, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
    n20380, n20381, n20382, n20383, n20384, n20385, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20415, n20416, n20417, n20418,
    n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
    n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20443, n20444, n20445, n20446, n20447,
    n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20457,
    n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
    n20467, n20468, n20469, n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
    n20496, n20497, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
    n20506, n20507, n20508, n20509, n20510, n20511, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20541, n20542, n20543, n20544,
    n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
    n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20583,
    n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
    n20593, n20594, n20595, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20622,
    n20623, n20624, n20625, n20626, n20627, n20628, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
    n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20662, n20663,
    n20664, n20665, n20666, n20667, n20668, n20670, n20671, n20672, n20673,
    n20674, n20675, n20676, n20678, n20679, n20680, n20681, n20683, n20684,
    n20685, n20686, n20688, n20689, n20690, n20691, n20693, n20694, n20695,
    n20696, n20698, n20699, n20700, n20701, n20703, n20704, n20705, n20706,
    n20708, n20709, n20710, n20711, n20713, n20714, n20715, n20716, n20718,
    n20719, n20720, n20722, n20723, n20724, n20726, n20727, n20728, n20730,
    n20731, n20732, n20734, n20735, n20736, n20738, n20739, n20740, n20742,
    n20743, n20744, n20746, n20747, n20748, n20750, n20751, n20752, n20754,
    n20755, n20756, n20758, n20759, n20760, n20762, n20763, n20764, n20766,
    n20767, n20768, n20770, n20771, n20772, n20774, n20775, n20776, n20778,
    n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
    n20788, n20789, n20790, n20791, n20792, n20794, n20795, n20796, n20797,
    n20799, n20800, n20801, n20802, n20804, n20805, n20806, n20807, n20809,
    n20810, n20811, n20812, n20814, n20815, n20816, n20817, n20819, n20820,
    n20821, n20822, n20824, n20825, n20826, n20827, n20829, n20830, n20831,
    n20832, n20834, n20835, n20836, n20837, n20839, n20840, n20841, n20842,
    n20844, n20845, n20846, n20847, n20849, n20850, n20851, n20852, n20854,
    n20855, n20856, n20857, n20859, n20860, n20861, n20862, n20864, n20865,
    n20866, n20867, n20869, n20870, n20871, n20872, n20873, n20875, n20876,
    n20877, n20878, n20880, n20881, n20882, n20883, n20885, n20886, n20887,
    n20888, n20890, n20891, n20892, n20893, n20895, n20896, n20897, n20898,
    n20900, n20901, n20902, n20903, n20905, n20906, n20907, n20908, n20910,
    n20911, n20912, n20913, n20915, n20916, n20917, n20918, n20920, n20921,
    n20922, n20923, n20925, n20926, n20927, n20928, n20930, n20931, n20932,
    n20933, n20935, n20936, n20937, n20938, n20940, n20941, n20942, n20943,
    n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960, n20962, n20963, n20964,
    n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
    n20974, n20975, n20976, n20977, n20978, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
    n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
    n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
    n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
    n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
    n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21092, n21093, n21094, n21095, n21096,
    n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
    n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
    n21115, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
    n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21161, n21162,
    n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
    n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
    n21181, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21208, n21209,
    n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21227, n21228,
    n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
    n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
    n21247, n21248, n21249, n21250, n21252, n21253, n21254, n21255, n21256,
    n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21299, n21300, n21301, n21302, n21303,
    n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
    n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
    n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
    n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
    n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
    n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
    n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
    n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
    n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
    n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
    n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
    n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
    n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
    n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
    n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
    n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
    n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
    n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
    n21550, n21551, n21552, n21553, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21669,
    n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
    n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
    n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
    n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
    n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
    n21724, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
    n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
    n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
    n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
    n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
    n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
    n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
    n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
    n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
    n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21832, n21833,
    n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
    n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
    n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
    n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21906,
    n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
    n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
    n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
    n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
    n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
    n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
    n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
    n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
    n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
    n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
    n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
    n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
    n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
    n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
    n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
    n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
    n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
    n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
    n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
    n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
    n22198, n22199, n22200, n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
    n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
    n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
    n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
    n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
    n22354, n22355, n22356, n22357, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22368, n22369, n22370, n22371, n22373, n22374,
    n22375, n22376, n22378, n22379, n22380, n22381, n22383, n22384, n22385,
    n22386, n22388, n22389, n22390, n22391, n22393, n22394, n22395, n22396,
    n22398, n22399, n22400, n22401, n22403, n22404, n22405, n22406, n22408,
    n22409, n22410, n22411, n22413, n22414, n22415, n22416, n22418, n22419,
    n22420, n22421, n22423, n22424, n22425, n22426, n22428, n22429, n22430,
    n22431, n22433, n22434, n22435, n22436, n22438, n22439, n22440, n22441,
    n22443, n22444, n22445, n22446, n22448, n22449, n22450, n22451, n22453,
    n22454, n22455, n22456, n22458, n22459, n22460, n22461, n22463, n22464,
    n22465, n22466, n22468, n22469, n22470, n22471, n22473, n22474, n22475,
    n22476, n22478, n22479, n22480, n22481, n22483, n22484, n22485, n22486,
    n22488, n22489, n22490, n22491, n22493, n22494, n22495, n22496, n22498,
    n22499, n22500, n22501, n22503, n22504, n22505, n22506, n22508, n22509,
    n22510, n22511, n22513, n22514, n22515, n22516, n22518, n22519, n22521,
    n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
    n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
    n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
    n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557,
    n22558, n22559, n22560, n22561, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
    n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22604, n22605,
    n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
    n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
    n22624, n22625, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
    n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
    n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22677, n22678, n22679, n22680,
    n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
    n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
    n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
    n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22743, n22744, n22745, n22746,
    n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
    n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
    n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
    n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
    n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22875, n22876, n22877, n22878,
    n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
    n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
    n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22941, n22942, n22943, n22944,
    n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
    n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
    n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
    n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
    n23020, n23021, n23022, n23023, n23024, n23025, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
    n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
    n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
    n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
    n23086, n23087, n23088, n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
    n23105, n23106, n23107, n23108, n23109, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
    n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23132, n23133,
    n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
    n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
    n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
    n23171, n23172, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
    n23190, n23191, n23192, n23193, n23195, n23196, n23197, n23198, n23199,
    n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
    n23209, n23210, n23211, n23212, n23213, n23214, n23216, n23217, n23218,
    n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23234, n23235, n23236, n23237,
    n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
    n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23273, n23274,
    n23275, n23276, n23277, n23278, n23279, n23281, n23282, n23284, n23285,
    n23286, n23288, n23289, n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23299, n23300, n23302, n23303, n23304, n23305, n23307, n23308,
    n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23326, n23327,
    n23328, n23330, n23331, n23333, n23334, n23335, n23337, n23339, n23340,
    n23341, n23342, n23343, n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23355, n23356, n23357, n23359, n23360, n23362,
    n23363, n23365, n23366, n23368, n23369, n23370, n23371, n23372, n23373,
    n23375, n23376, n23377, n23378, n23380, n23381, n23382, n23383, n23385,
    n23386, n23387, n23388, n23390, n23391, n23392, n23393, n23395, n23396,
    n23397, n23398, n23400, n23401, n23402, n23403, n23405, n23406, n23407,
    n23408, n23410, n23411, n23412, n23413, n23415, n23416, n23417, n23418,
    n23420, n23421, n23422, n23423, n23425, n23426, n23427, n23428, n23430,
    n23431, n23432, n23433, n23435, n23436, n23437, n23438, n23440, n23441,
    n23442, n23443, n23445, n23446, n23447, n23448, n23450, n23451, n23452,
    n23453, n23455, n23456, n23457, n23458, n23460, n23461, n23462, n23463,
    n23465, n23466, n23467, n23468, n23470, n23471, n23472, n23473, n23475,
    n23476, n23477, n23478, n23480, n23481, n23482, n23483, n23485, n23486,
    n23487, n23488, n23490, n23491, n23492, n23493, n23495, n23496, n23497,
    n23498, n23500, n23501, n23502, n23503, n23505, n23506, n23507, n23508,
    n23510, n23511, n23512, n23513, n23515, n23516, n23517, n23518, n23520,
    n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
    n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
    n23539, n23540, n23541, n23542, n23543, n23545, n23546, n23547, n23548,
    n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
    n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
    n23569, n23570, n23571, n23572, n23573, n23574, n23576, n23577, n23609,
    n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
    n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
    n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
    n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
    n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
    n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
    n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
    n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
    n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
    n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
    n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
    n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
    n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
    n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
    n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
    n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
    n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
    n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
    n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
    n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
    n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
    n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
    n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
    n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
    n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
    n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
    n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
    n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
    n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
    n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
    n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
    n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
    n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
    n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
    n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
    n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
    n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
    n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
    n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
    n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
    n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
    n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
    n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
    n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
    n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
    n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
    n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
    n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
    n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
    n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
    n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
    n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24568, n24569, n24570, n24571, n24572, n24573,
    n24574, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24620, n24621,
    n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
    n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
    n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
    n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
    n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
    n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
    n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
    n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
    n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
    n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
    n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
    n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
    n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
    n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
    n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
    n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
    n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
    n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
    n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
    n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
    n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
    n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
    n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
    n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837,
    n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
    n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
    n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
    n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
    n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
    n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
    n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
    n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909,
    n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
    n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
    n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
    n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
    n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
    n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
    n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
    n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
    n25059, n25060, n25061, n25062, n25064, n25065, n25066, n25067, n25068,
    n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
    n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
    n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25139, n25140, n25141, n25142, n25143,
    n25144, n25145, n25146, n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
    n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25193, n25194,
    n25195, n25196, n25197, n25198, n25199, n25200, n25202, n25203, n25204,
    n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
    n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
    n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25271, n25272,
    n25273, n25274, n25275, n25276, n25277, n25278, n25280, n25281, n25282,
    n25283, n25284, n25285, n25286, n25287, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
    n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
    n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
    n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25340,
    n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25349, n25350,
    n25351, n25352, n25353, n25354, n25355, n25356, n25358, n25359, n25360,
    n25361, n25362, n25363, n25364, n25365, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25376, n25377, n25378, n25379, n25380,
    n25381, n25382, n25383, n25385, n25386, n25387, n25388, n25389, n25390,
    n25391, n25392, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
    n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
    n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
    n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25445, n25446, n25447, n25448,
    n25449, n25450, n25451, n25452, n25454, n25455, n25456, n25457, n25458,
    n25459, n25460, n25461, n25463, n25464, n25465, n25466, n25467, n25468,
    n25469, n25470, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
    n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526,
    n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25546, n25547,
    n25548, n25549, n25550, n25551, n25552, n25553, n25555, n25556, n25557,
    n25558, n25559, n25560, n25561, n25562, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25582, n25583, n25584, n25585, n25586, n25587,
    n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
    n25606, n25607, n25608, n25609, n25610, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25621, n25622, n25623, n25624, n25625,
    n25626, n25627, n25628, n25630, n25631, n25632, n25633, n25634, n25635,
    n25636, n25637, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
    n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25666,
    n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25704,
    n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25713, n25714,
    n25715, n25716, n25717, n25718, n25719, n25720, n25722, n25723, n25724,
    n25725, n25726, n25727, n25728, n25729, n25731, n25732, n25733, n25734,
    n25735, n25736, n25737, n25738, n25740, n25741, n25742, n25743, n25744,
    n25745, n25746, n25747, n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
    n25765, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774,
    n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
    n25793, n25794, n25795, n25796, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25807, n25808, n25809, n25810, n25811, n25812,
    n25813, n25814, n25816, n25817, n25818, n25819, n25820, n25821, n25822,
    n25823, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
    n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25852, n25853,
    n25854, n25855, n25856, n25857, n25858, n25859, n25861, n25862, n25863,
    n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
    n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25908, n25909, n25910, n25911,
    n25912, n25913, n25914, n25915, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25935, n25936, n25937, n25938, n25939, n25940, n25941,
    n25942, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
    n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
    n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
    n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
    n25980, n25981, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
    n25990, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
    n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26010,
    n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26019, n26020,
    n26021, n26022, n26023, n26024, n26025, n26026, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26037, n26038, n26039, n26040,
    n26041, n26042, n26043, n26044, n26046, n26047, n26048, n26049, n26050,
    n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
    n26069, n26070, n26071, n26072, n26073, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26084, n26085, n26086, n26087, n26088,
    n26089, n26090, n26091, n26093, n26094, n26095, n26096, n26097, n26098,
    n26099, n26100, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
    n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26129,
    n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26138, n26139,
    n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
    n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
    n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
    n26167, n26168, n26169, n26170, n26171, n26173, n26174, n26175, n26176,
    n26177, n26178, n26179, n26180, n26182, n26183, n26184, n26185, n26186,
    n26187, n26188, n26189, n26191, n26192, n26193, n26194, n26195, n26196,
    n26197, n26198, n26200, n26201, n26202, n26203, n26204, n26205, n26206,
    n26207, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
    n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26236, n26237,
    n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246,
    n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
    n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26265,
    n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281, n26283, n26284, n26285,
    n26286, n26287, n26288, n26289, n26290, n26292, n26293, n26294, n26295,
    n26296, n26297, n26298, n26299, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26310, n26311, n26312, n26313, n26314, n26315,
    n26316, n26317, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
    n26326, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
    n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26358, n26359, n26360, n26361, n26362, n26363,
    n26364, n26365, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
    n26374, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
    n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26394,
    n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26403, n26404,
    n26405, n26406, n26407, n26408, n26409, n26410, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26421, n26422, n26423, n26424,
    n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
    n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
    n26443, n26444, n26445, n26446, n26447, n26448, n26450, n26451, n26452,
    n26453, n26454, n26455, n26456, n26457, n26459, n26460, n26461, n26462,
    n26463, n26464, n26465, n26466, n26468, n26469, n26470, n26471, n26472,
    n26473, n26474, n26475, n26477, n26478, n26479, n26480, n26481, n26482,
    n26483, n26484, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
    n26493, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
    n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26513,
    n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
    n26524, n26525, n26526, n26527, n26528, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26538, n26539, n26540, n26541, n26542, n26543,
    n26544, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26554,
    n26555, n26556, n26557, n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26567, n26568, n26569, n26571, n26572, n26573, n26574,
    n26575, n26576, n26577, n26578, n26579, n26580, n26582, n26583, n26584,
    n26585, n26586, n26587, n26588, n26589, n26591, n26592, n26593, n26594,
    n26595, n26596, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
    n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
    n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622,
    n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
    n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
    n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
    n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
    n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
    n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
    n26677, n26678, n26679, n26681, n26682, n26683, n26684, n26685, n26686,
    n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
    n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
    n26723, n26724, n26725, n26726, n26727, n26728, n26730, n26731, n26732,
    n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
    n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750,
    n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
    n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
    n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
    n26778, n26779, n26780, n26781, n26783, n26784, n26785, n26786, n26787,
    n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
    n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
    n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
    n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
    n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
    n26933, n26934, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
    n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
    n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
    n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
    n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
    n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
    n27042, n27043, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
    n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
    n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
    n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
    n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
    n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
    n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
    n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
    n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
    n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
    n27142, n27143, n27144, n27145, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
    n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
    n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
    n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214,
    n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27229, n27230, n27231, n27232, n27233,
    n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
    n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
    n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
    n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
    n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278,
    n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
    n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
    n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
    n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27348, n27349, n27350, n27351,
    n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
    n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
    n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
    n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
    n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
    n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
    n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
    n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
    n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
    n27433, n27434, n27435, n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
    n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
    n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
    n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
    n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
    n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
    n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
    n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
    n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
    n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
    n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614,
    n27615, n27616, n27617, n27618, n27619, n27621, n27622, n27623, n27624,
    n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
    n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
    n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
    n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
    n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
    n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678,
    n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
    n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
    n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
    n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27794, n27795, n27796, n27797,
    n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
    n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
    n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
    n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
    n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
    n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
    n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27882, n27883, n27884, n27885, n27886, n27887, n27888,
    n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
    n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
    n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
    n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
    n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
    n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
    n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
    n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960,
    n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
    n27970, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
    n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
    n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
    n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28033, n28034,
    n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
    n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
    n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061,
    n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070,
    n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28080,
    n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
    n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
    n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
    n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
    n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
    n28126, n28127, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
    n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
    n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177, n28179, n28180, n28181,
    n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190,
    n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
    n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
    n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
    n28218, n28219, n28220, n28221, n28222, n28224, n28225, n28226, n28227,
    n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
    n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245,
    n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254,
    n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263,
    n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
    n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
    n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318,
    n28319, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
    n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
    n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
    n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
    n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
    n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
    n28374, n28375, n28376, n28378, n28379, n28380, n28381, n28382, n28383,
    n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
    n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
    n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
    n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
    n28420, n28421, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
    n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
    n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28520, n28521,
    n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
    n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
    n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
    n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
    n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
    n28613, n28614, n28615, n28616, n28617, n28619, n28620, n28621, n28622,
    n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
    n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
    n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
    n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
    n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
    n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
    n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28685, n28686,
    n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
    n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
    n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
    n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
    n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
    n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750,
    n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
    n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
    n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
    n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28814,
    n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
    n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
    n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
    n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
    n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
    n28860, n28861, n28862, n28863, n28865, n28866, n28867, n28868, n28869,
    n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878,
    n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
    n28888, n28889, n28890, n28891, n28892, n28893, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
    n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
    n28925, n28926, n28927, n28928, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
    n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
    n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29003, n29004, n29005, n29006, n29007, n29008,
    n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
    n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29036,
    n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045,
    n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
    n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
    n29064, n29065, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
    n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
    n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
    n29092, n29093, n29094, n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
    n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
    n29129, n29130, n29131, n29132, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
    n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162, n29164, n29165, n29166,
    n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
    n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
    n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
    n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
    n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
    n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
    n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29265, n29266, n29267, n29268,
    n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277,
    n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
    n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333,
    n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
    n29352, n29353, n29354, n29356, n29357, n29358, n29359, n29360, n29361,
    n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
    n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
    n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388,
    n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397,
    n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
    n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
    n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
    n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
    n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
    n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
    n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29460, n29461,
    n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
    n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
    n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
    n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
    n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29524, n29525,
    n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
    n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
    n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
    n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
    n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
    n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607,
    n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616,
    n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
    n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
    n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
    n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652,
    n29653, n29654, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
    n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
    n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29782, n29783, n29785, n29786, n29787, n29788, n29789, n29790,
    n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
    n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
    n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
    n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
    n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844,
    n29845, n29846, n29847, n29848, n29849, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
    n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
    n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
    n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981,
    n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
    n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
    n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
    n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
    n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
    n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
    n30036, n30037, n30039, n30040, n30041, n30042, n30043, n30044, n30045,
    n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
    n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
    n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
    n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
    n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
    n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
    n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
    n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
    n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
    n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
    n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172,
    n30173, n30174, n30175, n30176, n30177, n30178, n30180, n30181, n30182,
    n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
    n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
    n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
    n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236,
    n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
    n30246, n30247, n30248, n30250, n30251, n30252, n30253, n30254, n30255,
    n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
    n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
    n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
    n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
    n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300,
    n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309,
    n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
    n30319, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
    n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
    n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364,
    n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
    n30383, n30384, n30385, n30386, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
    n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428,
    n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
    n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30455, n30456,
    n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
    n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474,
    n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
    n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30508, n30509, n30510, n30511, n30512,
    n30513, n30514, n30515, n30517, n30518, n30519, n30520, n30521, n30522,
    n30523, n30524, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
    n30533, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
    n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30553,
    n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569, n30571, n30572, n30573,
    n30574, n30575, n30577, n30578, n30579, n30580, n30581, n30583, n30584,
    n30585, n30586, n30587, n30589, n30590, n30591, n30592, n30593, n30595,
    n30596, n30597, n30598, n30599, n30601, n30602, n30603, n30604, n30605,
    n30607, n30608, n30609, n30610, n30611, n30613, n30614, n30615, n30616,
    n30617, n30619, n30620, n30621, n30622, n30624, n30625, n30626, n30627,
    n30629, n30630, n30631, n30632, n30634, n30635, n30636, n30637, n30639,
    n30640, n30641, n30642, n30644, n30645, n30646, n30647, n30649, n30650,
    n30651, n30652, n30654, n30655, n30656, n30657, n30659, n30660, n30661,
    n30662, n30664, n30665, n30666, n30667, n30669, n30670, n30671, n30672,
    n30674, n30675, n30676, n30677, n30679, n30680, n30681, n30682, n30684,
    n30685, n30686, n30687, n30689, n30690, n30691, n30692, n30694, n30695,
    n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
    n30705, n30706, n30708, n30709, n30710, n30711, n30713, n30714, n30715,
    n30716, n30718, n30719, n30720, n30721, n30723, n30724, n30725, n30726,
    n30728, n30729, n30730, n30731, n30733, n30734, n30735, n30736, n30738,
    n30739, n30740, n30741, n30743, n30744, n30745, n30746, n30748, n30749,
    n30750, n30751, n30753, n30754, n30755, n30756, n30758, n30759, n30760,
    n30761, n30763, n30764, n30765, n30766, n30768, n30769, n30770, n30771,
    n30773, n30774, n30775, n30776, n30778, n30779, n30780, n30781, n30783,
    n30784, n30785, n30786, n30787, n30789, n30790, n30791, n30792, n30794,
    n30795, n30796, n30797, n30799, n30800, n30801, n30802, n30804, n30805,
    n30806, n30807, n30809, n30810, n30811, n30812, n30814, n30815, n30816,
    n30817, n30819, n30820, n30821, n30822, n30824, n30825, n30826, n30827,
    n30829, n30830, n30831, n30832, n30834, n30835, n30836, n30837, n30839,
    n30840, n30841, n30842, n30844, n30845, n30846, n30847, n30849, n30850,
    n30851, n30852, n30854, n30855, n30856, n30857, n30860, n30861, n30862,
    n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30881,
    n30882, n30883, n30884, n30886, n30887, n30888, n30889, n30891, n30892,
    n30893, n30894, n30896, n30897, n30898, n30899, n30901, n30902, n30903,
    n30904, n30906, n30907, n30908, n30909, n30911, n30912, n30913, n30914,
    n30916, n30917, n30918, n30919, n30921, n30922, n30923, n30924, n30926,
    n30927, n30928, n30929, n30931, n30932, n30933, n30934, n30936, n30937,
    n30938, n30939, n30941, n30942, n30943, n30944, n30946, n30947, n30948,
    n30949, n30951, n30952, n30953, n30954, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30966, n30967, n30968, n30969,
    n30970, n30971, n30973, n30974, n30975, n30976, n30977, n30978, n30980,
    n30981, n30982, n30983, n30984, n30985, n30987, n30988, n30989, n30990,
    n30991, n30992, n30994, n30995, n30996, n30997, n30998, n30999, n31001,
    n31002, n31003, n31004, n31005, n31006, n31008, n31009, n31010, n31011,
    n31012, n31013, n31015, n31016, n31017, n31018, n31019, n31020, n31022,
    n31023, n31024, n31025, n31026, n31027, n31029, n31030, n31031, n31032,
    n31033, n31034, n31036, n31037, n31038, n31039, n31040, n31041, n31043,
    n31044, n31045, n31046, n31047, n31048, n31050, n31051, n31052, n31053,
    n31054, n31055, n31057, n31058, n31059, n31060, n31061, n31062, n31064,
    n31065, n31066, n31067, n31068, n31070, n31071, n31072, n31073, n31074,
    n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31084,
    n31085, n31086, n31087, n31089, n31090, n31091, n31092, n31094, n31095,
    n31096, n31097, n31099, n31100, n31101, n31102, n31104, n31105, n31106,
    n31107, n31109, n31110, n31111, n31112, n31114, n31115, n31116, n31117,
    n31119, n31120, n31121, n31122, n31124, n31125, n31126, n31127, n31129,
    n31130, n31131, n31132, n31134, n31135, n31136, n31137, n31139, n31140,
    n31141, n31142, n31144, n31145, n31146, n31147, n31149, n31150, n31151,
    n31152, n31154, n31155, n31156, n31157, n31159, n31160, n31161, n31162,
    n31164, n31165, n31166, n31167, n31169, n31170, n31171, n31172, n31174,
    n31175, n31176, n31177, n31179, n31180, n31181, n31182, n31184, n31185,
    n31186, n31187, n31189, n31190, n31191, n31192, n31194, n31195, n31196,
    n31197, n31199, n31200, n31201, n31202, n31204, n31205, n31206, n31207,
    n31209, n31210, n31211, n31212, n31214, n31215, n31216, n31217, n31219,
    n31220, n31221, n31222, n31224, n31225, n31226, n31227, n31229, n31230,
    n31231, n31232, n31234, n31235, n31237, n31238, n31239, n31240, n31241,
    n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
    n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
    n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
    n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277,
    n31278, n31279, n31280, n31281, n31282, n31283, n31285, n31286, n31287,
    n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
    n31297, n31298, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
    n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325,
    n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
    n31335, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
    n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
    n31354, n31355, n31356, n31357, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
    n31373, n31374, n31375, n31376, n31377, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
    n31392, n31393, n31394, n31395, n31396, n31398, n31399, n31400, n31401,
    n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
    n31411, n31412, n31413, n31414, n31416, n31417, n31418, n31419, n31420,
    n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31434, n31435, n31436, n31437, n31438, n31439,
    n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
    n31449, n31450, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
    n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
    n31468, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
    n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31506,
    n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
    n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31524, n31525,
    n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534,
    n31535, n31536, n31537, n31538, n31539, n31540, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
    n31554, n31555, n31556, n31557, n31558, n31560, n31561, n31562, n31563,
    n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
    n31573, n31574, n31575, n31576, n31578, n31579, n31580, n31581, n31582,
    n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31596, n31597, n31598, n31599, n31600, n31601,
    n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
    n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629,
    n31630, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31649,
    n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
    n31659, n31660, n31661, n31662, n31663, n31664, n31666, n31667, n31668,
    n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677,
    n31678, n31679, n31680, n31681, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
    n31697, n31698, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
    n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725,
    n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
    n31745, n31746, n31747, n31748, n31749, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
    n31764, n31765, n31766, n31768, n31769, n31770, n31771, n31772, n31773,
    n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
    n31783, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
    n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
    n31812, n31813, n31814, n31815, n31816, n31817, n31819, n31820, n31821,
    n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
    n31831, n31832, n31833, n31834, n31836, n31837, n31838, n31839, n31840,
    n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
    n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873, n31875, n31876, n31877,
    n31878, n31879, n31880, n31881, n31882, n31884, n31885, n31886, n31888,
    n31889, n31890, n31892, n31893, n31895, n31896, n31898, n31899, n31901,
    n31902, n31903, n31904, n31906, n31907, n31908, n31909, n31910, n31911,
    n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
    n31922, n31923, n31924, n31926, n31927, n31929, n31930, n31931, n31933,
    n31935, n31936, n31937, n31938, n31939, n31941, n31942, n31943, n31944,
    n31945, n270, n275, n280, n285, n290, n295, n300, n305, n310, n315,
    n320, n325, n330, n335, n340, n345, n350, n355, n360, n365, n370, n375,
    n380, n385, n390, n395, n400, n405, n410, n415, n420, n425, n430, n435,
    n440, n445, n450, n455, n460, n465, n470, n475, n480, n485, n490, n495,
    n500, n505, n510, n515, n520, n525, n530, n535, n540, n545, n550, n555,
    n560, n565, n570, n575, n580, n585, n590, n595, n600, n605, n610, n615,
    n620, n625, n630, n635, n640, n645, n650, n655, n660, n665, n670, n675,
    n680, n685, n690, n695, n700, n705, n710, n715, n720, n725, n730, n735,
    n740, n745, n750, n755, n760, n765, n770, n775, n780, n785, n790, n795,
    n800, n805, n810, n815, n820, n825, n830, n835, n840, n845, n850, n855,
    n860, n865, n870, n875, n880, n885, n890, n895, n900, n905, n910, n915,
    n920, n925, n930, n935, n940, n945, n950, n955, n960, n965, n970, n975,
    n980, n985, n990, n995, n1000, n1005, n1010, n1015, n1020, n1025,
    n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075,
    n1080, n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1120, n1125,
    n1130, n1135, n1140, n1145, n1150, n1155, n1160, n1165, n1170, n1175,
    n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225,
    n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275,
    n1280, n1285, n1290, n1295, n1300, n1305, n1310, n1315, n1320, n1325,
    n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365, n1370, n1375,
    n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415, n1420, n1425,
    n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465, n1470, n1475,
    n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515, n1520, n1525,
    n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575,
    n1580, n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625,
    n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675,
    n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725,
    n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775,
    n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820, n1825,
    n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875,
    n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920, n1925,
    n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970, n1975,
    n1980, n1985, n1990, n1995, n2000, n2005, n2010, n2015, n2020, n2025,
    n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070, n2075,
    n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120, n2125,
    n2130, n2135, n2140, n2144, n2148, n2152, n2156, n2160, n2164, n2168,
    n2172, n2176, n2180, n2184, n2188, n2192, n2196, n2200, n2204, n2208,
    n2212, n2216, n2220, n2224, n2228, n2232, n2236, n2240, n2244, n2248,
    n2252, n2256, n2260, n2264, n2268, n2273, n2278, n2283, n2288, n2293,
    n2298, n2303, n2308, n2313, n2318, n2323, n2328, n2333, n2338, n2343,
    n2348, n2353, n2358, n2363, n2368, n2373, n2378, n2383, n2388, n2393,
    n2398, n2403, n2408, n2413, n2418, n2423, n2428, n2433, n2438, n2443,
    n2448, n2453, n2458, n2463, n2468, n2473, n2478, n2483, n2488, n2493,
    n2498, n2503, n2508, n2513, n2518, n2523, n2528, n2533, n2538, n2543,
    n2548, n2553, n2558, n2563, n2568, n2573, n2578, n2583, n2588, n2593,
    n2598, n2603, n2608, n2613, n2618, n2623, n2628, n2633, n2638, n2643,
    n2648, n2653, n2658, n2663, n2668, n2673, n2678, n2683, n2688, n2693,
    n2698, n2703, n2708, n2713, n2718, n2723, n2728, n2733, n2738, n2743,
    n2748, n2753, n2758, n2763, n2768, n2772, n2777, n2782, n2787, n2792,
    n2796, n2800, n2805, n2809, n2814, n2819, n2824, n2829, n2834, n2839,
    n2844, n2849, n2854, n2859, n2864, n2869, n2874, n2879, n2884, n2889,
    n2894, n2899, n2904, n2909, n2914, n2919, n2924, n2929, n2934, n2939,
    n2944, n2949, n2954, n2959, n2964, n2969, n2974, n2979, n2984, n2989,
    n2994, n2999, n3004, n3009, n3014, n3019, n3024, n3029, n3034, n3039,
    n3044, n3049, n3054, n3059, n3064, n3069, n3074, n3079, n3084, n3089,
    n3094, n3099, n3104, n3109, n3114, n3119, n3124, n3129, n3134, n3139,
    n3144, n3149, n3154, n3159, n3164, n3169, n3174, n3179, n3184, n3189,
    n3194, n3199, n3204, n3209, n3214, n3219, n3224, n3229, n3234, n3239,
    n3244, n3249, n3254, n3259, n3264, n3269, n3274, n3279, n3284, n3289,
    n3294, n3299, n3304, n3309, n3314, n3319, n3324, n3329, n3334, n3339,
    n3344, n3349, n3354, n3359, n3364, n3369, n3374, n3379, n3384, n3389,
    n3394, n3399, n3404, n3409, n3414, n3419, n3424, n3429, n3434, n3439,
    n3444, n3449, n3454, n3459, n3464, n3469, n3474, n3479, n3484, n3489,
    n3494, n3499, n3504, n3509, n3514, n3519, n3524, n3529, n3534, n3539,
    n3544, n3549, n3554, n3559, n3564, n3569, n3574, n3579, n3584, n3589,
    n3594, n3599, n3604, n3609, n3614, n3619, n3624, n3629, n3634, n3639,
    n3644, n3649, n3654, n3659, n3664, n3669, n3674, n3679, n3684, n3689,
    n3694, n3699, n3704, n3709, n3714, n3719, n3724, n3729, n3734, n3739,
    n3744, n3749, n3754, n3759, n3764, n3769, n3774, n3779, n3784, n3789,
    n3794, n3799, n3804, n3809, n3814, n3819, n3824, n3829, n3834, n3839,
    n3844, n3849, n3854, n3859, n3864, n3869, n3874, n3879, n3884, n3889,
    n3894, n3899, n3904, n3909, n3914, n3919, n3924, n3929, n3934, n3939,
    n3944, n3949, n3954, n3959, n3964, n3969, n3974, n3979, n3984, n3989,
    n3994, n3999, n4004, n4009, n4014, n4019, n4024, n4029, n4034, n4039,
    n4044, n4049, n4054, n4059, n4064, n4069, n4074, n4079, n4084, n4089,
    n4094, n4099, n4104, n4109, n4114, n4119, n4124, n4129, n4134, n4139,
    n4144, n4149, n4154, n4159, n4164, n4169, n4174, n4179, n4184, n4189,
    n4194, n4199, n4204, n4209, n4214, n4219, n4224, n4229, n4234, n4239,
    n4244, n4249, n4254, n4259, n4264, n4269, n4274, n4279, n4284, n4289,
    n4294, n4299, n4304, n4309, n4314, n4319, n4324, n4329, n4334, n4339,
    n4344, n4349, n4354, n4359, n4364, n4369, n4374, n4379, n4384, n4389,
    n4394, n4399, n4404, n4409, n4414, n4419, n4424, n4429, n4434, n4439,
    n4444, n4449, n4454, n4459, n4464, n4469, n4474, n4479, n4484, n4489,
    n4494, n4499, n4504, n4509, n4514, n4519, n4524, n4529, n4534, n4539,
    n4544, n4549, n4554, n4559, n4564, n4569, n4574, n4579, n4584, n4589,
    n4594, n4599, n4604, n4609, n4614, n4619, n4624, n4629, n4634, n4639,
    n4644, n4649, n4654, n4659, n4664, n4669, n4674, n4679, n4684, n4689,
    n4694, n4699, n4704, n4709, n4714, n4719, n4724, n4729, n4734, n4739,
    n4744, n4749, n4754, n4759, n4764, n4769, n4774, n4779, n4784, n4789,
    n4794, n4799, n4804, n4809, n4814, n4819, n4824, n4829, n4834, n4839,
    n4844, n4849, n4854, n4859, n4864, n4869, n4874, n4879, n4884, n4889,
    n4894, n4899, n4904, n4909, n4914, n4919, n4924, n4929, n4934, n4939,
    n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979, n4984, n4989,
    n4994, n4999, n5004, n5009, n5014, n5019, n5024, n5029, n5034, n5039,
    n5044, n5049, n5054, n5059, n5064, n5069, n5074, n5079, n5084, n5088,
    n5092, n5096, n5100, n5104, n5108, n5112, n5116, n5120, n5124, n5128,
    n5132, n5136, n5140, n5144, n5148, n5152, n5156, n5160, n5164, n5168,
    n5172, n5176, n5180, n5184, n5188, n5192, n5196, n5200, n5204, n5209,
    n5214, n5219, n5224, n5229, n5234, n5239, n5244, n5249, n5254, n5259,
    n5264, n5269, n5274, n5279, n5284, n5289, n5294, n5299, n5304, n5309,
    n5314, n5319, n5324, n5329, n5334, n5339, n5344, n5349, n5354, n5359,
    n5364, n5369, n5374, n5379, n5384, n5389, n5394, n5399, n5404, n5409,
    n5414, n5419, n5424, n5429, n5434, n5439, n5444, n5449, n5454, n5459,
    n5464, n5469, n5474, n5479, n5484, n5489, n5494, n5499, n5504, n5509,
    n5514, n5519, n5524, n5529, n5534, n5539, n5544, n5549, n5554, n5559,
    n5564, n5569, n5574, n5579, n5584, n5589, n5594, n5599, n5604, n5609,
    n5614, n5619, n5624, n5629, n5634, n5639, n5644, n5649, n5654, n5659,
    n5664, n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709,
    n5714, n5719, n5724, n5729, n5734, n5739, n5744, n5749, n5754, n5759,
    n5764, n5769, n5774, n5779, n5784, n5789, n5794, n5799, n5804, n5809,
    n5814, n5819, n5824, n5829, n5834, n5839, n5844, n5849, n5854, n5859,
    n5864, n5869, n5874, n5879, n5884, n5889, n5894, n5899, n5904, n5909,
    n5914, n5919, n5924, n5929, n5934, n5939, n5944, n5949, n5954, n5959,
    n5964, n5969, n5974, n5979, n5984, n5989, n5994, n5999, n6004, n6009,
    n6014, n6019, n6024, n6029, n6034, n6039, n6044, n6049, n6054, n6059,
    n6064, n6069, n6074, n6079, n6084, n6089, n6094, n6099, n6104, n6109,
    n6114, n6119, n6124, n6129, n6134, n6139, n6144, n6149, n6154, n6159,
    n6164, n6169, n6174, n6179, n6184, n6189, n6194, n6199, n6204, n6209,
    n6214, n6219, n6224, n6229, n6234, n6239, n6244, n6249, n6254, n6259,
    n6264, n6269, n6274, n6279, n6284, n6289, n6294, n6299, n6304, n6309,
    n6314, n6319, n6324, n6329, n6334, n6339, n6344, n6349, n6354, n6359,
    n6364, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409,
    n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6454, n6459,
    n6464, n6469, n6474, n6479, n6484, n6489, n6494, n6499, n6504, n6509,
    n6514, n6519, n6524, n6529, n6534, n6539, n6544, n6549, n6554, n6559,
    n6564, n6569, n6574, n6579, n6584, n6589, n6594, n6599, n6604, n6609,
    n6614, n6619, n6624, n6629, n6634, n6639, n6644, n6649, n6654, n6659,
    n6664, n6669, n6674, n6679, n6684, n6689, n6694, n6699, n6704, n6709,
    n6714, n6719, n6724, n6729, n6734, n6739, n6744, n6749, n6754, n6759,
    n6764, n6769, n6774, n6779, n6784, n6789, n6794, n6799, n6804, n6809,
    n6814, n6819, n6824, n6829, n6834, n6839, n6844, n6849, n6854, n6859,
    n6864, n6869, n6874, n6879, n6884, n6889, n6894, n6899, n6904, n6909,
    n6914, n6919, n6924, n6929, n6934, n6939, n6944, n6949, n6954, n6959,
    n6964, n6969, n6974, n6979, n6984, n6989, n6994, n6999, n7004, n7009,
    n7014, n7019, n7024, n7029, n7034, n7039, n7044, n7049, n7054, n7059,
    n7064, n7069, n7074, n7079, n7084, n7089, n7094, n7099, n7104, n7109,
    n7114, n7119, n7124, n7129, n7134, n7139, n7144, n7149, n7154, n7159,
    n7164, n7169, n7174, n7179, n7184, n7189, n7194, n7199, n7204, n7209,
    n7214, n7219, n7224, n7229, n7234, n7239, n7244, n7249, n7254, n7259,
    n7264, n7268, n7273;
  assign n4380 = P3_DATAO_REG_30_ & ~P3_DATAO_REG_31_;
  assign n4381 = P1_DATAO_REG_30_ & ~P1_DATAO_REG_31_;
  assign n4382 = P2_DATAO_REG_30_ & ~P2_DATAO_REG_31_;
  assign n4383 = ~n4380 & ~n4381;
  assign n4384_1 = ~n4382 & n4383;
  assign n4385 = P3_ADDRESS_REG_29_ & n4384_1;
  assign n4386 = P2_ADDRESS_REG_29_ & ~n4384_1;
  assign U355 = n4385 | n4386;
  assign n4388 = P3_ADDRESS_REG_28_ & n4384_1;
  assign n4389_1 = P2_ADDRESS_REG_28_ & ~n4384_1;
  assign U356 = n4388 | n4389_1;
  assign n4391 = P3_ADDRESS_REG_27_ & n4384_1;
  assign n4392 = P2_ADDRESS_REG_27_ & ~n4384_1;
  assign U357 = n4391 | n4392;
  assign n4394_1 = P3_ADDRESS_REG_26_ & n4384_1;
  assign n4395 = P2_ADDRESS_REG_26_ & ~n4384_1;
  assign U358 = n4394_1 | n4395;
  assign n4397 = P3_ADDRESS_REG_25_ & n4384_1;
  assign n4398 = P2_ADDRESS_REG_25_ & ~n4384_1;
  assign U359 = n4397 | n4398;
  assign n4400 = P3_ADDRESS_REG_24_ & n4384_1;
  assign n4401 = P2_ADDRESS_REG_24_ & ~n4384_1;
  assign U360 = n4400 | n4401;
  assign n4403 = P3_ADDRESS_REG_23_ & n4384_1;
  assign n4404_1 = P2_ADDRESS_REG_23_ & ~n4384_1;
  assign U361 = n4403 | n4404_1;
  assign n4406 = P3_ADDRESS_REG_22_ & n4384_1;
  assign n4407 = P2_ADDRESS_REG_22_ & ~n4384_1;
  assign U362 = n4406 | n4407;
  assign n4409_1 = P3_ADDRESS_REG_21_ & n4384_1;
  assign n4410 = P2_ADDRESS_REG_21_ & ~n4384_1;
  assign U363 = n4409_1 | n4410;
  assign n4412 = P3_ADDRESS_REG_20_ & n4384_1;
  assign n4413 = P2_ADDRESS_REG_20_ & ~n4384_1;
  assign U364 = n4412 | n4413;
  assign n4415 = P3_ADDRESS_REG_19_ & n4384_1;
  assign n4416 = P2_ADDRESS_REG_19_ & ~n4384_1;
  assign U366 = n4415 | n4416;
  assign n4418 = P3_ADDRESS_REG_18_ & n4384_1;
  assign n4419_1 = P2_ADDRESS_REG_18_ & ~n4384_1;
  assign U367 = n4418 | n4419_1;
  assign n4421 = P3_ADDRESS_REG_17_ & n4384_1;
  assign n4422 = P2_ADDRESS_REG_17_ & ~n4384_1;
  assign U368 = n4421 | n4422;
  assign n4424_1 = P3_ADDRESS_REG_16_ & n4384_1;
  assign n4425 = P2_ADDRESS_REG_16_ & ~n4384_1;
  assign U369 = n4424_1 | n4425;
  assign n4427 = P3_ADDRESS_REG_15_ & n4384_1;
  assign n4428 = P2_ADDRESS_REG_15_ & ~n4384_1;
  assign U370 = n4427 | n4428;
  assign n4430 = P3_ADDRESS_REG_14_ & n4384_1;
  assign n4431 = P2_ADDRESS_REG_14_ & ~n4384_1;
  assign U371 = n4430 | n4431;
  assign n4433 = P3_ADDRESS_REG_13_ & n4384_1;
  assign n4434_1 = P2_ADDRESS_REG_13_ & ~n4384_1;
  assign U372 = n4433 | n4434_1;
  assign n4436 = P3_ADDRESS_REG_12_ & n4384_1;
  assign n4437 = P2_ADDRESS_REG_12_ & ~n4384_1;
  assign U373 = n4436 | n4437;
  assign n4439_1 = P3_ADDRESS_REG_11_ & n4384_1;
  assign n4440 = P2_ADDRESS_REG_11_ & ~n4384_1;
  assign U374 = n4439_1 | n4440;
  assign n4442 = P3_ADDRESS_REG_10_ & n4384_1;
  assign n4443 = P2_ADDRESS_REG_10_ & ~n4384_1;
  assign U375 = n4442 | n4443;
  assign n4445 = P3_ADDRESS_REG_9_ & n4384_1;
  assign n4446 = P2_ADDRESS_REG_9_ & ~n4384_1;
  assign U347 = n4445 | n4446;
  assign n4448 = P3_ADDRESS_REG_8_ & n4384_1;
  assign n4449_1 = P2_ADDRESS_REG_8_ & ~n4384_1;
  assign U348 = n4448 | n4449_1;
  assign n4451 = P3_ADDRESS_REG_7_ & n4384_1;
  assign n4452 = P2_ADDRESS_REG_7_ & ~n4384_1;
  assign U349 = n4451 | n4452;
  assign n4454_1 = P3_ADDRESS_REG_6_ & n4384_1;
  assign n4455 = P2_ADDRESS_REG_6_ & ~n4384_1;
  assign U350 = n4454_1 | n4455;
  assign n4457 = P3_ADDRESS_REG_5_ & n4384_1;
  assign n4458 = P2_ADDRESS_REG_5_ & ~n4384_1;
  assign U351 = n4457 | n4458;
  assign n4460 = P3_ADDRESS_REG_4_ & n4384_1;
  assign n4461 = P2_ADDRESS_REG_4_ & ~n4384_1;
  assign U352 = n4460 | n4461;
  assign n4463 = P3_ADDRESS_REG_3_ & n4384_1;
  assign n4464_1 = P2_ADDRESS_REG_3_ & ~n4384_1;
  assign U353 = n4463 | n4464_1;
  assign n4466 = P3_ADDRESS_REG_2_ & n4384_1;
  assign n4467 = P2_ADDRESS_REG_2_ & ~n4384_1;
  assign U354 = n4466 | n4467;
  assign n4469_1 = P3_ADDRESS_REG_1_ & n4384_1;
  assign n4470 = P2_ADDRESS_REG_1_ & ~n4384_1;
  assign U365 = n4469_1 | n4470;
  assign n4472 = P3_ADDRESS_REG_0_ & n4384_1;
  assign n4473 = P2_ADDRESS_REG_0_ & ~n4384_1;
  assign U376 = n4472 | n4473;
  assign n4475 = ~P1_BE_N_REG_3_ & ~P1_BE_N_REG_1_;
  assign n4476 = ~P1_D_C_N_REG & n4475;
  assign n4477 = ~P1_ADS_N_REG & n4476;
  assign n4478 = ~P1_BE_N_REG_0_ & n4477;
  assign n4479_1 = ~P1_ADDRESS_REG_20_ & ~P1_ADDRESS_REG_13_;
  assign n4480 = ~P1_ADDRESS_REG_3_ & n4479_1;
  assign n4481 = ~P1_ADDRESS_REG_27_ & n4480;
  assign n4482 = ~P1_ADDRESS_REG_2_ & n4481;
  assign n4483 = ~P1_ADDRESS_REG_5_ & n4482;
  assign n4484_1 = ~P1_ADDRESS_REG_15_ & n4483;
  assign n4485 = ~P1_ADDRESS_REG_26_ & ~P1_ADDRESS_REG_21_;
  assign n4486 = ~P1_ADDRESS_REG_28_ & n4485;
  assign n4487 = ~P1_ADDRESS_REG_6_ & n4486;
  assign n4488 = ~P1_ADDRESS_REG_12_ & n4487;
  assign n4489_1 = ~P1_ADDRESS_REG_14_ & n4488;
  assign n4490 = ~P1_ADDRESS_REG_4_ & n4489_1;
  assign n4491 = ~P1_ADDRESS_REG_16_ & ~P1_ADDRESS_REG_0_;
  assign n4492 = ~P1_ADDRESS_REG_18_ & n4491;
  assign n4493 = ~P1_ADDRESS_REG_8_ & n4492;
  assign n4494_1 = ~P1_ADDRESS_REG_23_ & n4493;
  assign n4495 = ~P1_ADDRESS_REG_1_ & n4494_1;
  assign n4496 = ~P1_ADDRESS_REG_11_ & n4495;
  assign n4497 = ~P1_ADDRESS_REG_17_ & ~P1_ADDRESS_REG_9_;
  assign n4498 = ~P1_ADDRESS_REG_7_ & n4497;
  assign n4499_1 = ~P1_ADDRESS_REG_22_ & n4498;
  assign n4500 = ~P1_ADDRESS_REG_10_ & n4499_1;
  assign n4501 = ~P1_ADDRESS_REG_19_ & n4500;
  assign n4502 = ~P1_ADDRESS_REG_25_ & n4501;
  assign n4503 = ~P1_ADDRESS_REG_24_ & n4502;
  assign n4504_1 = n4484_1 & n4490;
  assign n4505 = n4496 & n4504_1;
  assign n4506 = n4503 & n4505;
  assign n4507 = P1_ADDRESS_REG_29_ & ~n4506;
  assign n4508 = ~P1_BE_N_REG_2_ & P1_M_IO_N_REG;
  assign n4509_1 = P1_W_R_N_REG & n4508;
  assign n4510 = n4478 & n4509_1;
  assign n605 = ~n4507 | ~n4510;
  assign n4512 = P1_DATAO_REG_0_ & ~n605;
  assign n4513 = ~P2_ADDRESS_REG_20_ & ~P2_ADDRESS_REG_13_;
  assign n4514_1 = ~P2_ADDRESS_REG_3_ & n4513;
  assign n4515 = ~P2_ADDRESS_REG_27_ & n4514_1;
  assign n4516 = ~P2_ADDRESS_REG_2_ & n4515;
  assign n4517 = ~P2_ADDRESS_REG_5_ & n4516;
  assign n4518 = ~P2_ADDRESS_REG_15_ & n4517;
  assign n4519_1 = ~P2_ADDRESS_REG_26_ & ~P2_ADDRESS_REG_21_;
  assign n4520 = ~P2_ADDRESS_REG_28_ & n4519_1;
  assign n4521 = ~P2_ADDRESS_REG_6_ & n4520;
  assign n4522 = ~P2_ADDRESS_REG_12_ & n4521;
  assign n4523 = ~P2_ADDRESS_REG_14_ & n4522;
  assign n4524_1 = ~P2_ADDRESS_REG_4_ & n4523;
  assign n4525 = ~P2_ADDRESS_REG_16_ & ~P2_ADDRESS_REG_0_;
  assign n4526 = ~P2_ADDRESS_REG_18_ & n4525;
  assign n4527 = ~P2_ADDRESS_REG_8_ & n4526;
  assign n4528 = ~P2_ADDRESS_REG_23_ & n4527;
  assign n4529_1 = ~P2_ADDRESS_REG_1_ & n4528;
  assign n4530 = ~P2_ADDRESS_REG_11_ & n4529_1;
  assign n4531 = ~P2_ADDRESS_REG_17_ & ~P2_ADDRESS_REG_9_;
  assign n4532 = ~P2_ADDRESS_REG_7_ & n4531;
  assign n4533 = ~P2_ADDRESS_REG_22_ & n4532;
  assign n4534_1 = ~P2_ADDRESS_REG_10_ & n4533;
  assign n4535 = ~P2_ADDRESS_REG_19_ & n4534_1;
  assign n4536 = ~P2_ADDRESS_REG_25_ & n4535;
  assign n4537 = ~P2_ADDRESS_REG_24_ & n4536;
  assign n4538 = n4518 & n4524_1;
  assign n4539_1 = n4530 & n4538;
  assign n4540 = n4537 & n4539_1;
  assign n4541 = P2_ADDRESS_REG_29_ & ~n4540;
  assign n4542 = ~P2_BE_N_REG_3_ & ~P2_D_C_N_REG;
  assign n4543 = ~P2_BE_N_REG_0_ & ~P2_ADS_N_REG;
  assign n4544_1 = ~P2_BE_N_REG_2_ & n4543;
  assign n4545 = ~P2_BE_N_REG_1_ & n4544_1;
  assign n4546 = P2_W_R_N_REG & P2_M_IO_N_REG;
  assign n4547 = n4542 & n4546;
  assign n4548 = n4545 & n4547;
  assign n4549_1 = n4541 & n4548;
  assign n4550 = n605 & ~n4549_1;
  assign n4551 = BUF1_REG_0_ & n4550;
  assign n4552 = n605 & ~n4550;
  assign n4553 = P2_DATAO_REG_0_ & n4552;
  assign n4554_1 = ~n4512 & ~n4551;
  assign n270 = n4553 | ~n4554_1;
  assign n4556 = P1_DATAO_REG_1_ & ~n605;
  assign n4557 = BUF1_REG_1_ & n4550;
  assign n4558 = P2_DATAO_REG_1_ & n4552;
  assign n4559_1 = ~n4556 & ~n4557;
  assign n275 = n4558 | ~n4559_1;
  assign n4561 = P1_DATAO_REG_2_ & ~n605;
  assign n4562 = BUF1_REG_2_ & n4550;
  assign n4563 = P2_DATAO_REG_2_ & n4552;
  assign n4564_1 = ~n4561 & ~n4562;
  assign n280 = n4563 | ~n4564_1;
  assign n4566 = P1_DATAO_REG_3_ & ~n605;
  assign n4567 = BUF1_REG_3_ & n4550;
  assign n4568 = P2_DATAO_REG_3_ & n4552;
  assign n4569_1 = ~n4566 & ~n4567;
  assign n285 = n4568 | ~n4569_1;
  assign n4571 = P1_DATAO_REG_4_ & ~n605;
  assign n4572 = BUF1_REG_4_ & n4550;
  assign n4573 = P2_DATAO_REG_4_ & n4552;
  assign n4574_1 = ~n4571 & ~n4572;
  assign n290 = n4573 | ~n4574_1;
  assign n4576 = P1_DATAO_REG_5_ & ~n605;
  assign n4577 = BUF1_REG_5_ & n4550;
  assign n4578 = P2_DATAO_REG_5_ & n4552;
  assign n4579_1 = ~n4576 & ~n4577;
  assign n295 = n4578 | ~n4579_1;
  assign n4581 = P1_DATAO_REG_6_ & ~n605;
  assign n4582 = BUF1_REG_6_ & n4550;
  assign n4583 = P2_DATAO_REG_6_ & n4552;
  assign n4584_1 = ~n4581 & ~n4582;
  assign n300 = n4583 | ~n4584_1;
  assign n4586 = P1_DATAO_REG_7_ & ~n605;
  assign n4587 = BUF1_REG_7_ & n4550;
  assign n4588 = P2_DATAO_REG_7_ & n4552;
  assign n4589_1 = ~n4586 & ~n4587;
  assign n305 = n4588 | ~n4589_1;
  assign n4591 = P1_DATAO_REG_8_ & ~n605;
  assign n4592 = BUF1_REG_8_ & n4550;
  assign n4593 = P2_DATAO_REG_8_ & n4552;
  assign n4594_1 = ~n4591 & ~n4592;
  assign n310 = n4593 | ~n4594_1;
  assign n4596 = P1_DATAO_REG_9_ & ~n605;
  assign n4597 = BUF1_REG_9_ & n4550;
  assign n4598 = P2_DATAO_REG_9_ & n4552;
  assign n4599_1 = ~n4596 & ~n4597;
  assign n315 = n4598 | ~n4599_1;
  assign n4601 = P1_DATAO_REG_10_ & ~n605;
  assign n4602 = BUF1_REG_10_ & n4550;
  assign n4603 = P2_DATAO_REG_10_ & n4552;
  assign n4604_1 = ~n4601 & ~n4602;
  assign n320 = n4603 | ~n4604_1;
  assign n4606 = P1_DATAO_REG_11_ & ~n605;
  assign n4607 = BUF1_REG_11_ & n4550;
  assign n4608 = P2_DATAO_REG_11_ & n4552;
  assign n4609_1 = ~n4606 & ~n4607;
  assign n325 = n4608 | ~n4609_1;
  assign n4611 = P1_DATAO_REG_12_ & ~n605;
  assign n4612 = BUF1_REG_12_ & n4550;
  assign n4613 = P2_DATAO_REG_12_ & n4552;
  assign n4614_1 = ~n4611 & ~n4612;
  assign n330 = n4613 | ~n4614_1;
  assign n4616 = P1_DATAO_REG_13_ & ~n605;
  assign n4617 = BUF1_REG_13_ & n4550;
  assign n4618 = P2_DATAO_REG_13_ & n4552;
  assign n4619_1 = ~n4616 & ~n4617;
  assign n335 = n4618 | ~n4619_1;
  assign n4621 = P1_DATAO_REG_14_ & ~n605;
  assign n4622 = BUF1_REG_14_ & n4550;
  assign n4623 = P2_DATAO_REG_14_ & n4552;
  assign n4624_1 = ~n4621 & ~n4622;
  assign n340 = n4623 | ~n4624_1;
  assign n4626 = P1_DATAO_REG_15_ & ~n605;
  assign n4627 = BUF1_REG_15_ & n4550;
  assign n4628 = P2_DATAO_REG_15_ & n4552;
  assign n4629_1 = ~n4626 & ~n4627;
  assign n345 = n4628 | ~n4629_1;
  assign n4631 = P1_DATAO_REG_16_ & ~n605;
  assign n4632 = BUF1_REG_16_ & n4550;
  assign n4633 = P2_DATAO_REG_16_ & n4552;
  assign n4634_1 = ~n4631 & ~n4632;
  assign n350 = n4633 | ~n4634_1;
  assign n4636 = P1_DATAO_REG_17_ & ~n605;
  assign n4637 = BUF1_REG_17_ & n4550;
  assign n4638 = P2_DATAO_REG_17_ & n4552;
  assign n4639_1 = ~n4636 & ~n4637;
  assign n355 = n4638 | ~n4639_1;
  assign n4641 = P1_DATAO_REG_18_ & ~n605;
  assign n4642 = BUF1_REG_18_ & n4550;
  assign n4643 = P2_DATAO_REG_18_ & n4552;
  assign n4644_1 = ~n4641 & ~n4642;
  assign n360 = n4643 | ~n4644_1;
  assign n4646 = P1_DATAO_REG_19_ & ~n605;
  assign n4647 = BUF1_REG_19_ & n4550;
  assign n4648 = P2_DATAO_REG_19_ & n4552;
  assign n4649_1 = ~n4646 & ~n4647;
  assign n365 = n4648 | ~n4649_1;
  assign n4651 = P1_DATAO_REG_20_ & ~n605;
  assign n4652 = BUF1_REG_20_ & n4550;
  assign n4653 = P2_DATAO_REG_20_ & n4552;
  assign n4654_1 = ~n4651 & ~n4652;
  assign n370 = n4653 | ~n4654_1;
  assign n4656 = P1_DATAO_REG_21_ & ~n605;
  assign n4657 = BUF1_REG_21_ & n4550;
  assign n4658 = P2_DATAO_REG_21_ & n4552;
  assign n4659_1 = ~n4656 & ~n4657;
  assign n375 = n4658 | ~n4659_1;
  assign n4661 = P1_DATAO_REG_22_ & ~n605;
  assign n4662 = BUF1_REG_22_ & n4550;
  assign n4663 = P2_DATAO_REG_22_ & n4552;
  assign n4664_1 = ~n4661 & ~n4662;
  assign n380 = n4663 | ~n4664_1;
  assign n4666 = P1_DATAO_REG_23_ & ~n605;
  assign n4667 = BUF1_REG_23_ & n4550;
  assign n4668 = P2_DATAO_REG_23_ & n4552;
  assign n4669_1 = ~n4666 & ~n4667;
  assign n385 = n4668 | ~n4669_1;
  assign n4671 = P1_DATAO_REG_24_ & ~n605;
  assign n4672 = BUF1_REG_24_ & n4550;
  assign n4673 = P2_DATAO_REG_24_ & n4552;
  assign n4674_1 = ~n4671 & ~n4672;
  assign n390 = n4673 | ~n4674_1;
  assign n4676 = P1_DATAO_REG_25_ & ~n605;
  assign n4677 = BUF1_REG_25_ & n4550;
  assign n4678 = P2_DATAO_REG_25_ & n4552;
  assign n4679_1 = ~n4676 & ~n4677;
  assign n395 = n4678 | ~n4679_1;
  assign n4681 = P1_DATAO_REG_26_ & ~n605;
  assign n4682 = BUF1_REG_26_ & n4550;
  assign n4683 = P2_DATAO_REG_26_ & n4552;
  assign n4684_1 = ~n4681 & ~n4682;
  assign n400 = n4683 | ~n4684_1;
  assign n4686 = P1_DATAO_REG_27_ & ~n605;
  assign n4687 = BUF1_REG_27_ & n4550;
  assign n4688 = P2_DATAO_REG_27_ & n4552;
  assign n4689_1 = ~n4686 & ~n4687;
  assign n405 = n4688 | ~n4689_1;
  assign n4691 = P1_DATAO_REG_28_ & ~n605;
  assign n4692 = BUF1_REG_28_ & n4550;
  assign n4693 = P2_DATAO_REG_28_ & n4552;
  assign n4694_1 = ~n4691 & ~n4692;
  assign n410 = n4693 | ~n4694_1;
  assign n4696 = P1_DATAO_REG_29_ & ~n605;
  assign n4697 = BUF1_REG_29_ & n4550;
  assign n4698 = P2_DATAO_REG_29_ & n4552;
  assign n4699_1 = ~n4696 & ~n4697;
  assign n415 = n4698 | ~n4699_1;
  assign n4701 = P1_DATAO_REG_30_ & ~n605;
  assign n4702 = BUF1_REG_30_ & n4550;
  assign n4703 = P2_DATAO_REG_30_ & n4552;
  assign n4704_1 = ~n4701 & ~n4702;
  assign n420 = n4703 | ~n4704_1;
  assign n4706 = P1_DATAO_REG_31_ & ~n605;
  assign n4707 = BUF1_REG_31_ & n4550;
  assign n4708 = P2_DATAO_REG_31_ & n4552;
  assign n4709_1 = ~n4706 & ~n4707;
  assign n425 = n4708 | ~n4709_1;
  assign n595 = P2_ADDRESS_REG_29_ | ~n4548;
  assign n4712 = P2_DATAO_REG_0_ & ~n595;
  assign n4713 = BUF2_REG_0_ & n595;
  assign n430 = n4712 | n4713;
  assign n4715 = P2_DATAO_REG_1_ & ~n595;
  assign n4716 = BUF2_REG_1_ & n595;
  assign n435 = n4715 | n4716;
  assign n4718 = P2_DATAO_REG_2_ & ~n595;
  assign n4719_1 = BUF2_REG_2_ & n595;
  assign n440 = n4718 | n4719_1;
  assign n4721 = P2_DATAO_REG_3_ & ~n595;
  assign n4722 = BUF2_REG_3_ & n595;
  assign n445 = n4721 | n4722;
  assign n4724_1 = P2_DATAO_REG_4_ & ~n595;
  assign n4725 = BUF2_REG_4_ & n595;
  assign n450 = n4724_1 | n4725;
  assign n4727 = P2_DATAO_REG_5_ & ~n595;
  assign n4728 = BUF2_REG_5_ & n595;
  assign n455 = n4727 | n4728;
  assign n4730 = P2_DATAO_REG_6_ & ~n595;
  assign n4731 = BUF2_REG_6_ & n595;
  assign n460 = n4730 | n4731;
  assign n4733 = P2_DATAO_REG_7_ & ~n595;
  assign n4734_1 = BUF2_REG_7_ & n595;
  assign n465 = n4733 | n4734_1;
  assign n4736 = P2_DATAO_REG_8_ & ~n595;
  assign n4737 = BUF2_REG_8_ & n595;
  assign n470 = n4736 | n4737;
  assign n4739_1 = P2_DATAO_REG_9_ & ~n595;
  assign n4740 = BUF2_REG_9_ & n595;
  assign n475 = n4739_1 | n4740;
  assign n4742 = P2_DATAO_REG_10_ & ~n595;
  assign n4743 = BUF2_REG_10_ & n595;
  assign n480 = n4742 | n4743;
  assign n4745 = P2_DATAO_REG_11_ & ~n595;
  assign n4746 = BUF2_REG_11_ & n595;
  assign n485 = n4745 | n4746;
  assign n4748 = P2_DATAO_REG_12_ & ~n595;
  assign n4749_1 = BUF2_REG_12_ & n595;
  assign n490 = n4748 | n4749_1;
  assign n4751 = P2_DATAO_REG_13_ & ~n595;
  assign n4752 = BUF2_REG_13_ & n595;
  assign n495 = n4751 | n4752;
  assign n4754_1 = P2_DATAO_REG_14_ & ~n595;
  assign n4755 = BUF2_REG_14_ & n595;
  assign n500 = n4754_1 | n4755;
  assign n4757 = P2_DATAO_REG_15_ & ~n595;
  assign n4758 = BUF2_REG_15_ & n595;
  assign n505 = n4757 | n4758;
  assign n4760 = P2_DATAO_REG_16_ & ~n595;
  assign n4761 = BUF2_REG_16_ & n595;
  assign n510 = n4760 | n4761;
  assign n4763 = P2_DATAO_REG_17_ & ~n595;
  assign n4764_1 = BUF2_REG_17_ & n595;
  assign n515 = n4763 | n4764_1;
  assign n4766 = P2_DATAO_REG_18_ & ~n595;
  assign n4767 = BUF2_REG_18_ & n595;
  assign n520 = n4766 | n4767;
  assign n4769_1 = P2_DATAO_REG_19_ & ~n595;
  assign n4770 = BUF2_REG_19_ & n595;
  assign n525 = n4769_1 | n4770;
  assign n4772 = P2_DATAO_REG_20_ & ~n595;
  assign n4773 = BUF2_REG_20_ & n595;
  assign n530 = n4772 | n4773;
  assign n4775 = P2_DATAO_REG_21_ & ~n595;
  assign n4776 = BUF2_REG_21_ & n595;
  assign n535 = n4775 | n4776;
  assign n4778 = P2_DATAO_REG_22_ & ~n595;
  assign n4779_1 = BUF2_REG_22_ & n595;
  assign n540 = n4778 | n4779_1;
  assign n4781 = P2_DATAO_REG_23_ & ~n595;
  assign n4782 = BUF2_REG_23_ & n595;
  assign n545 = n4781 | n4782;
  assign n4784_1 = P2_DATAO_REG_24_ & ~n595;
  assign n4785 = BUF2_REG_24_ & n595;
  assign n550 = n4784_1 | n4785;
  assign n4787 = P2_DATAO_REG_25_ & ~n595;
  assign n4788 = BUF2_REG_25_ & n595;
  assign n555 = n4787 | n4788;
  assign n4790 = P2_DATAO_REG_26_ & ~n595;
  assign n4791 = BUF2_REG_26_ & n595;
  assign n560 = n4790 | n4791;
  assign n4793 = P2_DATAO_REG_27_ & ~n595;
  assign n4794_1 = BUF2_REG_27_ & n595;
  assign n565 = n4793 | n4794_1;
  assign n4796 = P2_DATAO_REG_28_ & ~n595;
  assign n4797 = BUF2_REG_28_ & n595;
  assign n570 = n4796 | n4797;
  assign n4799_1 = P2_DATAO_REG_29_ & ~n595;
  assign n4800 = BUF2_REG_29_ & n595;
  assign n575 = n4799_1 | n4800;
  assign n4802 = P2_DATAO_REG_30_ & ~n595;
  assign n4803 = BUF2_REG_30_ & n595;
  assign n580 = n4802 | n4803;
  assign n4805 = P2_DATAO_REG_31_ & ~n595;
  assign n4806 = BUF2_REG_31_ & n595;
  assign n585 = n4805 | n4806;
  assign n590 = ~n605 | ~n4549_1;
  assign n4809_1 = ~P3_BE_N_REG_3_ & ~P3_BE_N_REG_2_;
  assign n4810 = ~P3_BE_N_REG_1_ & ~P3_BE_N_REG_0_;
  assign n4811 = ~P3_ADS_N_REG & n4810;
  assign n4812 = ~P3_D_C_N_REG & n4811;
  assign n4813 = ~P3_W_R_N_REG & n4812;
  assign n4814_1 = P3_M_IO_N_REG & n4809_1;
  assign n4815 = n4813 & n4814_1;
  assign n600 = ~n595 | ~n4815;
  assign n4817 = P3_STATE_REG_1_ & ~P3_STATE_REG_0_;
  assign n4818 = P3_BYTEENABLE_REG_3_ & n4817;
  assign n4819_1 = P3_BE_N_REG_3_ & ~n4817;
  assign n610 = n4818 | n4819_1;
  assign n4821 = P3_BYTEENABLE_REG_2_ & n4817;
  assign n4822 = P3_BE_N_REG_2_ & ~n4817;
  assign n615 = n4821 | n4822;
  assign n4824_1 = P3_BYTEENABLE_REG_1_ & n4817;
  assign n4825 = P3_BE_N_REG_1_ & ~n4817;
  assign n620 = n4824_1 | n4825;
  assign n4827 = P3_BYTEENABLE_REG_0_ & n4817;
  assign n4828 = P3_BE_N_REG_0_ & ~n4817;
  assign n625 = n4827 | n4828;
  assign n4830 = P3_STATE_REG_2_ & n4817;
  assign n4831 = P3_REIP_REG_30_ & n4830;
  assign n4832 = ~P3_STATE_REG_2_ & n4817;
  assign n4833 = P3_REIP_REG_31_ & n4832;
  assign n4834_1 = P3_ADDRESS_REG_29_ & ~n4817;
  assign n4835 = ~n4831 & ~n4833;
  assign n630 = n4834_1 | ~n4835;
  assign n4837 = P3_REIP_REG_29_ & n4830;
  assign n4838 = P3_REIP_REG_30_ & n4832;
  assign n4839_1 = P3_ADDRESS_REG_28_ & ~n4817;
  assign n4840 = ~n4837 & ~n4838;
  assign n635 = n4839_1 | ~n4840;
  assign n4842 = P3_REIP_REG_28_ & n4830;
  assign n4843 = P3_REIP_REG_29_ & n4832;
  assign n4844_1 = P3_ADDRESS_REG_27_ & ~n4817;
  assign n4845 = ~n4842 & ~n4843;
  assign n640 = n4844_1 | ~n4845;
  assign n4847 = P3_REIP_REG_27_ & n4830;
  assign n4848 = P3_REIP_REG_28_ & n4832;
  assign n4849_1 = P3_ADDRESS_REG_26_ & ~n4817;
  assign n4850 = ~n4847 & ~n4848;
  assign n645 = n4849_1 | ~n4850;
  assign n4852 = P3_REIP_REG_26_ & n4830;
  assign n4853 = P3_REIP_REG_27_ & n4832;
  assign n4854_1 = P3_ADDRESS_REG_25_ & ~n4817;
  assign n4855 = ~n4852 & ~n4853;
  assign n650 = n4854_1 | ~n4855;
  assign n4857 = P3_REIP_REG_25_ & n4830;
  assign n4858 = P3_REIP_REG_26_ & n4832;
  assign n4859_1 = P3_ADDRESS_REG_24_ & ~n4817;
  assign n4860 = ~n4857 & ~n4858;
  assign n655 = n4859_1 | ~n4860;
  assign n4862 = P3_REIP_REG_24_ & n4830;
  assign n4863 = P3_REIP_REG_25_ & n4832;
  assign n4864_1 = P3_ADDRESS_REG_23_ & ~n4817;
  assign n4865 = ~n4862 & ~n4863;
  assign n660 = n4864_1 | ~n4865;
  assign n4867 = P3_REIP_REG_23_ & n4830;
  assign n4868 = P3_REIP_REG_24_ & n4832;
  assign n4869_1 = P3_ADDRESS_REG_22_ & ~n4817;
  assign n4870 = ~n4867 & ~n4868;
  assign n665 = n4869_1 | ~n4870;
  assign n4872 = P3_REIP_REG_22_ & n4830;
  assign n4873 = P3_REIP_REG_23_ & n4832;
  assign n4874_1 = P3_ADDRESS_REG_21_ & ~n4817;
  assign n4875 = ~n4872 & ~n4873;
  assign n670 = n4874_1 | ~n4875;
  assign n4877 = P3_REIP_REG_21_ & n4830;
  assign n4878 = P3_REIP_REG_22_ & n4832;
  assign n4879_1 = P3_ADDRESS_REG_20_ & ~n4817;
  assign n4880 = ~n4877 & ~n4878;
  assign n675 = n4879_1 | ~n4880;
  assign n4882 = P3_REIP_REG_20_ & n4830;
  assign n4883 = P3_REIP_REG_21_ & n4832;
  assign n4884_1 = P3_ADDRESS_REG_19_ & ~n4817;
  assign n4885 = ~n4882 & ~n4883;
  assign n680 = n4884_1 | ~n4885;
  assign n4887 = P3_REIP_REG_19_ & n4830;
  assign n4888 = P3_REIP_REG_20_ & n4832;
  assign n4889_1 = P3_ADDRESS_REG_18_ & ~n4817;
  assign n4890 = ~n4887 & ~n4888;
  assign n685 = n4889_1 | ~n4890;
  assign n4892 = P3_REIP_REG_18_ & n4830;
  assign n4893 = P3_REIP_REG_19_ & n4832;
  assign n4894_1 = P3_ADDRESS_REG_17_ & ~n4817;
  assign n4895 = ~n4892 & ~n4893;
  assign n690 = n4894_1 | ~n4895;
  assign n4897 = P3_REIP_REG_17_ & n4830;
  assign n4898 = P3_REIP_REG_18_ & n4832;
  assign n4899_1 = P3_ADDRESS_REG_16_ & ~n4817;
  assign n4900 = ~n4897 & ~n4898;
  assign n695 = n4899_1 | ~n4900;
  assign n4902 = P3_REIP_REG_16_ & n4830;
  assign n4903 = P3_REIP_REG_17_ & n4832;
  assign n4904_1 = P3_ADDRESS_REG_15_ & ~n4817;
  assign n4905 = ~n4902 & ~n4903;
  assign n700 = n4904_1 | ~n4905;
  assign n4907 = P3_REIP_REG_15_ & n4830;
  assign n4908 = P3_REIP_REG_16_ & n4832;
  assign n4909_1 = P3_ADDRESS_REG_14_ & ~n4817;
  assign n4910 = ~n4907 & ~n4908;
  assign n705 = n4909_1 | ~n4910;
  assign n4912 = P3_REIP_REG_14_ & n4830;
  assign n4913 = P3_REIP_REG_15_ & n4832;
  assign n4914_1 = P3_ADDRESS_REG_13_ & ~n4817;
  assign n4915 = ~n4912 & ~n4913;
  assign n710 = n4914_1 | ~n4915;
  assign n4917 = P3_REIP_REG_13_ & n4830;
  assign n4918 = P3_REIP_REG_14_ & n4832;
  assign n4919_1 = P3_ADDRESS_REG_12_ & ~n4817;
  assign n4920 = ~n4917 & ~n4918;
  assign n715 = n4919_1 | ~n4920;
  assign n4922 = P3_REIP_REG_12_ & n4830;
  assign n4923 = P3_REIP_REG_13_ & n4832;
  assign n4924_1 = P3_ADDRESS_REG_11_ & ~n4817;
  assign n4925 = ~n4922 & ~n4923;
  assign n720 = n4924_1 | ~n4925;
  assign n4927 = P3_REIP_REG_11_ & n4830;
  assign n4928 = P3_REIP_REG_12_ & n4832;
  assign n4929_1 = P3_ADDRESS_REG_10_ & ~n4817;
  assign n4930 = ~n4927 & ~n4928;
  assign n725 = n4929_1 | ~n4930;
  assign n4932 = P3_REIP_REG_10_ & n4830;
  assign n4933 = P3_REIP_REG_11_ & n4832;
  assign n4934_1 = P3_ADDRESS_REG_9_ & ~n4817;
  assign n4935 = ~n4932 & ~n4933;
  assign n730 = n4934_1 | ~n4935;
  assign n4937 = P3_REIP_REG_9_ & n4830;
  assign n4938 = P3_REIP_REG_10_ & n4832;
  assign n4939_1 = P3_ADDRESS_REG_8_ & ~n4817;
  assign n4940 = ~n4937 & ~n4938;
  assign n735 = n4939_1 | ~n4940;
  assign n4942 = P3_REIP_REG_8_ & n4830;
  assign n4943 = P3_REIP_REG_9_ & n4832;
  assign n4944_1 = P3_ADDRESS_REG_7_ & ~n4817;
  assign n4945 = ~n4942 & ~n4943;
  assign n740 = n4944_1 | ~n4945;
  assign n4947 = P3_REIP_REG_7_ & n4830;
  assign n4948 = P3_REIP_REG_8_ & n4832;
  assign n4949_1 = P3_ADDRESS_REG_6_ & ~n4817;
  assign n4950 = ~n4947 & ~n4948;
  assign n745 = n4949_1 | ~n4950;
  assign n4952 = P3_REIP_REG_6_ & n4830;
  assign n4953 = P3_REIP_REG_7_ & n4832;
  assign n4954_1 = P3_ADDRESS_REG_5_ & ~n4817;
  assign n4955 = ~n4952 & ~n4953;
  assign n750 = n4954_1 | ~n4955;
  assign n4957 = P3_REIP_REG_5_ & n4830;
  assign n4958 = P3_REIP_REG_6_ & n4832;
  assign n4959_1 = P3_ADDRESS_REG_4_ & ~n4817;
  assign n4960 = ~n4957 & ~n4958;
  assign n755 = n4959_1 | ~n4960;
  assign n4962 = P3_REIP_REG_4_ & n4830;
  assign n4963 = P3_REIP_REG_5_ & n4832;
  assign n4964_1 = P3_ADDRESS_REG_3_ & ~n4817;
  assign n4965 = ~n4962 & ~n4963;
  assign n760 = n4964_1 | ~n4965;
  assign n4967 = P3_REIP_REG_3_ & n4830;
  assign n4968 = P3_REIP_REG_4_ & n4832;
  assign n4969_1 = P3_ADDRESS_REG_2_ & ~n4817;
  assign n4970 = ~n4967 & ~n4968;
  assign n765 = n4969_1 | ~n4970;
  assign n4972 = P3_REIP_REG_2_ & n4830;
  assign n4973 = P3_REIP_REG_3_ & n4832;
  assign n4974_1 = P3_ADDRESS_REG_1_ & ~n4817;
  assign n4975 = ~n4972 & ~n4973;
  assign n770 = n4974_1 | ~n4975;
  assign n4977 = P3_REIP_REG_1_ & n4830;
  assign n4978 = P3_REIP_REG_2_ & n4832;
  assign n4979_1 = P3_ADDRESS_REG_0_ & ~n4817;
  assign n4980 = ~n4977 & ~n4978;
  assign n775 = n4979_1 | ~n4980;
  assign n4982 = ~P3_STATE_REG_2_ & P3_STATE_REG_1_;
  assign n4983 = NA & n4982;
  assign n4984_1 = P3_STATE_REG_0_ & ~n4983;
  assign n4985 = ~HOLD & ~P3_REQUESTPENDING_REG;
  assign n4986 = READY2 & READY22_REG;
  assign n4987 = ~n4985 & n4986;
  assign n4988 = n4982 & n4987;
  assign n4989_1 = ~P3_STATE_REG_2_ & ~P3_STATE_REG_1_;
  assign n4990 = HOLD & ~P3_REQUESTPENDING_REG;
  assign n4991 = n4989_1 & n4990;
  assign n4992 = ~n4988 & ~n4991;
  assign n4993 = n4984_1 & ~n4992;
  assign n4994_1 = ~n4830 & ~n4993;
  assign n4995 = ~HOLD & P3_REQUESTPENDING_REG;
  assign n4996 = P3_STATE_REG_0_ & ~n4995;
  assign n4997 = ~n4985 & n4996;
  assign n4998 = ~NA & ~P3_STATE_REG_0_;
  assign n4999_1 = n4985 & ~n4986;
  assign n5000 = ~n4986 & n4995;
  assign n5001 = P3_STATE_REG_1_ & ~n4999_1;
  assign n5002 = ~n5000 & n5001;
  assign n5003 = ~n4997 & ~n4998;
  assign n5004_1 = ~n5002 & n5003;
  assign n5005 = P3_STATE_REG_2_ & ~n5004_1;
  assign n780 = ~n4994_1 | n5005;
  assign n5007 = P3_STATE_REG_2_ & ~n4996;
  assign n5008 = P3_STATE_REG_0_ & P3_REQUESTPENDING_REG;
  assign n5009_1 = ~P3_STATE_REG_2_ & n5008;
  assign n5010 = ~n5007 & ~n5009_1;
  assign n5011 = ~P3_STATE_REG_1_ & ~n5010;
  assign n5012 = HOLD & ~n4986;
  assign n5013 = P3_STATE_REG_0_ & ~n5012;
  assign n5014_1 = P3_STATE_REG_2_ & ~n5013;
  assign n5015 = ~n4999_1 & ~n5014_1;
  assign n5016 = P3_STATE_REG_1_ & n5015;
  assign n5017 = n4817 & n4986;
  assign n5018 = ~n4832 & ~n5017;
  assign n5019_1 = ~n5011 & ~n5016;
  assign n785 = ~n5018 | ~n5019_1;
  assign n5021 = P3_STATE_REG_1_ & ~n5000;
  assign n5022 = n5008 & ~n5021;
  assign n5023 = ~P3_STATE_REG_2_ & ~n5022;
  assign n5024_1 = P3_STATE_REG_2_ & n4996;
  assign n5025 = NA & ~P3_STATE_REG_0_;
  assign n5026 = P3_STATE_REG_2_ & ~n4995;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~P3_STATE_REG_1_ & ~n5027;
  assign n5029_1 = ~n5023 & ~n5024_1;
  assign n790 = n5028 | ~n5029_1;
  assign n5031 = ~BS16 & ~n4989_1;
  assign n5032 = P3_STATE_REG_0_ & n4982;
  assign n5033 = ~P3_STATE_REG_1_ & ~P3_STATE_REG_0_;
  assign n5034_1 = ~n5032 & ~n5033;
  assign n5035 = n5031 & ~n5034_1;
  assign n5036 = P3_DATAWIDTH_REG_0_ & n5034_1;
  assign n795 = n5035 | n5036;
  assign n5038 = P3_DATAWIDTH_REG_1_ & n5034_1;
  assign n5039_1 = ~n5031 & ~n5034_1;
  assign n800 = n5038 | n5039_1;
  assign n805 = P3_DATAWIDTH_REG_2_ & n5034_1;
  assign n810 = P3_DATAWIDTH_REG_3_ & n5034_1;
  assign n815 = P3_DATAWIDTH_REG_4_ & n5034_1;
  assign n820 = P3_DATAWIDTH_REG_5_ & n5034_1;
  assign n825 = P3_DATAWIDTH_REG_6_ & n5034_1;
  assign n830 = P3_DATAWIDTH_REG_7_ & n5034_1;
  assign n835 = P3_DATAWIDTH_REG_8_ & n5034_1;
  assign n840 = P3_DATAWIDTH_REG_9_ & n5034_1;
  assign n845 = P3_DATAWIDTH_REG_10_ & n5034_1;
  assign n850 = P3_DATAWIDTH_REG_11_ & n5034_1;
  assign n855 = P3_DATAWIDTH_REG_12_ & n5034_1;
  assign n860 = P3_DATAWIDTH_REG_13_ & n5034_1;
  assign n865 = P3_DATAWIDTH_REG_14_ & n5034_1;
  assign n870 = P3_DATAWIDTH_REG_15_ & n5034_1;
  assign n875 = P3_DATAWIDTH_REG_16_ & n5034_1;
  assign n880 = P3_DATAWIDTH_REG_17_ & n5034_1;
  assign n885 = P3_DATAWIDTH_REG_18_ & n5034_1;
  assign n890 = P3_DATAWIDTH_REG_19_ & n5034_1;
  assign n895 = P3_DATAWIDTH_REG_20_ & n5034_1;
  assign n900 = P3_DATAWIDTH_REG_21_ & n5034_1;
  assign n905 = P3_DATAWIDTH_REG_22_ & n5034_1;
  assign n910 = P3_DATAWIDTH_REG_23_ & n5034_1;
  assign n915 = P3_DATAWIDTH_REG_24_ & n5034_1;
  assign n920 = P3_DATAWIDTH_REG_25_ & n5034_1;
  assign n925 = P3_DATAWIDTH_REG_26_ & n5034_1;
  assign n930 = P3_DATAWIDTH_REG_27_ & n5034_1;
  assign n935 = P3_DATAWIDTH_REG_28_ & n5034_1;
  assign n940 = P3_DATAWIDTH_REG_29_ & n5034_1;
  assign n945 = P3_DATAWIDTH_REG_30_ & n5034_1;
  assign n950 = P3_DATAWIDTH_REG_31_ & n5034_1;
  assign n5071 = P3_STATE2_REG_2_ & P3_STATE2_REG_1_;
  assign n5072 = P3_STATE2_REG_1_ & n4986;
  assign n5073 = ~P3_STATE2_REG_0_ & ~n5072;
  assign n5074_1 = ~P3_STATEBS16_REG & ~n4986;
  assign n5075 = P3_STATE_REG_2_ & ~P3_STATE_REG_1_;
  assign n5076 = ~n4982 & ~n5075;
  assign n5077 = ~P3_STATE_REG_0_ & ~n5076;
  assign n5078 = n5074_1 & n5077;
  assign n5079_1 = P3_INSTQUEUERD_ADDR_REG_1_ & P3_INSTQUEUERD_ADDR_REG_0_;
  assign n5080 = ~P3_INSTQUEUERD_ADDR_REG_2_ & n5079_1;
  assign n5081 = P3_INSTQUEUERD_ADDR_REG_3_ & n5080;
  assign n5082 = P3_INSTQUEUE_REG_11__5_ & n5081;
  assign n5083 = P3_INSTQUEUERD_ADDR_REG_1_ & ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign n5084_1 = ~P3_INSTQUEUERD_ADDR_REG_2_ & n5083;
  assign n5085 = P3_INSTQUEUERD_ADDR_REG_3_ & n5084_1;
  assign n5086 = P3_INSTQUEUE_REG_10__5_ & n5085;
  assign n5087 = ~n5082 & ~n5086;
  assign n5088_1 = ~P3_INSTQUEUERD_ADDR_REG_1_ & P3_INSTQUEUERD_ADDR_REG_0_;
  assign n5089 = ~P3_INSTQUEUERD_ADDR_REG_2_ & n5088_1;
  assign n5090 = P3_INSTQUEUERD_ADDR_REG_3_ & n5089;
  assign n5091 = P3_INSTQUEUE_REG_9__5_ & n5090;
  assign n5092_1 = ~P3_INSTQUEUERD_ADDR_REG_1_ & ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign n5093 = ~P3_INSTQUEUERD_ADDR_REG_2_ & n5092_1;
  assign n5094 = P3_INSTQUEUERD_ADDR_REG_3_ & n5093;
  assign n5095 = P3_INSTQUEUE_REG_8__5_ & n5094;
  assign n5096_1 = ~n5091 & ~n5095;
  assign n5097 = P3_INSTQUEUERD_ADDR_REG_3_ & P3_INSTQUEUERD_ADDR_REG_2_;
  assign n5098 = n5079_1 & n5097;
  assign n5099 = P3_INSTQUEUE_REG_15__5_ & n5098;
  assign n5100_1 = n5083 & n5097;
  assign n5101 = P3_INSTQUEUE_REG_14__5_ & n5100_1;
  assign n5102 = n5088_1 & n5097;
  assign n5103 = P3_INSTQUEUE_REG_13__5_ & n5102;
  assign n5104_1 = n5092_1 & n5097;
  assign n5105 = P3_INSTQUEUE_REG_12__5_ & n5104_1;
  assign n5106 = ~n5099 & ~n5101;
  assign n5107 = ~n5103 & n5106;
  assign n5108_1 = ~n5105 & n5107;
  assign n5109 = ~P3_INSTQUEUERD_ADDR_REG_3_ & P3_INSTQUEUERD_ADDR_REG_2_;
  assign n5110 = n5079_1 & n5109;
  assign n5111 = P3_INSTQUEUE_REG_7__5_ & n5110;
  assign n5112_1 = n5083 & n5109;
  assign n5113 = P3_INSTQUEUE_REG_6__5_ & n5112_1;
  assign n5114 = n5088_1 & n5109;
  assign n5115 = P3_INSTQUEUE_REG_5__5_ & n5114;
  assign n5116_1 = n5092_1 & n5109;
  assign n5117 = P3_INSTQUEUE_REG_4__5_ & n5116_1;
  assign n5118 = ~n5111 & ~n5113;
  assign n5119 = ~n5115 & n5118;
  assign n5120_1 = ~n5117 & n5119;
  assign n5121 = ~P3_INSTQUEUERD_ADDR_REG_3_ & n5080;
  assign n5122 = P3_INSTQUEUE_REG_3__5_ & n5121;
  assign n5123 = ~P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign n5124_1 = n5083 & n5123;
  assign n5125 = P3_INSTQUEUE_REG_2__5_ & n5124_1;
  assign n5126 = n5088_1 & n5123;
  assign n5127 = P3_INSTQUEUE_REG_1__5_ & n5126;
  assign n5128_1 = ~P3_INSTQUEUERD_ADDR_REG_3_ & n5093;
  assign n5129 = P3_INSTQUEUE_REG_0__5_ & n5128_1;
  assign n5130 = ~n5122 & ~n5125;
  assign n5131 = ~n5127 & n5130;
  assign n5132_1 = ~n5129 & n5131;
  assign n5133 = n5087 & n5096_1;
  assign n5134 = n5108_1 & n5133;
  assign n5135 = n5120_1 & n5134;
  assign n5136_1 = n5132_1 & n5135;
  assign n5137 = P3_INSTQUEUE_REG_11__6_ & n5081;
  assign n5138 = P3_INSTQUEUE_REG_10__6_ & n5085;
  assign n5139 = ~n5137 & ~n5138;
  assign n5140_1 = P3_INSTQUEUE_REG_9__6_ & n5090;
  assign n5141 = P3_INSTQUEUE_REG_8__6_ & n5094;
  assign n5142 = ~n5140_1 & ~n5141;
  assign n5143 = P3_INSTQUEUE_REG_15__6_ & n5098;
  assign n5144_1 = P3_INSTQUEUE_REG_14__6_ & n5100_1;
  assign n5145 = P3_INSTQUEUE_REG_13__6_ & n5102;
  assign n5146 = P3_INSTQUEUE_REG_12__6_ & n5104_1;
  assign n5147 = ~n5143 & ~n5144_1;
  assign n5148_1 = ~n5145 & n5147;
  assign n5149 = ~n5146 & n5148_1;
  assign n5150 = P3_INSTQUEUE_REG_7__6_ & n5110;
  assign n5151 = P3_INSTQUEUE_REG_6__6_ & n5112_1;
  assign n5152_1 = P3_INSTQUEUE_REG_5__6_ & n5114;
  assign n5153 = P3_INSTQUEUE_REG_4__6_ & n5116_1;
  assign n5154 = ~n5150 & ~n5151;
  assign n5155 = ~n5152_1 & n5154;
  assign n5156_1 = ~n5153 & n5155;
  assign n5157 = P3_INSTQUEUE_REG_3__6_ & n5121;
  assign n5158 = P3_INSTQUEUE_REG_2__6_ & n5124_1;
  assign n5159 = P3_INSTQUEUE_REG_1__6_ & n5126;
  assign n5160_1 = P3_INSTQUEUE_REG_0__6_ & n5128_1;
  assign n5161 = ~n5157 & ~n5158;
  assign n5162 = ~n5159 & n5161;
  assign n5163 = ~n5160_1 & n5162;
  assign n5164_1 = n5139 & n5142;
  assign n5165 = n5149 & n5164_1;
  assign n5166 = n5156_1 & n5165;
  assign n5167 = n5163 & n5166;
  assign n5168_1 = n5136_1 & n5167;
  assign n5169 = P3_INSTQUEUE_REG_11__4_ & n5081;
  assign n5170 = P3_INSTQUEUE_REG_10__4_ & n5085;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172_1 = P3_INSTQUEUE_REG_9__4_ & n5090;
  assign n5173 = P3_INSTQUEUE_REG_8__4_ & n5094;
  assign n5174 = ~n5172_1 & ~n5173;
  assign n5175 = P3_INSTQUEUE_REG_15__4_ & n5098;
  assign n5176_1 = P3_INSTQUEUE_REG_14__4_ & n5100_1;
  assign n5177 = P3_INSTQUEUE_REG_13__4_ & n5102;
  assign n5178 = P3_INSTQUEUE_REG_12__4_ & n5104_1;
  assign n5179 = ~n5175 & ~n5176_1;
  assign n5180_1 = ~n5177 & n5179;
  assign n5181 = ~n5178 & n5180_1;
  assign n5182 = P3_INSTQUEUE_REG_7__4_ & n5110;
  assign n5183 = P3_INSTQUEUE_REG_6__4_ & n5112_1;
  assign n5184_1 = P3_INSTQUEUE_REG_5__4_ & n5114;
  assign n5185 = P3_INSTQUEUE_REG_4__4_ & n5116_1;
  assign n5186 = ~n5182 & ~n5183;
  assign n5187 = ~n5184_1 & n5186;
  assign n5188_1 = ~n5185 & n5187;
  assign n5189 = P3_INSTQUEUE_REG_3__4_ & n5121;
  assign n5190 = P3_INSTQUEUE_REG_2__4_ & n5124_1;
  assign n5191 = P3_INSTQUEUE_REG_1__4_ & n5126;
  assign n5192_1 = P3_INSTQUEUE_REG_0__4_ & n5128_1;
  assign n5193 = ~n5189 & ~n5190;
  assign n5194 = ~n5191 & n5193;
  assign n5195 = ~n5192_1 & n5194;
  assign n5196_1 = n5171 & n5174;
  assign n5197 = n5181 & n5196_1;
  assign n5198 = n5188_1 & n5197;
  assign n5199 = n5195 & n5198;
  assign n5200_1 = P3_INSTQUEUE_REG_11__7_ & n5081;
  assign n5201 = P3_INSTQUEUE_REG_10__7_ & n5085;
  assign n5202 = ~n5200_1 & ~n5201;
  assign n5203 = P3_INSTQUEUE_REG_9__7_ & n5090;
  assign n5204_1 = P3_INSTQUEUE_REG_8__7_ & n5094;
  assign n5205 = ~n5203 & ~n5204_1;
  assign n5206 = P3_INSTQUEUE_REG_15__7_ & n5098;
  assign n5207 = P3_INSTQUEUE_REG_14__7_ & n5100_1;
  assign n5208 = P3_INSTQUEUE_REG_13__7_ & n5102;
  assign n5209_1 = P3_INSTQUEUE_REG_12__7_ & n5104_1;
  assign n5210 = ~n5206 & ~n5207;
  assign n5211 = ~n5208 & n5210;
  assign n5212 = ~n5209_1 & n5211;
  assign n5213 = P3_INSTQUEUE_REG_7__7_ & n5110;
  assign n5214_1 = P3_INSTQUEUE_REG_6__7_ & n5112_1;
  assign n5215 = P3_INSTQUEUE_REG_5__7_ & n5114;
  assign n5216 = P3_INSTQUEUE_REG_4__7_ & n5116_1;
  assign n5217 = ~n5213 & ~n5214_1;
  assign n5218 = ~n5215 & n5217;
  assign n5219_1 = ~n5216 & n5218;
  assign n5220 = P3_INSTQUEUE_REG_3__7_ & n5121;
  assign n5221 = P3_INSTQUEUE_REG_2__7_ & n5124_1;
  assign n5222 = P3_INSTQUEUE_REG_1__7_ & n5126;
  assign n5223 = P3_INSTQUEUE_REG_0__7_ & n5128_1;
  assign n5224_1 = ~n5220 & ~n5221;
  assign n5225 = ~n5222 & n5224_1;
  assign n5226 = ~n5223 & n5225;
  assign n5227 = n5202 & n5205;
  assign n5228 = n5212 & n5227;
  assign n5229_1 = n5219_1 & n5228;
  assign n5230 = n5226 & n5229_1;
  assign n5231 = P3_INSTQUEUE_REG_11__3_ & n5081;
  assign n5232 = P3_INSTQUEUE_REG_10__3_ & n5085;
  assign n5233 = ~n5231 & ~n5232;
  assign n5234_1 = P3_INSTQUEUE_REG_9__3_ & n5090;
  assign n5235 = P3_INSTQUEUE_REG_8__3_ & n5094;
  assign n5236 = ~n5234_1 & ~n5235;
  assign n5237 = P3_INSTQUEUE_REG_15__3_ & n5098;
  assign n5238 = P3_INSTQUEUE_REG_14__3_ & n5100_1;
  assign n5239_1 = P3_INSTQUEUE_REG_13__3_ & n5102;
  assign n5240 = P3_INSTQUEUE_REG_12__3_ & n5104_1;
  assign n5241 = ~n5237 & ~n5238;
  assign n5242 = ~n5239_1 & n5241;
  assign n5243 = ~n5240 & n5242;
  assign n5244_1 = P3_INSTQUEUE_REG_7__3_ & n5110;
  assign n5245 = P3_INSTQUEUE_REG_6__3_ & n5112_1;
  assign n5246 = P3_INSTQUEUE_REG_5__3_ & n5114;
  assign n5247 = P3_INSTQUEUE_REG_4__3_ & n5116_1;
  assign n5248 = ~n5244_1 & ~n5245;
  assign n5249_1 = ~n5246 & n5248;
  assign n5250 = ~n5247 & n5249_1;
  assign n5251 = P3_INSTQUEUE_REG_3__3_ & n5121;
  assign n5252 = P3_INSTQUEUE_REG_2__3_ & n5124_1;
  assign n5253 = P3_INSTQUEUE_REG_1__3_ & n5126;
  assign n5254_1 = P3_INSTQUEUE_REG_0__3_ & n5128_1;
  assign n5255 = ~n5251 & ~n5252;
  assign n5256 = ~n5253 & n5255;
  assign n5257 = ~n5254_1 & n5256;
  assign n5258 = n5233 & n5236;
  assign n5259_1 = n5243 & n5258;
  assign n5260 = n5250 & n5259_1;
  assign n5261 = n5257 & n5260;
  assign n5262 = P3_INSTQUEUE_REG_11__2_ & n5081;
  assign n5263 = P3_INSTQUEUE_REG_10__2_ & n5085;
  assign n5264_1 = ~n5262 & ~n5263;
  assign n5265 = P3_INSTQUEUE_REG_9__2_ & n5090;
  assign n5266 = P3_INSTQUEUE_REG_8__2_ & n5094;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = P3_INSTQUEUE_REG_15__2_ & n5098;
  assign n5269_1 = P3_INSTQUEUE_REG_14__2_ & n5100_1;
  assign n5270 = P3_INSTQUEUE_REG_13__2_ & n5102;
  assign n5271 = P3_INSTQUEUE_REG_12__2_ & n5104_1;
  assign n5272 = ~n5268 & ~n5269_1;
  assign n5273 = ~n5270 & n5272;
  assign n5274_1 = ~n5271 & n5273;
  assign n5275 = P3_INSTQUEUE_REG_7__2_ & n5110;
  assign n5276 = P3_INSTQUEUE_REG_6__2_ & n5112_1;
  assign n5277 = P3_INSTQUEUE_REG_5__2_ & n5114;
  assign n5278 = P3_INSTQUEUE_REG_4__2_ & n5116_1;
  assign n5279_1 = ~n5275 & ~n5276;
  assign n5280 = ~n5277 & n5279_1;
  assign n5281 = ~n5278 & n5280;
  assign n5282 = P3_INSTQUEUE_REG_3__2_ & n5121;
  assign n5283 = P3_INSTQUEUE_REG_2__2_ & n5124_1;
  assign n5284_1 = P3_INSTQUEUE_REG_1__2_ & n5126;
  assign n5285 = P3_INSTQUEUE_REG_0__2_ & n5128_1;
  assign n5286 = ~n5282 & ~n5283;
  assign n5287 = ~n5284_1 & n5286;
  assign n5288 = ~n5285 & n5287;
  assign n5289_1 = n5264_1 & n5267;
  assign n5290 = n5274_1 & n5289_1;
  assign n5291 = n5281 & n5290;
  assign n5292 = n5288 & n5291;
  assign n5293 = ~n5230 & ~n5261;
  assign n5294_1 = n5292 & n5293;
  assign n5295 = n5168_1 & n5199;
  assign n5296 = n5294_1 & n5295;
  assign n5297 = P3_INSTQUEUE_REG_11__1_ & n5081;
  assign n5298 = P3_INSTQUEUE_REG_10__1_ & n5085;
  assign n5299_1 = ~n5297 & ~n5298;
  assign n5300 = P3_INSTQUEUE_REG_9__1_ & n5090;
  assign n5301 = P3_INSTQUEUE_REG_8__1_ & n5094;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = P3_INSTQUEUE_REG_15__1_ & n5098;
  assign n5304_1 = P3_INSTQUEUE_REG_14__1_ & n5100_1;
  assign n5305 = P3_INSTQUEUE_REG_13__1_ & n5102;
  assign n5306 = P3_INSTQUEUE_REG_12__1_ & n5104_1;
  assign n5307 = ~n5303 & ~n5304_1;
  assign n5308 = ~n5305 & n5307;
  assign n5309_1 = ~n5306 & n5308;
  assign n5310 = P3_INSTQUEUE_REG_7__1_ & n5110;
  assign n5311 = P3_INSTQUEUE_REG_6__1_ & n5112_1;
  assign n5312 = P3_INSTQUEUE_REG_5__1_ & n5114;
  assign n5313 = P3_INSTQUEUE_REG_4__1_ & n5116_1;
  assign n5314_1 = ~n5310 & ~n5311;
  assign n5315 = ~n5312 & n5314_1;
  assign n5316 = ~n5313 & n5315;
  assign n5317 = P3_INSTQUEUE_REG_3__1_ & n5121;
  assign n5318 = P3_INSTQUEUE_REG_2__1_ & n5124_1;
  assign n5319_1 = P3_INSTQUEUE_REG_1__1_ & n5126;
  assign n5320 = P3_INSTQUEUE_REG_0__1_ & n5128_1;
  assign n5321 = ~n5317 & ~n5318;
  assign n5322 = ~n5319_1 & n5321;
  assign n5323 = ~n5320 & n5322;
  assign n5324_1 = n5299_1 & n5302;
  assign n5325 = n5309_1 & n5324_1;
  assign n5326 = n5316 & n5325;
  assign n5327 = n5323 & n5326;
  assign n5328 = P3_INSTQUEUE_REG_11__0_ & n5081;
  assign n5329_1 = P3_INSTQUEUE_REG_10__0_ & n5085;
  assign n5330 = ~n5328 & ~n5329_1;
  assign n5331 = P3_INSTQUEUE_REG_9__0_ & n5090;
  assign n5332 = P3_INSTQUEUE_REG_8__0_ & n5094;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334_1 = P3_INSTQUEUE_REG_15__0_ & n5098;
  assign n5335 = P3_INSTQUEUE_REG_14__0_ & n5100_1;
  assign n5336 = P3_INSTQUEUE_REG_13__0_ & n5102;
  assign n5337 = P3_INSTQUEUE_REG_12__0_ & n5104_1;
  assign n5338 = ~n5334_1 & ~n5335;
  assign n5339_1 = ~n5336 & n5338;
  assign n5340 = ~n5337 & n5339_1;
  assign n5341 = P3_INSTQUEUE_REG_7__0_ & n5110;
  assign n5342 = P3_INSTQUEUE_REG_6__0_ & n5112_1;
  assign n5343 = P3_INSTQUEUE_REG_5__0_ & n5114;
  assign n5344_1 = P3_INSTQUEUE_REG_4__0_ & n5116_1;
  assign n5345 = ~n5341 & ~n5342;
  assign n5346 = ~n5343 & n5345;
  assign n5347 = ~n5344_1 & n5346;
  assign n5348 = P3_INSTQUEUE_REG_3__0_ & n5121;
  assign n5349_1 = P3_INSTQUEUE_REG_2__0_ & n5124_1;
  assign n5350 = P3_INSTQUEUE_REG_1__0_ & n5126;
  assign n5351 = P3_INSTQUEUE_REG_0__0_ & n5128_1;
  assign n5352 = ~n5348 & ~n5349_1;
  assign n5353 = ~n5350 & n5352;
  assign n5354_1 = ~n5351 & n5353;
  assign n5355 = n5330 & n5333;
  assign n5356 = n5340 & n5355;
  assign n5357 = n5347 & n5356;
  assign n5358 = n5354_1 & n5357;
  assign n5359_1 = n5327 & ~n5358;
  assign n5360 = n5296 & n5359_1;
  assign n5361 = n5078 & n5360;
  assign n5362 = ~P3_STATE2_REG_1_ & ~n5361;
  assign n5363 = ~n4986 & n5077;
  assign n5364_1 = ~n5292 & ~n5327;
  assign n5365 = n5363 & n5364_1;
  assign n5366 = ~n4986 & ~n5292;
  assign n5367 = n5327 & n5366;
  assign n5368 = ~n4986 & n5292;
  assign n5369_1 = n5327 & ~n5363;
  assign n5370 = n5368 & ~n5369_1;
  assign n5371 = ~n5365 & ~n5367;
  assign n5372 = ~n5370 & n5371;
  assign n5373 = P3_INSTQUEUERD_ADDR_REG_4_ & ~P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n5374_1 = ~P3_INSTQUEUERD_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n5375 = P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_3_;
  assign n5376 = ~P3_INSTQUEUERD_ADDR_REG_2_ & P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n5377 = P3_INSTQUEUERD_ADDR_REG_2_ & ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n5378 = P3_INSTQUEUERD_ADDR_REG_0_ & ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5379_1 = P3_INSTQUEUEWR_ADDR_REG_1_ & ~n5378;
  assign n5380 = ~P3_INSTQUEUEWR_ADDR_REG_1_ & n5378;
  assign n5381 = ~P3_INSTQUEUERD_ADDR_REG_1_ & ~n5380;
  assign n5382 = ~n5379_1 & ~n5381;
  assign n5383 = ~n5377 & ~n5382;
  assign n5384_1 = ~n5376 & ~n5383;
  assign n5385 = ~n5375 & ~n5384_1;
  assign n5386 = ~n5374_1 & ~n5385;
  assign n5387 = ~P3_INSTQUEUERD_ADDR_REG_4_ & P3_INSTQUEUEWR_ADDR_REG_4_;
  assign n5388 = n5386 & ~n5387;
  assign n5389_1 = ~n5373 & ~n5388;
  assign n5390 = ~n5373 & ~n5387;
  assign n5391 = ~n5386 & ~n5390;
  assign n5392 = n5386 & n5390;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394_1 = ~n5374_1 & ~n5375;
  assign n5395 = ~n5384_1 & ~n5394_1;
  assign n5396 = n5384_1 & n5394_1;
  assign n5397 = ~n5395 & ~n5396;
  assign n5398 = ~P3_INSTQUEUERD_ADDR_REG_1_ & P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n5399_1 = P3_INSTQUEUERD_ADDR_REG_1_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n5400 = ~n5398 & ~n5399_1;
  assign n5401 = ~n5378 & ~n5400;
  assign n5402 = n5378 & n5400;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404_1 = ~n5376 & ~n5377;
  assign n5405 = ~n5382 & ~n5404_1;
  assign n5406 = n5382 & n5404_1;
  assign n5407 = ~n5405 & ~n5406;
  assign n5408 = n5393 & n5397;
  assign n5409_1 = n5403 & n5408;
  assign n5410 = n5407 & n5409_1;
  assign n5411 = n5389_1 & ~n5410;
  assign n5412 = ~n5327 & ~n5411;
  assign n5413 = n5327 & ~n5411;
  assign n5414_1 = ~n5412 & ~n5413;
  assign n5415 = ~n5230 & n5261;
  assign n5416 = ~n5136_1 & ~n5167;
  assign n5417 = n5199 & n5416;
  assign n5418 = n5415 & n5417;
  assign n5419_1 = n5358 & n5418;
  assign n5420 = n5414_1 & n5419_1;
  assign n5421 = ~n5292 & ~n5420;
  assign n5422 = ~n5261 & ~n5358;
  assign n5423 = ~n5230 & n5422;
  assign n5424_1 = n5295 & n5423;
  assign n5425 = ~n5412 & n5424_1;
  assign n5426 = ~n5413 & n5425;
  assign n5427 = n5292 & ~n5426;
  assign n5428 = ~n5421 & ~n5427;
  assign n5429_1 = n5372 & n5428;
  assign n5430 = ~P3_FLUSH_REG & ~P3_MORE_REG;
  assign n5431 = n5429_1 & ~n5430;
  assign n5432 = ~n5327 & n5358;
  assign n5433 = ~n5292 & n5432;
  assign n5434_1 = n5418 & n5433;
  assign n5435 = ~n5411 & n5434_1;
  assign n5436 = n5327 & n5358;
  assign n5437 = ~n5292 & n5436;
  assign n5438 = n5418 & n5437;
  assign n5439_1 = ~n5411 & n5438;
  assign n5440 = n5360 & ~n5411;
  assign n5441 = ~n5327 & ~n5358;
  assign n5442 = n5296 & n5441;
  assign n5443 = ~n5411 & n5442;
  assign n5444_1 = ~n5435 & ~n5439_1;
  assign n5445 = ~n5440 & n5444_1;
  assign n5446 = ~n5443 & n5445;
  assign n5447 = ~n5136_1 & n5167;
  assign n5448 = ~n5199 & n5447;
  assign n5449_1 = n5294_1 & n5448;
  assign n5450 = n5441 & n5449_1;
  assign n5451 = ~P3_INSTQUEUERD_ADDR_REG_0_ & P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5452 = ~n5378 & ~n5451;
  assign n5453 = n5403 & n5452;
  assign n5454_1 = ~n5407 & ~n5453;
  assign n5455 = n5408 & ~n5454_1;
  assign n5456 = n5389_1 & ~n5455;
  assign n5457 = n5450 & ~n5456;
  assign n5458 = n5436 & n5449_1;
  assign n5459_1 = ~n5456 & n5458;
  assign n5460 = n5294_1 & n5417;
  assign n5461 = n5359_1 & n5460;
  assign n5462 = n5393 & ~n5454_1;
  assign n5463 = n5397 & n5462;
  assign n5464_1 = n5389_1 & ~n5463;
  assign n5465 = n5461 & ~n5464_1;
  assign n5466 = n5441 & n5460;
  assign n5467 = ~n5403 & ~n5452;
  assign n5468 = n5408 & ~n5467;
  assign n5469_1 = n5407 & n5468;
  assign n5470 = n5389_1 & ~n5469_1;
  assign n5471 = n5466 & ~n5470;
  assign n5472 = ~n5457 & ~n5459_1;
  assign n5473 = ~n5465 & n5472;
  assign n5474_1 = ~n5471 & n5473;
  assign n5475 = n5446 & n5474_1;
  assign n5476 = ~n5429_1 & ~n5475;
  assign n5477 = ~n5327 & ~n5470;
  assign n5478 = n5327 & ~n5464_1;
  assign n5479_1 = ~n5477 & ~n5478;
  assign n5480 = ~n5358 & n5460;
  assign n5481 = n5479_1 & n5480;
  assign n5482 = n5261 & n5292;
  assign n5483 = n5136_1 & ~n5167;
  assign n5484_1 = n5482 & n5483;
  assign n5485 = n5436 & n5484_1;
  assign n5486 = ~n5230 & n5485;
  assign n5487 = n5296 & ~n5358;
  assign n5488 = ~n5434_1 & ~n5486;
  assign n5489_1 = ~n5487 & n5488;
  assign n5490 = n5167 & n5261;
  assign n5491 = ~n5199 & n5292;
  assign n5492 = ~n5230 & n5436;
  assign n5493 = n5491 & n5492;
  assign n5494_1 = n5136_1 & ~n5292;
  assign n5495 = n5199 & n5230;
  assign n5496 = n5494_1 & n5495;
  assign n5497 = ~n5493 & ~n5496;
  assign n5498 = n5490 & ~n5497;
  assign n5499_1 = n5441 & n5495;
  assign n5500 = n5484_1 & n5499_1;
  assign n5501 = n5261 & ~n5292;
  assign n5502 = n5230 & n5432;
  assign n5503 = n5417 & n5501;
  assign n5504_1 = n5502 & n5503;
  assign n5505 = ~n5327 & n5460;
  assign n5506 = ~n5504_1 & ~n5505;
  assign n5507 = ~n5498 & ~n5500;
  assign n5508 = n5506 & n5507;
  assign n5509_1 = n5167 & ~n5230;
  assign n5510 = ~n5483 & ~n5509_1;
  assign n5511 = n5261 & n5510;
  assign n5512 = ~n5292 & ~n5511;
  assign n5513 = ~n5230 & ~n5483;
  assign n5514_1 = ~n5447 & n5513;
  assign n5515 = ~n5261 & n5514_1;
  assign n5516 = n5359_1 & ~n5515;
  assign n5517 = n5416 & n5436;
  assign n5518 = n5136_1 & n5230;
  assign n5519_1 = ~n5293 & ~n5518;
  assign n5520 = ~n5327 & n5519_1;
  assign n5521 = n5167 & n5199;
  assign n5522 = n5358 & n5521;
  assign n5523 = ~n5517 & ~n5520;
  assign n5524_1 = ~n5522 & n5523;
  assign n5525 = ~n5516 & n5524_1;
  assign n5526 = n5292 & ~n5525;
  assign n5527 = ~n5261 & ~n5521;
  assign n5528 = n5136_1 & n5527;
  assign n5529_1 = n5230 & n5327;
  assign n5530 = n5358 & ~n5529_1;
  assign n5531 = n5261 & ~n5530;
  assign n5532 = ~n5136_1 & n5531;
  assign n5533 = ~n5230 & ~n5416;
  assign n5534_1 = ~n5359_1 & n5533;
  assign n5535 = ~n5199 & ~n5534_1;
  assign n5536 = n5167 & ~n5327;
  assign n5537 = n5230 & n5536;
  assign n5538 = n5199 & ~n5327;
  assign n5539_1 = n5447 & n5538;
  assign n5540 = ~n5416 & n5432;
  assign n5541 = ~n5537 & ~n5539_1;
  assign n5542 = ~n5540 & n5541;
  assign n5543 = ~n5528 & ~n5532;
  assign n5544_1 = ~n5535 & n5543;
  assign n5545 = n5542 & n5544_1;
  assign n5546 = ~n5512 & ~n5526;
  assign n5547 = n5545 & n5546;
  assign n5548 = n5508 & n5547;
  assign n5549_1 = ~n5485 & n5548;
  assign n5550 = P3_INSTQUEUERD_ADDR_REG_0_ & ~n5549_1;
  assign n5551 = n5489_1 & ~n5550;
  assign n5552 = ~P3_INSTQUEUERD_ADDR_REG_2_ & ~n5551;
  assign n5553 = P3_INSTQUEUERD_ADDR_REG_1_ & n5552;
  assign n5554_1 = P3_INSTQUEUERD_ADDR_REG_2_ & ~n5489_1;
  assign n5555 = ~P3_INSTQUEUERD_ADDR_REG_1_ & n5554_1;
  assign n5556 = ~P3_INSTQUEUERD_ADDR_REG_2_ & P3_INSTQUEUERD_ADDR_REG_1_;
  assign n5557 = P3_INSTQUEUERD_ADDR_REG_2_ & ~P3_INSTQUEUERD_ADDR_REG_1_;
  assign n5558 = ~n5556 & ~n5557;
  assign n5559_1 = n5438 & ~n5558;
  assign n5560 = P3_INSTQUEUERD_ADDR_REG_2_ & ~n5079_1;
  assign n5561 = ~n5080 & ~n5560;
  assign n5562 = ~n5436 & ~n5441;
  assign n5563 = n5561 & ~n5562;
  assign n5564_1 = n5449_1 & n5563;
  assign n5565 = ~n5559_1 & ~n5564_1;
  assign n5566 = n5327 & n5490;
  assign n5567 = ~n5491 & ~n5496;
  assign n5568 = n5566 & ~n5567;
  assign n5569_1 = n5495 & ~n5562;
  assign n5570 = n5484_1 & n5569_1;
  assign n5571 = ~n5568 & ~n5570;
  assign n5572 = n5506 & n5571;
  assign n5573 = n5547 & n5572;
  assign n5574_1 = n5560 & ~n5573;
  assign n5575 = n5565 & ~n5574_1;
  assign n5576 = ~n5553 & ~n5555;
  assign n5577 = n5575 & n5576;
  assign n5578 = n5199 & n5358;
  assign n5579_1 = ~n5261 & ~n5432;
  assign n5580 = n5513 & ~n5578;
  assign n5581 = n5579_1 & n5580;
  assign n5582 = ~n5539_1 & n5581;
  assign n5583 = n5292 & ~n5582;
  assign n5584_1 = ~n5292 & ~n5419_1;
  assign n5585 = n5359_1 & ~n5514_1;
  assign n5586 = ~n5583 & ~n5584_1;
  assign n5587 = ~n5585 & n5586;
  assign n5588 = n5456 & n5458;
  assign n5589_1 = n5411 & n5438;
  assign n5590 = n5411 & n5442;
  assign n5591 = ~n5589_1 & ~n5590;
  assign n5592 = ~n4986 & ~n5591;
  assign n5593 = ~n5588 & ~n5592;
  assign n5594_1 = n5450 & n5456;
  assign n5595 = ~n5447 & n5491;
  assign n5596 = ~n5594_1 & ~n5595;
  assign n5597 = n5411 & n5434_1;
  assign n5598 = n5360 & n5411;
  assign n5599_1 = ~n5597 & ~n5598;
  assign n5600 = n5363 & ~n5599_1;
  assign n5601 = n5596 & ~n5600;
  assign n5602 = n5587 & n5593;
  assign n5603 = n5601 & n5602;
  assign n5604_1 = ~n5577 & ~n5603;
  assign n5605 = P3_INSTQUEUERD_ADDR_REG_2_ & n5603;
  assign n5606 = ~n5604_1 & ~n5605;
  assign n5607 = P3_INSTQUEUERD_ADDR_REG_1_ & n5109;
  assign n5608 = ~n5551 & n5607;
  assign n5609_1 = P3_INSTQUEUERD_ADDR_REG_2_ & n5079_1;
  assign n5610 = P3_INSTQUEUERD_ADDR_REG_3_ & ~n5609_1;
  assign n5611 = ~n5572 & n5610;
  assign n5612 = P3_INSTQUEUERD_ADDR_REG_2_ & P3_INSTQUEUERD_ADDR_REG_1_;
  assign n5613 = ~P3_INSTQUEUERD_ADDR_REG_3_ & n5612;
  assign n5614_1 = P3_INSTQUEUERD_ADDR_REG_3_ & ~n5612;
  assign n5615 = ~n5613 & ~n5614_1;
  assign n5616 = n5438 & ~n5615;
  assign n5617 = ~n5611 & ~n5616;
  assign n5618 = ~n5199 & n5486;
  assign n5619_1 = n5199 & n5486;
  assign n5620 = ~n5360 & ~n5442;
  assign n5621 = ~n5434_1 & n5620;
  assign n5622 = ~n5618 & ~n5619_1;
  assign n5623 = n5621 & n5622;
  assign n5624_1 = n5547 & n5623;
  assign n5625 = n5614_1 & ~n5624_1;
  assign n5626 = P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_INSTQUEUERD_ADDR_REG_0_;
  assign n5627 = ~n5547 & n5626;
  assign n5628 = ~n5079_1 & n5123;
  assign n5629_1 = ~P3_INSTQUEUERD_ADDR_REG_2_ & ~n5079_1;
  assign n5630 = P3_INSTQUEUERD_ADDR_REG_3_ & ~n5629_1;
  assign n5631 = ~n5628 & ~n5630;
  assign n5632 = ~n5562 & n5631;
  assign n5633 = n5449_1 & n5632;
  assign n5634_1 = ~n5627 & ~n5633;
  assign n5635 = n5617 & ~n5625;
  assign n5636 = n5634_1 & n5635;
  assign n5637 = ~n5608 & n5636;
  assign n5638 = ~n5603 & ~n5637;
  assign n5639_1 = P3_INSTQUEUERD_ADDR_REG_3_ & n5603;
  assign n5640 = ~n5638 & ~n5639_1;
  assign n5641 = ~n5606 & ~n5640;
  assign n5642 = P3_INSTQUEUERD_ADDR_REG_4_ & n5603;
  assign n5643 = P3_INSTQUEUERD_ADDR_REG_3_ & n5612;
  assign n5644_1 = ~P3_INSTQUEUERD_ADDR_REG_4_ & n5643;
  assign n5645 = P3_INSTQUEUERD_ADDR_REG_4_ & ~n5643;
  assign n5646 = ~n5644_1 & ~n5645;
  assign n5647 = n5438 & ~n5646;
  assign n5648 = ~n5603 & n5647;
  assign n5649_1 = ~n5642 & ~n5648;
  assign n5650 = ~n5641 & n5649_1;
  assign n5651 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & ~n5640;
  assign n5652 = ~P3_INSTQUEUEWR_ADDR_REG_4_ & ~n5649_1;
  assign n5653 = P3_INSTQUEUEWR_ADDR_REG_2_ & n5606;
  assign n5654_1 = P3_INSTQUEUEWR_ADDR_REG_3_ & n5640;
  assign n5655 = n5447 & n5493;
  assign n5656 = ~n5450 & ~n5655;
  assign n5657 = n5485 & n5495;
  assign n5658 = n5548 & ~n5657;
  assign n5659_1 = n5656 & n5658;
  assign n5660 = ~P3_INSTQUEUERD_ADDR_REG_0_ & ~n5659_1;
  assign n5661 = P3_INSTQUEUERD_ADDR_REG_0_ & ~n5489_1;
  assign n5662 = P3_INSTQUEUERD_ADDR_REG_0_ & n5438;
  assign n5663 = ~n5660 & ~n5661;
  assign n5664_1 = ~n5662 & n5663;
  assign n5665 = ~n5603 & ~n5664_1;
  assign n5666 = P3_INSTQUEUERD_ADDR_REG_0_ & n5603;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = P3_INSTQUEUEWR_ADDR_REG_0_ & n5667;
  assign n5669_1 = ~P3_INSTQUEUEWR_ADDR_REG_1_ & ~n5668;
  assign n5670 = ~P3_INSTQUEUEWR_ADDR_REG_2_ & ~n5606;
  assign n5671 = ~P3_INSTQUEUERD_ADDR_REG_1_ & ~n5551;
  assign n5672 = ~P3_INSTQUEUERD_ADDR_REG_1_ & n5438;
  assign n5673 = ~n5079_1 & ~n5092_1;
  assign n5674_1 = ~n5656 & n5673;
  assign n5675 = ~n5672 & ~n5674_1;
  assign n5676 = n5083 & ~n5658;
  assign n5677 = n5675 & ~n5676;
  assign n5678 = ~n5671 & n5677;
  assign n5679_1 = ~n5603 & ~n5678;
  assign n5680 = P3_INSTQUEUERD_ADDR_REG_1_ & n5603;
  assign n5681 = ~n5679_1 & ~n5680;
  assign n5682 = P3_INSTQUEUEWR_ADDR_REG_1_ & n5668;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684_1 = ~n5669_1 & ~n5670;
  assign n5685 = ~n5683 & n5684_1;
  assign n5686 = ~n5653 & ~n5654_1;
  assign n5687 = ~n5685 & n5686;
  assign n5688 = ~n5651 & ~n5652;
  assign n5689_1 = ~n5687 & n5688;
  assign n5690 = P3_INSTQUEUEWR_ADDR_REG_4_ & n5649_1;
  assign n5691 = ~n5689_1 & ~n5690;
  assign n5692 = ~n5431 & ~n5476;
  assign n5693 = ~n5481 & n5692;
  assign n5694_1 = n5650 & n5693;
  assign n5695 = ~n5691 & n5694_1;
  assign n5696 = n5362 & n5695;
  assign n5697 = P3_STATE2_REG_0_ & ~n5696;
  assign n5698 = ~n5073 & ~n5697;
  assign n5699_1 = P3_STATE2_REG_2_ & n5698;
  assign n5700 = P3_STATE2_REG_0_ & ~n5699_1;
  assign n5701 = n5071 & n5700;
  assign n5702 = P3_STATE2_REG_3_ & ~n5700;
  assign n955 = n5701 | n5702;
  assign n5704_1 = ~P3_STATE2_REG_2_ & ~n4986;
  assign n5705 = P3_STATE2_REG_0_ & ~n5704_1;
  assign n5706 = ~P3_STATE2_REG_0_ & ~P3_STATEBS16_REG;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = P3_STATE2_REG_1_ & n5707;
  assign n5709_1 = P3_STATE2_REG_2_ & ~P3_STATE2_REG_1_;
  assign n5710 = ~n5708 & ~n5709_1;
  assign n5711 = P3_STATE2_REG_2_ & ~n5700;
  assign n960 = ~n5710 | n5711;
  assign n5713 = P3_STATE2_REG_0_ & n5709_1;
  assign n5714_1 = ~n5699_1 & n5713;
  assign n5715 = ~P3_STATE2_REG_2_ & P3_STATE2_REG_0_;
  assign n5716 = n4986 & n5715;
  assign n5717 = ~n5699_1 & ~n5716;
  assign n5718 = P3_STATE2_REG_1_ & ~n5717;
  assign n5719_1 = ~P3_STATE2_REG_3_ & ~P3_STATE2_REG_1_;
  assign n5720 = ~n4986 & n5719_1;
  assign n5721 = n5700 & n5720;
  assign n5722 = P3_STATE2_REG_1_ & ~P3_STATE2_REG_0_;
  assign n5723 = ~P3_STATE2_REG_2_ & n5722;
  assign n5724_1 = ~P3_STATEBS16_REG & n5723;
  assign n5725 = ~n5714_1 & ~n5718;
  assign n5726 = ~n5721 & n5725;
  assign n965 = n5724_1 | ~n5726;
  assign n5728 = P3_STATE2_REG_3_ & ~P3_INSTQUEUERD_ADDR_REG_4_;
  assign n5729_1 = ~P3_STATE2_REG_2_ & ~P3_STATE2_REG_1_;
  assign n5730 = n5728 & n5729_1;
  assign n5731 = ~n5699_1 & ~n5730;
  assign n5732 = ~P3_STATE2_REG_0_ & n5731;
  assign n5733 = P3_INSTADDRPOINTER_REG_0_ & P3_INSTADDRPOINTER_REG_31_;
  assign n5734_1 = P3_INSTADDRPOINTER_REG_0_ & ~P3_INSTADDRPOINTER_REG_31_;
  assign n5735 = ~n5733 & ~n5734_1;
  assign n5736 = P3_FLUSH_REG & n5735;
  assign n5737 = P3_INSTQUEUERD_ADDR_REG_0_ & ~P3_FLUSH_REG;
  assign n5738 = ~n5736 & ~n5737;
  assign n5739_1 = P3_INSTADDRPOINTER_REG_0_ & ~P3_INSTADDRPOINTER_REG_1_;
  assign n5740 = ~P3_INSTADDRPOINTER_REG_0_ & P3_INSTADDRPOINTER_REG_1_;
  assign n5741 = ~n5739_1 & ~n5740;
  assign n5742 = P3_INSTADDRPOINTER_REG_31_ & ~n5741;
  assign n5743 = P3_INSTADDRPOINTER_REG_1_ & ~P3_INSTADDRPOINTER_REG_31_;
  assign n5744_1 = ~n5742 & ~n5743;
  assign n5745 = ~n5735 & n5744_1;
  assign n5746 = P3_FLUSH_REG & n5745;
  assign n5747 = P3_INSTQUEUERD_ADDR_REG_1_ & ~P3_FLUSH_REG;
  assign n5748 = ~n5746 & ~n5747;
  assign n5749_1 = n5738 & n5748;
  assign n5750 = P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_FLUSH_REG;
  assign n5751 = ~n5735 & ~n5744_1;
  assign n5752 = P3_FLUSH_REG & n5751;
  assign n5753 = P3_INSTQUEUERD_ADDR_REG_2_ & ~P3_FLUSH_REG;
  assign n5754_1 = ~n5752 & ~n5753;
  assign n5755 = ~n5749_1 & n5750;
  assign n5756 = ~n5754_1 & n5755;
  assign n5757 = P3_INSTQUEUERD_ADDR_REG_4_ & ~P3_FLUSH_REG;
  assign n5758 = ~n5756 & ~n5757;
  assign n5759_1 = n5071 & n5758;
  assign n5760 = ~n5699_1 & ~n5759_1;
  assign n5761 = P3_STATE2_REG_0_ & ~n5760;
  assign n5762 = P3_STATE2_REG_3_ & P3_STATE2_REG_0_;
  assign n5763 = n5729_1 & n5762;
  assign n5764_1 = ~n5716 & ~n5763;
  assign n5765 = ~n5695 & n5713;
  assign n5766 = n5764_1 & ~n5765;
  assign n5767 = ~n5732 & ~n5761;
  assign n970 = ~n5766 | ~n5767;
  assign n5769_1 = P3_INSTQUEUEWR_ADDR_REG_1_ & P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5770 = P3_INSTQUEUEWR_ADDR_REG_2_ & n5769_1;
  assign n5771 = P3_INSTQUEUEWR_ADDR_REG_3_ & n5770;
  assign n5772 = P3_STATE2_REG_3_ & ~n5771;
  assign n5773 = ~P3_STATE2_REG_2_ & P3_STATE2_REG_1_;
  assign n5774_1 = ~n5709_1 & ~n5773;
  assign n5775 = ~n5728 & n5774_1;
  assign n5776 = ~P3_STATE2_REG_0_ & ~n5775;
  assign n5777 = ~n5772 & n5776;
  assign n5778 = ~P3_INSTQUEUEWR_ADDR_REG_2_ & n5769_1;
  assign n5779_1 = P3_INSTQUEUEWR_ADDR_REG_2_ & ~n5769_1;
  assign n5780 = ~n5778 & ~n5779_1;
  assign n5781 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & n5770;
  assign n5782 = P3_INSTQUEUEWR_ADDR_REG_3_ & ~n5770;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784_1 = ~n5780 & ~n5783;
  assign n5785 = ~P3_INSTQUEUEWR_ADDR_REG_1_ & P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5786 = P3_INSTQUEUEWR_ADDR_REG_1_ & ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5787 = ~n5785 & ~n5786;
  assign n5788 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5787;
  assign n5789_1 = n5784_1 & n5788;
  assign n5790 = ~n5771 & ~n5789_1;
  assign n5791 = ~P3_STATE2_REG_3_ & ~P3_STATE2_REG_2_;
  assign n5792 = ~P3_STATEBS16_REG & n5791;
  assign n5793 = ~P3_STATE2_REG_2_ & ~n5792;
  assign n5794_1 = P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5787;
  assign n5795 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & n5787;
  assign n5796 = ~n5794_1 & ~n5795;
  assign n5797 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5796;
  assign n5798 = P3_INSTQUEUEWR_ADDR_REG_0_ & n5796;
  assign n5799_1 = ~n5797 & ~n5798;
  assign n5800 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5799_1;
  assign n5801 = ~n5780 & ~n5788;
  assign n5802 = n5780 & n5788;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804_1 = P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5796;
  assign n5805 = ~n5803 & ~n5804_1;
  assign n5806 = n5803 & n5804_1;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = ~n5780 & n5783;
  assign n5809_1 = n5788 & n5808;
  assign n5810 = ~n5780 & n5788;
  assign n5811 = ~n5783 & ~n5810;
  assign n5812 = ~n5809_1 & ~n5811;
  assign n5813 = n5803 & ~n5812;
  assign n5814_1 = ~n5804_1 & ~n5812;
  assign n5815 = ~n5813 & ~n5814_1;
  assign n5816 = ~n5803 & n5812;
  assign n5817 = n5804_1 & n5816;
  assign n5818 = n5815 & ~n5817;
  assign n5819_1 = ~n5807 & ~n5818;
  assign n5820 = n5800 & n5819_1;
  assign n5821 = ~n5803 & ~n5812;
  assign n5822 = n5804_1 & n5821;
  assign n5823 = ~n5820 & ~n5822;
  assign n5824_1 = n5793 & ~n5823;
  assign n5825 = n5790 & ~n5824_1;
  assign n5826 = n5777 & ~n5825;
  assign n5827 = P3_INSTQUEUE_REG_15__7_ & ~n5826;
  assign n5828 = P3_STATEBS16_REG & n5791;
  assign n5829_1 = n5776 & n5828;
  assign n5830 = BUF2_REG_23_ & n5829_1;
  assign n5831 = n5822 & n5830;
  assign n5832 = P3_STATE2_REG_3_ & n5776;
  assign n5833 = ~n5230 & n5832;
  assign n5834_1 = n5771 & n5833;
  assign n5835 = ~n5831 & ~n5834_1;
  assign n5836 = BUF2_REG_31_ & n5829_1;
  assign n5837 = n5820 & n5836;
  assign n5838 = n5835 & ~n5837;
  assign n5839_1 = n5823 & n5828;
  assign n5840 = n5793 & ~n5839_1;
  assign n5841 = ~n5790 & ~n5840;
  assign n5842 = BUF2_REG_7_ & n5776;
  assign n5843 = n5841 & n5842;
  assign n5844_1 = ~n5827 & n5838;
  assign n975 = n5843 | ~n5844_1;
  assign n5846 = P3_INSTQUEUE_REG_15__6_ & ~n5826;
  assign n5847 = BUF2_REG_22_ & n5829_1;
  assign n5848 = n5822 & n5847;
  assign n5849_1 = ~n5167 & n5832;
  assign n5850 = n5771 & n5849_1;
  assign n5851 = ~n5848 & ~n5850;
  assign n5852 = BUF2_REG_30_ & n5829_1;
  assign n5853 = n5820 & n5852;
  assign n5854_1 = n5851 & ~n5853;
  assign n5855 = BUF2_REG_6_ & n5776;
  assign n5856 = n5841 & n5855;
  assign n5857 = ~n5846 & n5854_1;
  assign n980 = n5856 | ~n5857;
  assign n5859_1 = P3_INSTQUEUE_REG_15__5_ & ~n5826;
  assign n5860 = BUF2_REG_21_ & n5829_1;
  assign n5861 = n5822 & n5860;
  assign n5862 = ~n5136_1 & n5832;
  assign n5863 = n5771 & n5862;
  assign n5864_1 = ~n5861 & ~n5863;
  assign n5865 = BUF2_REG_29_ & n5829_1;
  assign n5866 = n5820 & n5865;
  assign n5867 = n5864_1 & ~n5866;
  assign n5868 = BUF2_REG_5_ & n5776;
  assign n5869_1 = n5841 & n5868;
  assign n5870 = ~n5859_1 & n5867;
  assign n985 = n5869_1 | ~n5870;
  assign n5872 = P3_INSTQUEUE_REG_15__4_ & ~n5826;
  assign n5873 = BUF2_REG_20_ & n5829_1;
  assign n5874_1 = n5822 & n5873;
  assign n5875 = ~n5199 & n5832;
  assign n5876 = n5771 & n5875;
  assign n5877 = ~n5874_1 & ~n5876;
  assign n5878 = BUF2_REG_28_ & n5829_1;
  assign n5879_1 = n5820 & n5878;
  assign n5880 = n5877 & ~n5879_1;
  assign n5881 = BUF2_REG_4_ & n5776;
  assign n5882 = n5841 & n5881;
  assign n5883 = ~n5872 & n5880;
  assign n990 = n5882 | ~n5883;
  assign n5885 = P3_INSTQUEUE_REG_15__3_ & ~n5826;
  assign n5886 = BUF2_REG_19_ & n5829_1;
  assign n5887 = n5822 & n5886;
  assign n5888 = ~n5261 & n5832;
  assign n5889_1 = n5771 & n5888;
  assign n5890 = ~n5887 & ~n5889_1;
  assign n5891 = BUF2_REG_27_ & n5829_1;
  assign n5892 = n5820 & n5891;
  assign n5893 = n5890 & ~n5892;
  assign n5894_1 = BUF2_REG_3_ & n5776;
  assign n5895 = n5841 & n5894_1;
  assign n5896 = ~n5885 & n5893;
  assign n995 = n5895 | ~n5896;
  assign n5898 = P3_INSTQUEUE_REG_15__2_ & ~n5826;
  assign n5899_1 = BUF2_REG_18_ & n5829_1;
  assign n5900 = n5822 & n5899_1;
  assign n5901 = ~n5292 & n5832;
  assign n5902 = n5771 & n5901;
  assign n5903 = ~n5900 & ~n5902;
  assign n5904_1 = BUF2_REG_26_ & n5829_1;
  assign n5905 = n5820 & n5904_1;
  assign n5906 = n5903 & ~n5905;
  assign n5907 = BUF2_REG_2_ & n5776;
  assign n5908 = n5841 & n5907;
  assign n5909_1 = ~n5898 & n5906;
  assign n1000 = n5908 | ~n5909_1;
  assign n5911 = P3_INSTQUEUE_REG_15__1_ & ~n5826;
  assign n5912 = BUF2_REG_17_ & n5829_1;
  assign n5913 = n5822 & n5912;
  assign n5914_1 = ~n5327 & n5832;
  assign n5915 = n5771 & n5914_1;
  assign n5916 = ~n5913 & ~n5915;
  assign n5917 = BUF2_REG_25_ & n5829_1;
  assign n5918 = n5820 & n5917;
  assign n5919_1 = n5916 & ~n5918;
  assign n5920 = BUF2_REG_1_ & n5776;
  assign n5921 = n5841 & n5920;
  assign n5922 = ~n5911 & n5919_1;
  assign n1005 = n5921 | ~n5922;
  assign n5924_1 = P3_INSTQUEUE_REG_15__0_ & ~n5826;
  assign n5925 = BUF2_REG_16_ & n5829_1;
  assign n5926 = n5822 & n5925;
  assign n5927 = ~n5358 & n5832;
  assign n5928 = n5771 & n5927;
  assign n5929_1 = ~n5926 & ~n5928;
  assign n5930 = BUF2_REG_24_ & n5829_1;
  assign n5931 = n5820 & n5930;
  assign n5932 = n5929_1 & ~n5931;
  assign n5933 = BUF2_REG_0_ & n5776;
  assign n5934_1 = n5841 & n5933;
  assign n5935 = ~n5924_1 & n5932;
  assign n1010 = n5934_1 | ~n5935;
  assign n5937 = P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n5938 = P3_INSTQUEUEWR_ADDR_REG_2_ & ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n5939_1 = n5937 & n5938;
  assign n5940 = P3_STATE2_REG_3_ & ~n5939_1;
  assign n5941 = n5776 & ~n5940;
  assign n5942 = n5784_1 & n5794_1;
  assign n5943 = ~n5939_1 & ~n5942;
  assign n5944_1 = P3_INSTQUEUEWR_ADDR_REG_0_ & ~n5799_1;
  assign n5945 = n5819_1 & n5944_1;
  assign n5946 = n5797 & n5821;
  assign n5947 = ~n5945 & ~n5946;
  assign n5948 = n5793 & ~n5947;
  assign n5949_1 = n5943 & ~n5948;
  assign n5950 = n5941 & ~n5949_1;
  assign n5951 = P3_INSTQUEUE_REG_14__7_ & ~n5950;
  assign n5952 = n5830 & n5946;
  assign n5953 = n5833 & n5939_1;
  assign n5954_1 = ~n5952 & ~n5953;
  assign n5955 = n5836 & n5945;
  assign n5956 = n5954_1 & ~n5955;
  assign n5957 = n5828 & n5947;
  assign n5958 = n5793 & ~n5957;
  assign n5959_1 = ~n5943 & ~n5958;
  assign n5960 = n5842 & n5959_1;
  assign n5961 = ~n5951 & n5956;
  assign n1015 = n5960 | ~n5961;
  assign n5963 = P3_INSTQUEUE_REG_14__6_ & ~n5950;
  assign n5964_1 = n5847 & n5946;
  assign n5965 = n5849_1 & n5939_1;
  assign n5966 = ~n5964_1 & ~n5965;
  assign n5967 = n5852 & n5945;
  assign n5968 = n5966 & ~n5967;
  assign n5969_1 = n5855 & n5959_1;
  assign n5970 = ~n5963 & n5968;
  assign n1020 = n5969_1 | ~n5970;
  assign n5972 = P3_INSTQUEUE_REG_14__5_ & ~n5950;
  assign n5973 = n5860 & n5946;
  assign n5974_1 = n5862 & n5939_1;
  assign n5975 = ~n5973 & ~n5974_1;
  assign n5976 = n5865 & n5945;
  assign n5977 = n5975 & ~n5976;
  assign n5978 = n5868 & n5959_1;
  assign n5979_1 = ~n5972 & n5977;
  assign n1025 = n5978 | ~n5979_1;
  assign n5981 = P3_INSTQUEUE_REG_14__4_ & ~n5950;
  assign n5982 = n5873 & n5946;
  assign n5983 = n5875 & n5939_1;
  assign n5984_1 = ~n5982 & ~n5983;
  assign n5985 = n5878 & n5945;
  assign n5986 = n5984_1 & ~n5985;
  assign n5987 = n5881 & n5959_1;
  assign n5988 = ~n5981 & n5986;
  assign n1030 = n5987 | ~n5988;
  assign n5990 = P3_INSTQUEUE_REG_14__3_ & ~n5950;
  assign n5991 = n5886 & n5946;
  assign n5992 = n5888 & n5939_1;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994_1 = n5891 & n5945;
  assign n5995 = n5993 & ~n5994_1;
  assign n5996 = n5894_1 & n5959_1;
  assign n5997 = ~n5990 & n5995;
  assign n1035 = n5996 | ~n5997;
  assign n5999_1 = P3_INSTQUEUE_REG_14__2_ & ~n5950;
  assign n6000 = n5899_1 & n5946;
  assign n6001 = n5901 & n5939_1;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = n5904_1 & n5945;
  assign n6004_1 = n6002 & ~n6003;
  assign n6005 = n5907 & n5959_1;
  assign n6006 = ~n5999_1 & n6004_1;
  assign n1040 = n6005 | ~n6006;
  assign n6008 = P3_INSTQUEUE_REG_14__1_ & ~n5950;
  assign n6009_1 = n5912 & n5946;
  assign n6010 = n5914_1 & n5939_1;
  assign n6011 = ~n6009_1 & ~n6010;
  assign n6012 = n5917 & n5945;
  assign n6013 = n6011 & ~n6012;
  assign n6014_1 = n5920 & n5959_1;
  assign n6015 = ~n6008 & n6013;
  assign n1045 = n6014_1 | ~n6015;
  assign n6017 = P3_INSTQUEUE_REG_14__0_ & ~n5950;
  assign n6018 = n5925 & n5946;
  assign n6019_1 = n5927 & n5939_1;
  assign n6020 = ~n6018 & ~n6019_1;
  assign n6021 = n5930 & n5945;
  assign n6022 = n6020 & ~n6021;
  assign n6023 = n5933 & n5959_1;
  assign n6024_1 = ~n6017 & n6022;
  assign n1050 = n6023 | ~n6024_1;
  assign n6026 = P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n6027 = n5785 & n6026;
  assign n6028 = P3_STATE2_REG_3_ & ~n6027;
  assign n6029_1 = n5776 & ~n6028;
  assign n6030 = n5784_1 & n5795;
  assign n6031 = ~n6027 & ~n6030;
  assign n6032 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & n5799_1;
  assign n6033 = n5819_1 & n6032;
  assign n6034_1 = n5798 & n5821;
  assign n6035 = ~n6033 & ~n6034_1;
  assign n6036 = n5793 & ~n6035;
  assign n6037 = n6031 & ~n6036;
  assign n6038 = n6029_1 & ~n6037;
  assign n6039_1 = P3_INSTQUEUE_REG_13__7_ & ~n6038;
  assign n6040 = n5830 & n6034_1;
  assign n6041 = n5833 & n6027;
  assign n6042 = ~n6040 & ~n6041;
  assign n6043 = n5836 & n6033;
  assign n6044_1 = n6042 & ~n6043;
  assign n6045 = n5828 & n6035;
  assign n6046 = n5793 & ~n6045;
  assign n6047 = ~n6031 & ~n6046;
  assign n6048 = n5842 & n6047;
  assign n6049_1 = ~n6039_1 & n6044_1;
  assign n1055 = n6048 | ~n6049_1;
  assign n6051 = P3_INSTQUEUE_REG_13__6_ & ~n6038;
  assign n6052 = n5847 & n6034_1;
  assign n6053 = n5849_1 & n6027;
  assign n6054_1 = ~n6052 & ~n6053;
  assign n6055 = n5852 & n6033;
  assign n6056 = n6054_1 & ~n6055;
  assign n6057 = n5855 & n6047;
  assign n6058 = ~n6051 & n6056;
  assign n1060 = n6057 | ~n6058;
  assign n6060 = P3_INSTQUEUE_REG_13__5_ & ~n6038;
  assign n6061 = n5860 & n6034_1;
  assign n6062 = n5862 & n6027;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064_1 = n5865 & n6033;
  assign n6065 = n6063 & ~n6064_1;
  assign n6066 = n5868 & n6047;
  assign n6067 = ~n6060 & n6065;
  assign n1065 = n6066 | ~n6067;
  assign n6069_1 = P3_INSTQUEUE_REG_13__4_ & ~n6038;
  assign n6070 = n5873 & n6034_1;
  assign n6071 = n5875 & n6027;
  assign n6072 = ~n6070 & ~n6071;
  assign n6073 = n5878 & n6033;
  assign n6074_1 = n6072 & ~n6073;
  assign n6075 = n5881 & n6047;
  assign n6076 = ~n6069_1 & n6074_1;
  assign n1070 = n6075 | ~n6076;
  assign n6078 = P3_INSTQUEUE_REG_13__3_ & ~n6038;
  assign n6079_1 = n5886 & n6034_1;
  assign n6080 = n5888 & n6027;
  assign n6081 = ~n6079_1 & ~n6080;
  assign n6082 = n5891 & n6033;
  assign n6083 = n6081 & ~n6082;
  assign n6084_1 = n5894_1 & n6047;
  assign n6085 = ~n6078 & n6083;
  assign n1075 = n6084_1 | ~n6085;
  assign n6087 = P3_INSTQUEUE_REG_13__2_ & ~n6038;
  assign n6088 = n5899_1 & n6034_1;
  assign n6089_1 = n5901 & n6027;
  assign n6090 = ~n6088 & ~n6089_1;
  assign n6091 = n5904_1 & n6033;
  assign n6092 = n6090 & ~n6091;
  assign n6093 = n5907 & n6047;
  assign n6094_1 = ~n6087 & n6092;
  assign n1080 = n6093 | ~n6094_1;
  assign n6096 = P3_INSTQUEUE_REG_13__1_ & ~n6038;
  assign n6097 = n5912 & n6034_1;
  assign n6098 = n5914_1 & n6027;
  assign n6099_1 = ~n6097 & ~n6098;
  assign n6100 = n5917 & n6033;
  assign n6101 = n6099_1 & ~n6100;
  assign n6102 = n5920 & n6047;
  assign n6103 = ~n6096 & n6101;
  assign n1085 = n6102 | ~n6103;
  assign n6105 = P3_INSTQUEUE_REG_13__0_ & ~n6038;
  assign n6106 = n5925 & n6034_1;
  assign n6107 = n5927 & n6027;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109_1 = n5930 & n6033;
  assign n6110 = n6108 & ~n6109_1;
  assign n6111 = n5933 & n6047;
  assign n6112 = ~n6105 & n6110;
  assign n1090 = n6111 | ~n6112;
  assign n6114_1 = P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n6115 = n5938 & n6114_1;
  assign n6116 = P3_STATE2_REG_3_ & ~n6115;
  assign n6117 = n5776 & ~n6116;
  assign n6118 = P3_INSTQUEUEWR_ADDR_REG_0_ & n5799_1;
  assign n6119_1 = n5819_1 & n6118;
  assign n6120 = ~P3_INSTQUEUEWR_ADDR_REG_0_ & n5796;
  assign n6121 = n5821 & n6120;
  assign n6122 = ~n6119_1 & ~n6121;
  assign n6123 = n5793 & ~n6122;
  assign n6124_1 = n5784_1 & n5787;
  assign n6125 = ~n6123 & ~n6124_1;
  assign n6126 = n6117 & ~n6125;
  assign n6127 = P3_INSTQUEUE_REG_12__7_ & ~n6126;
  assign n6128 = n5830 & n6121;
  assign n6129_1 = n5833 & n6115;
  assign n6130 = ~n6128 & ~n6129_1;
  assign n6131 = n5836 & n6119_1;
  assign n6132 = n6130 & ~n6131;
  assign n6133 = n5828 & n6122;
  assign n6134_1 = n5793 & ~n6133;
  assign n6135 = n6124_1 & ~n6134_1;
  assign n6136 = n5842 & n6135;
  assign n6137 = ~n6127 & n6132;
  assign n1095 = n6136 | ~n6137;
  assign n6139_1 = P3_INSTQUEUE_REG_12__6_ & ~n6126;
  assign n6140 = n5847 & n6121;
  assign n6141 = n5849_1 & n6115;
  assign n6142 = ~n6140 & ~n6141;
  assign n6143 = n5852 & n6119_1;
  assign n6144_1 = n6142 & ~n6143;
  assign n6145 = n5855 & n6135;
  assign n6146 = ~n6139_1 & n6144_1;
  assign n1100 = n6145 | ~n6146;
  assign n6148 = P3_INSTQUEUE_REG_12__5_ & ~n6126;
  assign n6149_1 = n5860 & n6121;
  assign n6150 = n5862 & n6115;
  assign n6151 = ~n6149_1 & ~n6150;
  assign n6152 = n5865 & n6119_1;
  assign n6153 = n6151 & ~n6152;
  assign n6154_1 = n5868 & n6135;
  assign n6155 = ~n6148 & n6153;
  assign n1105 = n6154_1 | ~n6155;
  assign n6157 = P3_INSTQUEUE_REG_12__4_ & ~n6126;
  assign n6158 = n5873 & n6121;
  assign n6159_1 = n5875 & n6115;
  assign n6160 = ~n6158 & ~n6159_1;
  assign n6161 = n5878 & n6119_1;
  assign n6162 = n6160 & ~n6161;
  assign n6163 = n5881 & n6135;
  assign n6164_1 = ~n6157 & n6162;
  assign n1110 = n6163 | ~n6164_1;
  assign n6166 = P3_INSTQUEUE_REG_12__3_ & ~n6126;
  assign n6167 = n5886 & n6121;
  assign n6168 = n5888 & n6115;
  assign n6169_1 = ~n6167 & ~n6168;
  assign n6170 = n5891 & n6119_1;
  assign n6171 = n6169_1 & ~n6170;
  assign n6172 = n5894_1 & n6135;
  assign n6173 = ~n6166 & n6171;
  assign n1115 = n6172 | ~n6173;
  assign n6175 = P3_INSTQUEUE_REG_12__2_ & ~n6126;
  assign n6176 = n5899_1 & n6121;
  assign n6177 = n5901 & n6115;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179_1 = n5904_1 & n6119_1;
  assign n6180 = n6178 & ~n6179_1;
  assign n6181 = n5907 & n6135;
  assign n6182 = ~n6175 & n6180;
  assign n1120 = n6181 | ~n6182;
  assign n6184_1 = P3_INSTQUEUE_REG_12__1_ & ~n6126;
  assign n6185 = n5912 & n6121;
  assign n6186 = n5914_1 & n6115;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = n5917 & n6119_1;
  assign n6189_1 = n6187 & ~n6188;
  assign n6190 = n5920 & n6135;
  assign n6191 = ~n6184_1 & n6189_1;
  assign n1125 = n6190 | ~n6191;
  assign n6193 = P3_INSTQUEUE_REG_12__0_ & ~n6126;
  assign n6194_1 = n5925 & n6121;
  assign n6195 = n5927 & n6115;
  assign n6196 = ~n6194_1 & ~n6195;
  assign n6197 = n5930 & n6119_1;
  assign n6198 = n6196 & ~n6197;
  assign n6199_1 = n5933 & n6135;
  assign n6200 = ~n6193 & n6198;
  assign n1130 = n6199_1 | ~n6200;
  assign n6202 = P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n6203 = n5769_1 & n6202;
  assign n6204_1 = P3_STATE2_REG_3_ & ~n6203;
  assign n6205 = n5776 & ~n6204_1;
  assign n6206 = n5780 & ~n5783;
  assign n6207 = n5788 & n6206;
  assign n6208 = ~n6203 & ~n6207;
  assign n6209_1 = n5807 & ~n5818;
  assign n6210 = n5800 & n6209_1;
  assign n6211 = n5804_1 & n5813;
  assign n6212 = ~n6210 & ~n6211;
  assign n6213 = n5793 & ~n6212;
  assign n6214_1 = n6208 & ~n6213;
  assign n6215 = n6205 & ~n6214_1;
  assign n6216 = P3_INSTQUEUE_REG_11__7_ & ~n6215;
  assign n6217 = n5830 & n6211;
  assign n6218 = n5833 & n6203;
  assign n6219_1 = ~n6217 & ~n6218;
  assign n6220 = n5836 & n6210;
  assign n6221 = n6219_1 & ~n6220;
  assign n6222 = n5828 & n6212;
  assign n6223 = n5793 & ~n6222;
  assign n6224_1 = ~n6208 & ~n6223;
  assign n6225 = n5842 & n6224_1;
  assign n6226 = ~n6216 & n6221;
  assign n1135 = n6225 | ~n6226;
  assign n6228 = P3_INSTQUEUE_REG_11__6_ & ~n6215;
  assign n6229_1 = n5847 & n6211;
  assign n6230 = n5849_1 & n6203;
  assign n6231 = ~n6229_1 & ~n6230;
  assign n6232 = n5852 & n6210;
  assign n6233 = n6231 & ~n6232;
  assign n6234_1 = n5855 & n6224_1;
  assign n6235 = ~n6228 & n6233;
  assign n1140 = n6234_1 | ~n6235;
  assign n6237 = P3_INSTQUEUE_REG_11__5_ & ~n6215;
  assign n6238 = n5860 & n6211;
  assign n6239_1 = n5862 & n6203;
  assign n6240 = ~n6238 & ~n6239_1;
  assign n6241 = n5865 & n6210;
  assign n6242 = n6240 & ~n6241;
  assign n6243 = n5868 & n6224_1;
  assign n6244_1 = ~n6237 & n6242;
  assign n1145 = n6243 | ~n6244_1;
  assign n6246 = P3_INSTQUEUE_REG_11__4_ & ~n6215;
  assign n6247 = n5873 & n6211;
  assign n6248 = n5875 & n6203;
  assign n6249_1 = ~n6247 & ~n6248;
  assign n6250 = n5878 & n6210;
  assign n6251 = n6249_1 & ~n6250;
  assign n6252 = n5881 & n6224_1;
  assign n6253 = ~n6246 & n6251;
  assign n1150 = n6252 | ~n6253;
  assign n6255 = P3_INSTQUEUE_REG_11__3_ & ~n6215;
  assign n6256 = n5886 & n6211;
  assign n6257 = n5888 & n6203;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259_1 = n5891 & n6210;
  assign n6260 = n6258 & ~n6259_1;
  assign n6261 = n5894_1 & n6224_1;
  assign n6262 = ~n6255 & n6260;
  assign n1155 = n6261 | ~n6262;
  assign n6264_1 = P3_INSTQUEUE_REG_11__2_ & ~n6215;
  assign n6265 = n5899_1 & n6211;
  assign n6266 = n5901 & n6203;
  assign n6267 = ~n6265 & ~n6266;
  assign n6268 = n5904_1 & n6210;
  assign n6269_1 = n6267 & ~n6268;
  assign n6270 = n5907 & n6224_1;
  assign n6271 = ~n6264_1 & n6269_1;
  assign n1160 = n6270 | ~n6271;
  assign n6273 = P3_INSTQUEUE_REG_11__1_ & ~n6215;
  assign n6274_1 = n5912 & n6211;
  assign n6275 = n5914_1 & n6203;
  assign n6276 = ~n6274_1 & ~n6275;
  assign n6277 = n5917 & n6210;
  assign n6278 = n6276 & ~n6277;
  assign n6279_1 = n5920 & n6224_1;
  assign n6280 = ~n6273 & n6278;
  assign n1165 = n6279_1 | ~n6280;
  assign n6282 = P3_INSTQUEUE_REG_11__0_ & ~n6215;
  assign n6283 = n5925 & n6211;
  assign n6284_1 = n5927 & n6203;
  assign n6285 = ~n6283 & ~n6284_1;
  assign n6286 = n5930 & n6210;
  assign n6287 = n6285 & ~n6286;
  assign n6288 = n5933 & n6224_1;
  assign n6289_1 = ~n6282 & n6287;
  assign n1170 = n6288 | ~n6289_1;
  assign n6291 = ~P3_INSTQUEUEWR_ADDR_REG_2_ & ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n6292 = n5937 & n6291;
  assign n6293 = P3_STATE2_REG_3_ & ~n6292;
  assign n6294_1 = n5776 & ~n6293;
  assign n6295 = n5794_1 & n6206;
  assign n6296 = ~n6292 & ~n6295;
  assign n6297 = n5944_1 & n6209_1;
  assign n6298 = n5797 & n5813;
  assign n6299_1 = ~n6297 & ~n6298;
  assign n6300 = n5793 & ~n6299_1;
  assign n6301 = n6296 & ~n6300;
  assign n6302 = n6294_1 & ~n6301;
  assign n6303 = P3_INSTQUEUE_REG_10__7_ & ~n6302;
  assign n6304_1 = n5830 & n6298;
  assign n6305 = n5833 & n6292;
  assign n6306 = ~n6304_1 & ~n6305;
  assign n6307 = n5836 & n6297;
  assign n6308 = n6306 & ~n6307;
  assign n6309_1 = n5828 & n6299_1;
  assign n6310 = n5793 & ~n6309_1;
  assign n6311 = ~n6296 & ~n6310;
  assign n6312 = n5842 & n6311;
  assign n6313 = ~n6303 & n6308;
  assign n1175 = n6312 | ~n6313;
  assign n6315 = P3_INSTQUEUE_REG_10__6_ & ~n6302;
  assign n6316 = n5847 & n6298;
  assign n6317 = n5849_1 & n6292;
  assign n6318 = ~n6316 & ~n6317;
  assign n6319_1 = n5852 & n6297;
  assign n6320 = n6318 & ~n6319_1;
  assign n6321 = n5855 & n6311;
  assign n6322 = ~n6315 & n6320;
  assign n1180 = n6321 | ~n6322;
  assign n6324_1 = P3_INSTQUEUE_REG_10__5_ & ~n6302;
  assign n6325 = n5860 & n6298;
  assign n6326 = n5862 & n6292;
  assign n6327 = ~n6325 & ~n6326;
  assign n6328 = n5865 & n6297;
  assign n6329_1 = n6327 & ~n6328;
  assign n6330 = n5868 & n6311;
  assign n6331 = ~n6324_1 & n6329_1;
  assign n1185 = n6330 | ~n6331;
  assign n6333 = P3_INSTQUEUE_REG_10__4_ & ~n6302;
  assign n6334_1 = n5873 & n6298;
  assign n6335 = n5875 & n6292;
  assign n6336 = ~n6334_1 & ~n6335;
  assign n6337 = n5878 & n6297;
  assign n6338 = n6336 & ~n6337;
  assign n6339_1 = n5881 & n6311;
  assign n6340 = ~n6333 & n6338;
  assign n1190 = n6339_1 | ~n6340;
  assign n6342 = P3_INSTQUEUE_REG_10__3_ & ~n6302;
  assign n6343 = n5886 & n6298;
  assign n6344_1 = n5888 & n6292;
  assign n6345 = ~n6343 & ~n6344_1;
  assign n6346 = n5891 & n6297;
  assign n6347 = n6345 & ~n6346;
  assign n6348 = n5894_1 & n6311;
  assign n6349_1 = ~n6342 & n6347;
  assign n1195 = n6348 | ~n6349_1;
  assign n6351 = P3_INSTQUEUE_REG_10__2_ & ~n6302;
  assign n6352 = n5899_1 & n6298;
  assign n6353 = n5901 & n6292;
  assign n6354_1 = ~n6352 & ~n6353;
  assign n6355 = n5904_1 & n6297;
  assign n6356 = n6354_1 & ~n6355;
  assign n6357 = n5907 & n6311;
  assign n6358 = ~n6351 & n6356;
  assign n1200 = n6357 | ~n6358;
  assign n6360 = P3_INSTQUEUE_REG_10__1_ & ~n6302;
  assign n6361 = n5912 & n6298;
  assign n6362 = n5914_1 & n6292;
  assign n6363 = ~n6361 & ~n6362;
  assign n6364_1 = n5917 & n6297;
  assign n6365 = n6363 & ~n6364_1;
  assign n6366 = n5920 & n6311;
  assign n6367 = ~n6360 & n6365;
  assign n1205 = n6366 | ~n6367;
  assign n6369_1 = P3_INSTQUEUE_REG_10__0_ & ~n6302;
  assign n6370 = n5925 & n6298;
  assign n6371 = n5927 & n6292;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = n5930 & n6297;
  assign n6374_1 = n6372 & ~n6373;
  assign n6375 = n5933 & n6311;
  assign n6376 = ~n6369_1 & n6374_1;
  assign n1210 = n6375 | ~n6376;
  assign n6378 = n5785 & n6202;
  assign n6379_1 = P3_STATE2_REG_3_ & ~n6378;
  assign n6380 = n5776 & ~n6379_1;
  assign n6381 = n5795 & n6206;
  assign n6382 = ~n6378 & ~n6381;
  assign n6383 = n6032 & n6209_1;
  assign n6384_1 = n5798 & n5813;
  assign n6385 = ~n6383 & ~n6384_1;
  assign n6386 = n5793 & ~n6385;
  assign n6387 = n6382 & ~n6386;
  assign n6388 = n6380 & ~n6387;
  assign n6389_1 = P3_INSTQUEUE_REG_9__7_ & ~n6388;
  assign n6390 = n5830 & n6384_1;
  assign n6391 = n5833 & n6378;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = n5836 & n6383;
  assign n6394_1 = n6392 & ~n6393;
  assign n6395 = n5828 & n6385;
  assign n6396 = n5793 & ~n6395;
  assign n6397 = ~n6382 & ~n6396;
  assign n6398 = n5842 & n6397;
  assign n6399_1 = ~n6389_1 & n6394_1;
  assign n1215 = n6398 | ~n6399_1;
  assign n6401 = P3_INSTQUEUE_REG_9__6_ & ~n6388;
  assign n6402 = n5847 & n6384_1;
  assign n6403 = n5849_1 & n6378;
  assign n6404_1 = ~n6402 & ~n6403;
  assign n6405 = n5852 & n6383;
  assign n6406 = n6404_1 & ~n6405;
  assign n6407 = n5855 & n6397;
  assign n6408 = ~n6401 & n6406;
  assign n1220 = n6407 | ~n6408;
  assign n6410 = P3_INSTQUEUE_REG_9__5_ & ~n6388;
  assign n6411 = n5860 & n6384_1;
  assign n6412 = n5862 & n6378;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414_1 = n5865 & n6383;
  assign n6415 = n6413 & ~n6414_1;
  assign n6416 = n5868 & n6397;
  assign n6417 = ~n6410 & n6415;
  assign n1225 = n6416 | ~n6417;
  assign n6419_1 = P3_INSTQUEUE_REG_9__4_ & ~n6388;
  assign n6420 = n5873 & n6384_1;
  assign n6421 = n5875 & n6378;
  assign n6422 = ~n6420 & ~n6421;
  assign n6423 = n5878 & n6383;
  assign n6424_1 = n6422 & ~n6423;
  assign n6425 = n5881 & n6397;
  assign n6426 = ~n6419_1 & n6424_1;
  assign n1230 = n6425 | ~n6426;
  assign n6428 = P3_INSTQUEUE_REG_9__3_ & ~n6388;
  assign n6429_1 = n5886 & n6384_1;
  assign n6430 = n5888 & n6378;
  assign n6431 = ~n6429_1 & ~n6430;
  assign n6432 = n5891 & n6383;
  assign n6433 = n6431 & ~n6432;
  assign n6434_1 = n5894_1 & n6397;
  assign n6435 = ~n6428 & n6433;
  assign n1235 = n6434_1 | ~n6435;
  assign n6437 = P3_INSTQUEUE_REG_9__2_ & ~n6388;
  assign n6438 = n5899_1 & n6384_1;
  assign n6439_1 = n5901 & n6378;
  assign n6440 = ~n6438 & ~n6439_1;
  assign n6441 = n5904_1 & n6383;
  assign n6442 = n6440 & ~n6441;
  assign n6443 = n5907 & n6397;
  assign n6444_1 = ~n6437 & n6442;
  assign n1240 = n6443 | ~n6444_1;
  assign n6446 = P3_INSTQUEUE_REG_9__1_ & ~n6388;
  assign n6447 = n5912 & n6384_1;
  assign n6448 = n5914_1 & n6378;
  assign n6449_1 = ~n6447 & ~n6448;
  assign n6450 = n5917 & n6383;
  assign n6451 = n6449_1 & ~n6450;
  assign n6452 = n5920 & n6397;
  assign n6453 = ~n6446 & n6451;
  assign n1245 = n6452 | ~n6453;
  assign n6455 = P3_INSTQUEUE_REG_9__0_ & ~n6388;
  assign n6456 = n5925 & n6384_1;
  assign n6457 = n5927 & n6378;
  assign n6458 = ~n6456 & ~n6457;
  assign n6459_1 = n5930 & n6383;
  assign n6460 = n6458 & ~n6459_1;
  assign n6461 = n5933 & n6397;
  assign n6462 = ~n6455 & n6460;
  assign n1250 = n6461 | ~n6462;
  assign n6464_1 = n6114_1 & n6291;
  assign n6465 = P3_STATE2_REG_3_ & ~n6464_1;
  assign n6466 = n5776 & ~n6465;
  assign n6467 = n6118 & n6209_1;
  assign n6468 = n5813 & n6120;
  assign n6469_1 = ~n6467 & ~n6468;
  assign n6470 = n5793 & ~n6469_1;
  assign n6471 = n5787 & n6206;
  assign n6472 = ~n6470 & ~n6471;
  assign n6473 = n6466 & ~n6472;
  assign n6474_1 = P3_INSTQUEUE_REG_8__7_ & ~n6473;
  assign n6475 = n5830 & n6468;
  assign n6476 = n5833 & n6464_1;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = n5836 & n6467;
  assign n6479_1 = n6477 & ~n6478;
  assign n6480 = n5828 & n6469_1;
  assign n6481 = n5793 & ~n6480;
  assign n6482 = n6471 & ~n6481;
  assign n6483 = n5842 & n6482;
  assign n6484_1 = ~n6474_1 & n6479_1;
  assign n1255 = n6483 | ~n6484_1;
  assign n6486 = P3_INSTQUEUE_REG_8__6_ & ~n6473;
  assign n6487 = n5847 & n6468;
  assign n6488 = n5849_1 & n6464_1;
  assign n6489_1 = ~n6487 & ~n6488;
  assign n6490 = n5852 & n6467;
  assign n6491 = n6489_1 & ~n6490;
  assign n6492 = n5855 & n6482;
  assign n6493 = ~n6486 & n6491;
  assign n1260 = n6492 | ~n6493;
  assign n6495 = P3_INSTQUEUE_REG_8__5_ & ~n6473;
  assign n6496 = n5860 & n6468;
  assign n6497 = n5862 & n6464_1;
  assign n6498 = ~n6496 & ~n6497;
  assign n6499_1 = n5865 & n6467;
  assign n6500 = n6498 & ~n6499_1;
  assign n6501 = n5868 & n6482;
  assign n6502 = ~n6495 & n6500;
  assign n1265 = n6501 | ~n6502;
  assign n6504_1 = P3_INSTQUEUE_REG_8__4_ & ~n6473;
  assign n6505 = n5873 & n6468;
  assign n6506 = n5875 & n6464_1;
  assign n6507 = ~n6505 & ~n6506;
  assign n6508 = n5878 & n6467;
  assign n6509_1 = n6507 & ~n6508;
  assign n6510 = n5881 & n6482;
  assign n6511 = ~n6504_1 & n6509_1;
  assign n1270 = n6510 | ~n6511;
  assign n6513 = P3_INSTQUEUE_REG_8__3_ & ~n6473;
  assign n6514_1 = n5886 & n6468;
  assign n6515 = n5888 & n6464_1;
  assign n6516 = ~n6514_1 & ~n6515;
  assign n6517 = n5891 & n6467;
  assign n6518 = n6516 & ~n6517;
  assign n6519_1 = n5894_1 & n6482;
  assign n6520 = ~n6513 & n6518;
  assign n1275 = n6519_1 | ~n6520;
  assign n6522 = P3_INSTQUEUE_REG_8__2_ & ~n6473;
  assign n6523 = n5899_1 & n6468;
  assign n6524_1 = n5901 & n6464_1;
  assign n6525 = ~n6523 & ~n6524_1;
  assign n6526 = n5904_1 & n6467;
  assign n6527 = n6525 & ~n6526;
  assign n6528 = n5907 & n6482;
  assign n6529_1 = ~n6522 & n6527;
  assign n1280 = n6528 | ~n6529_1;
  assign n6531 = P3_INSTQUEUE_REG_8__1_ & ~n6473;
  assign n6532 = n5912 & n6468;
  assign n6533 = n5914_1 & n6464_1;
  assign n6534_1 = ~n6532 & ~n6533;
  assign n6535 = n5917 & n6467;
  assign n6536 = n6534_1 & ~n6535;
  assign n6537 = n5920 & n6482;
  assign n6538 = ~n6531 & n6536;
  assign n1285 = n6537 | ~n6538;
  assign n6540 = P3_INSTQUEUE_REG_8__0_ & ~n6473;
  assign n6541 = n5925 & n6468;
  assign n6542 = n5927 & n6464_1;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544_1 = n5930 & n6467;
  assign n6545 = n6543 & ~n6544_1;
  assign n6546 = n5933 & n6482;
  assign n6547 = ~n6540 & n6545;
  assign n1290 = n6546 | ~n6547;
  assign n6549_1 = P3_STATE2_REG_3_ & ~n5781;
  assign n6550 = n5776 & ~n6549_1;
  assign n6551 = ~n5781 & ~n5809_1;
  assign n6552 = ~n5807 & n5818;
  assign n6553 = n5800 & n6552;
  assign n6554_1 = ~n5817 & ~n6553;
  assign n6555 = n5793 & ~n6554_1;
  assign n6556 = n6551 & ~n6555;
  assign n6557 = n6550 & ~n6556;
  assign n6558 = P3_INSTQUEUE_REG_7__7_ & ~n6557;
  assign n6559_1 = n5817 & n5830;
  assign n6560 = n5781 & n5833;
  assign n6561 = ~n6559_1 & ~n6560;
  assign n6562 = n5836 & n6553;
  assign n6563 = n6561 & ~n6562;
  assign n6564_1 = n5828 & n6554_1;
  assign n6565 = n5793 & ~n6564_1;
  assign n6566 = ~n6551 & ~n6565;
  assign n6567 = n5842 & n6566;
  assign n6568 = ~n6558 & n6563;
  assign n1295 = n6567 | ~n6568;
  assign n6570 = P3_INSTQUEUE_REG_7__6_ & ~n6557;
  assign n6571 = n5817 & n5847;
  assign n6572 = n5781 & n5849_1;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574_1 = n5852 & n6553;
  assign n6575 = n6573 & ~n6574_1;
  assign n6576 = n5855 & n6566;
  assign n6577 = ~n6570 & n6575;
  assign n1300 = n6576 | ~n6577;
  assign n6579_1 = P3_INSTQUEUE_REG_7__5_ & ~n6557;
  assign n6580 = n5817 & n5860;
  assign n6581 = n5781 & n5862;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = n5865 & n6553;
  assign n6584_1 = n6582 & ~n6583;
  assign n6585 = n5868 & n6566;
  assign n6586 = ~n6579_1 & n6584_1;
  assign n1305 = n6585 | ~n6586;
  assign n6588 = P3_INSTQUEUE_REG_7__4_ & ~n6557;
  assign n6589_1 = n5817 & n5873;
  assign n6590 = n5781 & n5875;
  assign n6591 = ~n6589_1 & ~n6590;
  assign n6592 = n5878 & n6553;
  assign n6593 = n6591 & ~n6592;
  assign n6594_1 = n5881 & n6566;
  assign n6595 = ~n6588 & n6593;
  assign n1310 = n6594_1 | ~n6595;
  assign n6597 = P3_INSTQUEUE_REG_7__3_ & ~n6557;
  assign n6598 = n5817 & n5886;
  assign n6599_1 = n5781 & n5888;
  assign n6600 = ~n6598 & ~n6599_1;
  assign n6601 = n5891 & n6553;
  assign n6602 = n6600 & ~n6601;
  assign n6603 = n5894_1 & n6566;
  assign n6604_1 = ~n6597 & n6602;
  assign n1315 = n6603 | ~n6604_1;
  assign n6606 = P3_INSTQUEUE_REG_7__2_ & ~n6557;
  assign n6607 = n5817 & n5899_1;
  assign n6608 = n5781 & n5901;
  assign n6609_1 = ~n6607 & ~n6608;
  assign n6610 = n5904_1 & n6553;
  assign n6611 = n6609_1 & ~n6610;
  assign n6612 = n5907 & n6566;
  assign n6613 = ~n6606 & n6611;
  assign n1320 = n6612 | ~n6613;
  assign n6615 = P3_INSTQUEUE_REG_7__1_ & ~n6557;
  assign n6616 = n5817 & n5912;
  assign n6617 = n5781 & n5914_1;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619_1 = n5917 & n6553;
  assign n6620 = n6618 & ~n6619_1;
  assign n6621 = n5920 & n6566;
  assign n6622 = ~n6615 & n6620;
  assign n1325 = n6621 | ~n6622;
  assign n6624_1 = P3_INSTQUEUE_REG_7__0_ & ~n6557;
  assign n6625 = n5817 & n5925;
  assign n6626 = n5781 & n5927;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = n5930 & n6553;
  assign n6629_1 = n6627 & ~n6628;
  assign n6630 = n5933 & n6566;
  assign n6631 = ~n6624_1 & n6629_1;
  assign n1330 = n6630 | ~n6631;
  assign n6633 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n6634_1 = n5938 & n6633;
  assign n6635 = P3_STATE2_REG_3_ & ~n6634_1;
  assign n6636 = n5776 & ~n6635;
  assign n6637 = n5794_1 & n5808;
  assign n6638 = ~n6634_1 & ~n6637;
  assign n6639_1 = n5944_1 & n6552;
  assign n6640 = n5797 & n5816;
  assign n6641 = ~n6639_1 & ~n6640;
  assign n6642 = n5793 & ~n6641;
  assign n6643 = n6638 & ~n6642;
  assign n6644_1 = n6636 & ~n6643;
  assign n6645 = P3_INSTQUEUE_REG_6__7_ & ~n6644_1;
  assign n6646 = n5830 & n6640;
  assign n6647 = n5833 & n6634_1;
  assign n6648 = ~n6646 & ~n6647;
  assign n6649_1 = n5836 & n6639_1;
  assign n6650 = n6648 & ~n6649_1;
  assign n6651 = n5828 & n6641;
  assign n6652 = n5793 & ~n6651;
  assign n6653 = ~n6638 & ~n6652;
  assign n6654_1 = n5842 & n6653;
  assign n6655 = ~n6645 & n6650;
  assign n1335 = n6654_1 | ~n6655;
  assign n6657 = P3_INSTQUEUE_REG_6__6_ & ~n6644_1;
  assign n6658 = n5847 & n6640;
  assign n6659_1 = n5849_1 & n6634_1;
  assign n6660 = ~n6658 & ~n6659_1;
  assign n6661 = n5852 & n6639_1;
  assign n6662 = n6660 & ~n6661;
  assign n6663 = n5855 & n6653;
  assign n6664_1 = ~n6657 & n6662;
  assign n1340 = n6663 | ~n6664_1;
  assign n6666 = P3_INSTQUEUE_REG_6__5_ & ~n6644_1;
  assign n6667 = n5860 & n6640;
  assign n6668 = n5862 & n6634_1;
  assign n6669_1 = ~n6667 & ~n6668;
  assign n6670 = n5865 & n6639_1;
  assign n6671 = n6669_1 & ~n6670;
  assign n6672 = n5868 & n6653;
  assign n6673 = ~n6666 & n6671;
  assign n1345 = n6672 | ~n6673;
  assign n6675 = P3_INSTQUEUE_REG_6__4_ & ~n6644_1;
  assign n6676 = n5873 & n6640;
  assign n6677 = n5875 & n6634_1;
  assign n6678 = ~n6676 & ~n6677;
  assign n6679_1 = n5878 & n6639_1;
  assign n6680 = n6678 & ~n6679_1;
  assign n6681 = n5881 & n6653;
  assign n6682 = ~n6675 & n6680;
  assign n1350 = n6681 | ~n6682;
  assign n6684_1 = P3_INSTQUEUE_REG_6__3_ & ~n6644_1;
  assign n6685 = n5886 & n6640;
  assign n6686 = n5888 & n6634_1;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = n5891 & n6639_1;
  assign n6689_1 = n6687 & ~n6688;
  assign n6690 = n5894_1 & n6653;
  assign n6691 = ~n6684_1 & n6689_1;
  assign n1355 = n6690 | ~n6691;
  assign n6693 = P3_INSTQUEUE_REG_6__2_ & ~n6644_1;
  assign n6694_1 = n5899_1 & n6640;
  assign n6695 = n5901 & n6634_1;
  assign n6696 = ~n6694_1 & ~n6695;
  assign n6697 = n5904_1 & n6639_1;
  assign n6698 = n6696 & ~n6697;
  assign n6699_1 = n5907 & n6653;
  assign n6700 = ~n6693 & n6698;
  assign n1360 = n6699_1 | ~n6700;
  assign n6702 = P3_INSTQUEUE_REG_6__1_ & ~n6644_1;
  assign n6703 = n5912 & n6640;
  assign n6704_1 = n5914_1 & n6634_1;
  assign n6705 = ~n6703 & ~n6704_1;
  assign n6706 = n5917 & n6639_1;
  assign n6707 = n6705 & ~n6706;
  assign n6708 = n5920 & n6653;
  assign n6709_1 = ~n6702 & n6707;
  assign n1365 = n6708 | ~n6709_1;
  assign n6711 = P3_INSTQUEUE_REG_6__0_ & ~n6644_1;
  assign n6712 = n5925 & n6640;
  assign n6713 = n5927 & n6634_1;
  assign n6714_1 = ~n6712 & ~n6713;
  assign n6715 = n5930 & n6639_1;
  assign n6716 = n6714_1 & ~n6715;
  assign n6717 = n5933 & n6653;
  assign n6718 = ~n6711 & n6716;
  assign n1370 = n6717 | ~n6718;
  assign n6720 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n6721 = n5785 & n6720;
  assign n6722 = P3_STATE2_REG_3_ & ~n6721;
  assign n6723 = n5776 & ~n6722;
  assign n6724_1 = n5795 & n5808;
  assign n6725 = ~n6721 & ~n6724_1;
  assign n6726 = n6032 & n6552;
  assign n6727 = n5798 & n5816;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729_1 = n5793 & ~n6728;
  assign n6730 = n6725 & ~n6729_1;
  assign n6731 = n6723 & ~n6730;
  assign n6732 = P3_INSTQUEUE_REG_5__7_ & ~n6731;
  assign n6733 = n5830 & n6727;
  assign n6734_1 = n5833 & n6721;
  assign n6735 = ~n6733 & ~n6734_1;
  assign n6736 = n5836 & n6726;
  assign n6737 = n6735 & ~n6736;
  assign n6738 = n5828 & n6728;
  assign n6739_1 = n5793 & ~n6738;
  assign n6740 = ~n6725 & ~n6739_1;
  assign n6741 = n5842 & n6740;
  assign n6742 = ~n6732 & n6737;
  assign n1375 = n6741 | ~n6742;
  assign n6744_1 = P3_INSTQUEUE_REG_5__6_ & ~n6731;
  assign n6745 = n5847 & n6727;
  assign n6746 = n5849_1 & n6721;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = n5852 & n6726;
  assign n6749_1 = n6747 & ~n6748;
  assign n6750 = n5855 & n6740;
  assign n6751 = ~n6744_1 & n6749_1;
  assign n1380 = n6750 | ~n6751;
  assign n6753 = P3_INSTQUEUE_REG_5__5_ & ~n6731;
  assign n6754_1 = n5860 & n6727;
  assign n6755 = n5862 & n6721;
  assign n6756 = ~n6754_1 & ~n6755;
  assign n6757 = n5865 & n6726;
  assign n6758 = n6756 & ~n6757;
  assign n6759_1 = n5868 & n6740;
  assign n6760 = ~n6753 & n6758;
  assign n1385 = n6759_1 | ~n6760;
  assign n6762 = P3_INSTQUEUE_REG_5__4_ & ~n6731;
  assign n6763 = n5873 & n6727;
  assign n6764_1 = n5875 & n6721;
  assign n6765 = ~n6763 & ~n6764_1;
  assign n6766 = n5878 & n6726;
  assign n6767 = n6765 & ~n6766;
  assign n6768 = n5881 & n6740;
  assign n6769_1 = ~n6762 & n6767;
  assign n1390 = n6768 | ~n6769_1;
  assign n6771 = P3_INSTQUEUE_REG_5__3_ & ~n6731;
  assign n6772 = n5886 & n6727;
  assign n6773 = n5888 & n6721;
  assign n6774_1 = ~n6772 & ~n6773;
  assign n6775 = n5891 & n6726;
  assign n6776 = n6774_1 & ~n6775;
  assign n6777 = n5894_1 & n6740;
  assign n6778 = ~n6771 & n6776;
  assign n1395 = n6777 | ~n6778;
  assign n6780 = P3_INSTQUEUE_REG_5__2_ & ~n6731;
  assign n6781 = n5899_1 & n6727;
  assign n6782 = n5901 & n6721;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784_1 = n5904_1 & n6726;
  assign n6785 = n6783 & ~n6784_1;
  assign n6786 = n5907 & n6740;
  assign n6787 = ~n6780 & n6785;
  assign n1400 = n6786 | ~n6787;
  assign n6789_1 = P3_INSTQUEUE_REG_5__1_ & ~n6731;
  assign n6790 = n5912 & n6727;
  assign n6791 = n5914_1 & n6721;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = n5917 & n6726;
  assign n6794_1 = n6792 & ~n6793;
  assign n6795 = n5920 & n6740;
  assign n6796 = ~n6789_1 & n6794_1;
  assign n1405 = n6795 | ~n6796;
  assign n6798 = P3_INSTQUEUE_REG_5__0_ & ~n6731;
  assign n6799_1 = n5925 & n6727;
  assign n6800 = n5927 & n6721;
  assign n6801 = ~n6799_1 & ~n6800;
  assign n6802 = n5930 & n6726;
  assign n6803 = n6801 & ~n6802;
  assign n6804_1 = n5933 & n6740;
  assign n6805 = ~n6798 & n6803;
  assign n1410 = n6804_1 | ~n6805;
  assign n6807 = n5816 & n6120;
  assign n6808 = n5830 & n6807;
  assign n6809_1 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n6810 = n5938 & n6809_1;
  assign n6811 = n5833 & n6810;
  assign n6812 = n5793 & ~n5828;
  assign n6813 = n5787 & n5808;
  assign n6814_1 = ~n6812 & n6813;
  assign n6815 = n5842 & n6814_1;
  assign n6816 = ~n6808 & ~n6811;
  assign n6817 = ~n6815 & n6816;
  assign n6818 = n6118 & n6552;
  assign n6819_1 = n5836 & n6818;
  assign n6820 = n6817 & ~n6819_1;
  assign n6821 = P3_STATE2_REG_3_ & ~n6810;
  assign n6822 = n5776 & ~n6821;
  assign n6823 = ~n6807 & ~n6818;
  assign n6824_1 = n5793 & ~n6823;
  assign n6825 = ~n6813 & ~n6824_1;
  assign n6826 = n6822 & ~n6825;
  assign n6827 = P3_INSTQUEUE_REG_4__7_ & ~n6826;
  assign n1415 = ~n6820 | n6827;
  assign n6829_1 = n5847 & n6807;
  assign n6830 = n5849_1 & n6810;
  assign n6831 = n5855 & n6814_1;
  assign n6832 = ~n6829_1 & ~n6830;
  assign n6833 = ~n6831 & n6832;
  assign n6834_1 = n5852 & n6818;
  assign n6835 = n6833 & ~n6834_1;
  assign n6836 = P3_INSTQUEUE_REG_4__6_ & ~n6826;
  assign n1420 = ~n6835 | n6836;
  assign n6838 = n5860 & n6807;
  assign n6839_1 = n5862 & n6810;
  assign n6840 = n5868 & n6814_1;
  assign n6841 = ~n6838 & ~n6839_1;
  assign n6842 = ~n6840 & n6841;
  assign n6843 = n5865 & n6818;
  assign n6844_1 = n6842 & ~n6843;
  assign n6845 = P3_INSTQUEUE_REG_4__5_ & ~n6826;
  assign n1425 = ~n6844_1 | n6845;
  assign n6847 = n5873 & n6807;
  assign n6848 = n5875 & n6810;
  assign n6849_1 = n5881 & n6814_1;
  assign n6850 = ~n6847 & ~n6848;
  assign n6851 = ~n6849_1 & n6850;
  assign n6852 = n5878 & n6818;
  assign n6853 = n6851 & ~n6852;
  assign n6854_1 = P3_INSTQUEUE_REG_4__4_ & ~n6826;
  assign n1430 = ~n6853 | n6854_1;
  assign n6856 = n5886 & n6807;
  assign n6857 = n5888 & n6810;
  assign n6858 = n5894_1 & n6814_1;
  assign n6859_1 = ~n6856 & ~n6857;
  assign n6860 = ~n6858 & n6859_1;
  assign n6861 = n5891 & n6818;
  assign n6862 = n6860 & ~n6861;
  assign n6863 = P3_INSTQUEUE_REG_4__3_ & ~n6826;
  assign n1435 = ~n6862 | n6863;
  assign n6865 = n5899_1 & n6807;
  assign n6866 = n5901 & n6810;
  assign n6867 = n5907 & n6814_1;
  assign n6868 = ~n6865 & ~n6866;
  assign n6869_1 = ~n6867 & n6868;
  assign n6870 = n5904_1 & n6818;
  assign n6871 = n6869_1 & ~n6870;
  assign n6872 = P3_INSTQUEUE_REG_4__2_ & ~n6826;
  assign n1440 = ~n6871 | n6872;
  assign n6874_1 = n5912 & n6807;
  assign n6875 = n5914_1 & n6810;
  assign n6876 = n5920 & n6814_1;
  assign n6877 = ~n6874_1 & ~n6875;
  assign n6878 = ~n6876 & n6877;
  assign n6879_1 = n5917 & n6818;
  assign n6880 = n6878 & ~n6879_1;
  assign n6881 = P3_INSTQUEUE_REG_4__1_ & ~n6826;
  assign n1445 = ~n6880 | n6881;
  assign n6883 = n5925 & n6807;
  assign n6884_1 = n5927 & n6810;
  assign n6885 = n5933 & n6814_1;
  assign n6886 = ~n6883 & ~n6884_1;
  assign n6887 = ~n6885 & n6886;
  assign n6888 = n5930 & n6818;
  assign n6889_1 = n6887 & ~n6888;
  assign n6890 = P3_INSTQUEUE_REG_4__0_ & ~n6826;
  assign n1450 = ~n6889_1 | n6890;
  assign n6892 = n5803 & n5812;
  assign n6893 = n5804_1 & n6892;
  assign n6894_1 = n5830 & n6893;
  assign n6895 = ~P3_INSTQUEUEWR_ADDR_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n6896 = n5769_1 & n6895;
  assign n6897 = n5833 & n6896;
  assign n6898 = n5780 & n5783;
  assign n6899_1 = n5788 & n6898;
  assign n6900 = ~n6896 & ~n6899_1;
  assign n6901 = ~n6812 & ~n6900;
  assign n6902 = n5842 & n6901;
  assign n6903 = ~n6894_1 & ~n6897;
  assign n6904_1 = ~n6902 & n6903;
  assign n6905 = n5807 & n5818;
  assign n6906 = n5800 & n6905;
  assign n6907 = n5836 & n6906;
  assign n6908 = n6904_1 & ~n6907;
  assign n6909_1 = P3_STATE2_REG_3_ & ~n6896;
  assign n6910 = n5776 & ~n6909_1;
  assign n6911 = ~n6893 & ~n6906;
  assign n6912 = n5793 & ~n6911;
  assign n6913 = n6900 & ~n6912;
  assign n6914_1 = n6910 & ~n6913;
  assign n6915 = P3_INSTQUEUE_REG_3__7_ & ~n6914_1;
  assign n1455 = ~n6908 | n6915;
  assign n6917 = n5847 & n6893;
  assign n6918 = n5849_1 & n6896;
  assign n6919_1 = n5855 & n6901;
  assign n6920 = ~n6917 & ~n6918;
  assign n6921 = ~n6919_1 & n6920;
  assign n6922 = n5852 & n6906;
  assign n6923 = n6921 & ~n6922;
  assign n6924_1 = P3_INSTQUEUE_REG_3__6_ & ~n6914_1;
  assign n1460 = ~n6923 | n6924_1;
  assign n6926 = n5860 & n6893;
  assign n6927 = n5862 & n6896;
  assign n6928 = n5868 & n6901;
  assign n6929_1 = ~n6926 & ~n6927;
  assign n6930 = ~n6928 & n6929_1;
  assign n6931 = n5865 & n6906;
  assign n6932 = n6930 & ~n6931;
  assign n6933 = P3_INSTQUEUE_REG_3__5_ & ~n6914_1;
  assign n1465 = ~n6932 | n6933;
  assign n6935 = n5873 & n6893;
  assign n6936 = n5875 & n6896;
  assign n6937 = n5881 & n6901;
  assign n6938 = ~n6935 & ~n6936;
  assign n6939_1 = ~n6937 & n6938;
  assign n6940 = n5878 & n6906;
  assign n6941 = n6939_1 & ~n6940;
  assign n6942 = P3_INSTQUEUE_REG_3__4_ & ~n6914_1;
  assign n1470 = ~n6941 | n6942;
  assign n6944_1 = n5886 & n6893;
  assign n6945 = n5888 & n6896;
  assign n6946 = n5894_1 & n6901;
  assign n6947 = ~n6944_1 & ~n6945;
  assign n6948 = ~n6946 & n6947;
  assign n6949_1 = n5891 & n6906;
  assign n6950 = n6948 & ~n6949_1;
  assign n6951 = P3_INSTQUEUE_REG_3__3_ & ~n6914_1;
  assign n1475 = ~n6950 | n6951;
  assign n6953 = n5899_1 & n6893;
  assign n6954_1 = n5901 & n6896;
  assign n6955 = n5907 & n6901;
  assign n6956 = ~n6953 & ~n6954_1;
  assign n6957 = ~n6955 & n6956;
  assign n6958 = n5904_1 & n6906;
  assign n6959_1 = n6957 & ~n6958;
  assign n6960 = P3_INSTQUEUE_REG_3__2_ & ~n6914_1;
  assign n1480 = ~n6959_1 | n6960;
  assign n6962 = n5912 & n6893;
  assign n6963 = n5914_1 & n6896;
  assign n6964_1 = n5920 & n6901;
  assign n6965 = ~n6962 & ~n6963;
  assign n6966 = ~n6964_1 & n6965;
  assign n6967 = n5917 & n6906;
  assign n6968 = n6966 & ~n6967;
  assign n6969_1 = P3_INSTQUEUE_REG_3__1_ & ~n6914_1;
  assign n1485 = ~n6968 | n6969_1;
  assign n6971 = n5925 & n6893;
  assign n6972 = n5927 & n6896;
  assign n6973 = n5933 & n6901;
  assign n6974_1 = ~n6971 & ~n6972;
  assign n6975 = ~n6973 & n6974_1;
  assign n6976 = n5930 & n6906;
  assign n6977 = n6975 & ~n6976;
  assign n6978 = P3_INSTQUEUE_REG_3__0_ & ~n6914_1;
  assign n1490 = ~n6977 | n6978;
  assign n6980 = n5797 & n6892;
  assign n6981 = n5830 & n6980;
  assign n6982 = n6291 & n6633;
  assign n6983 = n5833 & n6982;
  assign n6984_1 = n5794_1 & n6898;
  assign n6985 = ~n6982 & ~n6984_1;
  assign n6986 = ~n6812 & ~n6985;
  assign n6987 = n5842 & n6986;
  assign n6988 = ~n6981 & ~n6983;
  assign n6989_1 = ~n6987 & n6988;
  assign n6990 = n5944_1 & n6905;
  assign n6991 = n5836 & n6990;
  assign n6992 = n6989_1 & ~n6991;
  assign n6993 = P3_STATE2_REG_3_ & ~n6982;
  assign n6994_1 = n5776 & ~n6993;
  assign n6995 = ~n6980 & ~n6990;
  assign n6996 = n5793 & ~n6995;
  assign n6997 = n6985 & ~n6996;
  assign n6998 = n6994_1 & ~n6997;
  assign n6999_1 = P3_INSTQUEUE_REG_2__7_ & ~n6998;
  assign n1495 = ~n6992 | n6999_1;
  assign n7001 = n5847 & n6980;
  assign n7002 = n5849_1 & n6982;
  assign n7003 = n5855 & n6986;
  assign n7004_1 = ~n7001 & ~n7002;
  assign n7005 = ~n7003 & n7004_1;
  assign n7006 = n5852 & n6990;
  assign n7007 = n7005 & ~n7006;
  assign n7008 = P3_INSTQUEUE_REG_2__6_ & ~n6998;
  assign n1500 = ~n7007 | n7008;
  assign n7010 = n5860 & n6980;
  assign n7011 = n5862 & n6982;
  assign n7012 = n5868 & n6986;
  assign n7013 = ~n7010 & ~n7011;
  assign n7014_1 = ~n7012 & n7013;
  assign n7015 = n5865 & n6990;
  assign n7016 = n7014_1 & ~n7015;
  assign n7017 = P3_INSTQUEUE_REG_2__5_ & ~n6998;
  assign n1505 = ~n7016 | n7017;
  assign n7019_1 = n5873 & n6980;
  assign n7020 = n5875 & n6982;
  assign n7021 = n5881 & n6986;
  assign n7022 = ~n7019_1 & ~n7020;
  assign n7023 = ~n7021 & n7022;
  assign n7024_1 = n5878 & n6990;
  assign n7025 = n7023 & ~n7024_1;
  assign n7026 = P3_INSTQUEUE_REG_2__4_ & ~n6998;
  assign n1510 = ~n7025 | n7026;
  assign n7028 = n5886 & n6980;
  assign n7029_1 = n5888 & n6982;
  assign n7030 = n5894_1 & n6986;
  assign n7031 = ~n7028 & ~n7029_1;
  assign n7032 = ~n7030 & n7031;
  assign n7033 = n5891 & n6990;
  assign n7034_1 = n7032 & ~n7033;
  assign n7035 = P3_INSTQUEUE_REG_2__3_ & ~n6998;
  assign n1515 = ~n7034_1 | n7035;
  assign n7037 = n5899_1 & n6980;
  assign n7038 = n5901 & n6982;
  assign n7039_1 = n5907 & n6986;
  assign n7040 = ~n7037 & ~n7038;
  assign n7041 = ~n7039_1 & n7040;
  assign n7042 = n5904_1 & n6990;
  assign n7043 = n7041 & ~n7042;
  assign n7044_1 = P3_INSTQUEUE_REG_2__2_ & ~n6998;
  assign n1520 = ~n7043 | n7044_1;
  assign n7046 = n5912 & n6980;
  assign n7047 = n5914_1 & n6982;
  assign n7048 = n5920 & n6986;
  assign n7049_1 = ~n7046 & ~n7047;
  assign n7050 = ~n7048 & n7049_1;
  assign n7051 = n5917 & n6990;
  assign n7052 = n7050 & ~n7051;
  assign n7053 = P3_INSTQUEUE_REG_2__1_ & ~n6998;
  assign n1525 = ~n7052 | n7053;
  assign n7055 = n5925 & n6980;
  assign n7056 = n5927 & n6982;
  assign n7057 = n5933 & n6986;
  assign n7058 = ~n7055 & ~n7056;
  assign n7059_1 = ~n7057 & n7058;
  assign n7060 = n5930 & n6990;
  assign n7061 = n7059_1 & ~n7060;
  assign n7062 = P3_INSTQUEUE_REG_2__0_ & ~n6998;
  assign n1530 = ~n7061 | n7062;
  assign n7064_1 = n5798 & n6892;
  assign n7065 = n5830 & n7064_1;
  assign n7066 = n5785 & n6895;
  assign n7067 = n5833 & n7066;
  assign n7068 = n5795 & n6898;
  assign n7069_1 = ~n7066 & ~n7068;
  assign n7070 = ~n6812 & ~n7069_1;
  assign n7071 = n5842 & n7070;
  assign n7072 = ~n7065 & ~n7067;
  assign n7073 = ~n7071 & n7072;
  assign n7074_1 = n6032 & n6905;
  assign n7075 = n5836 & n7074_1;
  assign n7076 = n7073 & ~n7075;
  assign n7077 = P3_STATE2_REG_3_ & ~n7066;
  assign n7078 = n5776 & ~n7077;
  assign n7079_1 = ~n7064_1 & ~n7074_1;
  assign n7080 = n5793 & ~n7079_1;
  assign n7081 = n7069_1 & ~n7080;
  assign n7082 = n7078 & ~n7081;
  assign n7083 = P3_INSTQUEUE_REG_1__7_ & ~n7082;
  assign n1535 = ~n7076 | n7083;
  assign n7085 = n5847 & n7064_1;
  assign n7086 = n5849_1 & n7066;
  assign n7087 = n5855 & n7070;
  assign n7088 = ~n7085 & ~n7086;
  assign n7089_1 = ~n7087 & n7088;
  assign n7090 = n5852 & n7074_1;
  assign n7091 = n7089_1 & ~n7090;
  assign n7092 = P3_INSTQUEUE_REG_1__6_ & ~n7082;
  assign n1540 = ~n7091 | n7092;
  assign n7094_1 = n5860 & n7064_1;
  assign n7095 = n5862 & n7066;
  assign n7096 = n5868 & n7070;
  assign n7097 = ~n7094_1 & ~n7095;
  assign n7098 = ~n7096 & n7097;
  assign n7099_1 = n5865 & n7074_1;
  assign n7100 = n7098 & ~n7099_1;
  assign n7101 = P3_INSTQUEUE_REG_1__5_ & ~n7082;
  assign n1545 = ~n7100 | n7101;
  assign n7103 = n5873 & n7064_1;
  assign n7104_1 = n5875 & n7066;
  assign n7105 = n5881 & n7070;
  assign n7106 = ~n7103 & ~n7104_1;
  assign n7107 = ~n7105 & n7106;
  assign n7108 = n5878 & n7074_1;
  assign n7109_1 = n7107 & ~n7108;
  assign n7110 = P3_INSTQUEUE_REG_1__4_ & ~n7082;
  assign n1550 = ~n7109_1 | n7110;
  assign n7112 = n5886 & n7064_1;
  assign n7113 = n5888 & n7066;
  assign n7114_1 = n5894_1 & n7070;
  assign n7115 = ~n7112 & ~n7113;
  assign n7116 = ~n7114_1 & n7115;
  assign n7117 = n5891 & n7074_1;
  assign n7118 = n7116 & ~n7117;
  assign n7119_1 = P3_INSTQUEUE_REG_1__3_ & ~n7082;
  assign n1555 = ~n7118 | n7119_1;
  assign n7121 = n5899_1 & n7064_1;
  assign n7122 = n5901 & n7066;
  assign n7123 = n5907 & n7070;
  assign n7124_1 = ~n7121 & ~n7122;
  assign n7125 = ~n7123 & n7124_1;
  assign n7126 = n5904_1 & n7074_1;
  assign n7127 = n7125 & ~n7126;
  assign n7128 = P3_INSTQUEUE_REG_1__2_ & ~n7082;
  assign n1560 = ~n7127 | n7128;
  assign n7130 = n5912 & n7064_1;
  assign n7131 = n5914_1 & n7066;
  assign n7132 = n5920 & n7070;
  assign n7133 = ~n7130 & ~n7131;
  assign n7134_1 = ~n7132 & n7133;
  assign n7135 = n5917 & n7074_1;
  assign n7136 = n7134_1 & ~n7135;
  assign n7137 = P3_INSTQUEUE_REG_1__1_ & ~n7082;
  assign n1565 = ~n7136 | n7137;
  assign n7139_1 = n5925 & n7064_1;
  assign n7140 = n5927 & n7066;
  assign n7141 = n5933 & n7070;
  assign n7142 = ~n7139_1 & ~n7140;
  assign n7143 = ~n7141 & n7142;
  assign n7144_1 = n5930 & n7074_1;
  assign n7145 = n7143 & ~n7144_1;
  assign n7146 = P3_INSTQUEUE_REG_1__0_ & ~n7082;
  assign n1570 = ~n7145 | n7146;
  assign n7148 = n6120 & n6892;
  assign n7149_1 = n5830 & n7148;
  assign n7150 = n6291 & n6809_1;
  assign n7151 = n5833 & n7150;
  assign n7152 = n5787 & n6898;
  assign n7153 = ~n6812 & n7152;
  assign n7154_1 = n5842 & n7153;
  assign n7155 = ~n7149_1 & ~n7151;
  assign n7156 = ~n7154_1 & n7155;
  assign n7157 = n6118 & n6905;
  assign n7158 = n5836 & n7157;
  assign n7159_1 = n7156 & ~n7158;
  assign n7160 = P3_STATE2_REG_3_ & ~n7150;
  assign n7161 = n5776 & ~n7160;
  assign n7162 = ~n7148 & ~n7157;
  assign n7163 = n5793 & ~n7162;
  assign n7164_1 = ~n7152 & ~n7163;
  assign n7165 = n7161 & ~n7164_1;
  assign n7166 = P3_INSTQUEUE_REG_0__7_ & ~n7165;
  assign n1575 = ~n7159_1 | n7166;
  assign n7168 = n5847 & n7148;
  assign n7169_1 = n5849_1 & n7150;
  assign n7170 = n5855 & n7153;
  assign n7171 = ~n7168 & ~n7169_1;
  assign n7172 = ~n7170 & n7171;
  assign n7173 = n5852 & n7157;
  assign n7174_1 = n7172 & ~n7173;
  assign n7175 = P3_INSTQUEUE_REG_0__6_ & ~n7165;
  assign n1580 = ~n7174_1 | n7175;
  assign n7177 = n5860 & n7148;
  assign n7178 = n5862 & n7150;
  assign n7179_1 = n5868 & n7153;
  assign n7180 = ~n7177 & ~n7178;
  assign n7181 = ~n7179_1 & n7180;
  assign n7182 = n5865 & n7157;
  assign n7183 = n7181 & ~n7182;
  assign n7184_1 = P3_INSTQUEUE_REG_0__5_ & ~n7165;
  assign n1585 = ~n7183 | n7184_1;
  assign n7186 = n5873 & n7148;
  assign n7187 = n5875 & n7150;
  assign n7188 = n5881 & n7153;
  assign n7189_1 = ~n7186 & ~n7187;
  assign n7190 = ~n7188 & n7189_1;
  assign n7191 = n5878 & n7157;
  assign n7192 = n7190 & ~n7191;
  assign n7193 = P3_INSTQUEUE_REG_0__4_ & ~n7165;
  assign n1590 = ~n7192 | n7193;
  assign n7195 = n5886 & n7148;
  assign n7196 = n5888 & n7150;
  assign n7197 = n5894_1 & n7153;
  assign n7198 = ~n7195 & ~n7196;
  assign n7199_1 = ~n7197 & n7198;
  assign n7200 = n5891 & n7157;
  assign n7201 = n7199_1 & ~n7200;
  assign n7202 = P3_INSTQUEUE_REG_0__3_ & ~n7165;
  assign n1595 = ~n7201 | n7202;
  assign n7204_1 = n5899_1 & n7148;
  assign n7205 = n5901 & n7150;
  assign n7206 = n5907 & n7153;
  assign n7207 = ~n7204_1 & ~n7205;
  assign n7208 = ~n7206 & n7207;
  assign n7209_1 = n5904_1 & n7157;
  assign n7210 = n7208 & ~n7209_1;
  assign n7211 = P3_INSTQUEUE_REG_0__2_ & ~n7165;
  assign n1600 = ~n7210 | n7211;
  assign n7213 = n5912 & n7148;
  assign n7214_1 = n5914_1 & n7150;
  assign n7215 = n5920 & n7153;
  assign n7216 = ~n7213 & ~n7214_1;
  assign n7217 = ~n7215 & n7216;
  assign n7218 = n5917 & n7157;
  assign n7219_1 = n7217 & ~n7218;
  assign n7220 = P3_INSTQUEUE_REG_0__1_ & ~n7165;
  assign n1605 = ~n7219_1 | n7220;
  assign n7222 = n5925 & n7148;
  assign n7223 = n5927 & n7150;
  assign n7224_1 = n5933 & n7153;
  assign n7225 = ~n7222 & ~n7223;
  assign n7226 = ~n7224_1 & n7225;
  assign n7227 = n5930 & n7157;
  assign n7228 = n7226 & ~n7227;
  assign n7229_1 = P3_INSTQUEUE_REG_0__0_ & ~n7165;
  assign n1610 = ~n7228 | n7229_1;
  assign n7231 = P3_STATE2_REG_3_ & ~P3_STATE2_REG_0_;
  assign n7232 = P3_STATE2_REG_0_ & P3_FLUSH_REG;
  assign n7233 = n5071 & n7232;
  assign n7234_1 = ~n7231 & ~n7233;
  assign n7235 = ~n5603 & n5713;
  assign n7236 = n7234_1 & ~n7235;
  assign n7237 = P3_INSTQUEUERD_ADDR_REG_4_ & n7236;
  assign n7238 = ~n5646 & n5719_1;
  assign n7239_1 = n5438 & n7238;
  assign n7240 = ~n7236 & n7239_1;
  assign n1615 = n7237 | n7240;
  assign n7242 = ~n5637 & n5719_1;
  assign n7243 = ~n5110 & ~n5610;
  assign n7244_1 = n5728 & ~n7243;
  assign n7245 = ~n7242 & ~n7244_1;
  assign n7246 = ~n7236 & ~n7245;
  assign n7247 = P3_INSTQUEUERD_ADDR_REG_3_ & n7236;
  assign n1620 = n7246 | n7247;
  assign n7249_1 = ~n5561 & n5728;
  assign n7250 = P3_STATE2_REG_1_ & ~n5735;
  assign n7251 = ~n5744_1 & n7250;
  assign n7252 = ~n7249_1 & ~n7251;
  assign n7253 = ~n5577 & n5719_1;
  assign n7254_1 = n7252 & ~n7253;
  assign n7255 = ~n7236 & ~n7254_1;
  assign n7256 = P3_INSTQUEUERD_ADDR_REG_2_ & n7236;
  assign n1625 = n7255 | n7256;
  assign n7258 = n5673 & n5728;
  assign n7259_1 = n5744_1 & n7250;
  assign n7260 = ~n7258 & ~n7259_1;
  assign n7261 = ~n5678 & n5719_1;
  assign n7262 = n7260 & ~n7261;
  assign n7263 = ~n7236 & ~n7262;
  assign n7264_1 = P3_INSTQUEUERD_ADDR_REG_1_ & n7236;
  assign n1630 = n7263 | n7264_1;
  assign n7266 = P3_STATE2_REG_1_ & n5735;
  assign n7267 = ~P3_INSTQUEUERD_ADDR_REG_0_ & n5728;
  assign n7268_1 = ~n7266 & ~n7267;
  assign n7269 = ~n5664_1 & n5719_1;
  assign n7270 = n7268_1 & ~n7269;
  assign n7271 = ~n7236 & ~n7270;
  assign n7272 = P3_INSTQUEUERD_ADDR_REG_0_ & n7236;
  assign n1635 = n7271 | n7272;
  assign n7274 = P3_STATE2_REG_0_ & n5071;
  assign n7275 = ~n5758 & n7274;
  assign n7276 = ~n5776 & ~n7233;
  assign n7277 = ~n7275 & n7276;
  assign n1640 = P3_INSTQUEUEWR_ADDR_REG_4_ & n7277;
  assign n7279 = P3_STATE2_REG_3_ & ~n5770;
  assign n7280 = ~n7277 & ~n7279;
  assign n7281 = P3_INSTQUEUEWR_ADDR_REG_3_ & ~n7280;
  assign n7282 = ~n5719_1 & ~n5792;
  assign n7283 = ~n5812 & ~n7282;
  assign n7284 = P3_STATE2_REG_3_ & n5781;
  assign n7285 = ~n7283 & ~n7284;
  assign n7286 = n5800 & ~n5807;
  assign n7287 = ~n5818 & ~n7286;
  assign n7288 = ~n6553 & ~n7287;
  assign n7289 = n5828 & ~n7288;
  assign n7290 = n7285 & ~n7289;
  assign n7291 = ~n7277 & ~n7290;
  assign n1645 = n7281 | n7291;
  assign n7293 = ~n5803 & ~n7282;
  assign n7294 = P3_STATE2_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_2_;
  assign n7295 = n5769_1 & n7294;
  assign n7296 = ~n7293 & ~n7295;
  assign n7297 = ~n5800 & ~n5807;
  assign n7298 = n5800 & n5807;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = n5828 & ~n7299;
  assign n7301 = n7296 & ~n7300;
  assign n7302 = ~n7277 & ~n7301;
  assign n7303 = P3_STATE2_REG_3_ & ~n5769_1;
  assign n7304 = ~n7277 & ~n7303;
  assign n7305 = P3_INSTQUEUEWR_ADDR_REG_2_ & ~n7304;
  assign n1650 = n7302 | n7305;
  assign n7307 = ~n5796 & ~n7282;
  assign n7308 = P3_STATE2_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_1_;
  assign n7309 = ~n5799_1 & n5828;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = P3_INSTQUEUEWR_ADDR_REG_0_ & ~n7310;
  assign n7312 = n5828 & n6032;
  assign n7313 = ~n7307 & ~n7311;
  assign n7314 = ~n7312 & n7313;
  assign n7315 = ~n7277 & ~n7314;
  assign n7316 = P3_STATE2_REG_3_ & ~P3_INSTQUEUEWR_ADDR_REG_0_;
  assign n7317 = ~n7277 & ~n7316;
  assign n7318 = P3_INSTQUEUEWR_ADDR_REG_1_ & ~n7317;
  assign n1655 = n7315 | n7318;
  assign n7320 = ~n5719_1 & ~n5791;
  assign n7321 = ~n7277 & n7320;
  assign n7322 = P3_INSTQUEUEWR_ADDR_REG_0_ & ~n7321;
  assign n7323 = ~n5759_1 & ~n7316;
  assign n7324 = ~n7277 & ~n7323;
  assign n1660 = n7322 | n7324;
  assign n7326 = ~P3_STATE2_REG_1_ & n5791;
  assign n7327 = ~P3_STATE2_REG_0_ & n7326;
  assign n7328 = n5367 & n5411;
  assign n7329 = ~n5199 & ~n5358;
  assign n7330 = n5456 & n7329;
  assign n7331 = n5365 & n5411;
  assign n7332 = ~n5595 & ~n7330;
  assign n7333 = ~n7331 & n7332;
  assign n7334 = n5416 & n5464_1;
  assign n7335 = n5168_1 & n5363;
  assign n7336 = n5411 & n7335;
  assign n7337 = ~n7334 & ~n7336;
  assign n7338 = n5327 & ~n7337;
  assign n7339 = ~n5167 & n5470;
  assign n7340 = ~n4986 & n5136_1;
  assign n7341 = n5411 & n7340;
  assign n7342 = ~n7339 & ~n7341;
  assign n7343 = ~n5327 & ~n7342;
  assign n7344 = n5358 & n5456;
  assign n7345 = ~n7338 & ~n7343;
  assign n7346 = ~n7344 & n7345;
  assign n7347 = n5292 & ~n7346;
  assign n7348 = n5587 & ~n7328;
  assign n7349 = n7333 & n7348;
  assign n7350 = ~n7347 & n7349;
  assign n7351 = n5713 & ~n7350;
  assign n7352 = ~n7327 & ~n7351;
  assign n7353 = P3_STATE2_REG_2_ & ~n7352;
  assign n7354 = ~P3_INSTADDRPOINTER_REG_0_ & n5657;
  assign n7355 = ~P3_INSTADDRPOINTER_REG_0_ & n5500;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = ~P3_INSTADDRPOINTER_REG_0_ & ~n5547;
  assign n7358 = P3_INSTADDRPOINTER_REG_0_ & n5618;
  assign n7359 = P3_INSTADDRPOINTER_REG_0_ & n5619_1;
  assign n7360 = n5359_1 & n5490;
  assign n7361 = n5496 & n7360;
  assign n7362 = ~P3_INSTADDRPOINTER_REG_0_ & n7361;
  assign n7363 = n5436 & n5490;
  assign n7364 = n5496 & n7363;
  assign n7365 = ~P3_INSTADDRPOINTER_REG_0_ & n7364;
  assign n7366 = ~n7362 & ~n7365;
  assign n7367 = P3_INSTADDRPOINTER_REG_0_ & n5434_1;
  assign n7368 = n7366 & ~n7367;
  assign n7369 = n5561 & n7243;
  assign n7370 = P3_INSTQUEUERD_ADDR_REG_0_ & ~n5673;
  assign n7371 = n7369 & n7370;
  assign n7372 = P3_INSTQUEUE_REG_0__0_ & n7371;
  assign n7373 = ~P3_INSTQUEUERD_ADDR_REG_0_ & ~n5673;
  assign n7374 = n7369 & n7373;
  assign n7375 = P3_INSTQUEUE_REG_1__0_ & n7374;
  assign n7376 = P3_INSTQUEUERD_ADDR_REG_0_ & n5673;
  assign n7377 = n7369 & n7376;
  assign n7378 = P3_INSTQUEUE_REG_2__0_ & n7377;
  assign n7379 = ~P3_INSTQUEUERD_ADDR_REG_0_ & n5673;
  assign n7380 = n7369 & n7379;
  assign n7381 = P3_INSTQUEUE_REG_3__0_ & n7380;
  assign n7382 = ~n7372 & ~n7375;
  assign n7383 = ~n7378 & n7382;
  assign n7384 = ~n7381 & n7383;
  assign n7385 = ~n5561 & n7243;
  assign n7386 = n7370 & n7385;
  assign n7387 = P3_INSTQUEUE_REG_4__0_ & n7386;
  assign n7388 = n7373 & n7385;
  assign n7389 = P3_INSTQUEUE_REG_5__0_ & n7388;
  assign n7390 = n7376 & n7385;
  assign n7391 = P3_INSTQUEUE_REG_6__0_ & n7390;
  assign n7392 = n7379 & n7385;
  assign n7393 = P3_INSTQUEUE_REG_7__0_ & n7392;
  assign n7394 = ~n7387 & ~n7389;
  assign n7395 = ~n7391 & n7394;
  assign n7396 = ~n7393 & n7395;
  assign n7397 = n5561 & ~n7243;
  assign n7398 = n7370 & n7397;
  assign n7399 = P3_INSTQUEUE_REG_8__0_ & n7398;
  assign n7400 = n7373 & n7397;
  assign n7401 = P3_INSTQUEUE_REG_9__0_ & n7400;
  assign n7402 = n7376 & n7397;
  assign n7403 = P3_INSTQUEUE_REG_10__0_ & n7402;
  assign n7404 = n7379 & n7397;
  assign n7405 = P3_INSTQUEUE_REG_11__0_ & n7404;
  assign n7406 = ~n7399 & ~n7401;
  assign n7407 = ~n7403 & n7406;
  assign n7408 = ~n7405 & n7407;
  assign n7409 = ~n5561 & ~n7243;
  assign n7410 = n7370 & n7409;
  assign n7411 = P3_INSTQUEUE_REG_12__0_ & n7410;
  assign n7412 = n7373 & n7409;
  assign n7413 = P3_INSTQUEUE_REG_13__0_ & n7412;
  assign n7414 = n7376 & n7409;
  assign n7415 = P3_INSTQUEUE_REG_14__0_ & n7414;
  assign n7416 = n7379 & n7409;
  assign n7417 = P3_INSTQUEUE_REG_15__0_ & n7416;
  assign n7418 = ~n7411 & ~n7413;
  assign n7419 = ~n7415 & n7418;
  assign n7420 = ~n7417 & n7419;
  assign n7421 = n7384 & n7396;
  assign n7422 = n7408 & n7421;
  assign n7423 = n7420 & n7422;
  assign n7424 = ~P3_INSTADDRPOINTER_REG_0_ & ~n7423;
  assign n7425 = P3_INSTADDRPOINTER_REG_0_ & n7423;
  assign n7426 = ~n7424 & ~n7425;
  assign n7427 = P3_INSTQUEUE_REG_0__7_ & n7371;
  assign n7428 = P3_INSTQUEUE_REG_1__7_ & n7374;
  assign n7429 = P3_INSTQUEUE_REG_2__7_ & n7377;
  assign n7430 = P3_INSTQUEUE_REG_3__7_ & n7380;
  assign n7431 = ~n7427 & ~n7428;
  assign n7432 = ~n7429 & n7431;
  assign n7433 = ~n7430 & n7432;
  assign n7434 = P3_INSTQUEUE_REG_4__7_ & n7386;
  assign n7435 = P3_INSTQUEUE_REG_5__7_ & n7388;
  assign n7436 = P3_INSTQUEUE_REG_6__7_ & n7390;
  assign n7437 = P3_INSTQUEUE_REG_7__7_ & n7392;
  assign n7438 = ~n7434 & ~n7435;
  assign n7439 = ~n7436 & n7438;
  assign n7440 = ~n7437 & n7439;
  assign n7441 = P3_INSTQUEUE_REG_8__7_ & n7398;
  assign n7442 = P3_INSTQUEUE_REG_9__7_ & n7400;
  assign n7443 = P3_INSTQUEUE_REG_10__7_ & n7402;
  assign n7444 = P3_INSTQUEUE_REG_11__7_ & n7404;
  assign n7445 = ~n7441 & ~n7442;
  assign n7446 = ~n7443 & n7445;
  assign n7447 = ~n7444 & n7446;
  assign n7448 = P3_INSTQUEUE_REG_12__7_ & n7410;
  assign n7449 = P3_INSTQUEUE_REG_13__7_ & n7412;
  assign n7450 = P3_INSTQUEUE_REG_14__7_ & n7414;
  assign n7451 = P3_INSTQUEUE_REG_15__7_ & n7416;
  assign n7452 = ~n7448 & ~n7449;
  assign n7453 = ~n7450 & n7452;
  assign n7454 = ~n7451 & n7453;
  assign n7455 = n7433 & n7440;
  assign n7456 = n7447 & n7455;
  assign n7457 = n7454 & n7456;
  assign n7458 = n5466 & ~n7457;
  assign n7459 = ~n7426 & n7458;
  assign n7460 = n5466 & n7457;
  assign n7461 = ~n7426 & n7460;
  assign n7462 = ~n7358 & ~n7359;
  assign n7463 = n7368 & n7462;
  assign n7464 = ~n7459 & n7463;
  assign n7465 = ~n7461 & n7464;
  assign n7466 = n5432 & n5460;
  assign n7467 = ~P3_INSTADDRPOINTER_REG_0_ & n7466;
  assign n7468 = ~P3_INSTADDRPOINTER_REG_0_ & n5504_1;
  assign n7469 = n5261 & n5447;
  assign n7470 = n5493 & n7469;
  assign n7471 = ~P3_INSTADDRPOINTER_REG_0_ & n7470;
  assign n7472 = ~P3_INSTADDRPOINTER_REG_0_ & n7423;
  assign n7473 = P3_INSTADDRPOINTER_REG_0_ & ~n7423;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n5461 & ~n7474;
  assign n7476 = n5136_1 & n5490;
  assign n7477 = n5493 & n7476;
  assign n7478 = ~P3_INSTADDRPOINTER_REG_0_ & n7477;
  assign n7479 = ~n7467 & ~n7468;
  assign n7480 = ~n7471 & n7479;
  assign n7481 = ~n7475 & n7480;
  assign n7482 = ~n7478 & n7481;
  assign n7483 = P3_INSTADDRPOINTER_REG_0_ & n5360;
  assign n7484 = P3_INSTADDRPOINTER_REG_0_ & n5438;
  assign n7485 = P3_INSTADDRPOINTER_REG_0_ & n5442;
  assign n7486 = ~P3_INSTADDRPOINTER_REG_0_ & n5458;
  assign n7487 = ~P3_INSTADDRPOINTER_REG_0_ & n5450;
  assign n7488 = ~n7483 & ~n7484;
  assign n7489 = ~n7485 & n7488;
  assign n7490 = ~n7486 & n7489;
  assign n7491 = ~n7487 & n7490;
  assign n7492 = n7482 & n7491;
  assign n7493 = n7356 & ~n7357;
  assign n7494 = n7465 & n7493;
  assign n7495 = n7492 & n7494;
  assign n7496 = n7353 & ~n7495;
  assign n7497 = ~P3_STATE2_REG_2_ & ~n7352;
  assign n7498 = P3_REIP_REG_0_ & n7497;
  assign n7499 = P3_INSTADDRPOINTER_REG_0_ & n7352;
  assign n7500 = ~n7496 & ~n7498;
  assign n1665 = n7499 | ~n7500;
  assign n7502 = P3_INSTADDRPOINTER_REG_1_ & n7352;
  assign n7503 = P3_REIP_REG_1_ & n7497;
  assign n7504 = ~n5547 & ~n5741;
  assign n7505 = n5657 & ~n5741;
  assign n7506 = n5500 & ~n5741;
  assign n7507 = ~n7505 & ~n7506;
  assign n7508 = ~P3_INSTADDRPOINTER_REG_1_ & n7473;
  assign n7509 = P3_INSTADDRPOINTER_REG_1_ & ~n7473;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = P3_INSTQUEUE_REG_0__1_ & n7371;
  assign n7512 = P3_INSTQUEUE_REG_1__1_ & n7374;
  assign n7513 = P3_INSTQUEUE_REG_2__1_ & n7377;
  assign n7514 = P3_INSTQUEUE_REG_3__1_ & n7380;
  assign n7515 = ~n7511 & ~n7512;
  assign n7516 = ~n7513 & n7515;
  assign n7517 = ~n7514 & n7516;
  assign n7518 = P3_INSTQUEUE_REG_4__1_ & n7386;
  assign n7519 = P3_INSTQUEUE_REG_5__1_ & n7388;
  assign n7520 = P3_INSTQUEUE_REG_6__1_ & n7390;
  assign n7521 = P3_INSTQUEUE_REG_7__1_ & n7392;
  assign n7522 = ~n7518 & ~n7519;
  assign n7523 = ~n7520 & n7522;
  assign n7524 = ~n7521 & n7523;
  assign n7525 = P3_INSTQUEUE_REG_8__1_ & n7398;
  assign n7526 = P3_INSTQUEUE_REG_9__1_ & n7400;
  assign n7527 = P3_INSTQUEUE_REG_10__1_ & n7402;
  assign n7528 = P3_INSTQUEUE_REG_11__1_ & n7404;
  assign n7529 = ~n7525 & ~n7526;
  assign n7530 = ~n7527 & n7529;
  assign n7531 = ~n7528 & n7530;
  assign n7532 = P3_INSTQUEUE_REG_12__1_ & n7410;
  assign n7533 = P3_INSTQUEUE_REG_13__1_ & n7412;
  assign n7534 = P3_INSTQUEUE_REG_14__1_ & n7414;
  assign n7535 = P3_INSTQUEUE_REG_15__1_ & n7416;
  assign n7536 = ~n7532 & ~n7533;
  assign n7537 = ~n7534 & n7536;
  assign n7538 = ~n7535 & n7537;
  assign n7539 = n7517 & n7524;
  assign n7540 = n7531 & n7539;
  assign n7541 = n7538 & n7540;
  assign n7542 = ~n7510 & ~n7541;
  assign n7543 = ~P3_INSTADDRPOINTER_REG_1_ & ~n7473;
  assign n7544 = n7541 & n7543;
  assign n7545 = n7473 & n7541;
  assign n7546 = P3_INSTADDRPOINTER_REG_1_ & n7545;
  assign n7547 = ~n7542 & ~n7544;
  assign n7548 = ~n7546 & n7547;
  assign n7549 = n7460 & ~n7548;
  assign n7550 = ~n5741 & n7477;
  assign n7551 = ~n5741 & n7470;
  assign n7552 = ~n5741 & n7466;
  assign n7553 = n5504_1 & ~n5741;
  assign n7554 = ~n7550 & ~n7551;
  assign n7555 = ~n7552 & n7554;
  assign n7556 = ~n7553 & n7555;
  assign n7557 = ~P3_INSTADDRPOINTER_REG_1_ & n5360;
  assign n7558 = ~P3_INSTADDRPOINTER_REG_1_ & n5438;
  assign n7559 = ~P3_INSTADDRPOINTER_REG_1_ & n5442;
  assign n7560 = n5458 & ~n5741;
  assign n7561 = n5450 & ~n5741;
  assign n7562 = ~n7557 & ~n7558;
  assign n7563 = ~n7559 & n7562;
  assign n7564 = ~n7560 & n7563;
  assign n7565 = ~n7561 & n7564;
  assign n7566 = ~P3_INSTADDRPOINTER_REG_1_ & n7425;
  assign n7567 = P3_INSTADDRPOINTER_REG_1_ & ~n7425;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = ~n7423 & n7541;
  assign n7570 = n7423 & ~n7541;
  assign n7571 = ~n7569 & ~n7570;
  assign n7572 = ~n7568 & n7571;
  assign n7573 = ~P3_INSTADDRPOINTER_REG_1_ & ~n7425;
  assign n7574 = ~n7571 & n7573;
  assign n7575 = n7425 & ~n7571;
  assign n7576 = P3_INSTADDRPOINTER_REG_1_ & n7575;
  assign n7577 = ~n7572 & ~n7574;
  assign n7578 = ~n7576 & n7577;
  assign n7579 = n5461 & ~n7578;
  assign n7580 = n7556 & n7565;
  assign n7581 = ~n7579 & n7580;
  assign n7582 = ~P3_INSTADDRPOINTER_REG_1_ & n5618;
  assign n7583 = ~P3_INSTADDRPOINTER_REG_1_ & n5619_1;
  assign n7584 = ~n5741 & n7361;
  assign n7585 = ~n5741 & n7364;
  assign n7586 = ~n7584 & ~n7585;
  assign n7587 = ~P3_INSTADDRPOINTER_REG_1_ & n5434_1;
  assign n7588 = n7586 & ~n7587;
  assign n7589 = n7458 & ~n7548;
  assign n7590 = ~n7582 & ~n7583;
  assign n7591 = n7588 & n7590;
  assign n7592 = ~n7589 & n7591;
  assign n7593 = ~n7504 & n7507;
  assign n7594 = ~n7549 & n7593;
  assign n7595 = n7581 & n7594;
  assign n7596 = n7592 & n7595;
  assign n7597 = n7353 & ~n7596;
  assign n7598 = ~n7502 & ~n7503;
  assign n1670 = n7597 | ~n7598;
  assign n7600 = P3_INSTADDRPOINTER_REG_2_ & n7352;
  assign n7601 = P3_REIP_REG_2_ & n7497;
  assign n7602 = P3_INSTADDRPOINTER_REG_0_ & P3_INSTADDRPOINTER_REG_1_;
  assign n7603 = ~P3_INSTADDRPOINTER_REG_2_ & n7602;
  assign n7604 = P3_INSTADDRPOINTER_REG_2_ & ~n7602;
  assign n7605 = ~n7603 & ~n7604;
  assign n7606 = ~n5547 & ~n7605;
  assign n7607 = P3_INSTADDRPOINTER_REG_1_ & ~P3_INSTADDRPOINTER_REG_2_;
  assign n7608 = ~P3_INSTADDRPOINTER_REG_1_ & P3_INSTADDRPOINTER_REG_2_;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = n5618 & ~n7609;
  assign n7611 = n5619_1 & ~n7609;
  assign n7612 = n7361 & ~n7605;
  assign n7613 = n7364 & ~n7605;
  assign n7614 = ~n7612 & ~n7613;
  assign n7615 = n5434_1 & ~n7609;
  assign n7616 = n7614 & ~n7615;
  assign n7617 = ~n7610 & ~n7611;
  assign n7618 = n7616 & n7617;
  assign n7619 = ~n7473 & ~n7541;
  assign n7620 = P3_INSTADDRPOINTER_REG_1_ & ~n7619;
  assign n7621 = ~n7545 & ~n7620;
  assign n7622 = P3_INSTQUEUE_REG_0__2_ & n7371;
  assign n7623 = P3_INSTQUEUE_REG_1__2_ & n7374;
  assign n7624 = P3_INSTQUEUE_REG_2__2_ & n7377;
  assign n7625 = P3_INSTQUEUE_REG_3__2_ & n7380;
  assign n7626 = ~n7622 & ~n7623;
  assign n7627 = ~n7624 & n7626;
  assign n7628 = ~n7625 & n7627;
  assign n7629 = P3_INSTQUEUE_REG_4__2_ & n7386;
  assign n7630 = P3_INSTQUEUE_REG_5__2_ & n7388;
  assign n7631 = P3_INSTQUEUE_REG_6__2_ & n7390;
  assign n7632 = P3_INSTQUEUE_REG_7__2_ & n7392;
  assign n7633 = ~n7629 & ~n7630;
  assign n7634 = ~n7631 & n7633;
  assign n7635 = ~n7632 & n7634;
  assign n7636 = P3_INSTQUEUE_REG_8__2_ & n7398;
  assign n7637 = P3_INSTQUEUE_REG_9__2_ & n7400;
  assign n7638 = P3_INSTQUEUE_REG_10__2_ & n7402;
  assign n7639 = P3_INSTQUEUE_REG_11__2_ & n7404;
  assign n7640 = ~n7636 & ~n7637;
  assign n7641 = ~n7638 & n7640;
  assign n7642 = ~n7639 & n7641;
  assign n7643 = P3_INSTQUEUE_REG_12__2_ & n7410;
  assign n7644 = P3_INSTQUEUE_REG_13__2_ & n7412;
  assign n7645 = P3_INSTQUEUE_REG_14__2_ & n7414;
  assign n7646 = P3_INSTQUEUE_REG_15__2_ & n7416;
  assign n7647 = ~n7643 & ~n7644;
  assign n7648 = ~n7645 & n7647;
  assign n7649 = ~n7646 & n7648;
  assign n7650 = n7628 & n7635;
  assign n7651 = n7642 & n7650;
  assign n7652 = n7649 & n7651;
  assign n7653 = ~n7541 & n7652;
  assign n7654 = n7541 & ~n7652;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = ~P3_INSTADDRPOINTER_REG_2_ & ~n7655;
  assign n7657 = P3_INSTADDRPOINTER_REG_2_ & n7655;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = n7621 & ~n7658;
  assign n7660 = ~n7621 & n7658;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = n7460 & ~n7661;
  assign n7663 = n5657 & ~n7605;
  assign n7664 = n5500 & ~n7605;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = P3_INSTADDRPOINTER_REG_1_ & n7473;
  assign n7667 = P3_INSTADDRPOINTER_REG_1_ & n7541;
  assign n7668 = ~n7545 & ~n7666;
  assign n7669 = ~n7667 & n7668;
  assign n7670 = ~n7658 & n7669;
  assign n7671 = ~P3_INSTADDRPOINTER_REG_2_ & n7655;
  assign n7672 = P3_INSTADDRPOINTER_REG_2_ & ~n7655;
  assign n7673 = ~n7671 & ~n7672;
  assign n7674 = ~n7669 & ~n7673;
  assign n7675 = ~n7670 & ~n7674;
  assign n7676 = n7458 & ~n7675;
  assign n7677 = n7665 & ~n7676;
  assign n7678 = n7477 & ~n7605;
  assign n7679 = n7470 & ~n7605;
  assign n7680 = n7466 & ~n7605;
  assign n7681 = n5504_1 & ~n7605;
  assign n7682 = ~n7678 & ~n7679;
  assign n7683 = ~n7680 & n7682;
  assign n7684 = ~n7681 & n7683;
  assign n7685 = n5360 & ~n7609;
  assign n7686 = n5438 & ~n7609;
  assign n7687 = n5442 & ~n7609;
  assign n7688 = ~P3_INSTADDRPOINTER_REG_2_ & ~n7602;
  assign n7689 = P3_INSTADDRPOINTER_REG_2_ & n7602;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 = n5458 & ~n7690;
  assign n7692 = n5450 & ~n7690;
  assign n7693 = ~n7685 & ~n7686;
  assign n7694 = ~n7687 & n7693;
  assign n7695 = ~n7691 & n7694;
  assign n7696 = ~n7692 & n7695;
  assign n7697 = ~n7423 & ~n7541;
  assign n7698 = n7652 & ~n7697;
  assign n7699 = ~n7652 & n7697;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = ~P3_INSTADDRPOINTER_REG_2_ & ~n7700;
  assign n7702 = P3_INSTADDRPOINTER_REG_2_ & n7700;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = ~n7425 & n7571;
  assign n7705 = P3_INSTADDRPOINTER_REG_1_ & ~n7704;
  assign n7706 = ~n7575 & ~n7705;
  assign n7707 = ~n7703 & n7706;
  assign n7708 = ~P3_INSTADDRPOINTER_REG_2_ & n7700;
  assign n7709 = P3_INSTADDRPOINTER_REG_2_ & ~n7700;
  assign n7710 = ~n7708 & ~n7709;
  assign n7711 = ~n7706 & ~n7710;
  assign n7712 = ~n7707 & ~n7711;
  assign n7713 = n5461 & ~n7712;
  assign n7714 = n7684 & n7696;
  assign n7715 = ~n7713 & n7714;
  assign n7716 = ~n7606 & n7618;
  assign n7717 = ~n7662 & n7716;
  assign n7718 = n7677 & n7717;
  assign n7719 = n7715 & n7718;
  assign n7720 = n7353 & ~n7719;
  assign n7721 = ~n7600 & ~n7601;
  assign n1675 = n7720 | ~n7721;
  assign n7723 = P3_INSTADDRPOINTER_REG_3_ & n7352;
  assign n7724 = P3_REIP_REG_3_ & n7497;
  assign n7725 = ~P3_INSTADDRPOINTER_REG_3_ & n7689;
  assign n7726 = P3_INSTADDRPOINTER_REG_3_ & ~n7689;
  assign n7727 = ~n7725 & ~n7726;
  assign n7728 = n5657 & ~n7727;
  assign n7729 = n5500 & ~n7727;
  assign n7730 = ~n7728 & ~n7729;
  assign n7731 = ~n5547 & ~n7727;
  assign n7732 = P3_INSTADDRPOINTER_REG_1_ & P3_INSTADDRPOINTER_REG_2_;
  assign n7733 = ~P3_INSTADDRPOINTER_REG_3_ & n7732;
  assign n7734 = P3_INSTADDRPOINTER_REG_3_ & ~n7732;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = n5618 & ~n7735;
  assign n7737 = n5619_1 & ~n7735;
  assign n7738 = n7361 & ~n7727;
  assign n7739 = P3_INSTADDRPOINTER_REG_0_ & P3_INSTADDRPOINTER_REG_2_;
  assign n7740 = P3_INSTADDRPOINTER_REG_1_ & n7739;
  assign n7741 = P3_INSTADDRPOINTER_REG_3_ & ~n7740;
  assign n7742 = ~P3_INSTADDRPOINTER_REG_3_ & n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = n7364 & ~n7743;
  assign n7745 = ~n7738 & ~n7744;
  assign n7746 = n5434_1 & ~n7735;
  assign n7747 = n7745 & ~n7746;
  assign n7748 = ~n7736 & ~n7737;
  assign n7749 = n7747 & n7748;
  assign n7750 = ~n7669 & ~n7671;
  assign n7751 = ~n7672 & ~n7750;
  assign n7752 = P3_INSTQUEUE_REG_0__3_ & n7371;
  assign n7753 = P3_INSTQUEUE_REG_1__3_ & n7374;
  assign n7754 = P3_INSTQUEUE_REG_2__3_ & n7377;
  assign n7755 = P3_INSTQUEUE_REG_3__3_ & n7380;
  assign n7756 = ~n7752 & ~n7753;
  assign n7757 = ~n7754 & n7756;
  assign n7758 = ~n7755 & n7757;
  assign n7759 = P3_INSTQUEUE_REG_4__3_ & n7386;
  assign n7760 = P3_INSTQUEUE_REG_5__3_ & n7388;
  assign n7761 = P3_INSTQUEUE_REG_6__3_ & n7390;
  assign n7762 = P3_INSTQUEUE_REG_7__3_ & n7392;
  assign n7763 = ~n7759 & ~n7760;
  assign n7764 = ~n7761 & n7763;
  assign n7765 = ~n7762 & n7764;
  assign n7766 = P3_INSTQUEUE_REG_8__3_ & n7398;
  assign n7767 = P3_INSTQUEUE_REG_9__3_ & n7400;
  assign n7768 = P3_INSTQUEUE_REG_10__3_ & n7402;
  assign n7769 = P3_INSTQUEUE_REG_11__3_ & n7404;
  assign n7770 = ~n7766 & ~n7767;
  assign n7771 = ~n7768 & n7770;
  assign n7772 = ~n7769 & n7771;
  assign n7773 = P3_INSTQUEUE_REG_12__3_ & n7410;
  assign n7774 = P3_INSTQUEUE_REG_13__3_ & n7412;
  assign n7775 = P3_INSTQUEUE_REG_14__3_ & n7414;
  assign n7776 = P3_INSTQUEUE_REG_15__3_ & n7416;
  assign n7777 = ~n7773 & ~n7774;
  assign n7778 = ~n7775 & n7777;
  assign n7779 = ~n7776 & n7778;
  assign n7780 = n7758 & n7765;
  assign n7781 = n7772 & n7780;
  assign n7782 = n7779 & n7781;
  assign n7783 = ~n7541 & ~n7652;
  assign n7784 = n7782 & ~n7783;
  assign n7785 = ~n7782 & n7783;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = ~P3_INSTADDRPOINTER_REG_3_ & n7786;
  assign n7788 = P3_INSTADDRPOINTER_REG_3_ & ~n7786;
  assign n7789 = ~n7787 & ~n7788;
  assign n7790 = n7751 & ~n7789;
  assign n7791 = P3_INSTADDRPOINTER_REG_3_ & n7786;
  assign n7792 = ~P3_INSTADDRPOINTER_REG_3_ & ~n7786;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = ~n7751 & ~n7793;
  assign n7795 = ~n7790 & ~n7794;
  assign n7796 = n7458 & ~n7795;
  assign n7797 = ~n7621 & ~n7671;
  assign n7798 = ~n7672 & ~n7797;
  assign n7799 = n7782 & n7783;
  assign n7800 = ~n7782 & ~n7783;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~P3_INSTADDRPOINTER_REG_3_ & n7801;
  assign n7803 = ~n7798 & ~n7802;
  assign n7804 = P3_INSTADDRPOINTER_REG_3_ & ~n7801;
  assign n7805 = n7803 & ~n7804;
  assign n7806 = ~P3_INSTADDRPOINTER_REG_3_ & ~n7801;
  assign n7807 = P3_INSTADDRPOINTER_REG_3_ & n7801;
  assign n7808 = ~n7806 & ~n7807;
  assign n7809 = n7798 & n7808;
  assign n7810 = ~n7805 & ~n7809;
  assign n7811 = n7460 & n7810;
  assign n7812 = ~n7796 & ~n7811;
  assign n7813 = n7477 & ~n7727;
  assign n7814 = n7470 & ~n7727;
  assign n7815 = n7466 & ~n7727;
  assign n7816 = n5504_1 & ~n7727;
  assign n7817 = ~n7813 & ~n7814;
  assign n7818 = ~n7815 & n7817;
  assign n7819 = ~n7816 & n7818;
  assign n7820 = n5360 & ~n7735;
  assign n7821 = n5438 & ~n7735;
  assign n7822 = n5442 & ~n7735;
  assign n7823 = ~P3_INSTADDRPOINTER_REG_3_ & n7688;
  assign n7824 = P3_INSTADDRPOINTER_REG_3_ & ~n7688;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = n5458 & n7825;
  assign n7827 = n5450 & n7825;
  assign n7828 = ~n7820 & ~n7821;
  assign n7829 = ~n7822 & n7828;
  assign n7830 = ~n7826 & n7829;
  assign n7831 = ~n7827 & n7830;
  assign n7832 = n7706 & ~n7709;
  assign n7833 = n7698 & n7782;
  assign n7834 = ~n7698 & ~n7782;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = P3_INSTADDRPOINTER_REG_3_ & n7835;
  assign n7837 = ~n7708 & n7835;
  assign n7838 = P3_INSTADDRPOINTER_REG_3_ & ~n7708;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~n7832 & ~n7836;
  assign n7841 = ~n7839 & n7840;
  assign n7842 = ~P3_INSTADDRPOINTER_REG_3_ & n7835;
  assign n7843 = P3_INSTADDRPOINTER_REG_3_ & ~n7835;
  assign n7844 = ~n7842 & ~n7843;
  assign n7845 = ~n7709 & n7844;
  assign n7846 = ~n7706 & ~n7708;
  assign n7847 = n7845 & ~n7846;
  assign n7848 = ~n7841 & ~n7847;
  assign n7849 = n5461 & n7848;
  assign n7850 = n7819 & n7831;
  assign n7851 = ~n7849 & n7850;
  assign n7852 = n7730 & ~n7731;
  assign n7853 = n7749 & n7852;
  assign n7854 = n7812 & n7853;
  assign n7855 = n7851 & n7854;
  assign n7856 = n7353 & ~n7855;
  assign n7857 = ~n7723 & ~n7724;
  assign n1680 = n7856 | ~n7857;
  assign n7859 = P3_INSTADDRPOINTER_REG_4_ & n7352;
  assign n7860 = P3_REIP_REG_4_ & n7497;
  assign n7861 = P3_INSTADDRPOINTER_REG_3_ & n7689;
  assign n7862 = ~P3_INSTADDRPOINTER_REG_4_ & n7861;
  assign n7863 = P3_INSTADDRPOINTER_REG_4_ & ~n7861;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~n5547 & ~n7864;
  assign n7866 = P3_INSTADDRPOINTER_REG_3_ & n7732;
  assign n7867 = ~P3_INSTADDRPOINTER_REG_4_ & n7866;
  assign n7868 = P3_INSTADDRPOINTER_REG_4_ & ~n7866;
  assign n7869 = ~n7867 & ~n7868;
  assign n7870 = n5618 & ~n7869;
  assign n7871 = n5619_1 & ~n7869;
  assign n7872 = n7361 & ~n7864;
  assign n7873 = P3_INSTADDRPOINTER_REG_3_ & n7740;
  assign n7874 = ~P3_INSTADDRPOINTER_REG_4_ & n7873;
  assign n7875 = P3_INSTADDRPOINTER_REG_4_ & ~n7873;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = n7364 & ~n7876;
  assign n7878 = ~n7872 & ~n7877;
  assign n7879 = n5434_1 & ~n7869;
  assign n7880 = n7878 & ~n7879;
  assign n7881 = ~n7870 & ~n7871;
  assign n7882 = n7880 & n7881;
  assign n7883 = P3_INSTQUEUE_REG_0__4_ & n7371;
  assign n7884 = P3_INSTQUEUE_REG_1__4_ & n7374;
  assign n7885 = P3_INSTQUEUE_REG_2__4_ & n7377;
  assign n7886 = P3_INSTQUEUE_REG_3__4_ & n7380;
  assign n7887 = ~n7883 & ~n7884;
  assign n7888 = ~n7885 & n7887;
  assign n7889 = ~n7886 & n7888;
  assign n7890 = P3_INSTQUEUE_REG_4__4_ & n7386;
  assign n7891 = P3_INSTQUEUE_REG_5__4_ & n7388;
  assign n7892 = P3_INSTQUEUE_REG_6__4_ & n7390;
  assign n7893 = P3_INSTQUEUE_REG_7__4_ & n7392;
  assign n7894 = ~n7890 & ~n7891;
  assign n7895 = ~n7892 & n7894;
  assign n7896 = ~n7893 & n7895;
  assign n7897 = P3_INSTQUEUE_REG_8__4_ & n7398;
  assign n7898 = P3_INSTQUEUE_REG_9__4_ & n7400;
  assign n7899 = P3_INSTQUEUE_REG_10__4_ & n7402;
  assign n7900 = P3_INSTQUEUE_REG_11__4_ & n7404;
  assign n7901 = ~n7897 & ~n7898;
  assign n7902 = ~n7899 & n7901;
  assign n7903 = ~n7900 & n7902;
  assign n7904 = P3_INSTQUEUE_REG_12__4_ & n7410;
  assign n7905 = P3_INSTQUEUE_REG_13__4_ & n7412;
  assign n7906 = P3_INSTQUEUE_REG_14__4_ & n7414;
  assign n7907 = P3_INSTQUEUE_REG_15__4_ & n7416;
  assign n7908 = ~n7904 & ~n7905;
  assign n7909 = ~n7906 & n7908;
  assign n7910 = ~n7907 & n7909;
  assign n7911 = n7889 & n7896;
  assign n7912 = n7903 & n7911;
  assign n7913 = n7910 & n7912;
  assign n7914 = n7785 & n7913;
  assign n7915 = ~n7785 & ~n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = P3_INSTADDRPOINTER_REG_4_ & ~n7916;
  assign n7918 = ~P3_INSTADDRPOINTER_REG_4_ & n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7803 & ~n7804;
  assign n7921 = n7919 & ~n7920;
  assign n7922 = ~P3_INSTADDRPOINTER_REG_4_ & ~n7916;
  assign n7923 = P3_INSTADDRPOINTER_REG_4_ & n7916;
  assign n7924 = ~n7922 & ~n7923;
  assign n7925 = ~n7804 & n7924;
  assign n7926 = ~n7803 & n7925;
  assign n7927 = ~n7921 & ~n7926;
  assign n7928 = n7460 & n7927;
  assign n7929 = n5657 & ~n7864;
  assign n7930 = n5500 & ~n7864;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = ~n7671 & ~n7792;
  assign n7933 = ~n7666 & ~n7667;
  assign n7934 = ~n7672 & n7933;
  assign n7935 = ~n7545 & n7934;
  assign n7936 = n7932 & ~n7935;
  assign n7937 = ~n7791 & ~n7936;
  assign n7938 = n7785 & ~n7913;
  assign n7939 = ~n7785 & n7913;
  assign n7940 = ~n7938 & ~n7939;
  assign n7941 = ~P3_INSTADDRPOINTER_REG_4_ & n7940;
  assign n7942 = P3_INSTADDRPOINTER_REG_4_ & ~n7940;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = n7937 & ~n7943;
  assign n7945 = P3_INSTADDRPOINTER_REG_4_ & n7940;
  assign n7946 = ~P3_INSTADDRPOINTER_REG_4_ & ~n7940;
  assign n7947 = ~n7945 & ~n7946;
  assign n7948 = ~n7937 & ~n7947;
  assign n7949 = ~n7944 & ~n7948;
  assign n7950 = n7458 & ~n7949;
  assign n7951 = n7931 & ~n7950;
  assign n7952 = n7477 & ~n7864;
  assign n7953 = n7470 & ~n7864;
  assign n7954 = n7466 & ~n7864;
  assign n7955 = n5504_1 & ~n7864;
  assign n7956 = ~n7952 & ~n7953;
  assign n7957 = ~n7954 & n7956;
  assign n7958 = ~n7955 & n7957;
  assign n7959 = n5360 & ~n7869;
  assign n7960 = n5438 & ~n7869;
  assign n7961 = n5442 & ~n7869;
  assign n7962 = ~P3_INSTADDRPOINTER_REG_4_ & n7824;
  assign n7963 = P3_INSTADDRPOINTER_REG_4_ & ~n7824;
  assign n7964 = ~n7962 & ~n7963;
  assign n7965 = n5458 & ~n7964;
  assign n7966 = n5450 & ~n7964;
  assign n7967 = ~n7959 & ~n7960;
  assign n7968 = ~n7961 & n7967;
  assign n7969 = ~n7965 & n7968;
  assign n7970 = ~n7966 & n7969;
  assign n7971 = n7834 & n7913;
  assign n7972 = ~n7834 & ~n7913;
  assign n7973 = ~n7971 & ~n7972;
  assign n7974 = ~P3_INSTADDRPOINTER_REG_4_ & ~n7973;
  assign n7975 = P3_INSTADDRPOINTER_REG_4_ & n7973;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = n7709 & n7835;
  assign n7978 = ~n7709 & ~n7835;
  assign n7979 = P3_INSTADDRPOINTER_REG_3_ & ~n7978;
  assign n7980 = ~n7977 & ~n7979;
  assign n7981 = ~n7706 & ~n7839;
  assign n7982 = n7980 & ~n7981;
  assign n7983 = ~n7976 & n7982;
  assign n7984 = ~P3_INSTADDRPOINTER_REG_4_ & n7973;
  assign n7985 = P3_INSTADDRPOINTER_REG_4_ & ~n7973;
  assign n7986 = ~n7984 & ~n7985;
  assign n7987 = ~n7982 & ~n7986;
  assign n7988 = ~n7983 & ~n7987;
  assign n7989 = n5461 & ~n7988;
  assign n7990 = n7958 & n7970;
  assign n7991 = ~n7989 & n7990;
  assign n7992 = ~n7865 & n7882;
  assign n7993 = ~n7928 & n7992;
  assign n7994 = n7951 & n7993;
  assign n7995 = n7991 & n7994;
  assign n7996 = n7353 & ~n7995;
  assign n7997 = ~n7859 & ~n7860;
  assign n1685 = n7996 | ~n7997;
  assign n7999 = P3_INSTADDRPOINTER_REG_5_ & n7352;
  assign n8000 = P3_REIP_REG_5_ & n7497;
  assign n8001 = P3_INSTADDRPOINTER_REG_4_ & n7866;
  assign n8002 = ~P3_INSTADDRPOINTER_REG_5_ & n8001;
  assign n8003 = P3_INSTADDRPOINTER_REG_5_ & ~n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = n5618 & ~n8004;
  assign n8006 = n5619_1 & ~n8004;
  assign n8007 = P3_INSTADDRPOINTER_REG_4_ & n7861;
  assign n8008 = ~P3_INSTADDRPOINTER_REG_5_ & n8007;
  assign n8009 = P3_INSTADDRPOINTER_REG_5_ & ~n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = n7361 & ~n8010;
  assign n8012 = P3_INSTADDRPOINTER_REG_3_ & P3_INSTADDRPOINTER_REG_4_;
  assign n8013 = n7740 & n8012;
  assign n8014 = P3_INSTADDRPOINTER_REG_5_ & ~n8013;
  assign n8015 = ~P3_INSTADDRPOINTER_REG_5_ & n8013;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = n7364 & ~n8016;
  assign n8018 = ~n8011 & ~n8017;
  assign n8019 = n5434_1 & ~n8004;
  assign n8020 = n8018 & ~n8019;
  assign n8021 = ~n8005 & ~n8006;
  assign n8022 = n8020 & n8021;
  assign n8023 = ~n5547 & ~n8010;
  assign n8024 = n7791 & ~n7946;
  assign n8025 = ~n7945 & ~n8024;
  assign n8026 = n7932 & ~n7946;
  assign n8027 = ~n7935 & n8026;
  assign n8028 = n8025 & ~n8027;
  assign n8029 = P3_INSTQUEUE_REG_0__5_ & n7371;
  assign n8030 = P3_INSTQUEUE_REG_1__5_ & n7374;
  assign n8031 = P3_INSTQUEUE_REG_2__5_ & n7377;
  assign n8032 = P3_INSTQUEUE_REG_3__5_ & n7380;
  assign n8033 = ~n8029 & ~n8030;
  assign n8034 = ~n8031 & n8033;
  assign n8035 = ~n8032 & n8034;
  assign n8036 = P3_INSTQUEUE_REG_4__5_ & n7386;
  assign n8037 = P3_INSTQUEUE_REG_5__5_ & n7388;
  assign n8038 = P3_INSTQUEUE_REG_6__5_ & n7390;
  assign n8039 = P3_INSTQUEUE_REG_7__5_ & n7392;
  assign n8040 = ~n8036 & ~n8037;
  assign n8041 = ~n8038 & n8040;
  assign n8042 = ~n8039 & n8041;
  assign n8043 = P3_INSTQUEUE_REG_8__5_ & n7398;
  assign n8044 = P3_INSTQUEUE_REG_9__5_ & n7400;
  assign n8045 = P3_INSTQUEUE_REG_10__5_ & n7402;
  assign n8046 = P3_INSTQUEUE_REG_11__5_ & n7404;
  assign n8047 = ~n8043 & ~n8044;
  assign n8048 = ~n8045 & n8047;
  assign n8049 = ~n8046 & n8048;
  assign n8050 = P3_INSTQUEUE_REG_12__5_ & n7410;
  assign n8051 = P3_INSTQUEUE_REG_13__5_ & n7412;
  assign n8052 = P3_INSTQUEUE_REG_14__5_ & n7414;
  assign n8053 = P3_INSTQUEUE_REG_15__5_ & n7416;
  assign n8054 = ~n8050 & ~n8051;
  assign n8055 = ~n8052 & n8054;
  assign n8056 = ~n8053 & n8055;
  assign n8057 = n8035 & n8042;
  assign n8058 = n8049 & n8057;
  assign n8059 = n8056 & n8058;
  assign n8060 = ~n7938 & n8059;
  assign n8061 = ~n7913 & ~n8059;
  assign n8062 = n7785 & n8061;
  assign n8063 = ~n8060 & ~n8062;
  assign n8064 = ~P3_INSTADDRPOINTER_REG_5_ & n8063;
  assign n8065 = P3_INSTADDRPOINTER_REG_5_ & ~n8063;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = n8028 & ~n8066;
  assign n8068 = ~n8028 & n8066;
  assign n8069 = ~n8067 & ~n8068;
  assign n8070 = n7458 & ~n8069;
  assign n8071 = n5657 & ~n8010;
  assign n8072 = n5500 & ~n8010;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = n7804 & ~n7918;
  assign n8075 = ~n7917 & ~n8074;
  assign n8076 = ~n7802 & ~n7918;
  assign n8077 = ~n7798 & n8076;
  assign n8078 = n8075 & ~n8077;
  assign n8079 = n7938 & n8059;
  assign n8080 = ~n7938 & ~n8059;
  assign n8081 = ~n8079 & ~n8080;
  assign n8082 = ~P3_INSTADDRPOINTER_REG_5_ & ~n8081;
  assign n8083 = P3_INSTADDRPOINTER_REG_5_ & n8081;
  assign n8084 = ~n8082 & ~n8083;
  assign n8085 = n8078 & ~n8084;
  assign n8086 = ~n8078 & n8084;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = n7460 & ~n8087;
  assign n8089 = n8073 & ~n8088;
  assign n8090 = n7477 & ~n8010;
  assign n8091 = n7470 & ~n8010;
  assign n8092 = n7466 & ~n8010;
  assign n8093 = n5504_1 & ~n8010;
  assign n8094 = ~n8090 & ~n8091;
  assign n8095 = ~n8092 & n8094;
  assign n8096 = ~n8093 & n8095;
  assign n8097 = n5360 & ~n8004;
  assign n8098 = n5438 & ~n8004;
  assign n8099 = n5442 & ~n8004;
  assign n8100 = P3_INSTADDRPOINTER_REG_4_ & n7824;
  assign n8101 = ~P3_INSTADDRPOINTER_REG_5_ & n8100;
  assign n8102 = P3_INSTADDRPOINTER_REG_5_ & ~n8100;
  assign n8103 = ~n8101 & ~n8102;
  assign n8104 = n5458 & ~n8103;
  assign n8105 = n5450 & ~n8103;
  assign n8106 = ~n8097 & ~n8098;
  assign n8107 = ~n8099 & n8106;
  assign n8108 = ~n8104 & n8107;
  assign n8109 = ~n8105 & n8108;
  assign n8110 = n7834 & ~n7913;
  assign n8111 = n8059 & n8110;
  assign n8112 = ~n8059 & ~n8110;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = P3_INSTADDRPOINTER_REG_5_ & ~n8113;
  assign n8115 = ~P3_INSTADDRPOINTER_REG_5_ & n8113;
  assign n8116 = ~n7984 & ~n8115;
  assign n8117 = ~n8114 & n8116;
  assign n8118 = n7982 & ~n7985;
  assign n8119 = n8117 & ~n8118;
  assign n8120 = ~P3_INSTADDRPOINTER_REG_5_ & ~n8113;
  assign n8121 = P3_INSTADDRPOINTER_REG_5_ & n8113;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n7985 & n8122;
  assign n8124 = ~n7982 & ~n7984;
  assign n8125 = n8123 & ~n8124;
  assign n8126 = ~n8119 & ~n8125;
  assign n8127 = n5461 & n8126;
  assign n8128 = n8096 & n8109;
  assign n8129 = ~n8127 & n8128;
  assign n8130 = n8022 & ~n8023;
  assign n8131 = ~n8070 & n8130;
  assign n8132 = n8089 & n8131;
  assign n8133 = n8129 & n8132;
  assign n8134 = n7353 & ~n8133;
  assign n8135 = ~n7999 & ~n8000;
  assign n1690 = n8134 | ~n8135;
  assign n8137 = P3_INSTADDRPOINTER_REG_6_ & n7352;
  assign n8138 = P3_REIP_REG_6_ & n7497;
  assign n8139 = P3_INSTADDRPOINTER_REG_5_ & n8001;
  assign n8140 = ~P3_INSTADDRPOINTER_REG_6_ & n8139;
  assign n8141 = P3_INSTADDRPOINTER_REG_6_ & ~n8139;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = n5618 & ~n8142;
  assign n8144 = n5619_1 & ~n8142;
  assign n8145 = P3_INSTADDRPOINTER_REG_5_ & n8007;
  assign n8146 = ~P3_INSTADDRPOINTER_REG_6_ & n8145;
  assign n8147 = P3_INSTADDRPOINTER_REG_6_ & ~n8145;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = n7361 & ~n8148;
  assign n8150 = P3_INSTADDRPOINTER_REG_5_ & n8013;
  assign n8151 = ~P3_INSTADDRPOINTER_REG_6_ & n8150;
  assign n8152 = P3_INSTADDRPOINTER_REG_6_ & ~n8150;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n7364 & ~n8153;
  assign n8155 = ~n8149 & ~n8154;
  assign n8156 = n5434_1 & ~n8142;
  assign n8157 = n8155 & ~n8156;
  assign n8158 = ~n8143 & ~n8144;
  assign n8159 = n8157 & n8158;
  assign n8160 = ~n5547 & ~n8148;
  assign n8161 = ~P3_INSTADDRPOINTER_REG_5_ & ~n8063;
  assign n8162 = ~n8028 & ~n8161;
  assign n8163 = P3_INSTADDRPOINTER_REG_5_ & n8063;
  assign n8164 = ~n8162 & ~n8163;
  assign n8165 = P3_INSTQUEUE_REG_0__6_ & n7371;
  assign n8166 = P3_INSTQUEUE_REG_1__6_ & n7374;
  assign n8167 = P3_INSTQUEUE_REG_2__6_ & n7377;
  assign n8168 = P3_INSTQUEUE_REG_3__6_ & n7380;
  assign n8169 = ~n8165 & ~n8166;
  assign n8170 = ~n8167 & n8169;
  assign n8171 = ~n8168 & n8170;
  assign n8172 = P3_INSTQUEUE_REG_4__6_ & n7386;
  assign n8173 = P3_INSTQUEUE_REG_5__6_ & n7388;
  assign n8174 = P3_INSTQUEUE_REG_6__6_ & n7390;
  assign n8175 = P3_INSTQUEUE_REG_7__6_ & n7392;
  assign n8176 = ~n8172 & ~n8173;
  assign n8177 = ~n8174 & n8176;
  assign n8178 = ~n8175 & n8177;
  assign n8179 = P3_INSTQUEUE_REG_8__6_ & n7398;
  assign n8180 = P3_INSTQUEUE_REG_9__6_ & n7400;
  assign n8181 = P3_INSTQUEUE_REG_10__6_ & n7402;
  assign n8182 = P3_INSTQUEUE_REG_11__6_ & n7404;
  assign n8183 = ~n8179 & ~n8180;
  assign n8184 = ~n8181 & n8183;
  assign n8185 = ~n8182 & n8184;
  assign n8186 = P3_INSTQUEUE_REG_12__6_ & n7410;
  assign n8187 = P3_INSTQUEUE_REG_13__6_ & n7412;
  assign n8188 = P3_INSTQUEUE_REG_14__6_ & n7414;
  assign n8189 = P3_INSTQUEUE_REG_15__6_ & n7416;
  assign n8190 = ~n8186 & ~n8187;
  assign n8191 = ~n8188 & n8190;
  assign n8192 = ~n8189 & n8191;
  assign n8193 = n8171 & n8178;
  assign n8194 = n8185 & n8193;
  assign n8195 = n8192 & n8194;
  assign n8196 = n8062 & ~n8195;
  assign n8197 = ~n8062 & n8195;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = ~P3_INSTADDRPOINTER_REG_6_ & n8198;
  assign n8200 = P3_INSTADDRPOINTER_REG_6_ & ~n8198;
  assign n8201 = ~n8199 & ~n8200;
  assign n8202 = n8164 & ~n8201;
  assign n8203 = ~n8164 & n8201;
  assign n8204 = ~n8202 & ~n8203;
  assign n8205 = n7458 & ~n8204;
  assign n8206 = n5657 & ~n8148;
  assign n8207 = n5500 & ~n8148;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = ~n8078 & ~n8081;
  assign n8210 = P3_INSTADDRPOINTER_REG_5_ & ~n8078;
  assign n8211 = P3_INSTADDRPOINTER_REG_5_ & ~n8081;
  assign n8212 = ~n8209 & ~n8210;
  assign n8213 = ~n8211 & n8212;
  assign n8214 = n7938 & ~n8059;
  assign n8215 = n8195 & n8214;
  assign n8216 = ~n8195 & ~n8214;
  assign n8217 = ~n8215 & ~n8216;
  assign n8218 = ~P3_INSTADDRPOINTER_REG_6_ & ~n8217;
  assign n8219 = P3_INSTADDRPOINTER_REG_6_ & n8217;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = n8213 & ~n8220;
  assign n8222 = ~n8213 & n8220;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = n7460 & ~n8223;
  assign n8225 = n8208 & ~n8224;
  assign n8226 = n7477 & ~n8148;
  assign n8227 = n7470 & ~n8148;
  assign n8228 = n7466 & ~n8148;
  assign n8229 = n5504_1 & ~n8148;
  assign n8230 = ~n8226 & ~n8227;
  assign n8231 = ~n8228 & n8230;
  assign n8232 = ~n8229 & n8231;
  assign n8233 = n5360 & ~n8142;
  assign n8234 = n5438 & ~n8142;
  assign n8235 = n5442 & ~n8142;
  assign n8236 = P3_INSTADDRPOINTER_REG_5_ & n8100;
  assign n8237 = ~P3_INSTADDRPOINTER_REG_6_ & n8236;
  assign n8238 = P3_INSTADDRPOINTER_REG_6_ & ~n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = n5458 & ~n8239;
  assign n8241 = n5450 & ~n8239;
  assign n8242 = ~n8233 & ~n8234;
  assign n8243 = ~n8235 & n8242;
  assign n8244 = ~n8240 & n8243;
  assign n8245 = ~n8241 & n8244;
  assign n8246 = n7985 & ~n8113;
  assign n8247 = ~n7985 & n8113;
  assign n8248 = P3_INSTADDRPOINTER_REG_5_ & ~n8247;
  assign n8249 = ~n8246 & ~n8248;
  assign n8250 = ~n7982 & n8116;
  assign n8251 = n8249 & ~n8250;
  assign n8252 = ~n8059 & n8110;
  assign n8253 = n8195 & n8252;
  assign n8254 = ~n8195 & ~n8252;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = ~P3_INSTADDRPOINTER_REG_6_ & ~n8255;
  assign n8257 = P3_INSTADDRPOINTER_REG_6_ & n8255;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = n8251 & ~n8258;
  assign n8260 = ~n8251 & n8258;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = n5461 & ~n8261;
  assign n8263 = n8232 & n8245;
  assign n8264 = ~n8262 & n8263;
  assign n8265 = n8159 & ~n8160;
  assign n8266 = ~n8205 & n8265;
  assign n8267 = n8225 & n8266;
  assign n8268 = n8264 & n8267;
  assign n8269 = n7353 & ~n8268;
  assign n8270 = ~n8137 & ~n8138;
  assign n1695 = n8269 | ~n8270;
  assign n8272 = P3_INSTADDRPOINTER_REG_7_ & n7352;
  assign n8273 = P3_REIP_REG_7_ & n7497;
  assign n8274 = P3_INSTADDRPOINTER_REG_6_ & n8139;
  assign n8275 = ~P3_INSTADDRPOINTER_REG_7_ & n8274;
  assign n8276 = P3_INSTADDRPOINTER_REG_7_ & ~n8274;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = n5618 & ~n8277;
  assign n8279 = n5619_1 & ~n8277;
  assign n8280 = P3_INSTADDRPOINTER_REG_6_ & n8145;
  assign n8281 = ~P3_INSTADDRPOINTER_REG_7_ & n8280;
  assign n8282 = P3_INSTADDRPOINTER_REG_7_ & ~n8280;
  assign n8283 = ~n8281 & ~n8282;
  assign n8284 = n7361 & ~n8283;
  assign n8285 = P3_INSTADDRPOINTER_REG_5_ & P3_INSTADDRPOINTER_REG_6_;
  assign n8286 = n8013 & n8285;
  assign n8287 = P3_INSTADDRPOINTER_REG_7_ & ~n8286;
  assign n8288 = ~P3_INSTADDRPOINTER_REG_7_ & n8286;
  assign n8289 = ~n8287 & ~n8288;
  assign n8290 = n7364 & ~n8289;
  assign n8291 = ~n8284 & ~n8290;
  assign n8292 = n5434_1 & ~n8277;
  assign n8293 = n8291 & ~n8292;
  assign n8294 = ~n8278 & ~n8279;
  assign n8295 = n8293 & n8294;
  assign n8296 = ~n5547 & ~n8283;
  assign n8297 = P3_INSTADDRPOINTER_REG_6_ & n8198;
  assign n8298 = ~P3_INSTADDRPOINTER_REG_6_ & ~n8198;
  assign n8299 = ~n8164 & ~n8298;
  assign n8300 = ~n8297 & ~n8299;
  assign n8301 = n7457 & ~n8196;
  assign n8302 = ~n7457 & ~n8195;
  assign n8303 = n8062 & n8302;
  assign n8304 = ~n8301 & ~n8303;
  assign n8305 = ~P3_INSTADDRPOINTER_REG_7_ & n8304;
  assign n8306 = P3_INSTADDRPOINTER_REG_7_ & ~n8304;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = n8300 & ~n8307;
  assign n8309 = ~n8300 & n8307;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = n7458 & ~n8310;
  assign n8312 = n5657 & ~n8283;
  assign n8313 = n5500 & ~n8283;
  assign n8314 = ~n8312 & ~n8313;
  assign n8315 = P3_INSTADDRPOINTER_REG_6_ & ~n8217;
  assign n8316 = ~P3_INSTADDRPOINTER_REG_6_ & n8217;
  assign n8317 = ~n8213 & ~n8316;
  assign n8318 = ~n8315 & ~n8317;
  assign n8319 = ~n8195 & n8214;
  assign n8320 = n7457 & n8319;
  assign n8321 = ~n7457 & ~n8319;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = ~P3_INSTADDRPOINTER_REG_7_ & ~n8322;
  assign n8324 = P3_INSTADDRPOINTER_REG_7_ & n8322;
  assign n8325 = ~n8323 & ~n8324;
  assign n8326 = n8318 & ~n8325;
  assign n8327 = ~n8318 & n8325;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = n7460 & ~n8328;
  assign n8330 = n8314 & ~n8329;
  assign n8331 = n7477 & ~n8283;
  assign n8332 = n7470 & ~n8283;
  assign n8333 = n7466 & ~n8283;
  assign n8334 = n5504_1 & ~n8283;
  assign n8335 = ~n8331 & ~n8332;
  assign n8336 = ~n8333 & n8335;
  assign n8337 = ~n8334 & n8336;
  assign n8338 = n5360 & ~n8277;
  assign n8339 = n5438 & ~n8277;
  assign n8340 = n5442 & ~n8277;
  assign n8341 = P3_INSTADDRPOINTER_REG_6_ & n8236;
  assign n8342 = ~P3_INSTADDRPOINTER_REG_7_ & n8341;
  assign n8343 = P3_INSTADDRPOINTER_REG_7_ & ~n8341;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = n5458 & ~n8344;
  assign n8346 = n5450 & ~n8344;
  assign n8347 = ~n8338 & ~n8339;
  assign n8348 = ~n8340 & n8347;
  assign n8349 = ~n8345 & n8348;
  assign n8350 = ~n8346 & n8349;
  assign n8351 = P3_INSTADDRPOINTER_REG_6_ & ~n8255;
  assign n8352 = ~P3_INSTADDRPOINTER_REG_6_ & n8255;
  assign n8353 = ~n8251 & ~n8352;
  assign n8354 = ~n8351 & ~n8353;
  assign n8355 = ~n8195 & n8252;
  assign n8356 = n7457 & n8355;
  assign n8357 = ~n7457 & ~n8355;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = ~P3_INSTADDRPOINTER_REG_7_ & ~n8358;
  assign n8360 = P3_INSTADDRPOINTER_REG_7_ & n8358;
  assign n8361 = ~n8359 & ~n8360;
  assign n8362 = n8354 & ~n8361;
  assign n8363 = ~n8354 & n8361;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n5461 & ~n8364;
  assign n8366 = n8337 & n8350;
  assign n8367 = ~n8365 & n8366;
  assign n8368 = n8295 & ~n8296;
  assign n8369 = ~n8311 & n8368;
  assign n8370 = n8330 & n8369;
  assign n8371 = n8367 & n8370;
  assign n8372 = n7353 & ~n8371;
  assign n8373 = ~n8272 & ~n8273;
  assign n1700 = n8372 | ~n8373;
  assign n8375 = P3_INSTADDRPOINTER_REG_8_ & n7352;
  assign n8376 = P3_REIP_REG_8_ & n7497;
  assign n8377 = P3_INSTADDRPOINTER_REG_7_ & n8274;
  assign n8378 = ~P3_INSTADDRPOINTER_REG_8_ & n8377;
  assign n8379 = P3_INSTADDRPOINTER_REG_8_ & ~n8377;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = n5618 & ~n8380;
  assign n8382 = n5619_1 & ~n8380;
  assign n8383 = n5434_1 & ~n8380;
  assign n8384 = P3_INSTADDRPOINTER_REG_7_ & n8286;
  assign n8385 = ~P3_INSTADDRPOINTER_REG_8_ & n8384;
  assign n8386 = P3_INSTADDRPOINTER_REG_8_ & ~n8384;
  assign n8387 = ~n8385 & ~n8386;
  assign n8388 = n7364 & ~n8387;
  assign n8389 = P3_INSTADDRPOINTER_REG_7_ & n8280;
  assign n8390 = ~P3_INSTADDRPOINTER_REG_8_ & n8389;
  assign n8391 = P3_INSTADDRPOINTER_REG_8_ & ~n8389;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = n7361 & ~n8392;
  assign n8394 = ~n8383 & ~n8388;
  assign n8395 = ~n8393 & n8394;
  assign n8396 = ~n8381 & ~n8382;
  assign n8397 = n8395 & n8396;
  assign n8398 = ~n5547 & ~n8392;
  assign n8399 = ~P3_INSTADDRPOINTER_REG_7_ & ~n8304;
  assign n8400 = ~n8300 & ~n8399;
  assign n8401 = P3_INSTADDRPOINTER_REG_7_ & n8304;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = P3_INSTADDRPOINTER_REG_8_ & n8303;
  assign n8404 = ~P3_INSTADDRPOINTER_REG_8_ & ~n8303;
  assign n8405 = ~n8403 & ~n8404;
  assign n8406 = n8402 & ~n8405;
  assign n8407 = ~n8402 & n8405;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = n7458 & ~n8408;
  assign n8410 = n5657 & ~n8392;
  assign n8411 = n5500 & ~n8392;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = ~n8318 & ~n8322;
  assign n8414 = P3_INSTADDRPOINTER_REG_7_ & ~n8318;
  assign n8415 = P3_INSTADDRPOINTER_REG_7_ & ~n8322;
  assign n8416 = ~n8413 & ~n8414;
  assign n8417 = ~n8415 & n8416;
  assign n8418 = n8214 & n8302;
  assign n8419 = ~P3_INSTADDRPOINTER_REG_8_ & n8418;
  assign n8420 = P3_INSTADDRPOINTER_REG_8_ & ~n8418;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = n8417 & ~n8421;
  assign n8423 = ~n8417 & n8421;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = n7460 & ~n8424;
  assign n8426 = n8412 & ~n8425;
  assign n8427 = n7477 & ~n8392;
  assign n8428 = n5504_1 & ~n8392;
  assign n8429 = n7466 & ~n8392;
  assign n8430 = n7470 & ~n8392;
  assign n8431 = ~n8427 & ~n8428;
  assign n8432 = ~n8429 & n8431;
  assign n8433 = ~n8430 & n8432;
  assign n8434 = n5360 & ~n8380;
  assign n8435 = n5438 & ~n8380;
  assign n8436 = n5442 & ~n8380;
  assign n8437 = P3_INSTADDRPOINTER_REG_7_ & n8341;
  assign n8438 = ~P3_INSTADDRPOINTER_REG_8_ & n8437;
  assign n8439 = P3_INSTADDRPOINTER_REG_8_ & ~n8437;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = n5458 & ~n8440;
  assign n8442 = n5450 & ~n8440;
  assign n8443 = ~n8434 & ~n8435;
  assign n8444 = ~n8436 & n8443;
  assign n8445 = ~n8441 & n8444;
  assign n8446 = ~n8442 & n8445;
  assign n8447 = ~n8354 & ~n8358;
  assign n8448 = P3_INSTADDRPOINTER_REG_7_ & ~n8354;
  assign n8449 = P3_INSTADDRPOINTER_REG_7_ & ~n8358;
  assign n8450 = ~n8447 & ~n8448;
  assign n8451 = ~n8449 & n8450;
  assign n8452 = n8252 & n8302;
  assign n8453 = ~P3_INSTADDRPOINTER_REG_8_ & n8452;
  assign n8454 = P3_INSTADDRPOINTER_REG_8_ & ~n8452;
  assign n8455 = ~n8453 & ~n8454;
  assign n8456 = n8451 & ~n8455;
  assign n8457 = ~n8451 & n8455;
  assign n8458 = ~n8456 & ~n8457;
  assign n8459 = n5461 & ~n8458;
  assign n8460 = n8433 & n8446;
  assign n8461 = ~n8459 & n8460;
  assign n8462 = n8397 & ~n8398;
  assign n8463 = ~n8409 & n8462;
  assign n8464 = n8426 & n8463;
  assign n8465 = n8461 & n8464;
  assign n8466 = n7353 & ~n8465;
  assign n8467 = ~n8375 & ~n8376;
  assign n1705 = n8466 | ~n8467;
  assign n8469 = P3_INSTADDRPOINTER_REG_9_ & n7352;
  assign n8470 = P3_REIP_REG_9_ & n7497;
  assign n8471 = P3_INSTADDRPOINTER_REG_8_ & n8377;
  assign n8472 = ~P3_INSTADDRPOINTER_REG_9_ & n8471;
  assign n8473 = P3_INSTADDRPOINTER_REG_9_ & ~n8471;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = n5618 & ~n8474;
  assign n8476 = n5619_1 & ~n8474;
  assign n8477 = P3_INSTADDRPOINTER_REG_8_ & n8389;
  assign n8478 = ~P3_INSTADDRPOINTER_REG_9_ & n8477;
  assign n8479 = P3_INSTADDRPOINTER_REG_9_ & ~n8477;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = n7361 & ~n8480;
  assign n8482 = n5434_1 & ~n8474;
  assign n8483 = P3_INSTADDRPOINTER_REG_7_ & P3_INSTADDRPOINTER_REG_8_;
  assign n8484 = n8286 & n8483;
  assign n8485 = P3_INSTADDRPOINTER_REG_9_ & ~n8484;
  assign n8486 = ~P3_INSTADDRPOINTER_REG_9_ & n8484;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = n7364 & ~n8487;
  assign n8489 = ~n8482 & ~n8488;
  assign n8490 = ~n8475 & ~n8476;
  assign n8491 = ~n8481 & n8490;
  assign n8492 = n8489 & n8491;
  assign n8493 = ~n5547 & ~n8480;
  assign n8494 = P3_INSTADDRPOINTER_REG_8_ & ~n8402;
  assign n8495 = ~n8303 & ~n8402;
  assign n8496 = P3_INSTADDRPOINTER_REG_8_ & ~n8303;
  assign n8497 = ~n8494 & ~n8495;
  assign n8498 = ~n8496 & n8497;
  assign n8499 = P3_INSTADDRPOINTER_REG_9_ & n8303;
  assign n8500 = ~P3_INSTADDRPOINTER_REG_9_ & ~n8303;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = n8498 & ~n8501;
  assign n8503 = P3_INSTADDRPOINTER_REG_9_ & ~n8303;
  assign n8504 = ~P3_INSTADDRPOINTER_REG_9_ & n8303;
  assign n8505 = ~n8503 & ~n8504;
  assign n8506 = ~n8498 & ~n8505;
  assign n8507 = ~n8502 & ~n8506;
  assign n8508 = n7458 & ~n8507;
  assign n8509 = n5657 & ~n8480;
  assign n8510 = n5500 & ~n8480;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = P3_INSTADDRPOINTER_REG_8_ & n8418;
  assign n8513 = ~P3_INSTADDRPOINTER_REG_8_ & ~n8418;
  assign n8514 = ~n8417 & ~n8513;
  assign n8515 = ~n8512 & ~n8514;
  assign n8516 = ~P3_INSTADDRPOINTER_REG_9_ & n8515;
  assign n8517 = P3_INSTADDRPOINTER_REG_9_ & ~n8515;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = n7460 & n8518;
  assign n8520 = n8511 & ~n8519;
  assign n8521 = n7477 & ~n8480;
  assign n8522 = n5504_1 & ~n8480;
  assign n8523 = n7466 & ~n8480;
  assign n8524 = n7470 & ~n8480;
  assign n8525 = ~n8521 & ~n8522;
  assign n8526 = ~n8523 & n8525;
  assign n8527 = ~n8524 & n8526;
  assign n8528 = n5360 & ~n8474;
  assign n8529 = n5438 & ~n8474;
  assign n8530 = n5442 & ~n8474;
  assign n8531 = P3_INSTADDRPOINTER_REG_8_ & n8437;
  assign n8532 = ~P3_INSTADDRPOINTER_REG_9_ & n8531;
  assign n8533 = P3_INSTADDRPOINTER_REG_9_ & ~n8531;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = n5458 & ~n8534;
  assign n8536 = n5450 & ~n8534;
  assign n8537 = ~n8528 & ~n8529;
  assign n8538 = ~n8530 & n8537;
  assign n8539 = ~n8535 & n8538;
  assign n8540 = ~n8536 & n8539;
  assign n8541 = P3_INSTADDRPOINTER_REG_8_ & n8452;
  assign n8542 = ~P3_INSTADDRPOINTER_REG_8_ & ~n8452;
  assign n8543 = ~n8451 & ~n8542;
  assign n8544 = ~n8541 & ~n8543;
  assign n8545 = ~P3_INSTADDRPOINTER_REG_9_ & n8544;
  assign n8546 = P3_INSTADDRPOINTER_REG_9_ & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n5461 & n8547;
  assign n8549 = n8527 & n8540;
  assign n8550 = ~n8548 & n8549;
  assign n8551 = n8492 & ~n8493;
  assign n8552 = ~n8508 & n8551;
  assign n8553 = n8520 & n8552;
  assign n8554 = n8550 & n8553;
  assign n8555 = n7353 & ~n8554;
  assign n8556 = ~n8469 & ~n8470;
  assign n1710 = n8555 | ~n8556;
  assign n8558 = P3_INSTADDRPOINTER_REG_10_ & n7352;
  assign n8559 = P3_REIP_REG_10_ & n7497;
  assign n8560 = P3_INSTADDRPOINTER_REG_9_ & n8477;
  assign n8561 = ~P3_INSTADDRPOINTER_REG_10_ & n8560;
  assign n8562 = P3_INSTADDRPOINTER_REG_10_ & ~n8560;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = ~n5547 & ~n8563;
  assign n8565 = P3_INSTADDRPOINTER_REG_9_ & n8471;
  assign n8566 = ~P3_INSTADDRPOINTER_REG_10_ & n8565;
  assign n8567 = P3_INSTADDRPOINTER_REG_10_ & ~n8565;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = n5618 & ~n8568;
  assign n8570 = n5619_1 & ~n8568;
  assign n8571 = n7361 & ~n8563;
  assign n8572 = n5434_1 & ~n8568;
  assign n8573 = P3_INSTADDRPOINTER_REG_9_ & n8484;
  assign n8574 = ~P3_INSTADDRPOINTER_REG_10_ & n8573;
  assign n8575 = P3_INSTADDRPOINTER_REG_10_ & ~n8573;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = n7364 & ~n8576;
  assign n8578 = ~n8572 & ~n8577;
  assign n8579 = ~n8569 & ~n8570;
  assign n8580 = ~n8571 & n8579;
  assign n8581 = n8578 & n8580;
  assign n8582 = ~P3_INSTADDRPOINTER_REG_10_ & ~n8517;
  assign n8583 = P3_INSTADDRPOINTER_REG_9_ & P3_INSTADDRPOINTER_REG_10_;
  assign n8584 = ~n8515 & n8583;
  assign n8585 = ~n8582 & ~n8584;
  assign n8586 = n7460 & n8585;
  assign n8587 = n7477 & ~n8563;
  assign n8588 = n5504_1 & ~n8563;
  assign n8589 = n7466 & ~n8563;
  assign n8590 = n7470 & ~n8563;
  assign n8591 = ~n8587 & ~n8588;
  assign n8592 = ~n8589 & n8591;
  assign n8593 = ~n8590 & n8592;
  assign n8594 = n5360 & ~n8568;
  assign n8595 = n5438 & ~n8568;
  assign n8596 = n5442 & ~n8568;
  assign n8597 = P3_INSTADDRPOINTER_REG_9_ & n8531;
  assign n8598 = ~P3_INSTADDRPOINTER_REG_10_ & n8597;
  assign n8599 = P3_INSTADDRPOINTER_REG_10_ & ~n8597;
  assign n8600 = ~n8598 & ~n8599;
  assign n8601 = n5458 & ~n8600;
  assign n8602 = n5450 & ~n8600;
  assign n8603 = ~n8594 & ~n8595;
  assign n8604 = ~n8596 & n8603;
  assign n8605 = ~n8601 & n8604;
  assign n8606 = ~n8602 & n8605;
  assign n8607 = ~P3_INSTADDRPOINTER_REG_10_ & ~n8546;
  assign n8608 = ~n8544 & n8583;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = n5461 & n8609;
  assign n8611 = n8593 & n8606;
  assign n8612 = ~n8610 & n8611;
  assign n8613 = n5657 & ~n8563;
  assign n8614 = n5500 & ~n8563;
  assign n8615 = ~n8613 & ~n8614;
  assign n8616 = ~n8498 & ~n8504;
  assign n8617 = ~n8503 & ~n8616;
  assign n8618 = ~P3_INSTADDRPOINTER_REG_10_ & ~n8303;
  assign n8619 = P3_INSTADDRPOINTER_REG_10_ & n8303;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = n8617 & ~n8620;
  assign n8622 = P3_INSTADDRPOINTER_REG_10_ & ~n8303;
  assign n8623 = ~P3_INSTADDRPOINTER_REG_10_ & n8303;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~n8617 & ~n8624;
  assign n8626 = ~n8621 & ~n8625;
  assign n8627 = n7458 & ~n8626;
  assign n8628 = n8615 & ~n8627;
  assign n8629 = ~n8564 & n8581;
  assign n8630 = ~n8586 & n8629;
  assign n8631 = n8612 & n8630;
  assign n8632 = n8628 & n8631;
  assign n8633 = n7353 & ~n8632;
  assign n8634 = ~n8558 & ~n8559;
  assign n1715 = n8633 | ~n8634;
  assign n8636 = P3_INSTADDRPOINTER_REG_11_ & n7352;
  assign n8637 = P3_REIP_REG_11_ & n7497;
  assign n8638 = P3_INSTADDRPOINTER_REG_10_ & n8560;
  assign n8639 = ~P3_INSTADDRPOINTER_REG_11_ & n8638;
  assign n8640 = P3_INSTADDRPOINTER_REG_11_ & ~n8638;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = ~n5547 & ~n8641;
  assign n8643 = P3_INSTADDRPOINTER_REG_10_ & n8565;
  assign n8644 = ~P3_INSTADDRPOINTER_REG_11_ & n8643;
  assign n8645 = P3_INSTADDRPOINTER_REG_11_ & ~n8643;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = n5618 & ~n8646;
  assign n8648 = n5619_1 & ~n8646;
  assign n8649 = n7361 & ~n8641;
  assign n8650 = n5434_1 & ~n8646;
  assign n8651 = n8484 & n8583;
  assign n8652 = P3_INSTADDRPOINTER_REG_11_ & ~n8651;
  assign n8653 = ~P3_INSTADDRPOINTER_REG_11_ & n8651;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = n7364 & ~n8654;
  assign n8656 = ~n8650 & ~n8655;
  assign n8657 = ~n8647 & ~n8648;
  assign n8658 = ~n8649 & n8657;
  assign n8659 = n8656 & n8658;
  assign n8660 = P3_INSTADDRPOINTER_REG_11_ & ~n8584;
  assign n8661 = ~P3_INSTADDRPOINTER_REG_11_ & n8584;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = n7460 & ~n8662;
  assign n8664 = n5657 & ~n8641;
  assign n8665 = n5500 & ~n8641;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~n8504 & ~n8623;
  assign n8668 = ~n8498 & n8667;
  assign n8669 = ~n8503 & ~n8622;
  assign n8670 = ~n8668 & n8669;
  assign n8671 = ~P3_INSTADDRPOINTER_REG_11_ & ~n8303;
  assign n8672 = P3_INSTADDRPOINTER_REG_11_ & n8303;
  assign n8673 = ~n8671 & ~n8672;
  assign n8674 = n8670 & ~n8673;
  assign n8675 = ~n8670 & n8673;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = n7458 & ~n8676;
  assign n8678 = n8666 & ~n8677;
  assign n8679 = n7477 & ~n8641;
  assign n8680 = n5504_1 & ~n8641;
  assign n8681 = n7466 & ~n8641;
  assign n8682 = n7470 & ~n8641;
  assign n8683 = ~n8679 & ~n8680;
  assign n8684 = ~n8681 & n8683;
  assign n8685 = ~n8682 & n8684;
  assign n8686 = n5360 & ~n8646;
  assign n8687 = n5438 & ~n8646;
  assign n8688 = n5442 & ~n8646;
  assign n8689 = P3_INSTADDRPOINTER_REG_10_ & n8597;
  assign n8690 = ~P3_INSTADDRPOINTER_REG_11_ & n8689;
  assign n8691 = P3_INSTADDRPOINTER_REG_11_ & ~n8689;
  assign n8692 = ~n8690 & ~n8691;
  assign n8693 = n5458 & ~n8692;
  assign n8694 = n5450 & ~n8692;
  assign n8695 = ~n8686 & ~n8687;
  assign n8696 = ~n8688 & n8695;
  assign n8697 = ~n8693 & n8696;
  assign n8698 = ~n8694 & n8697;
  assign n8699 = P3_INSTADDRPOINTER_REG_11_ & ~n8608;
  assign n8700 = ~P3_INSTADDRPOINTER_REG_11_ & n8608;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = n5461 & ~n8701;
  assign n8703 = n8685 & n8698;
  assign n8704 = ~n8702 & n8703;
  assign n8705 = ~n8642 & n8659;
  assign n8706 = ~n8663 & n8705;
  assign n8707 = n8678 & n8706;
  assign n8708 = n8704 & n8707;
  assign n8709 = n7353 & ~n8708;
  assign n8710 = ~n8636 & ~n8637;
  assign n1720 = n8709 | ~n8710;
  assign n8712 = P3_INSTADDRPOINTER_REG_12_ & n7352;
  assign n8713 = P3_REIP_REG_12_ & n7497;
  assign n8714 = P3_INSTADDRPOINTER_REG_11_ & n8643;
  assign n8715 = ~P3_INSTADDRPOINTER_REG_12_ & n8714;
  assign n8716 = P3_INSTADDRPOINTER_REG_12_ & ~n8714;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = n5618 & ~n8717;
  assign n8719 = n5619_1 & ~n8717;
  assign n8720 = P3_INSTADDRPOINTER_REG_11_ & n8638;
  assign n8721 = ~P3_INSTADDRPOINTER_REG_12_ & n8720;
  assign n8722 = P3_INSTADDRPOINTER_REG_12_ & ~n8720;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = n7361 & ~n8723;
  assign n8725 = n5434_1 & ~n8717;
  assign n8726 = P3_INSTADDRPOINTER_REG_11_ & n8651;
  assign n8727 = ~P3_INSTADDRPOINTER_REG_12_ & n8726;
  assign n8728 = P3_INSTADDRPOINTER_REG_12_ & ~n8726;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = n7364 & ~n8729;
  assign n8731 = ~n8725 & ~n8730;
  assign n8732 = ~n8718 & ~n8719;
  assign n8733 = ~n8724 & n8732;
  assign n8734 = n8731 & n8733;
  assign n8735 = ~n5547 & ~n8723;
  assign n8736 = ~P3_INSTADDRPOINTER_REG_12_ & ~n8303;
  assign n8737 = P3_INSTADDRPOINTER_REG_12_ & n8303;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = ~P3_INSTADDRPOINTER_REG_11_ & n8303;
  assign n8740 = n8667 & ~n8739;
  assign n8741 = ~n8498 & n8740;
  assign n8742 = P3_INSTADDRPOINTER_REG_11_ & ~n8303;
  assign n8743 = n8669 & ~n8742;
  assign n8744 = ~n8741 & n8743;
  assign n8745 = ~n8738 & n8744;
  assign n8746 = ~P3_INSTADDRPOINTER_REG_12_ & n8303;
  assign n8747 = P3_INSTADDRPOINTER_REG_12_ & ~n8303;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~n8744 & ~n8748;
  assign n8750 = ~n8745 & ~n8749;
  assign n8751 = n7458 & ~n8750;
  assign n8752 = n5657 & ~n8723;
  assign n8753 = n5500 & ~n8723;
  assign n8754 = ~n8752 & ~n8753;
  assign n8755 = P3_INSTADDRPOINTER_REG_11_ & n8584;
  assign n8756 = ~P3_INSTADDRPOINTER_REG_12_ & ~n8755;
  assign n8757 = P3_INSTADDRPOINTER_REG_11_ & P3_INSTADDRPOINTER_REG_12_;
  assign n8758 = n8584 & n8757;
  assign n8759 = ~n8756 & ~n8758;
  assign n8760 = n7460 & n8759;
  assign n8761 = n8754 & ~n8760;
  assign n8762 = n7477 & ~n8723;
  assign n8763 = n5504_1 & ~n8723;
  assign n8764 = n7466 & ~n8723;
  assign n8765 = n7470 & ~n8723;
  assign n8766 = ~n8762 & ~n8763;
  assign n8767 = ~n8764 & n8766;
  assign n8768 = ~n8765 & n8767;
  assign n8769 = n5360 & ~n8717;
  assign n8770 = n5438 & ~n8717;
  assign n8771 = n5442 & ~n8717;
  assign n8772 = P3_INSTADDRPOINTER_REG_11_ & n8689;
  assign n8773 = ~P3_INSTADDRPOINTER_REG_12_ & n8772;
  assign n8774 = P3_INSTADDRPOINTER_REG_12_ & ~n8772;
  assign n8775 = ~n8773 & ~n8774;
  assign n8776 = n5458 & ~n8775;
  assign n8777 = n5450 & ~n8775;
  assign n8778 = ~n8769 & ~n8770;
  assign n8779 = ~n8771 & n8778;
  assign n8780 = ~n8776 & n8779;
  assign n8781 = ~n8777 & n8780;
  assign n8782 = P3_INSTADDRPOINTER_REG_11_ & n8608;
  assign n8783 = ~P3_INSTADDRPOINTER_REG_12_ & ~n8782;
  assign n8784 = n8608 & n8757;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = n5461 & n8785;
  assign n8787 = n8768 & n8781;
  assign n8788 = ~n8786 & n8787;
  assign n8789 = n8734 & ~n8735;
  assign n8790 = ~n8751 & n8789;
  assign n8791 = n8761 & n8790;
  assign n8792 = n8788 & n8791;
  assign n8793 = n7353 & ~n8792;
  assign n8794 = ~n8712 & ~n8713;
  assign n1725 = n8793 | ~n8794;
  assign n8796 = P3_INSTADDRPOINTER_REG_13_ & n7352;
  assign n8797 = P3_REIP_REG_13_ & n7497;
  assign n8798 = P3_INSTADDRPOINTER_REG_12_ & n8714;
  assign n8799 = ~P3_INSTADDRPOINTER_REG_13_ & n8798;
  assign n8800 = P3_INSTADDRPOINTER_REG_13_ & ~n8798;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = n5618 & ~n8801;
  assign n8803 = n5619_1 & ~n8801;
  assign n8804 = P3_INSTADDRPOINTER_REG_12_ & n8720;
  assign n8805 = ~P3_INSTADDRPOINTER_REG_13_ & n8804;
  assign n8806 = P3_INSTADDRPOINTER_REG_13_ & ~n8804;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = n7361 & ~n8807;
  assign n8809 = n5434_1 & ~n8801;
  assign n8810 = n8651 & n8757;
  assign n8811 = P3_INSTADDRPOINTER_REG_13_ & ~n8810;
  assign n8812 = ~P3_INSTADDRPOINTER_REG_13_ & n8810;
  assign n8813 = ~n8811 & ~n8812;
  assign n8814 = n7364 & ~n8813;
  assign n8815 = ~n8809 & ~n8814;
  assign n8816 = ~n8802 & ~n8803;
  assign n8817 = ~n8808 & n8816;
  assign n8818 = n8815 & n8817;
  assign n8819 = ~n5547 & ~n8807;
  assign n8820 = P3_INSTADDRPOINTER_REG_13_ & ~n8303;
  assign n8821 = P3_INSTADDRPOINTER_REG_12_ & P3_INSTADDRPOINTER_REG_13_;
  assign n8822 = n8303 & ~n8821;
  assign n8823 = ~n8820 & ~n8822;
  assign n8824 = n8744 & ~n8747;
  assign n8825 = n8823 & ~n8824;
  assign n8826 = ~P3_INSTADDRPOINTER_REG_13_ & ~n8303;
  assign n8827 = P3_INSTADDRPOINTER_REG_13_ & n8303;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = ~n8747 & n8828;
  assign n8830 = ~n8744 & ~n8746;
  assign n8831 = n8829 & ~n8830;
  assign n8832 = ~n8825 & ~n8831;
  assign n8833 = n7458 & n8832;
  assign n8834 = n5657 & ~n8807;
  assign n8835 = n5500 & ~n8807;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = ~P3_INSTADDRPOINTER_REG_13_ & ~n8758;
  assign n8838 = P3_INSTADDRPOINTER_REG_13_ & n8758;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = n7460 & n8839;
  assign n8841 = n8836 & ~n8840;
  assign n8842 = n7477 & ~n8807;
  assign n8843 = n5504_1 & ~n8807;
  assign n8844 = n7466 & ~n8807;
  assign n8845 = n7470 & ~n8807;
  assign n8846 = ~n8842 & ~n8843;
  assign n8847 = ~n8844 & n8846;
  assign n8848 = ~n8845 & n8847;
  assign n8849 = n5360 & ~n8801;
  assign n8850 = n5438 & ~n8801;
  assign n8851 = n5442 & ~n8801;
  assign n8852 = P3_INSTADDRPOINTER_REG_12_ & n8772;
  assign n8853 = ~P3_INSTADDRPOINTER_REG_13_ & n8852;
  assign n8854 = P3_INSTADDRPOINTER_REG_13_ & ~n8852;
  assign n8855 = ~n8853 & ~n8854;
  assign n8856 = n5458 & ~n8855;
  assign n8857 = n5450 & ~n8855;
  assign n8858 = ~n8849 & ~n8850;
  assign n8859 = ~n8851 & n8858;
  assign n8860 = ~n8856 & n8859;
  assign n8861 = ~n8857 & n8860;
  assign n8862 = ~P3_INSTADDRPOINTER_REG_13_ & ~n8784;
  assign n8863 = P3_INSTADDRPOINTER_REG_13_ & n8784;
  assign n8864 = ~n8862 & ~n8863;
  assign n8865 = n5461 & n8864;
  assign n8866 = n8848 & n8861;
  assign n8867 = ~n8865 & n8866;
  assign n8868 = n8818 & ~n8819;
  assign n8869 = ~n8833 & n8868;
  assign n8870 = n8841 & n8869;
  assign n8871 = n8867 & n8870;
  assign n8872 = n7353 & ~n8871;
  assign n8873 = ~n8796 & ~n8797;
  assign n1730 = n8872 | ~n8873;
  assign n8875 = P3_INSTADDRPOINTER_REG_14_ & n7352;
  assign n8876 = P3_REIP_REG_14_ & n7497;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = P3_INSTADDRPOINTER_REG_13_ & n8804;
  assign n8879 = ~P3_INSTADDRPOINTER_REG_14_ & n8878;
  assign n8880 = P3_INSTADDRPOINTER_REG_14_ & ~n8878;
  assign n8881 = ~n8879 & ~n8880;
  assign n8882 = n7477 & ~n8881;
  assign n8883 = n5504_1 & ~n8881;
  assign n8884 = n7466 & ~n8881;
  assign n8885 = n7470 & ~n8881;
  assign n8886 = ~n8882 & ~n8883;
  assign n8887 = ~n8884 & n8886;
  assign n8888 = ~n8885 & n8887;
  assign n8889 = P3_INSTADDRPOINTER_REG_13_ & n8798;
  assign n8890 = ~P3_INSTADDRPOINTER_REG_14_ & n8889;
  assign n8891 = P3_INSTADDRPOINTER_REG_14_ & ~n8889;
  assign n8892 = ~n8890 & ~n8891;
  assign n8893 = n5360 & ~n8892;
  assign n8894 = n5438 & ~n8892;
  assign n8895 = n5442 & ~n8892;
  assign n8896 = P3_INSTADDRPOINTER_REG_13_ & n8852;
  assign n8897 = ~P3_INSTADDRPOINTER_REG_14_ & n8896;
  assign n8898 = P3_INSTADDRPOINTER_REG_14_ & ~n8896;
  assign n8899 = ~n8897 & ~n8898;
  assign n8900 = n5458 & ~n8899;
  assign n8901 = n5450 & ~n8899;
  assign n8902 = ~n8893 & ~n8894;
  assign n8903 = ~n8895 & n8902;
  assign n8904 = ~n8900 & n8903;
  assign n8905 = ~n8901 & n8904;
  assign n8906 = ~P3_INSTADDRPOINTER_REG_14_ & n8863;
  assign n8907 = P3_INSTADDRPOINTER_REG_14_ & ~n8863;
  assign n8908 = ~n8906 & ~n8907;
  assign n8909 = n5461 & ~n8908;
  assign n8910 = n8888 & n8905;
  assign n8911 = ~n8909 & n8910;
  assign n8912 = n5657 & ~n8881;
  assign n8913 = n5500 & ~n8881;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = ~n5547 & ~n8881;
  assign n8916 = n5618 & ~n8892;
  assign n8917 = n5619_1 & ~n8892;
  assign n8918 = n7361 & ~n8881;
  assign n8919 = n5434_1 & ~n8892;
  assign n8920 = P3_INSTADDRPOINTER_REG_13_ & n8810;
  assign n8921 = ~P3_INSTADDRPOINTER_REG_14_ & n8920;
  assign n8922 = P3_INSTADDRPOINTER_REG_14_ & ~n8920;
  assign n8923 = ~n8921 & ~n8922;
  assign n8924 = n7364 & ~n8923;
  assign n8925 = ~n8919 & ~n8924;
  assign n8926 = ~n8916 & ~n8917;
  assign n8927 = ~n8918 & n8926;
  assign n8928 = n8925 & n8927;
  assign n8929 = ~n8747 & ~n8820;
  assign n8930 = n8743 & n8929;
  assign n8931 = n8740 & ~n8822;
  assign n8932 = ~n8498 & n8931;
  assign n8933 = n8930 & ~n8932;
  assign n8934 = ~P3_INSTADDRPOINTER_REG_14_ & ~n8303;
  assign n8935 = P3_INSTADDRPOINTER_REG_14_ & n8303;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = n8933 & ~n8936;
  assign n8938 = ~n8933 & n8936;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = n7458 & ~n8939;
  assign n8941 = ~P3_INSTADDRPOINTER_REG_14_ & n8838;
  assign n8942 = P3_INSTADDRPOINTER_REG_14_ & ~n8838;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = n7460 & ~n8943;
  assign n8945 = n8914 & ~n8915;
  assign n8946 = n8928 & n8945;
  assign n8947 = ~n8940 & n8946;
  assign n8948 = ~n8944 & n8947;
  assign n8949 = n8911 & n8948;
  assign n8950 = n7353 & ~n8949;
  assign n1735 = ~n8877 | n8950;
  assign n8952 = P3_INSTADDRPOINTER_REG_15_ & n7352;
  assign n8953 = P3_REIP_REG_15_ & n7497;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = P3_INSTADDRPOINTER_REG_14_ & n8878;
  assign n8956 = ~P3_INSTADDRPOINTER_REG_15_ & n8955;
  assign n8957 = P3_INSTADDRPOINTER_REG_15_ & ~n8955;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = n7477 & ~n8958;
  assign n8960 = n5504_1 & ~n8958;
  assign n8961 = n7466 & ~n8958;
  assign n8962 = n7470 & ~n8958;
  assign n8963 = ~n8959 & ~n8960;
  assign n8964 = ~n8961 & n8963;
  assign n8965 = ~n8962 & n8964;
  assign n8966 = P3_INSTADDRPOINTER_REG_14_ & n8889;
  assign n8967 = ~P3_INSTADDRPOINTER_REG_15_ & n8966;
  assign n8968 = P3_INSTADDRPOINTER_REG_15_ & ~n8966;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = n5360 & ~n8969;
  assign n8971 = n5438 & ~n8969;
  assign n8972 = n5442 & ~n8969;
  assign n8973 = P3_INSTADDRPOINTER_REG_14_ & n8896;
  assign n8974 = ~P3_INSTADDRPOINTER_REG_15_ & n8973;
  assign n8975 = P3_INSTADDRPOINTER_REG_15_ & ~n8973;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = n5458 & ~n8976;
  assign n8978 = n5450 & ~n8976;
  assign n8979 = ~n8970 & ~n8971;
  assign n8980 = ~n8972 & n8979;
  assign n8981 = ~n8977 & n8980;
  assign n8982 = ~n8978 & n8981;
  assign n8983 = P3_INSTADDRPOINTER_REG_14_ & n8863;
  assign n8984 = ~P3_INSTADDRPOINTER_REG_15_ & ~n8983;
  assign n8985 = P3_INSTADDRPOINTER_REG_14_ & P3_INSTADDRPOINTER_REG_15_;
  assign n8986 = P3_INSTADDRPOINTER_REG_13_ & n8985;
  assign n8987 = n8784 & n8986;
  assign n8988 = ~n8984 & ~n8987;
  assign n8989 = n5461 & n8988;
  assign n8990 = n8965 & n8982;
  assign n8991 = ~n8989 & n8990;
  assign n8992 = n5657 & ~n8958;
  assign n8993 = n5500 & ~n8958;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = ~n5547 & ~n8958;
  assign n8996 = n5618 & ~n8969;
  assign n8997 = n5619_1 & ~n8969;
  assign n8998 = n7361 & ~n8958;
  assign n8999 = n5434_1 & ~n8969;
  assign n9000 = P3_INSTADDRPOINTER_REG_13_ & P3_INSTADDRPOINTER_REG_14_;
  assign n9001 = n8810 & n9000;
  assign n9002 = P3_INSTADDRPOINTER_REG_15_ & ~n9001;
  assign n9003 = ~P3_INSTADDRPOINTER_REG_15_ & n9001;
  assign n9004 = ~n9002 & ~n9003;
  assign n9005 = n7364 & ~n9004;
  assign n9006 = ~n8999 & ~n9005;
  assign n9007 = ~n8996 & ~n8997;
  assign n9008 = ~n8998 & n9007;
  assign n9009 = n9006 & n9008;
  assign n9010 = P3_INSTADDRPOINTER_REG_14_ & ~n8303;
  assign n9011 = ~P3_INSTADDRPOINTER_REG_14_ & n8303;
  assign n9012 = ~n8933 & ~n9011;
  assign n9013 = ~n9010 & ~n9012;
  assign n9014 = ~P3_INSTADDRPOINTER_REG_15_ & ~n8303;
  assign n9015 = P3_INSTADDRPOINTER_REG_15_ & n8303;
  assign n9016 = ~n9014 & ~n9015;
  assign n9017 = n9013 & ~n9016;
  assign n9018 = ~n9013 & n9016;
  assign n9019 = ~n9017 & ~n9018;
  assign n9020 = n7458 & ~n9019;
  assign n9021 = P3_INSTADDRPOINTER_REG_14_ & n8838;
  assign n9022 = ~P3_INSTADDRPOINTER_REG_15_ & ~n9021;
  assign n9023 = n8758 & n8986;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = n7460 & n9024;
  assign n9026 = n8994 & ~n8995;
  assign n9027 = n9009 & n9026;
  assign n9028 = ~n9020 & n9027;
  assign n9029 = ~n9025 & n9028;
  assign n9030 = n8991 & n9029;
  assign n9031 = n7353 & ~n9030;
  assign n1740 = ~n8954 | n9031;
  assign n9033 = P3_INSTADDRPOINTER_REG_16_ & n7352;
  assign n9034 = P3_REIP_REG_16_ & n7497;
  assign n9035 = P3_INSTADDRPOINTER_REG_15_ & n8955;
  assign n9036 = ~P3_INSTADDRPOINTER_REG_16_ & n9035;
  assign n9037 = P3_INSTADDRPOINTER_REG_16_ & ~n9035;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~n5547 & ~n9038;
  assign n9040 = P3_INSTADDRPOINTER_REG_15_ & n8966;
  assign n9041 = ~P3_INSTADDRPOINTER_REG_16_ & n9040;
  assign n9042 = P3_INSTADDRPOINTER_REG_16_ & ~n9040;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = n5618 & ~n9043;
  assign n9045 = n5619_1 & ~n9043;
  assign n9046 = n7361 & ~n9038;
  assign n9047 = n5434_1 & ~n9043;
  assign n9048 = P3_INSTADDRPOINTER_REG_15_ & n9001;
  assign n9049 = ~P3_INSTADDRPOINTER_REG_16_ & n9048;
  assign n9050 = P3_INSTADDRPOINTER_REG_16_ & ~n9048;
  assign n9051 = ~n9049 & ~n9050;
  assign n9052 = n7364 & ~n9051;
  assign n9053 = ~n9047 & ~n9052;
  assign n9054 = ~n9044 & ~n9045;
  assign n9055 = ~n9046 & n9054;
  assign n9056 = n9053 & n9055;
  assign n9057 = ~P3_INSTADDRPOINTER_REG_16_ & n9023;
  assign n9058 = P3_INSTADDRPOINTER_REG_16_ & ~n9023;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = n7460 & ~n9059;
  assign n9061 = n5657 & ~n9038;
  assign n9062 = n5500 & ~n9038;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = P3_INSTADDRPOINTER_REG_15_ & ~n8303;
  assign n9065 = ~P3_INSTADDRPOINTER_REG_15_ & n8303;
  assign n9066 = ~n9013 & ~n9065;
  assign n9067 = ~n9064 & ~n9066;
  assign n9068 = ~P3_INSTADDRPOINTER_REG_16_ & ~n8303;
  assign n9069 = P3_INSTADDRPOINTER_REG_16_ & n8303;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = n9067 & ~n9070;
  assign n9072 = ~n9067 & n9070;
  assign n9073 = ~n9071 & ~n9072;
  assign n9074 = n7458 & ~n9073;
  assign n9075 = n9063 & ~n9074;
  assign n9076 = n7477 & ~n9038;
  assign n9077 = n5504_1 & ~n9038;
  assign n9078 = n7466 & ~n9038;
  assign n9079 = n7470 & ~n9038;
  assign n9080 = ~n9076 & ~n9077;
  assign n9081 = ~n9078 & n9080;
  assign n9082 = ~n9079 & n9081;
  assign n9083 = n5360 & ~n9043;
  assign n9084 = n5438 & ~n9043;
  assign n9085 = n5442 & ~n9043;
  assign n9086 = P3_INSTADDRPOINTER_REG_15_ & n8973;
  assign n9087 = ~P3_INSTADDRPOINTER_REG_16_ & n9086;
  assign n9088 = P3_INSTADDRPOINTER_REG_16_ & ~n9086;
  assign n9089 = ~n9087 & ~n9088;
  assign n9090 = n5458 & ~n9089;
  assign n9091 = n5450 & ~n9089;
  assign n9092 = ~n9083 & ~n9084;
  assign n9093 = ~n9085 & n9092;
  assign n9094 = ~n9090 & n9093;
  assign n9095 = ~n9091 & n9094;
  assign n9096 = ~P3_INSTADDRPOINTER_REG_16_ & n8987;
  assign n9097 = P3_INSTADDRPOINTER_REG_16_ & ~n8987;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = n5461 & ~n9098;
  assign n9100 = n9082 & n9095;
  assign n9101 = ~n9099 & n9100;
  assign n9102 = ~n9039 & n9056;
  assign n9103 = ~n9060 & n9102;
  assign n9104 = n9075 & n9103;
  assign n9105 = n9101 & n9104;
  assign n9106 = n7353 & ~n9105;
  assign n9107 = ~n9033 & ~n9034;
  assign n1745 = n9106 | ~n9107;
  assign n9109 = P3_INSTADDRPOINTER_REG_17_ & n7352;
  assign n9110 = P3_REIP_REG_17_ & n7497;
  assign n9111 = P3_INSTADDRPOINTER_REG_16_ & n9035;
  assign n9112 = ~P3_INSTADDRPOINTER_REG_17_ & n9111;
  assign n9113 = P3_INSTADDRPOINTER_REG_17_ & ~n9111;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = ~n5547 & ~n9114;
  assign n9116 = n5657 & ~n9114;
  assign n9117 = n5500 & ~n9114;
  assign n9118 = ~n9116 & ~n9117;
  assign n9119 = P3_INSTADDRPOINTER_REG_16_ & n9023;
  assign n9120 = ~P3_INSTADDRPOINTER_REG_17_ & ~n9119;
  assign n9121 = P3_INSTADDRPOINTER_REG_16_ & P3_INSTADDRPOINTER_REG_17_;
  assign n9122 = n9023 & n9121;
  assign n9123 = ~n9120 & ~n9122;
  assign n9124 = n7460 & n9123;
  assign n9125 = n7477 & ~n9114;
  assign n9126 = n5504_1 & ~n9114;
  assign n9127 = n7466 & ~n9114;
  assign n9128 = n7470 & ~n9114;
  assign n9129 = ~n9125 & ~n9126;
  assign n9130 = ~n9127 & n9129;
  assign n9131 = ~n9128 & n9130;
  assign n9132 = P3_INSTADDRPOINTER_REG_16_ & n9040;
  assign n9133 = ~P3_INSTADDRPOINTER_REG_17_ & n9132;
  assign n9134 = P3_INSTADDRPOINTER_REG_17_ & ~n9132;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = n5360 & ~n9135;
  assign n9137 = n5438 & ~n9135;
  assign n9138 = n5442 & ~n9135;
  assign n9139 = P3_INSTADDRPOINTER_REG_16_ & n9086;
  assign n9140 = ~P3_INSTADDRPOINTER_REG_17_ & n9139;
  assign n9141 = P3_INSTADDRPOINTER_REG_17_ & ~n9139;
  assign n9142 = ~n9140 & ~n9141;
  assign n9143 = n5458 & ~n9142;
  assign n9144 = n5450 & ~n9142;
  assign n9145 = ~n9136 & ~n9137;
  assign n9146 = ~n9138 & n9145;
  assign n9147 = ~n9143 & n9146;
  assign n9148 = ~n9144 & n9147;
  assign n9149 = P3_INSTADDRPOINTER_REG_16_ & n8987;
  assign n9150 = ~P3_INSTADDRPOINTER_REG_17_ & ~n9149;
  assign n9151 = n8987 & n9121;
  assign n9152 = ~n9150 & ~n9151;
  assign n9153 = n5461 & n9152;
  assign n9154 = n9131 & n9148;
  assign n9155 = ~n9153 & n9154;
  assign n9156 = n5618 & ~n9135;
  assign n9157 = n5619_1 & ~n9135;
  assign n9158 = n7361 & ~n9114;
  assign n9159 = n5434_1 & ~n9135;
  assign n9160 = P3_INSTADDRPOINTER_REG_15_ & P3_INSTADDRPOINTER_REG_16_;
  assign n9161 = n9001 & n9160;
  assign n9162 = P3_INSTADDRPOINTER_REG_17_ & ~n9161;
  assign n9163 = ~P3_INSTADDRPOINTER_REG_17_ & n9161;
  assign n9164 = ~n9162 & ~n9163;
  assign n9165 = n7364 & ~n9164;
  assign n9166 = ~n9159 & ~n9165;
  assign n9167 = ~n9067 & n9121;
  assign n9168 = n8303 & ~n9167;
  assign n9169 = P3_INSTADDRPOINTER_REG_17_ & ~n8303;
  assign n9170 = ~P3_INSTADDRPOINTER_REG_16_ & ~n9064;
  assign n9171 = ~n9066 & n9170;
  assign n9172 = ~n9168 & ~n9169;
  assign n9173 = ~n9171 & n9172;
  assign n9174 = P3_INSTADDRPOINTER_REG_17_ & n9171;
  assign n9175 = ~n8303 & ~n9174;
  assign n9176 = P3_INSTADDRPOINTER_REG_17_ & n8303;
  assign n9177 = P3_INSTADDRPOINTER_REG_16_ & ~n9067;
  assign n9178 = ~n9175 & ~n9176;
  assign n9179 = ~n9177 & n9178;
  assign n9180 = ~n9173 & ~n9179;
  assign n9181 = n7458 & n9180;
  assign n9182 = ~n9156 & ~n9157;
  assign n9183 = ~n9158 & n9182;
  assign n9184 = n9166 & n9183;
  assign n9185 = ~n9181 & n9184;
  assign n9186 = ~n9115 & n9118;
  assign n9187 = ~n9124 & n9186;
  assign n9188 = n9155 & n9187;
  assign n9189 = n9185 & n9188;
  assign n9190 = n7353 & ~n9189;
  assign n9191 = ~n9109 & ~n9110;
  assign n1750 = n9190 | ~n9191;
  assign n9193 = P3_INSTADDRPOINTER_REG_18_ & n7352;
  assign n9194 = P3_REIP_REG_18_ & n7497;
  assign n9195 = P3_INSTADDRPOINTER_REG_17_ & n9111;
  assign n9196 = ~P3_INSTADDRPOINTER_REG_18_ & n9195;
  assign n9197 = P3_INSTADDRPOINTER_REG_18_ & ~n9195;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n5547 & ~n9198;
  assign n9200 = P3_INSTADDRPOINTER_REG_17_ & n9132;
  assign n9201 = ~P3_INSTADDRPOINTER_REG_18_ & n9200;
  assign n9202 = P3_INSTADDRPOINTER_REG_18_ & ~n9200;
  assign n9203 = ~n9201 & ~n9202;
  assign n9204 = n5618 & ~n9203;
  assign n9205 = n5619_1 & ~n9203;
  assign n9206 = n7361 & ~n9198;
  assign n9207 = n5434_1 & ~n9203;
  assign n9208 = P3_INSTADDRPOINTER_REG_17_ & n9161;
  assign n9209 = ~P3_INSTADDRPOINTER_REG_18_ & n9208;
  assign n9210 = P3_INSTADDRPOINTER_REG_18_ & ~n9208;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = n7364 & ~n9211;
  assign n9213 = ~n9207 & ~n9212;
  assign n9214 = ~n9204 & ~n9205;
  assign n9215 = ~n9206 & n9214;
  assign n9216 = n9213 & n9215;
  assign n9217 = ~P3_INSTADDRPOINTER_REG_18_ & n9122;
  assign n9218 = P3_INSTADDRPOINTER_REG_18_ & ~n9122;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = n7460 & ~n9219;
  assign n9221 = n5657 & ~n9198;
  assign n9222 = n5500 & ~n9198;
  assign n9223 = ~n9221 & ~n9222;
  assign n9224 = ~n8303 & ~n9171;
  assign n9225 = ~n9167 & ~n9224;
  assign n9226 = ~n9169 & n9225;
  assign n9227 = ~P3_INSTADDRPOINTER_REG_18_ & ~n8303;
  assign n9228 = P3_INSTADDRPOINTER_REG_18_ & n8303;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = n9226 & ~n9229;
  assign n9231 = ~n9226 & n9229;
  assign n9232 = ~n9230 & ~n9231;
  assign n9233 = n7458 & ~n9232;
  assign n9234 = n9223 & ~n9233;
  assign n9235 = n7477 & ~n9198;
  assign n9236 = n5504_1 & ~n9198;
  assign n9237 = n7466 & ~n9198;
  assign n9238 = n7470 & ~n9198;
  assign n9239 = ~n9235 & ~n9236;
  assign n9240 = ~n9237 & n9239;
  assign n9241 = ~n9238 & n9240;
  assign n9242 = n5360 & ~n9203;
  assign n9243 = n5438 & ~n9203;
  assign n9244 = n5442 & ~n9203;
  assign n9245 = P3_INSTADDRPOINTER_REG_17_ & n9139;
  assign n9246 = ~P3_INSTADDRPOINTER_REG_18_ & n9245;
  assign n9247 = P3_INSTADDRPOINTER_REG_18_ & ~n9245;
  assign n9248 = ~n9246 & ~n9247;
  assign n9249 = n5458 & ~n9248;
  assign n9250 = n5450 & ~n9248;
  assign n9251 = ~n9242 & ~n9243;
  assign n9252 = ~n9244 & n9251;
  assign n9253 = ~n9249 & n9252;
  assign n9254 = ~n9250 & n9253;
  assign n9255 = ~P3_INSTADDRPOINTER_REG_18_ & n9151;
  assign n9256 = P3_INSTADDRPOINTER_REG_18_ & ~n9151;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = n5461 & ~n9257;
  assign n9259 = n9241 & n9254;
  assign n9260 = ~n9258 & n9259;
  assign n9261 = ~n9199 & n9216;
  assign n9262 = ~n9220 & n9261;
  assign n9263 = n9234 & n9262;
  assign n9264 = n9260 & n9263;
  assign n9265 = n7353 & ~n9264;
  assign n9266 = ~n9193 & ~n9194;
  assign n1755 = n9265 | ~n9266;
  assign n9268 = P3_INSTADDRPOINTER_REG_19_ & n7352;
  assign n9269 = P3_REIP_REG_19_ & n7497;
  assign n9270 = P3_INSTADDRPOINTER_REG_18_ & n9195;
  assign n9271 = ~P3_INSTADDRPOINTER_REG_19_ & n9270;
  assign n9272 = P3_INSTADDRPOINTER_REG_19_ & ~n9270;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = ~n5547 & ~n9273;
  assign n9275 = n5657 & ~n9273;
  assign n9276 = n5500 & ~n9273;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = P3_INSTADDRPOINTER_REG_18_ & n9122;
  assign n9279 = ~P3_INSTADDRPOINTER_REG_19_ & ~n9278;
  assign n9280 = P3_INSTADDRPOINTER_REG_18_ & P3_INSTADDRPOINTER_REG_19_;
  assign n9281 = n9122 & n9280;
  assign n9282 = ~n9279 & ~n9281;
  assign n9283 = n7460 & n9282;
  assign n9284 = n7477 & ~n9273;
  assign n9285 = n5504_1 & ~n9273;
  assign n9286 = n7466 & ~n9273;
  assign n9287 = n7470 & ~n9273;
  assign n9288 = ~n9284 & ~n9285;
  assign n9289 = ~n9286 & n9288;
  assign n9290 = ~n9287 & n9289;
  assign n9291 = P3_INSTADDRPOINTER_REG_18_ & n9200;
  assign n9292 = ~P3_INSTADDRPOINTER_REG_19_ & n9291;
  assign n9293 = P3_INSTADDRPOINTER_REG_19_ & ~n9291;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = n5360 & ~n9294;
  assign n9296 = n5438 & ~n9294;
  assign n9297 = n5442 & ~n9294;
  assign n9298 = P3_INSTADDRPOINTER_REG_18_ & n9245;
  assign n9299 = ~P3_INSTADDRPOINTER_REG_19_ & n9298;
  assign n9300 = P3_INSTADDRPOINTER_REG_19_ & ~n9298;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = n5458 & ~n9301;
  assign n9303 = n5450 & ~n9301;
  assign n9304 = ~n9295 & ~n9296;
  assign n9305 = ~n9297 & n9304;
  assign n9306 = ~n9302 & n9305;
  assign n9307 = ~n9303 & n9306;
  assign n9308 = P3_INSTADDRPOINTER_REG_18_ & n9151;
  assign n9309 = ~P3_INSTADDRPOINTER_REG_19_ & ~n9308;
  assign n9310 = n9151 & n9280;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = n5461 & n9311;
  assign n9313 = n9290 & n9307;
  assign n9314 = ~n9312 & n9313;
  assign n9315 = n5618 & ~n9294;
  assign n9316 = n5619_1 & ~n9294;
  assign n9317 = n7361 & ~n9273;
  assign n9318 = n5434_1 & ~n9294;
  assign n9319 = P3_INSTADDRPOINTER_REG_17_ & P3_INSTADDRPOINTER_REG_18_;
  assign n9320 = n9161 & n9319;
  assign n9321 = P3_INSTADDRPOINTER_REG_19_ & ~n9320;
  assign n9322 = ~P3_INSTADDRPOINTER_REG_19_ & n9320;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = n7364 & ~n9323;
  assign n9325 = ~n9318 & ~n9324;
  assign n9326 = ~P3_INSTADDRPOINTER_REG_19_ & ~n8303;
  assign n9327 = P3_INSTADDRPOINTER_REG_19_ & n8303;
  assign n9328 = ~n9326 & ~n9327;
  assign n9329 = ~P3_INSTADDRPOINTER_REG_18_ & n8303;
  assign n9330 = ~n9226 & ~n9329;
  assign n9331 = P3_INSTADDRPOINTER_REG_18_ & ~n8303;
  assign n9332 = ~n9330 & ~n9331;
  assign n9333 = ~n9328 & n9332;
  assign n9334 = ~P3_INSTADDRPOINTER_REG_19_ & n8303;
  assign n9335 = P3_INSTADDRPOINTER_REG_19_ & ~n8303;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = ~n9332 & ~n9336;
  assign n9338 = ~n9333 & ~n9337;
  assign n9339 = n7458 & ~n9338;
  assign n9340 = ~n9315 & ~n9316;
  assign n9341 = ~n9317 & n9340;
  assign n9342 = n9325 & n9341;
  assign n9343 = ~n9339 & n9342;
  assign n9344 = ~n9274 & n9277;
  assign n9345 = ~n9283 & n9344;
  assign n9346 = n9314 & n9345;
  assign n9347 = n9343 & n9346;
  assign n9348 = n7353 & ~n9347;
  assign n9349 = ~n9268 & ~n9269;
  assign n1760 = n9348 | ~n9349;
  assign n9351 = P3_INSTADDRPOINTER_REG_20_ & n7352;
  assign n9352 = P3_REIP_REG_20_ & n7497;
  assign n9353 = ~n9351 & ~n9352;
  assign n9354 = P3_INSTADDRPOINTER_REG_19_ & P3_INSTADDRPOINTER_REG_20_;
  assign n9355 = n8303 & ~n9354;
  assign n9356 = P3_INSTADDRPOINTER_REG_20_ & ~n8303;
  assign n9357 = ~n9355 & ~n9356;
  assign n9358 = n9332 & ~n9335;
  assign n9359 = n9357 & ~n9358;
  assign n9360 = ~P3_INSTADDRPOINTER_REG_19_ & n9332;
  assign n9361 = P3_INSTADDRPOINTER_REG_20_ & n9360;
  assign n9362 = ~n8303 & ~n9361;
  assign n9363 = P3_INSTADDRPOINTER_REG_20_ & n8303;
  assign n9364 = P3_INSTADDRPOINTER_REG_19_ & ~n9332;
  assign n9365 = ~n9362 & ~n9363;
  assign n9366 = ~n9364 & n9365;
  assign n9367 = ~n9359 & ~n9366;
  assign n9368 = n7458 & n9367;
  assign n9369 = P3_INSTADDRPOINTER_REG_19_ & n9270;
  assign n9370 = ~P3_INSTADDRPOINTER_REG_20_ & n9369;
  assign n9371 = P3_INSTADDRPOINTER_REG_20_ & ~n9369;
  assign n9372 = ~n9370 & ~n9371;
  assign n9373 = ~n5547 & ~n9372;
  assign n9374 = n5657 & ~n9372;
  assign n9375 = n5500 & ~n9372;
  assign n9376 = ~n9374 & ~n9375;
  assign n9377 = P3_INSTADDRPOINTER_REG_19_ & n9291;
  assign n9378 = ~P3_INSTADDRPOINTER_REG_20_ & n9377;
  assign n9379 = P3_INSTADDRPOINTER_REG_20_ & ~n9377;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = n5618 & ~n9380;
  assign n9382 = n5619_1 & ~n9380;
  assign n9383 = n7361 & ~n9372;
  assign n9384 = n5434_1 & ~n9380;
  assign n9385 = P3_INSTADDRPOINTER_REG_19_ & n9320;
  assign n9386 = ~P3_INSTADDRPOINTER_REG_20_ & n9385;
  assign n9387 = P3_INSTADDRPOINTER_REG_20_ & ~n9385;
  assign n9388 = ~n9386 & ~n9387;
  assign n9389 = n7364 & ~n9388;
  assign n9390 = ~n9384 & ~n9389;
  assign n9391 = ~n9381 & ~n9382;
  assign n9392 = ~n9383 & n9391;
  assign n9393 = n9390 & n9392;
  assign n9394 = ~P3_INSTADDRPOINTER_REG_20_ & ~n9281;
  assign n9395 = P3_INSTADDRPOINTER_REG_20_ & n9281;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = n7460 & n9396;
  assign n9398 = n7477 & ~n9372;
  assign n9399 = n5504_1 & ~n9372;
  assign n9400 = n7466 & ~n9372;
  assign n9401 = n7470 & ~n9372;
  assign n9402 = ~n9398 & ~n9399;
  assign n9403 = ~n9400 & n9402;
  assign n9404 = ~n9401 & n9403;
  assign n9405 = n5360 & ~n9380;
  assign n9406 = n5438 & ~n9380;
  assign n9407 = n5442 & ~n9380;
  assign n9408 = P3_INSTADDRPOINTER_REG_19_ & n9298;
  assign n9409 = ~P3_INSTADDRPOINTER_REG_20_ & n9408;
  assign n9410 = P3_INSTADDRPOINTER_REG_20_ & ~n9408;
  assign n9411 = ~n9409 & ~n9410;
  assign n9412 = n5458 & ~n9411;
  assign n9413 = n5450 & ~n9411;
  assign n9414 = ~n9405 & ~n9406;
  assign n9415 = ~n9407 & n9414;
  assign n9416 = ~n9412 & n9415;
  assign n9417 = ~n9413 & n9416;
  assign n9418 = ~P3_INSTADDRPOINTER_REG_20_ & ~n9310;
  assign n9419 = P3_INSTADDRPOINTER_REG_20_ & n9310;
  assign n9420 = ~n9418 & ~n9419;
  assign n9421 = n5461 & n9420;
  assign n9422 = n9404 & n9417;
  assign n9423 = ~n9421 & n9422;
  assign n9424 = ~n9373 & n9376;
  assign n9425 = n9393 & n9424;
  assign n9426 = ~n9397 & n9425;
  assign n9427 = n9423 & n9426;
  assign n9428 = ~n9368 & n9427;
  assign n9429 = n7353 & ~n9428;
  assign n1765 = ~n9353 | n9429;
  assign n9431 = P3_INSTADDRPOINTER_REG_21_ & n7352;
  assign n9432 = P3_REIP_REG_21_ & n7497;
  assign n9433 = ~n9431 & ~n9432;
  assign n9434 = ~n9332 & n9354;
  assign n9435 = ~n9356 & ~n9434;
  assign n9436 = ~n8303 & ~n9360;
  assign n9437 = n9435 & ~n9436;
  assign n9438 = ~P3_INSTADDRPOINTER_REG_21_ & ~n8303;
  assign n9439 = P3_INSTADDRPOINTER_REG_21_ & n8303;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = n9437 & ~n9440;
  assign n9442 = ~n9437 & n9440;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = n7458 & ~n9443;
  assign n9445 = P3_INSTADDRPOINTER_REG_20_ & n9369;
  assign n9446 = ~P3_INSTADDRPOINTER_REG_21_ & n9445;
  assign n9447 = P3_INSTADDRPOINTER_REG_21_ & ~n9445;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n5547 & ~n9448;
  assign n9450 = n5657 & ~n9448;
  assign n9451 = n5500 & ~n9448;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = P3_INSTADDRPOINTER_REG_20_ & n9377;
  assign n9454 = ~P3_INSTADDRPOINTER_REG_21_ & n9453;
  assign n9455 = P3_INSTADDRPOINTER_REG_21_ & ~n9453;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = n5618 & ~n9456;
  assign n9458 = n5619_1 & ~n9456;
  assign n9459 = n7361 & ~n9448;
  assign n9460 = n5434_1 & ~n9456;
  assign n9461 = n9320 & n9354;
  assign n9462 = P3_INSTADDRPOINTER_REG_21_ & ~n9461;
  assign n9463 = ~P3_INSTADDRPOINTER_REG_21_ & n9461;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = n7364 & ~n9464;
  assign n9466 = ~n9460 & ~n9465;
  assign n9467 = ~n9457 & ~n9458;
  assign n9468 = ~n9459 & n9467;
  assign n9469 = n9466 & n9468;
  assign n9470 = ~P3_INSTADDRPOINTER_REG_21_ & ~n9395;
  assign n9471 = P3_INSTADDRPOINTER_REG_21_ & n9395;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = n7460 & n9472;
  assign n9474 = n5360 & ~n9456;
  assign n9475 = n5438 & ~n9456;
  assign n9476 = n5442 & ~n9456;
  assign n9477 = P3_INSTADDRPOINTER_REG_20_ & n9408;
  assign n9478 = ~P3_INSTADDRPOINTER_REG_21_ & n9477;
  assign n9479 = P3_INSTADDRPOINTER_REG_21_ & ~n9477;
  assign n9480 = ~n9478 & ~n9479;
  assign n9481 = n5458 & ~n9480;
  assign n9482 = n5450 & ~n9480;
  assign n9483 = ~n9474 & ~n9475;
  assign n9484 = ~n9476 & n9483;
  assign n9485 = ~n9481 & n9484;
  assign n9486 = ~n9482 & n9485;
  assign n9487 = n7477 & ~n9448;
  assign n9488 = n5504_1 & ~n9448;
  assign n9489 = n7466 & ~n9448;
  assign n9490 = n7470 & ~n9448;
  assign n9491 = ~n9487 & ~n9488;
  assign n9492 = ~n9489 & n9491;
  assign n9493 = ~n9490 & n9492;
  assign n9494 = ~P3_INSTADDRPOINTER_REG_21_ & ~n9419;
  assign n9495 = P3_INSTADDRPOINTER_REG_20_ & P3_INSTADDRPOINTER_REG_21_;
  assign n9496 = n9310 & n9495;
  assign n9497 = ~n9494 & ~n9496;
  assign n9498 = n5461 & n9497;
  assign n9499 = n9486 & n9493;
  assign n9500 = ~n9498 & n9499;
  assign n9501 = ~n9449 & n9452;
  assign n9502 = n9469 & n9501;
  assign n9503 = ~n9473 & n9502;
  assign n9504 = n9500 & n9503;
  assign n9505 = ~n9444 & n9504;
  assign n9506 = n7353 & ~n9505;
  assign n1770 = ~n9433 | n9506;
  assign n9508 = P3_INSTADDRPOINTER_REG_22_ & n7352;
  assign n9509 = P3_REIP_REG_22_ & n7497;
  assign n9510 = ~n9508 & ~n9509;
  assign n9511 = P3_INSTADDRPOINTER_REG_21_ & n9477;
  assign n9512 = ~P3_INSTADDRPOINTER_REG_22_ & n9511;
  assign n9513 = P3_INSTADDRPOINTER_REG_22_ & ~n9511;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = n5458 & ~n9514;
  assign n9516 = n5450 & ~n9514;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = P3_INSTADDRPOINTER_REG_21_ & n9453;
  assign n9519 = ~P3_INSTADDRPOINTER_REG_22_ & n9518;
  assign n9520 = P3_INSTADDRPOINTER_REG_22_ & ~n9518;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = n5360 & ~n9521;
  assign n9523 = n5438 & ~n9521;
  assign n9524 = n5442 & ~n9521;
  assign n9525 = ~n9522 & ~n9523;
  assign n9526 = ~n9524 & n9525;
  assign n9527 = P3_INSTADDRPOINTER_REG_21_ & n9445;
  assign n9528 = ~P3_INSTADDRPOINTER_REG_22_ & n9527;
  assign n9529 = P3_INSTADDRPOINTER_REG_22_ & ~n9527;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = n7466 & ~n9530;
  assign n9532 = n7470 & ~n9530;
  assign n9533 = n5504_1 & ~n9530;
  assign n9534 = ~n9531 & ~n9532;
  assign n9535 = ~n9533 & n9534;
  assign n9536 = ~P3_INSTADDRPOINTER_REG_22_ & n9496;
  assign n9537 = P3_INSTADDRPOINTER_REG_22_ & ~n9496;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = n5461 & ~n9538;
  assign n9540 = n7477 & ~n9530;
  assign n9541 = ~n9539 & ~n9540;
  assign n9542 = n9517 & n9526;
  assign n9543 = n9535 & n9542;
  assign n9544 = n9541 & n9543;
  assign n9545 = P3_INSTADDRPOINTER_REG_21_ & n9354;
  assign n9546 = n8303 & ~n9545;
  assign n9547 = ~n9329 & ~n9546;
  assign n9548 = ~n9226 & n9547;
  assign n9549 = P3_INSTADDRPOINTER_REG_21_ & ~n8303;
  assign n9550 = ~n9331 & ~n9549;
  assign n9551 = ~n9335 & n9550;
  assign n9552 = ~n9356 & n9551;
  assign n9553 = ~n9548 & n9552;
  assign n9554 = ~P3_INSTADDRPOINTER_REG_22_ & ~n8303;
  assign n9555 = P3_INSTADDRPOINTER_REG_22_ & n8303;
  assign n9556 = ~n9554 & ~n9555;
  assign n9557 = n9553 & ~n9556;
  assign n9558 = ~n9553 & n9556;
  assign n9559 = ~n9557 & ~n9558;
  assign n9560 = n7458 & ~n9559;
  assign n9561 = ~n5547 & ~n9530;
  assign n9562 = n5657 & ~n9530;
  assign n9563 = n5500 & ~n9530;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = n5618 & ~n9521;
  assign n9566 = n5619_1 & ~n9521;
  assign n9567 = n7361 & ~n9530;
  assign n9568 = n5434_1 & ~n9521;
  assign n9569 = P3_INSTADDRPOINTER_REG_21_ & n9461;
  assign n9570 = ~P3_INSTADDRPOINTER_REG_22_ & n9569;
  assign n9571 = P3_INSTADDRPOINTER_REG_22_ & ~n9569;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = n7364 & ~n9572;
  assign n9574 = ~n9568 & ~n9573;
  assign n9575 = ~n9565 & ~n9566;
  assign n9576 = ~n9567 & n9575;
  assign n9577 = n9574 & n9576;
  assign n9578 = ~P3_INSTADDRPOINTER_REG_22_ & n9471;
  assign n9579 = P3_INSTADDRPOINTER_REG_22_ & ~n9471;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = n7460 & ~n9580;
  assign n9582 = ~n9560 & ~n9561;
  assign n9583 = n9564 & n9582;
  assign n9584 = n9577 & n9583;
  assign n9585 = ~n9581 & n9584;
  assign n9586 = n9544 & n9585;
  assign n9587 = n7353 & ~n9586;
  assign n1775 = ~n9510 | n9587;
  assign n9589 = P3_INSTADDRPOINTER_REG_23_ & n7352;
  assign n9590 = P3_REIP_REG_23_ & n7497;
  assign n9591 = ~n9589 & ~n9590;
  assign n9592 = P3_INSTADDRPOINTER_REG_22_ & n9511;
  assign n9593 = ~P3_INSTADDRPOINTER_REG_23_ & n9592;
  assign n9594 = P3_INSTADDRPOINTER_REG_23_ & ~n9592;
  assign n9595 = ~n9593 & ~n9594;
  assign n9596 = n5458 & ~n9595;
  assign n9597 = n5450 & ~n9595;
  assign n9598 = ~n9596 & ~n9597;
  assign n9599 = P3_INSTADDRPOINTER_REG_22_ & n9518;
  assign n9600 = ~P3_INSTADDRPOINTER_REG_23_ & n9599;
  assign n9601 = P3_INSTADDRPOINTER_REG_23_ & ~n9599;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = n5360 & ~n9602;
  assign n9604 = n5438 & ~n9602;
  assign n9605 = n5442 & ~n9602;
  assign n9606 = ~n9603 & ~n9604;
  assign n9607 = ~n9605 & n9606;
  assign n9608 = P3_INSTADDRPOINTER_REG_22_ & n9527;
  assign n9609 = ~P3_INSTADDRPOINTER_REG_23_ & n9608;
  assign n9610 = P3_INSTADDRPOINTER_REG_23_ & ~n9608;
  assign n9611 = ~n9609 & ~n9610;
  assign n9612 = n7466 & ~n9611;
  assign n9613 = n7470 & ~n9611;
  assign n9614 = n5504_1 & ~n9611;
  assign n9615 = ~n9612 & ~n9613;
  assign n9616 = ~n9614 & n9615;
  assign n9617 = P3_INSTADDRPOINTER_REG_22_ & n9496;
  assign n9618 = ~P3_INSTADDRPOINTER_REG_23_ & ~n9617;
  assign n9619 = P3_INSTADDRPOINTER_REG_22_ & P3_INSTADDRPOINTER_REG_23_;
  assign n9620 = n9496 & n9619;
  assign n9621 = ~n9618 & ~n9620;
  assign n9622 = n5461 & n9621;
  assign n9623 = n7477 & ~n9611;
  assign n9624 = ~n9622 & ~n9623;
  assign n9625 = n9598 & n9607;
  assign n9626 = n9616 & n9625;
  assign n9627 = n9624 & n9626;
  assign n9628 = ~P3_INSTADDRPOINTER_REG_22_ & n8303;
  assign n9629 = n9547 & ~n9628;
  assign n9630 = ~n9226 & n9629;
  assign n9631 = P3_INSTADDRPOINTER_REG_22_ & ~n8303;
  assign n9632 = n9552 & ~n9631;
  assign n9633 = ~n9630 & n9632;
  assign n9634 = ~P3_INSTADDRPOINTER_REG_23_ & ~n8303;
  assign n9635 = P3_INSTADDRPOINTER_REG_23_ & n8303;
  assign n9636 = ~n9634 & ~n9635;
  assign n9637 = n9633 & ~n9636;
  assign n9638 = ~n9633 & n9636;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = n7458 & ~n9639;
  assign n9641 = ~n5547 & ~n9611;
  assign n9642 = n5657 & ~n9611;
  assign n9643 = n5500 & ~n9611;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = n5618 & ~n9602;
  assign n9646 = n5619_1 & ~n9602;
  assign n9647 = n7361 & ~n9611;
  assign n9648 = n5434_1 & ~n9602;
  assign n9649 = P3_INSTADDRPOINTER_REG_21_ & P3_INSTADDRPOINTER_REG_22_;
  assign n9650 = n9461 & n9649;
  assign n9651 = P3_INSTADDRPOINTER_REG_23_ & ~n9650;
  assign n9652 = ~P3_INSTADDRPOINTER_REG_23_ & n9650;
  assign n9653 = ~n9651 & ~n9652;
  assign n9654 = n7364 & ~n9653;
  assign n9655 = ~n9648 & ~n9654;
  assign n9656 = ~n9645 & ~n9646;
  assign n9657 = ~n9647 & n9656;
  assign n9658 = n9655 & n9657;
  assign n9659 = P3_INSTADDRPOINTER_REG_22_ & n9471;
  assign n9660 = ~P3_INSTADDRPOINTER_REG_23_ & ~n9659;
  assign n9661 = n9471 & n9619;
  assign n9662 = ~n9660 & ~n9661;
  assign n9663 = n7460 & n9662;
  assign n9664 = ~n9640 & ~n9641;
  assign n9665 = n9644 & n9664;
  assign n9666 = n9658 & n9665;
  assign n9667 = ~n9663 & n9666;
  assign n9668 = n9627 & n9667;
  assign n9669 = n7353 & ~n9668;
  assign n1780 = ~n9591 | n9669;
  assign n9671 = P3_INSTADDRPOINTER_REG_24_ & n7352;
  assign n9672 = P3_REIP_REG_24_ & n7497;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = P3_INSTADDRPOINTER_REG_23_ & n9592;
  assign n9675 = ~P3_INSTADDRPOINTER_REG_24_ & n9674;
  assign n9676 = P3_INSTADDRPOINTER_REG_24_ & ~n9674;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = n5458 & ~n9677;
  assign n9679 = n5450 & ~n9677;
  assign n9680 = ~n9678 & ~n9679;
  assign n9681 = P3_INSTADDRPOINTER_REG_23_ & n9599;
  assign n9682 = ~P3_INSTADDRPOINTER_REG_24_ & n9681;
  assign n9683 = P3_INSTADDRPOINTER_REG_24_ & ~n9681;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = n5360 & ~n9684;
  assign n9686 = n5438 & ~n9684;
  assign n9687 = n5442 & ~n9684;
  assign n9688 = ~n9685 & ~n9686;
  assign n9689 = ~n9687 & n9688;
  assign n9690 = ~P3_INSTADDRPOINTER_REG_24_ & n9620;
  assign n9691 = P3_INSTADDRPOINTER_REG_24_ & ~n9620;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = n5461 & ~n9692;
  assign n9694 = P3_INSTADDRPOINTER_REG_23_ & n9608;
  assign n9695 = ~P3_INSTADDRPOINTER_REG_24_ & n9694;
  assign n9696 = P3_INSTADDRPOINTER_REG_24_ & ~n9694;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = n7477 & ~n9697;
  assign n9699 = ~n9693 & ~n9698;
  assign n9700 = n7466 & ~n9697;
  assign n9701 = n7470 & ~n9697;
  assign n9702 = n5504_1 & ~n9697;
  assign n9703 = ~n9700 & ~n9701;
  assign n9704 = ~n9702 & n9703;
  assign n9705 = n9680 & n9689;
  assign n9706 = n9699 & n9705;
  assign n9707 = n9704 & n9706;
  assign n9708 = ~P3_INSTADDRPOINTER_REG_23_ & n8303;
  assign n9709 = n9629 & ~n9708;
  assign n9710 = ~n9226 & n9709;
  assign n9711 = P3_INSTADDRPOINTER_REG_23_ & ~n8303;
  assign n9712 = n9632 & ~n9711;
  assign n9713 = ~n9710 & n9712;
  assign n9714 = ~P3_INSTADDRPOINTER_REG_24_ & ~n8303;
  assign n9715 = P3_INSTADDRPOINTER_REG_24_ & n8303;
  assign n9716 = ~n9714 & ~n9715;
  assign n9717 = n9713 & ~n9716;
  assign n9718 = ~n9713 & n9716;
  assign n9719 = ~n9717 & ~n9718;
  assign n9720 = n7458 & ~n9719;
  assign n9721 = ~n5547 & ~n9697;
  assign n9722 = n5657 & ~n9697;
  assign n9723 = n5500 & ~n9697;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = ~P3_INSTADDRPOINTER_REG_24_ & n9661;
  assign n9726 = P3_INSTADDRPOINTER_REG_24_ & ~n9661;
  assign n9727 = ~n9725 & ~n9726;
  assign n9728 = n7460 & ~n9727;
  assign n9729 = n5618 & ~n9684;
  assign n9730 = n5619_1 & ~n9684;
  assign n9731 = n7361 & ~n9697;
  assign n9732 = n5434_1 & ~n9684;
  assign n9733 = P3_INSTADDRPOINTER_REG_23_ & n9650;
  assign n9734 = ~P3_INSTADDRPOINTER_REG_24_ & n9733;
  assign n9735 = P3_INSTADDRPOINTER_REG_24_ & ~n9733;
  assign n9736 = ~n9734 & ~n9735;
  assign n9737 = n7364 & ~n9736;
  assign n9738 = ~n9732 & ~n9737;
  assign n9739 = ~n9729 & ~n9730;
  assign n9740 = ~n9731 & n9739;
  assign n9741 = n9738 & n9740;
  assign n9742 = ~n9720 & ~n9721;
  assign n9743 = n9724 & n9742;
  assign n9744 = ~n9728 & n9743;
  assign n9745 = n9741 & n9744;
  assign n9746 = n9707 & n9745;
  assign n9747 = n7353 & ~n9746;
  assign n1785 = ~n9673 | n9747;
  assign n9749 = P3_INSTADDRPOINTER_REG_25_ & n7352;
  assign n9750 = P3_REIP_REG_25_ & n7497;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = P3_INSTADDRPOINTER_REG_24_ & n9674;
  assign n9753 = ~P3_INSTADDRPOINTER_REG_25_ & n9752;
  assign n9754 = P3_INSTADDRPOINTER_REG_25_ & ~n9752;
  assign n9755 = ~n9753 & ~n9754;
  assign n9756 = n5458 & ~n9755;
  assign n9757 = n5450 & ~n9755;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = P3_INSTADDRPOINTER_REG_24_ & n9681;
  assign n9760 = ~P3_INSTADDRPOINTER_REG_25_ & n9759;
  assign n9761 = P3_INSTADDRPOINTER_REG_25_ & ~n9759;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = n5360 & ~n9762;
  assign n9764 = n5438 & ~n9762;
  assign n9765 = n5442 & ~n9762;
  assign n9766 = ~n9763 & ~n9764;
  assign n9767 = ~n9765 & n9766;
  assign n9768 = P3_INSTADDRPOINTER_REG_24_ & n9620;
  assign n9769 = ~P3_INSTADDRPOINTER_REG_25_ & ~n9768;
  assign n9770 = P3_INSTADDRPOINTER_REG_24_ & P3_INSTADDRPOINTER_REG_25_;
  assign n9771 = n9620 & n9770;
  assign n9772 = ~n9769 & ~n9771;
  assign n9773 = n5461 & n9772;
  assign n9774 = P3_INSTADDRPOINTER_REG_24_ & n9694;
  assign n9775 = ~P3_INSTADDRPOINTER_REG_25_ & n9774;
  assign n9776 = P3_INSTADDRPOINTER_REG_25_ & ~n9774;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = n7477 & ~n9777;
  assign n9779 = ~n9773 & ~n9778;
  assign n9780 = n7466 & ~n9777;
  assign n9781 = n7470 & ~n9777;
  assign n9782 = n5504_1 & ~n9777;
  assign n9783 = ~n9780 & ~n9781;
  assign n9784 = ~n9782 & n9783;
  assign n9785 = n9758 & n9767;
  assign n9786 = n9779 & n9785;
  assign n9787 = n9784 & n9786;
  assign n9788 = ~P3_INSTADDRPOINTER_REG_25_ & ~n8303;
  assign n9789 = P3_INSTADDRPOINTER_REG_25_ & n8303;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = P3_INSTADDRPOINTER_REG_24_ & ~n8303;
  assign n9792 = n9712 & ~n9791;
  assign n9793 = ~P3_INSTADDRPOINTER_REG_24_ & n8303;
  assign n9794 = n9709 & ~n9793;
  assign n9795 = ~n9226 & n9794;
  assign n9796 = n9792 & ~n9795;
  assign n9797 = ~n9790 & n9796;
  assign n9798 = ~P3_INSTADDRPOINTER_REG_25_ & n8303;
  assign n9799 = P3_INSTADDRPOINTER_REG_25_ & ~n8303;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = ~n9796 & ~n9800;
  assign n9802 = ~n9797 & ~n9801;
  assign n9803 = n7458 & ~n9802;
  assign n9804 = ~n5547 & ~n9777;
  assign n9805 = P3_INSTADDRPOINTER_REG_24_ & n9661;
  assign n9806 = ~P3_INSTADDRPOINTER_REG_25_ & ~n9805;
  assign n9807 = n9661 & n9770;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = n7460 & n9808;
  assign n9810 = n5657 & ~n9777;
  assign n9811 = n5500 & ~n9777;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = n5618 & ~n9762;
  assign n9814 = n5619_1 & ~n9762;
  assign n9815 = n7361 & ~n9777;
  assign n9816 = n5434_1 & ~n9762;
  assign n9817 = P3_INSTADDRPOINTER_REG_23_ & P3_INSTADDRPOINTER_REG_24_;
  assign n9818 = n9650 & n9817;
  assign n9819 = P3_INSTADDRPOINTER_REG_25_ & ~n9818;
  assign n9820 = ~P3_INSTADDRPOINTER_REG_25_ & n9818;
  assign n9821 = ~n9819 & ~n9820;
  assign n9822 = n7364 & ~n9821;
  assign n9823 = ~n9816 & ~n9822;
  assign n9824 = ~n9813 & ~n9814;
  assign n9825 = ~n9815 & n9824;
  assign n9826 = n9823 & n9825;
  assign n9827 = ~n9803 & ~n9804;
  assign n9828 = ~n9809 & n9827;
  assign n9829 = n9812 & n9828;
  assign n9830 = n9826 & n9829;
  assign n9831 = n9787 & n9830;
  assign n9832 = n7353 & ~n9831;
  assign n1790 = ~n9751 | n9832;
  assign n9834 = P3_INSTADDRPOINTER_REG_26_ & n7352;
  assign n9835 = P3_REIP_REG_26_ & n7497;
  assign n9836 = P3_INSTADDRPOINTER_REG_26_ & ~n8303;
  assign n9837 = P3_INSTADDRPOINTER_REG_25_ & P3_INSTADDRPOINTER_REG_26_;
  assign n9838 = n8303 & ~n9837;
  assign n9839 = ~n9836 & ~n9838;
  assign n9840 = n9796 & ~n9799;
  assign n9841 = n9839 & ~n9840;
  assign n9842 = ~P3_INSTADDRPOINTER_REG_26_ & ~n8303;
  assign n9843 = P3_INSTADDRPOINTER_REG_26_ & n8303;
  assign n9844 = ~n9842 & ~n9843;
  assign n9845 = ~n9799 & n9844;
  assign n9846 = ~n9796 & ~n9798;
  assign n9847 = n9845 & ~n9846;
  assign n9848 = ~n9841 & ~n9847;
  assign n9849 = n7458 & n9848;
  assign n9850 = ~P3_INSTADDRPOINTER_REG_26_ & ~n9807;
  assign n9851 = P3_INSTADDRPOINTER_REG_26_ & n9807;
  assign n9852 = ~n9850 & ~n9851;
  assign n9853 = n7460 & n9852;
  assign n9854 = ~n9849 & ~n9853;
  assign n9855 = P3_INSTADDRPOINTER_REG_25_ & n9774;
  assign n9856 = ~P3_INSTADDRPOINTER_REG_26_ & n9855;
  assign n9857 = P3_INSTADDRPOINTER_REG_26_ & ~n9855;
  assign n9858 = ~n9856 & ~n9857;
  assign n9859 = ~n5547 & ~n9858;
  assign n9860 = n5657 & ~n9858;
  assign n9861 = n5500 & ~n9858;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = P3_INSTADDRPOINTER_REG_25_ & n9759;
  assign n9864 = ~P3_INSTADDRPOINTER_REG_26_ & n9863;
  assign n9865 = P3_INSTADDRPOINTER_REG_26_ & ~n9863;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n5618 & ~n9866;
  assign n9868 = n5619_1 & ~n9866;
  assign n9869 = n7361 & ~n9858;
  assign n9870 = n5434_1 & ~n9866;
  assign n9871 = P3_INSTADDRPOINTER_REG_25_ & n9818;
  assign n9872 = ~P3_INSTADDRPOINTER_REG_26_ & n9871;
  assign n9873 = P3_INSTADDRPOINTER_REG_26_ & ~n9871;
  assign n9874 = ~n9872 & ~n9873;
  assign n9875 = n7364 & ~n9874;
  assign n9876 = ~n9870 & ~n9875;
  assign n9877 = ~n9867 & ~n9868;
  assign n9878 = ~n9869 & n9877;
  assign n9879 = n9876 & n9878;
  assign n9880 = P3_INSTADDRPOINTER_REG_25_ & n9752;
  assign n9881 = ~P3_INSTADDRPOINTER_REG_26_ & n9880;
  assign n9882 = P3_INSTADDRPOINTER_REG_26_ & ~n9880;
  assign n9883 = ~n9881 & ~n9882;
  assign n9884 = n5458 & ~n9883;
  assign n9885 = n5450 & ~n9883;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = n5360 & ~n9866;
  assign n9888 = n5438 & ~n9866;
  assign n9889 = n5442 & ~n9866;
  assign n9890 = ~n9887 & ~n9888;
  assign n9891 = ~n9889 & n9890;
  assign n9892 = ~P3_INSTADDRPOINTER_REG_26_ & ~n9771;
  assign n9893 = P3_INSTADDRPOINTER_REG_26_ & n9771;
  assign n9894 = ~n9892 & ~n9893;
  assign n9895 = n5461 & n9894;
  assign n9896 = n7477 & ~n9858;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = n7466 & ~n9858;
  assign n9899 = n7470 & ~n9858;
  assign n9900 = n5504_1 & ~n9858;
  assign n9901 = ~n9898 & ~n9899;
  assign n9902 = ~n9900 & n9901;
  assign n9903 = n9886 & n9891;
  assign n9904 = n9897 & n9903;
  assign n9905 = n9902 & n9904;
  assign n9906 = n9854 & ~n9859;
  assign n9907 = n9862 & n9906;
  assign n9908 = n9879 & n9907;
  assign n9909 = n9905 & n9908;
  assign n9910 = n7353 & ~n9909;
  assign n9911 = ~n9834 & ~n9835;
  assign n1795 = n9910 | ~n9911;
  assign n9913 = P3_INSTADDRPOINTER_REG_27_ & n7352;
  assign n9914 = P3_REIP_REG_27_ & n7497;
  assign n9915 = ~n9799 & ~n9836;
  assign n9916 = ~n9796 & ~n9838;
  assign n9917 = n9915 & ~n9916;
  assign n9918 = ~P3_INSTADDRPOINTER_REG_27_ & ~n8303;
  assign n9919 = P3_INSTADDRPOINTER_REG_27_ & n8303;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = n9917 & ~n9920;
  assign n9922 = ~n9917 & n9920;
  assign n9923 = ~n9921 & ~n9922;
  assign n9924 = n7458 & ~n9923;
  assign n9925 = ~P3_INSTADDRPOINTER_REG_27_ & n9851;
  assign n9926 = P3_INSTADDRPOINTER_REG_27_ & ~n9851;
  assign n9927 = ~n9925 & ~n9926;
  assign n9928 = n7460 & ~n9927;
  assign n9929 = ~n9924 & ~n9928;
  assign n9930 = P3_INSTADDRPOINTER_REG_26_ & n9855;
  assign n9931 = ~P3_INSTADDRPOINTER_REG_27_ & n9930;
  assign n9932 = P3_INSTADDRPOINTER_REG_27_ & ~n9930;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = ~n5547 & ~n9933;
  assign n9935 = n5657 & ~n9933;
  assign n9936 = n5500 & ~n9933;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = P3_INSTADDRPOINTER_REG_26_ & n9863;
  assign n9939 = ~P3_INSTADDRPOINTER_REG_27_ & n9938;
  assign n9940 = P3_INSTADDRPOINTER_REG_27_ & ~n9938;
  assign n9941 = ~n9939 & ~n9940;
  assign n9942 = n5618 & ~n9941;
  assign n9943 = n5619_1 & ~n9941;
  assign n9944 = n7361 & ~n9933;
  assign n9945 = n5434_1 & ~n9941;
  assign n9946 = n9818 & n9837;
  assign n9947 = P3_INSTADDRPOINTER_REG_27_ & ~n9946;
  assign n9948 = ~P3_INSTADDRPOINTER_REG_27_ & n9946;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = n7364 & ~n9949;
  assign n9951 = ~n9945 & ~n9950;
  assign n9952 = ~n9942 & ~n9943;
  assign n9953 = ~n9944 & n9952;
  assign n9954 = n9951 & n9953;
  assign n9955 = P3_INSTADDRPOINTER_REG_26_ & n9880;
  assign n9956 = ~P3_INSTADDRPOINTER_REG_27_ & n9955;
  assign n9957 = P3_INSTADDRPOINTER_REG_27_ & ~n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = n5458 & ~n9958;
  assign n9960 = n5450 & ~n9958;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = n5360 & ~n9941;
  assign n9963 = n5438 & ~n9941;
  assign n9964 = n5442 & ~n9941;
  assign n9965 = ~n9962 & ~n9963;
  assign n9966 = ~n9964 & n9965;
  assign n9967 = ~P3_INSTADDRPOINTER_REG_27_ & n9893;
  assign n9968 = P3_INSTADDRPOINTER_REG_27_ & ~n9893;
  assign n9969 = ~n9967 & ~n9968;
  assign n9970 = n5461 & ~n9969;
  assign n9971 = n7477 & ~n9933;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = n7466 & ~n9933;
  assign n9974 = n7470 & ~n9933;
  assign n9975 = n5504_1 & ~n9933;
  assign n9976 = ~n9973 & ~n9974;
  assign n9977 = ~n9975 & n9976;
  assign n9978 = n9961 & n9966;
  assign n9979 = n9972 & n9978;
  assign n9980 = n9977 & n9979;
  assign n9981 = n9929 & ~n9934;
  assign n9982 = n9937 & n9981;
  assign n9983 = n9954 & n9982;
  assign n9984 = n9980 & n9983;
  assign n9985 = n7353 & ~n9984;
  assign n9986 = ~n9913 & ~n9914;
  assign n1800 = n9985 | ~n9986;
  assign n9988 = P3_INSTADDRPOINTER_REG_28_ & n7352;
  assign n9989 = P3_REIP_REG_28_ & n7497;
  assign n9990 = P3_INSTADDRPOINTER_REG_27_ & P3_INSTADDRPOINTER_REG_28_;
  assign n9991 = ~n9917 & n9990;
  assign n9992 = n8303 & ~n9991;
  assign n9993 = P3_INSTADDRPOINTER_REG_28_ & ~n8303;
  assign n9994 = ~P3_INSTADDRPOINTER_REG_27_ & ~n9799;
  assign n9995 = ~n9836 & n9994;
  assign n9996 = ~n9916 & n9995;
  assign n9997 = ~n9992 & ~n9993;
  assign n9998 = ~n9996 & n9997;
  assign n9999 = P3_INSTADDRPOINTER_REG_28_ & n9996;
  assign n10000 = ~n8303 & ~n9999;
  assign n10001 = P3_INSTADDRPOINTER_REG_28_ & n8303;
  assign n10002 = P3_INSTADDRPOINTER_REG_27_ & ~n9917;
  assign n10003 = ~n10000 & ~n10001;
  assign n10004 = ~n10002 & n10003;
  assign n10005 = ~n9998 & ~n10004;
  assign n10006 = n7458 & n10005;
  assign n10007 = P3_INSTADDRPOINTER_REG_27_ & n9851;
  assign n10008 = ~P3_INSTADDRPOINTER_REG_28_ & ~n10007;
  assign n10009 = n9851 & n9990;
  assign n10010 = ~n10008 & ~n10009;
  assign n10011 = n7460 & n10010;
  assign n10012 = ~n10006 & ~n10011;
  assign n10013 = P3_INSTADDRPOINTER_REG_27_ & n9930;
  assign n10014 = ~P3_INSTADDRPOINTER_REG_28_ & n10013;
  assign n10015 = P3_INSTADDRPOINTER_REG_28_ & ~n10013;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = ~n5547 & ~n10016;
  assign n10018 = n5657 & ~n10016;
  assign n10019 = n5500 & ~n10016;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = P3_INSTADDRPOINTER_REG_27_ & n9938;
  assign n10022 = ~P3_INSTADDRPOINTER_REG_28_ & n10021;
  assign n10023 = P3_INSTADDRPOINTER_REG_28_ & ~n10021;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n5618 & ~n10024;
  assign n10026 = n5619_1 & ~n10024;
  assign n10027 = n7361 & ~n10016;
  assign n10028 = n5434_1 & ~n10024;
  assign n10029 = P3_INSTADDRPOINTER_REG_27_ & n9946;
  assign n10030 = ~P3_INSTADDRPOINTER_REG_28_ & n10029;
  assign n10031 = P3_INSTADDRPOINTER_REG_28_ & ~n10029;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = n7364 & ~n10032;
  assign n10034 = ~n10028 & ~n10033;
  assign n10035 = ~n10025 & ~n10026;
  assign n10036 = ~n10027 & n10035;
  assign n10037 = n10034 & n10036;
  assign n10038 = P3_INSTADDRPOINTER_REG_27_ & n9955;
  assign n10039 = ~P3_INSTADDRPOINTER_REG_28_ & n10038;
  assign n10040 = P3_INSTADDRPOINTER_REG_28_ & ~n10038;
  assign n10041 = ~n10039 & ~n10040;
  assign n10042 = n5458 & ~n10041;
  assign n10043 = n5450 & ~n10041;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = n5360 & ~n10024;
  assign n10046 = n5438 & ~n10024;
  assign n10047 = n5442 & ~n10024;
  assign n10048 = ~n10045 & ~n10046;
  assign n10049 = ~n10047 & n10048;
  assign n10050 = P3_INSTADDRPOINTER_REG_27_ & n9893;
  assign n10051 = ~P3_INSTADDRPOINTER_REG_28_ & ~n10050;
  assign n10052 = n9893 & n9990;
  assign n10053 = ~n10051 & ~n10052;
  assign n10054 = n5461 & n10053;
  assign n10055 = n7477 & ~n10016;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = n7466 & ~n10016;
  assign n10058 = n7470 & ~n10016;
  assign n10059 = n5504_1 & ~n10016;
  assign n10060 = ~n10057 & ~n10058;
  assign n10061 = ~n10059 & n10060;
  assign n10062 = n10044 & n10049;
  assign n10063 = n10056 & n10062;
  assign n10064 = n10061 & n10063;
  assign n10065 = n10012 & ~n10017;
  assign n10066 = n10020 & n10065;
  assign n10067 = n10037 & n10066;
  assign n10068 = n10064 & n10067;
  assign n10069 = n7353 & ~n10068;
  assign n10070 = ~n9988 & ~n9989;
  assign n1805 = n10069 | ~n10070;
  assign n10072 = P3_INSTADDRPOINTER_REG_29_ & n7352;
  assign n10073 = P3_REIP_REG_29_ & n7497;
  assign n10074 = ~n8303 & ~n9996;
  assign n10075 = ~n9993 & ~n10074;
  assign n10076 = ~n9991 & n10075;
  assign n10077 = P3_INSTADDRPOINTER_REG_29_ & n8303;
  assign n10078 = ~P3_INSTADDRPOINTER_REG_29_ & ~n8303;
  assign n10079 = ~n10077 & ~n10078;
  assign n10080 = n10076 & ~n10079;
  assign n10081 = ~n10076 & n10079;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = n7458 & ~n10082;
  assign n10084 = ~P3_INSTADDRPOINTER_REG_29_ & ~n10009;
  assign n10085 = P3_INSTADDRPOINTER_REG_29_ & n10009;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = n7460 & n10086;
  assign n10088 = ~n10083 & ~n10087;
  assign n10089 = P3_INSTADDRPOINTER_REG_28_ & n10013;
  assign n10090 = ~P3_INSTADDRPOINTER_REG_29_ & n10089;
  assign n10091 = P3_INSTADDRPOINTER_REG_29_ & ~n10089;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = ~n5547 & ~n10092;
  assign n10094 = n5657 & ~n10092;
  assign n10095 = n5500 & ~n10092;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = P3_INSTADDRPOINTER_REG_28_ & n10021;
  assign n10098 = ~P3_INSTADDRPOINTER_REG_29_ & n10097;
  assign n10099 = P3_INSTADDRPOINTER_REG_29_ & ~n10097;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = n5618 & ~n10100;
  assign n10102 = n5619_1 & ~n10100;
  assign n10103 = n7361 & ~n10092;
  assign n10104 = n5434_1 & ~n10100;
  assign n10105 = n9946 & n9990;
  assign n10106 = P3_INSTADDRPOINTER_REG_29_ & ~n10105;
  assign n10107 = ~P3_INSTADDRPOINTER_REG_29_ & n10105;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = n7364 & ~n10108;
  assign n10110 = ~n10104 & ~n10109;
  assign n10111 = ~n10101 & ~n10102;
  assign n10112 = ~n10103 & n10111;
  assign n10113 = n10110 & n10112;
  assign n10114 = P3_INSTADDRPOINTER_REG_28_ & n10038;
  assign n10115 = ~P3_INSTADDRPOINTER_REG_29_ & n10114;
  assign n10116 = P3_INSTADDRPOINTER_REG_29_ & ~n10114;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = n5458 & ~n10117;
  assign n10119 = n5450 & ~n10117;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = n5360 & ~n10100;
  assign n10122 = n5438 & ~n10100;
  assign n10123 = n5442 & ~n10100;
  assign n10124 = ~n10121 & ~n10122;
  assign n10125 = ~n10123 & n10124;
  assign n10126 = ~P3_INSTADDRPOINTER_REG_29_ & ~n10052;
  assign n10127 = P3_INSTADDRPOINTER_REG_29_ & n10052;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = n5461 & n10128;
  assign n10130 = n7477 & ~n10092;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = n7466 & ~n10092;
  assign n10133 = n7470 & ~n10092;
  assign n10134 = n5504_1 & ~n10092;
  assign n10135 = ~n10132 & ~n10133;
  assign n10136 = ~n10134 & n10135;
  assign n10137 = n10120 & n10125;
  assign n10138 = n10131 & n10137;
  assign n10139 = n10136 & n10138;
  assign n10140 = n10088 & ~n10093;
  assign n10141 = n10096 & n10140;
  assign n10142 = n10113 & n10141;
  assign n10143 = n10139 & n10142;
  assign n10144 = n7353 & ~n10143;
  assign n10145 = ~n10072 & ~n10073;
  assign n1810 = n10144 | ~n10145;
  assign n10147 = P3_INSTADDRPOINTER_REG_30_ & n7352;
  assign n10148 = P3_REIP_REG_30_ & n7497;
  assign n10149 = P3_INSTADDRPOINTER_REG_30_ & n8303;
  assign n10150 = ~P3_INSTADDRPOINTER_REG_30_ & ~n8303;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = P3_INSTADDRPOINTER_REG_29_ & ~n10076;
  assign n10153 = ~n8303 & ~n10076;
  assign n10154 = P3_INSTADDRPOINTER_REG_29_ & ~n8303;
  assign n10155 = ~n10152 & ~n10153;
  assign n10156 = ~n10154 & n10155;
  assign n10157 = ~n10151 & n10156;
  assign n10158 = n10151 & ~n10156;
  assign n10159 = ~n10157 & ~n10158;
  assign n10160 = n7458 & ~n10159;
  assign n10161 = ~P3_INSTADDRPOINTER_REG_30_ & n10085;
  assign n10162 = P3_INSTADDRPOINTER_REG_30_ & ~n10085;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = n7460 & ~n10163;
  assign n10165 = ~n10160 & ~n10164;
  assign n10166 = P3_INSTADDRPOINTER_REG_29_ & n10089;
  assign n10167 = ~P3_INSTADDRPOINTER_REG_30_ & n10166;
  assign n10168 = P3_INSTADDRPOINTER_REG_30_ & ~n10166;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~n5547 & ~n10169;
  assign n10171 = n5657 & ~n10169;
  assign n10172 = n5500 & ~n10169;
  assign n10173 = ~n10171 & ~n10172;
  assign n10174 = P3_INSTADDRPOINTER_REG_29_ & n10097;
  assign n10175 = ~P3_INSTADDRPOINTER_REG_30_ & n10174;
  assign n10176 = P3_INSTADDRPOINTER_REG_30_ & ~n10174;
  assign n10177 = ~n10175 & ~n10176;
  assign n10178 = n5618 & ~n10177;
  assign n10179 = n5619_1 & ~n10177;
  assign n10180 = n7361 & ~n10169;
  assign n10181 = n5434_1 & ~n10177;
  assign n10182 = P3_INSTADDRPOINTER_REG_29_ & n10105;
  assign n10183 = ~P3_INSTADDRPOINTER_REG_30_ & n10182;
  assign n10184 = P3_INSTADDRPOINTER_REG_30_ & ~n10182;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = n7364 & ~n10185;
  assign n10187 = ~n10181 & ~n10186;
  assign n10188 = ~n10178 & ~n10179;
  assign n10189 = ~n10180 & n10188;
  assign n10190 = n10187 & n10189;
  assign n10191 = P3_INSTADDRPOINTER_REG_29_ & n10114;
  assign n10192 = ~P3_INSTADDRPOINTER_REG_30_ & n10191;
  assign n10193 = P3_INSTADDRPOINTER_REG_30_ & ~n10191;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = n5458 & ~n10194;
  assign n10196 = n5450 & ~n10194;
  assign n10197 = ~n10195 & ~n10196;
  assign n10198 = n5360 & ~n10177;
  assign n10199 = n5438 & ~n10177;
  assign n10200 = n5442 & ~n10177;
  assign n10201 = ~n10198 & ~n10199;
  assign n10202 = ~n10200 & n10201;
  assign n10203 = ~P3_INSTADDRPOINTER_REG_30_ & n10127;
  assign n10204 = P3_INSTADDRPOINTER_REG_30_ & ~n10127;
  assign n10205 = ~n10203 & ~n10204;
  assign n10206 = n5461 & ~n10205;
  assign n10207 = n7477 & ~n10169;
  assign n10208 = ~n10206 & ~n10207;
  assign n10209 = n7466 & ~n10169;
  assign n10210 = n7470 & ~n10169;
  assign n10211 = n5504_1 & ~n10169;
  assign n10212 = ~n10209 & ~n10210;
  assign n10213 = ~n10211 & n10212;
  assign n10214 = n10197 & n10202;
  assign n10215 = n10208 & n10214;
  assign n10216 = n10213 & n10215;
  assign n10217 = n10165 & ~n10170;
  assign n10218 = n10173 & n10217;
  assign n10219 = n10190 & n10218;
  assign n10220 = n10216 & n10219;
  assign n10221 = n7353 & ~n10220;
  assign n10222 = ~n10147 & ~n10148;
  assign n1815 = n10221 | ~n10222;
  assign n10224 = P3_INSTADDRPOINTER_REG_31_ & n7352;
  assign n10225 = P3_REIP_REG_31_ & n7497;
  assign n10226 = P3_INSTADDRPOINTER_REG_30_ & n10127;
  assign n10227 = ~P3_INSTADDRPOINTER_REG_31_ & n10226;
  assign n10228 = P3_INSTADDRPOINTER_REG_31_ & ~n10226;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = n5461 & ~n10229;
  assign n10231 = P3_INSTADDRPOINTER_REG_30_ & n10166;
  assign n10232 = ~P3_INSTADDRPOINTER_REG_31_ & n10231;
  assign n10233 = P3_INSTADDRPOINTER_REG_31_ & ~n10231;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = n7477 & ~n10234;
  assign n10236 = n5504_1 & ~n10234;
  assign n10237 = ~n10235 & ~n10236;
  assign n10238 = P3_INSTADDRPOINTER_REG_30_ & n10174;
  assign n10239 = ~P3_INSTADDRPOINTER_REG_31_ & n10238;
  assign n10240 = P3_INSTADDRPOINTER_REG_31_ & ~n10238;
  assign n10241 = ~n10239 & ~n10240;
  assign n10242 = n5442 & ~n10241;
  assign n10243 = n5360 & ~n10241;
  assign n10244 = P3_INSTADDRPOINTER_REG_30_ & n10191;
  assign n10245 = ~P3_INSTADDRPOINTER_REG_31_ & n10244;
  assign n10246 = P3_INSTADDRPOINTER_REG_31_ & ~n10244;
  assign n10247 = ~n10245 & ~n10246;
  assign n10248 = n5450 & ~n10247;
  assign n10249 = ~n10242 & ~n10243;
  assign n10250 = ~n10248 & n10249;
  assign n10251 = n7466 & ~n10234;
  assign n10252 = n7470 & ~n10234;
  assign n10253 = n5458 & ~n10247;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = n10250 & ~n10251;
  assign n10256 = n10254 & n10255;
  assign n10257 = ~n10224 & ~n10225;
  assign n10258 = ~n10230 & n10257;
  assign n10259 = n10237 & n10258;
  assign n10260 = n10256 & n10259;
  assign n10261 = P3_INSTADDRPOINTER_REG_30_ & P3_INSTADDRPOINTER_REG_31_;
  assign n10262 = ~n10156 & n10261;
  assign n10263 = n8303 & ~n10262;
  assign n10264 = P3_INSTADDRPOINTER_REG_31_ & ~n8303;
  assign n10265 = ~P3_INSTADDRPOINTER_REG_30_ & n10156;
  assign n10266 = ~n10263 & ~n10264;
  assign n10267 = ~n10265 & n10266;
  assign n10268 = ~P3_INSTADDRPOINTER_REG_30_ & P3_INSTADDRPOINTER_REG_31_;
  assign n10269 = ~n10154 & n10268;
  assign n10270 = ~n10153 & n10269;
  assign n10271 = ~n8303 & ~n10270;
  assign n10272 = P3_INSTADDRPOINTER_REG_31_ & n8303;
  assign n10273 = P3_INSTADDRPOINTER_REG_30_ & ~n10156;
  assign n10274 = ~n10271 & ~n10272;
  assign n10275 = ~n10273 & n10274;
  assign n10276 = ~n10267 & ~n10275;
  assign n10277 = n7458 & n10276;
  assign n10278 = P3_INSTADDRPOINTER_REG_30_ & n10085;
  assign n10279 = ~P3_INSTADDRPOINTER_REG_31_ & n10278;
  assign n10280 = P3_INSTADDRPOINTER_REG_31_ & ~n10278;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n7460 & ~n10281;
  assign n10283 = ~n10277 & ~n10282;
  assign n10284 = ~n5547 & ~n10234;
  assign n10285 = n5657 & ~n10234;
  assign n10286 = n5500 & ~n10234;
  assign n10287 = ~n10285 & ~n10286;
  assign n10288 = n5619_1 & ~n10241;
  assign n10289 = n10287 & ~n10288;
  assign n10290 = n7361 & ~n10234;
  assign n10291 = n5618 & ~n10241;
  assign n10292 = n5438 & ~n10241;
  assign n10293 = n5434_1 & ~n10241;
  assign n10294 = P3_INSTADDRPOINTER_REG_30_ & n10182;
  assign n10295 = ~P3_INSTADDRPOINTER_REG_31_ & n10294;
  assign n10296 = P3_INSTADDRPOINTER_REG_31_ & ~n10294;
  assign n10297 = ~n10295 & ~n10296;
  assign n10298 = n7364 & ~n10297;
  assign n10299 = ~n10292 & ~n10293;
  assign n10300 = ~n10298 & n10299;
  assign n10301 = ~n10290 & ~n10291;
  assign n10302 = n10300 & n10301;
  assign n10303 = n10283 & ~n10284;
  assign n10304 = n10289 & n10303;
  assign n10305 = n10302 & n10304;
  assign n10306 = n10260 & n10305;
  assign n10307 = ~n7353 & ~n10224;
  assign n10308 = ~n10225 & n10307;
  assign n1820 = ~n10306 & ~n10308;
  assign n10310 = P3_STATE2_REG_0_ & ~n5327;
  assign n10311 = ~P3_STATE2_REG_0_ & ~n7320;
  assign n10312 = n5461 & n5464_1;
  assign n10313 = n5466 & n5470;
  assign n10314 = ~n10312 & ~n10313;
  assign n10315 = n5713 & ~n10314;
  assign n10316 = ~n10311 & ~n10315;
  assign n10317 = n10310 & ~n10316;
  assign n10318 = ~n7457 & n10317;
  assign n10319 = ~n7426 & n10318;
  assign n10320 = n7457 & n10317;
  assign n10321 = ~n7426 & n10320;
  assign n10322 = P3_STATE2_REG_1_ & ~n10316;
  assign n10323 = P3_STATEBS16_REG & n10322;
  assign n10324 = P3_PHYADDRPOINTER_REG_0_ & n10323;
  assign n10325 = ~P3_STATEBS16_REG & n10322;
  assign n10326 = P3_PHYADDRPOINTER_REG_0_ & n10325;
  assign n10327 = P3_PHYADDRPOINTER_REG_0_ & n10316;
  assign n10328 = P3_STATE2_REG_0_ & n5327;
  assign n10329 = ~n10316 & n10328;
  assign n10330 = ~n7474 & n10329;
  assign n10331 = P3_STATE2_REG_2_ & ~P3_STATE2_REG_0_;
  assign n10332 = ~n10316 & n10331;
  assign n10333 = P3_PHYADDRPOINTER_REG_0_ & n10332;
  assign n10334 = n5729_1 & ~n10316;
  assign n10335 = P3_REIP_REG_0_ & n10334;
  assign n10336 = ~n10327 & ~n10330;
  assign n10337 = ~n10333 & n10336;
  assign n10338 = ~n10335 & n10337;
  assign n10339 = ~n10319 & ~n10321;
  assign n10340 = ~n10324 & n10339;
  assign n10341 = ~n10326 & n10340;
  assign n1825 = ~n10338 | ~n10341;
  assign n10343 = ~n7548 & n10318;
  assign n10344 = ~n7548 & n10320;
  assign n10345 = P3_PHYADDRPOINTER_REG_1_ & n10323;
  assign n10346 = ~P3_PHYADDRPOINTER_REG_1_ & n10325;
  assign n10347 = P3_PHYADDRPOINTER_REG_1_ & n10316;
  assign n10348 = ~n7578 & n10329;
  assign n10349 = ~P3_PHYADDRPOINTER_REG_1_ & n10332;
  assign n10350 = P3_REIP_REG_1_ & n10334;
  assign n10351 = ~n10347 & ~n10348;
  assign n10352 = ~n10349 & n10351;
  assign n10353 = ~n10350 & n10352;
  assign n10354 = ~n10343 & ~n10344;
  assign n10355 = ~n10345 & n10354;
  assign n10356 = ~n10346 & n10355;
  assign n1830 = ~n10353 | ~n10356;
  assign n10358 = ~n7675 & n10318;
  assign n10359 = ~n7661 & n10320;
  assign n10360 = ~P3_PHYADDRPOINTER_REG_2_ & n10323;
  assign n10361 = P3_PHYADDRPOINTER_REG_1_ & ~P3_PHYADDRPOINTER_REG_2_;
  assign n10362 = ~P3_PHYADDRPOINTER_REG_1_ & P3_PHYADDRPOINTER_REG_2_;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = n10325 & ~n10363;
  assign n10365 = n10332 & ~n10363;
  assign n10366 = P3_REIP_REG_2_ & n10334;
  assign n10367 = P3_PHYADDRPOINTER_REG_2_ & n10316;
  assign n10368 = ~n7712 & n10329;
  assign n10369 = ~n10365 & ~n10366;
  assign n10370 = ~n10367 & n10369;
  assign n10371 = ~n10368 & n10370;
  assign n10372 = ~n10358 & ~n10359;
  assign n10373 = ~n10360 & n10372;
  assign n10374 = ~n10364 & n10373;
  assign n1835 = ~n10371 | ~n10374;
  assign n10376 = ~n7795 & n10318;
  assign n10377 = n7810 & n10320;
  assign n10378 = P3_PHYADDRPOINTER_REG_2_ & ~P3_PHYADDRPOINTER_REG_3_;
  assign n10379 = ~P3_PHYADDRPOINTER_REG_2_ & P3_PHYADDRPOINTER_REG_3_;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = n10323 & ~n10380;
  assign n10382 = P3_PHYADDRPOINTER_REG_1_ & P3_PHYADDRPOINTER_REG_2_;
  assign n10383 = ~P3_PHYADDRPOINTER_REG_3_ & n10382;
  assign n10384 = P3_PHYADDRPOINTER_REG_3_ & ~n10382;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = n10325 & ~n10385;
  assign n10387 = n10332 & ~n10385;
  assign n10388 = P3_REIP_REG_3_ & n10334;
  assign n10389 = P3_PHYADDRPOINTER_REG_3_ & n10316;
  assign n10390 = n7848 & n10329;
  assign n10391 = ~n10387 & ~n10388;
  assign n10392 = ~n10389 & n10391;
  assign n10393 = ~n10390 & n10392;
  assign n10394 = ~n10376 & ~n10377;
  assign n10395 = ~n10381 & n10394;
  assign n10396 = ~n10386 & n10395;
  assign n1840 = ~n10393 | ~n10396;
  assign n10398 = P3_PHYADDRPOINTER_REG_2_ & P3_PHYADDRPOINTER_REG_3_;
  assign n10399 = ~P3_PHYADDRPOINTER_REG_4_ & n10398;
  assign n10400 = P3_PHYADDRPOINTER_REG_4_ & ~n10398;
  assign n10401 = ~n10399 & ~n10400;
  assign n10402 = n10323 & ~n10401;
  assign n10403 = P3_PHYADDRPOINTER_REG_3_ & n10382;
  assign n10404 = ~P3_PHYADDRPOINTER_REG_4_ & n10403;
  assign n10405 = P3_PHYADDRPOINTER_REG_4_ & ~n10403;
  assign n10406 = ~n10404 & ~n10405;
  assign n10407 = n10325 & ~n10406;
  assign n10408 = n7927 & n10320;
  assign n10409 = ~n7949 & n10318;
  assign n10410 = n10332 & ~n10406;
  assign n10411 = P3_REIP_REG_4_ & n10334;
  assign n10412 = P3_PHYADDRPOINTER_REG_4_ & n10316;
  assign n10413 = ~n7988 & n10329;
  assign n10414 = ~n10410 & ~n10411;
  assign n10415 = ~n10412 & n10414;
  assign n10416 = ~n10413 & n10415;
  assign n10417 = ~n10402 & ~n10407;
  assign n10418 = ~n10408 & n10417;
  assign n10419 = ~n10409 & n10418;
  assign n1845 = ~n10416 | ~n10419;
  assign n10421 = P3_PHYADDRPOINTER_REG_4_ & n10398;
  assign n10422 = ~P3_PHYADDRPOINTER_REG_5_ & n10421;
  assign n10423 = P3_PHYADDRPOINTER_REG_5_ & ~n10421;
  assign n10424 = ~n10422 & ~n10423;
  assign n10425 = n10323 & ~n10424;
  assign n10426 = P3_PHYADDRPOINTER_REG_4_ & n10403;
  assign n10427 = ~P3_PHYADDRPOINTER_REG_5_ & n10426;
  assign n10428 = P3_PHYADDRPOINTER_REG_5_ & ~n10426;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = n10325 & ~n10429;
  assign n10431 = ~n8069 & n10318;
  assign n10432 = ~n8087 & n10320;
  assign n10433 = n10332 & ~n10429;
  assign n10434 = P3_REIP_REG_5_ & n10334;
  assign n10435 = P3_PHYADDRPOINTER_REG_5_ & n10316;
  assign n10436 = n8126 & n10329;
  assign n10437 = ~n10433 & ~n10434;
  assign n10438 = ~n10435 & n10437;
  assign n10439 = ~n10436 & n10438;
  assign n10440 = ~n10425 & ~n10430;
  assign n10441 = ~n10431 & n10440;
  assign n10442 = ~n10432 & n10441;
  assign n1850 = ~n10439 | ~n10442;
  assign n10444 = P3_PHYADDRPOINTER_REG_5_ & n10421;
  assign n10445 = ~P3_PHYADDRPOINTER_REG_6_ & n10444;
  assign n10446 = P3_PHYADDRPOINTER_REG_6_ & ~n10444;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = n10323 & ~n10447;
  assign n10449 = P3_PHYADDRPOINTER_REG_5_ & n10426;
  assign n10450 = ~P3_PHYADDRPOINTER_REG_6_ & n10449;
  assign n10451 = P3_PHYADDRPOINTER_REG_6_ & ~n10449;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = n10325 & ~n10452;
  assign n10454 = ~n8204 & n10318;
  assign n10455 = ~n8223 & n10320;
  assign n10456 = n10332 & ~n10452;
  assign n10457 = P3_REIP_REG_6_ & n10334;
  assign n10458 = P3_PHYADDRPOINTER_REG_6_ & n10316;
  assign n10459 = ~n8261 & n10329;
  assign n10460 = ~n10456 & ~n10457;
  assign n10461 = ~n10458 & n10460;
  assign n10462 = ~n10459 & n10461;
  assign n10463 = ~n10448 & ~n10453;
  assign n10464 = ~n10454 & n10463;
  assign n10465 = ~n10455 & n10464;
  assign n1855 = ~n10462 | ~n10465;
  assign n10467 = P3_PHYADDRPOINTER_REG_6_ & n10444;
  assign n10468 = ~P3_PHYADDRPOINTER_REG_7_ & n10467;
  assign n10469 = P3_PHYADDRPOINTER_REG_7_ & ~n10467;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = n10323 & ~n10470;
  assign n10472 = P3_PHYADDRPOINTER_REG_6_ & n10449;
  assign n10473 = ~P3_PHYADDRPOINTER_REG_7_ & n10472;
  assign n10474 = P3_PHYADDRPOINTER_REG_7_ & ~n10472;
  assign n10475 = ~n10473 & ~n10474;
  assign n10476 = n10325 & ~n10475;
  assign n10477 = ~n8310 & n10318;
  assign n10478 = ~n8328 & n10320;
  assign n10479 = n10332 & ~n10475;
  assign n10480 = P3_REIP_REG_7_ & n10334;
  assign n10481 = P3_PHYADDRPOINTER_REG_7_ & n10316;
  assign n10482 = ~n8364 & n10329;
  assign n10483 = ~n10479 & ~n10480;
  assign n10484 = ~n10481 & n10483;
  assign n10485 = ~n10482 & n10484;
  assign n10486 = ~n10471 & ~n10476;
  assign n10487 = ~n10477 & n10486;
  assign n10488 = ~n10478 & n10487;
  assign n1860 = ~n10485 | ~n10488;
  assign n10490 = P3_PHYADDRPOINTER_REG_7_ & n10467;
  assign n10491 = ~P3_PHYADDRPOINTER_REG_8_ & n10490;
  assign n10492 = P3_PHYADDRPOINTER_REG_8_ & ~n10490;
  assign n10493 = ~n10491 & ~n10492;
  assign n10494 = n10323 & ~n10493;
  assign n10495 = P3_PHYADDRPOINTER_REG_7_ & n10472;
  assign n10496 = ~P3_PHYADDRPOINTER_REG_8_ & n10495;
  assign n10497 = P3_PHYADDRPOINTER_REG_8_ & ~n10495;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = n10325 & ~n10498;
  assign n10500 = ~n8408 & n10318;
  assign n10501 = ~n8424 & n10320;
  assign n10502 = n10332 & ~n10498;
  assign n10503 = P3_REIP_REG_8_ & n10334;
  assign n10504 = P3_PHYADDRPOINTER_REG_8_ & n10316;
  assign n10505 = ~n8458 & n10329;
  assign n10506 = ~n10502 & ~n10503;
  assign n10507 = ~n10504 & n10506;
  assign n10508 = ~n10505 & n10507;
  assign n10509 = ~n10494 & ~n10499;
  assign n10510 = ~n10500 & n10509;
  assign n10511 = ~n10501 & n10510;
  assign n1865 = ~n10508 | ~n10511;
  assign n10513 = P3_PHYADDRPOINTER_REG_8_ & n10490;
  assign n10514 = ~P3_PHYADDRPOINTER_REG_9_ & n10513;
  assign n10515 = P3_PHYADDRPOINTER_REG_9_ & ~n10513;
  assign n10516 = ~n10514 & ~n10515;
  assign n10517 = n10323 & ~n10516;
  assign n10518 = P3_PHYADDRPOINTER_REG_8_ & n10495;
  assign n10519 = ~P3_PHYADDRPOINTER_REG_9_ & n10518;
  assign n10520 = P3_PHYADDRPOINTER_REG_9_ & ~n10518;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = n10325 & ~n10521;
  assign n10523 = ~n8507 & n10318;
  assign n10524 = n8518 & n10320;
  assign n10525 = n10332 & ~n10521;
  assign n10526 = P3_REIP_REG_9_ & n10334;
  assign n10527 = P3_PHYADDRPOINTER_REG_9_ & n10316;
  assign n10528 = n8547 & n10329;
  assign n10529 = ~n10525 & ~n10526;
  assign n10530 = ~n10527 & n10529;
  assign n10531 = ~n10528 & n10530;
  assign n10532 = ~n10517 & ~n10522;
  assign n10533 = ~n10523 & n10532;
  assign n10534 = ~n10524 & n10533;
  assign n1870 = ~n10531 | ~n10534;
  assign n10536 = P3_PHYADDRPOINTER_REG_9_ & n10513;
  assign n10537 = ~P3_PHYADDRPOINTER_REG_10_ & n10536;
  assign n10538 = P3_PHYADDRPOINTER_REG_10_ & ~n10536;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = n10323 & ~n10539;
  assign n10541 = P3_PHYADDRPOINTER_REG_9_ & n10518;
  assign n10542 = ~P3_PHYADDRPOINTER_REG_10_ & n10541;
  assign n10543 = P3_PHYADDRPOINTER_REG_10_ & ~n10541;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = n10325 & ~n10544;
  assign n10546 = n8585 & n10320;
  assign n10547 = ~n8626 & n10318;
  assign n10548 = n10332 & ~n10544;
  assign n10549 = P3_REIP_REG_10_ & n10334;
  assign n10550 = P3_PHYADDRPOINTER_REG_10_ & n10316;
  assign n10551 = n8609 & n10329;
  assign n10552 = ~n10548 & ~n10549;
  assign n10553 = ~n10550 & n10552;
  assign n10554 = ~n10551 & n10553;
  assign n10555 = ~n10540 & ~n10545;
  assign n10556 = ~n10546 & n10555;
  assign n10557 = ~n10547 & n10556;
  assign n1875 = ~n10554 | ~n10557;
  assign n10559 = P3_PHYADDRPOINTER_REG_10_ & n10536;
  assign n10560 = ~P3_PHYADDRPOINTER_REG_11_ & n10559;
  assign n10561 = P3_PHYADDRPOINTER_REG_11_ & ~n10559;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = n10323 & ~n10562;
  assign n10564 = P3_PHYADDRPOINTER_REG_10_ & n10541;
  assign n10565 = ~P3_PHYADDRPOINTER_REG_11_ & n10564;
  assign n10566 = P3_PHYADDRPOINTER_REG_11_ & ~n10564;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = n10325 & ~n10567;
  assign n10569 = ~n8662 & n10320;
  assign n10570 = ~n8676 & n10318;
  assign n10571 = n10332 & ~n10567;
  assign n10572 = P3_REIP_REG_11_ & n10334;
  assign n10573 = P3_PHYADDRPOINTER_REG_11_ & n10316;
  assign n10574 = ~n8701 & n10329;
  assign n10575 = ~n10571 & ~n10572;
  assign n10576 = ~n10573 & n10575;
  assign n10577 = ~n10574 & n10576;
  assign n10578 = ~n10563 & ~n10568;
  assign n10579 = ~n10569 & n10578;
  assign n10580 = ~n10570 & n10579;
  assign n1880 = ~n10577 | ~n10580;
  assign n10582 = P3_PHYADDRPOINTER_REG_11_ & n10559;
  assign n10583 = ~P3_PHYADDRPOINTER_REG_12_ & n10582;
  assign n10584 = P3_PHYADDRPOINTER_REG_12_ & ~n10582;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = n10323 & ~n10585;
  assign n10587 = P3_PHYADDRPOINTER_REG_11_ & n10564;
  assign n10588 = ~P3_PHYADDRPOINTER_REG_12_ & n10587;
  assign n10589 = P3_PHYADDRPOINTER_REG_12_ & ~n10587;
  assign n10590 = ~n10588 & ~n10589;
  assign n10591 = n10325 & ~n10590;
  assign n10592 = ~n8750 & n10318;
  assign n10593 = n8759 & n10320;
  assign n10594 = P3_PHYADDRPOINTER_REG_12_ & n10316;
  assign n10595 = P3_REIP_REG_12_ & n10334;
  assign n10596 = n10332 & ~n10590;
  assign n10597 = n8785 & n10329;
  assign n10598 = ~n10594 & ~n10595;
  assign n10599 = ~n10596 & n10598;
  assign n10600 = ~n10597 & n10599;
  assign n10601 = ~n10586 & ~n10591;
  assign n10602 = ~n10592 & n10601;
  assign n10603 = ~n10593 & n10602;
  assign n1885 = ~n10600 | ~n10603;
  assign n10605 = P3_PHYADDRPOINTER_REG_12_ & n10582;
  assign n10606 = ~P3_PHYADDRPOINTER_REG_13_ & n10605;
  assign n10607 = P3_PHYADDRPOINTER_REG_13_ & ~n10605;
  assign n10608 = ~n10606 & ~n10607;
  assign n10609 = n10323 & ~n10608;
  assign n10610 = P3_PHYADDRPOINTER_REG_12_ & n10587;
  assign n10611 = ~P3_PHYADDRPOINTER_REG_13_ & n10610;
  assign n10612 = P3_PHYADDRPOINTER_REG_13_ & ~n10610;
  assign n10613 = ~n10611 & ~n10612;
  assign n10614 = n10325 & ~n10613;
  assign n10615 = n8832 & n10318;
  assign n10616 = n8839 & n10320;
  assign n10617 = P3_PHYADDRPOINTER_REG_13_ & n10316;
  assign n10618 = P3_REIP_REG_13_ & n10334;
  assign n10619 = n10332 & ~n10613;
  assign n10620 = n8864 & n10329;
  assign n10621 = ~n10617 & ~n10618;
  assign n10622 = ~n10619 & n10621;
  assign n10623 = ~n10620 & n10622;
  assign n10624 = ~n10609 & ~n10614;
  assign n10625 = ~n10615 & n10624;
  assign n10626 = ~n10616 & n10625;
  assign n1890 = ~n10623 | ~n10626;
  assign n10628 = P3_PHYADDRPOINTER_REG_13_ & n10605;
  assign n10629 = ~P3_PHYADDRPOINTER_REG_14_ & n10628;
  assign n10630 = P3_PHYADDRPOINTER_REG_14_ & ~n10628;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = n10323 & ~n10631;
  assign n10633 = P3_PHYADDRPOINTER_REG_13_ & n10610;
  assign n10634 = ~P3_PHYADDRPOINTER_REG_14_ & n10633;
  assign n10635 = P3_PHYADDRPOINTER_REG_14_ & ~n10633;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = n10325 & ~n10636;
  assign n10638 = ~n8939 & n10318;
  assign n10639 = ~n8943 & n10320;
  assign n10640 = P3_PHYADDRPOINTER_REG_14_ & n10316;
  assign n10641 = P3_REIP_REG_14_ & n10334;
  assign n10642 = n10332 & ~n10636;
  assign n10643 = ~n8908 & n10329;
  assign n10644 = ~n10640 & ~n10641;
  assign n10645 = ~n10642 & n10644;
  assign n10646 = ~n10643 & n10645;
  assign n10647 = ~n10632 & ~n10637;
  assign n10648 = ~n10638 & n10647;
  assign n10649 = ~n10639 & n10648;
  assign n1895 = ~n10646 | ~n10649;
  assign n10651 = P3_PHYADDRPOINTER_REG_14_ & n10628;
  assign n10652 = ~P3_PHYADDRPOINTER_REG_15_ & n10651;
  assign n10653 = P3_PHYADDRPOINTER_REG_15_ & ~n10651;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = n10323 & ~n10654;
  assign n10656 = P3_PHYADDRPOINTER_REG_14_ & n10633;
  assign n10657 = ~P3_PHYADDRPOINTER_REG_15_ & n10656;
  assign n10658 = P3_PHYADDRPOINTER_REG_15_ & ~n10656;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = n10325 & ~n10659;
  assign n10661 = ~n9019 & n10318;
  assign n10662 = n9024 & n10320;
  assign n10663 = P3_PHYADDRPOINTER_REG_15_ & n10316;
  assign n10664 = P3_REIP_REG_15_ & n10334;
  assign n10665 = n10332 & ~n10659;
  assign n10666 = n8988 & n10329;
  assign n10667 = ~n10663 & ~n10664;
  assign n10668 = ~n10665 & n10667;
  assign n10669 = ~n10666 & n10668;
  assign n10670 = ~n10655 & ~n10660;
  assign n10671 = ~n10661 & n10670;
  assign n10672 = ~n10662 & n10671;
  assign n1900 = ~n10669 | ~n10672;
  assign n10674 = P3_PHYADDRPOINTER_REG_15_ & n10651;
  assign n10675 = ~P3_PHYADDRPOINTER_REG_16_ & n10674;
  assign n10676 = P3_PHYADDRPOINTER_REG_16_ & ~n10674;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = n10323 & ~n10677;
  assign n10679 = P3_PHYADDRPOINTER_REG_15_ & n10656;
  assign n10680 = ~P3_PHYADDRPOINTER_REG_16_ & n10679;
  assign n10681 = P3_PHYADDRPOINTER_REG_16_ & ~n10679;
  assign n10682 = ~n10680 & ~n10681;
  assign n10683 = n10325 & ~n10682;
  assign n10684 = ~n9059 & n10320;
  assign n10685 = ~n9073 & n10318;
  assign n10686 = P3_PHYADDRPOINTER_REG_16_ & n10316;
  assign n10687 = P3_REIP_REG_16_ & n10334;
  assign n10688 = n10332 & ~n10682;
  assign n10689 = ~n9098 & n10329;
  assign n10690 = ~n10686 & ~n10687;
  assign n10691 = ~n10688 & n10690;
  assign n10692 = ~n10689 & n10691;
  assign n10693 = ~n10678 & ~n10683;
  assign n10694 = ~n10684 & n10693;
  assign n10695 = ~n10685 & n10694;
  assign n1905 = ~n10692 | ~n10695;
  assign n10697 = P3_PHYADDRPOINTER_REG_16_ & n10674;
  assign n10698 = ~P3_PHYADDRPOINTER_REG_17_ & n10697;
  assign n10699 = P3_PHYADDRPOINTER_REG_17_ & ~n10697;
  assign n10700 = ~n10698 & ~n10699;
  assign n10701 = n10323 & ~n10700;
  assign n10702 = P3_PHYADDRPOINTER_REG_16_ & n10679;
  assign n10703 = ~P3_PHYADDRPOINTER_REG_17_ & n10702;
  assign n10704 = P3_PHYADDRPOINTER_REG_17_ & ~n10702;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = n10325 & ~n10705;
  assign n10707 = n9123 & n10320;
  assign n10708 = n9180 & n10318;
  assign n10709 = P3_PHYADDRPOINTER_REG_17_ & n10316;
  assign n10710 = P3_REIP_REG_17_ & n10334;
  assign n10711 = n10332 & ~n10705;
  assign n10712 = n9152 & n10329;
  assign n10713 = ~n10709 & ~n10710;
  assign n10714 = ~n10711 & n10713;
  assign n10715 = ~n10712 & n10714;
  assign n10716 = ~n10701 & ~n10706;
  assign n10717 = ~n10707 & n10716;
  assign n10718 = ~n10708 & n10717;
  assign n1910 = ~n10715 | ~n10718;
  assign n10720 = P3_PHYADDRPOINTER_REG_17_ & n10697;
  assign n10721 = ~P3_PHYADDRPOINTER_REG_18_ & n10720;
  assign n10722 = P3_PHYADDRPOINTER_REG_18_ & ~n10720;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = n10323 & ~n10723;
  assign n10725 = P3_PHYADDRPOINTER_REG_17_ & n10702;
  assign n10726 = ~P3_PHYADDRPOINTER_REG_18_ & n10725;
  assign n10727 = P3_PHYADDRPOINTER_REG_18_ & ~n10725;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = n10325 & ~n10728;
  assign n10730 = ~n9219 & n10320;
  assign n10731 = ~n9232 & n10318;
  assign n10732 = P3_PHYADDRPOINTER_REG_18_ & n10316;
  assign n10733 = P3_REIP_REG_18_ & n10334;
  assign n10734 = n10332 & ~n10728;
  assign n10735 = ~n9257 & n10329;
  assign n10736 = ~n10732 & ~n10733;
  assign n10737 = ~n10734 & n10736;
  assign n10738 = ~n10735 & n10737;
  assign n10739 = ~n10724 & ~n10729;
  assign n10740 = ~n10730 & n10739;
  assign n10741 = ~n10731 & n10740;
  assign n1915 = ~n10738 | ~n10741;
  assign n10743 = P3_PHYADDRPOINTER_REG_18_ & n10720;
  assign n10744 = ~P3_PHYADDRPOINTER_REG_19_ & n10743;
  assign n10745 = P3_PHYADDRPOINTER_REG_19_ & ~n10743;
  assign n10746 = ~n10744 & ~n10745;
  assign n10747 = n10323 & ~n10746;
  assign n10748 = P3_PHYADDRPOINTER_REG_18_ & n10725;
  assign n10749 = ~P3_PHYADDRPOINTER_REG_19_ & n10748;
  assign n10750 = P3_PHYADDRPOINTER_REG_19_ & ~n10748;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = n10325 & ~n10751;
  assign n10753 = n9282 & n10320;
  assign n10754 = ~n9338 & n10318;
  assign n10755 = P3_PHYADDRPOINTER_REG_19_ & n10316;
  assign n10756 = P3_REIP_REG_19_ & n10334;
  assign n10757 = n10332 & ~n10751;
  assign n10758 = n9311 & n10329;
  assign n10759 = ~n10755 & ~n10756;
  assign n10760 = ~n10757 & n10759;
  assign n10761 = ~n10758 & n10760;
  assign n10762 = ~n10747 & ~n10752;
  assign n10763 = ~n10753 & n10762;
  assign n10764 = ~n10754 & n10763;
  assign n1920 = ~n10761 | ~n10764;
  assign n10766 = P3_PHYADDRPOINTER_REG_19_ & n10743;
  assign n10767 = ~P3_PHYADDRPOINTER_REG_20_ & n10766;
  assign n10768 = P3_PHYADDRPOINTER_REG_20_ & ~n10766;
  assign n10769 = ~n10767 & ~n10768;
  assign n10770 = n10323 & ~n10769;
  assign n10771 = P3_PHYADDRPOINTER_REG_19_ & n10748;
  assign n10772 = ~P3_PHYADDRPOINTER_REG_20_ & n10771;
  assign n10773 = P3_PHYADDRPOINTER_REG_20_ & ~n10771;
  assign n10774 = ~n10772 & ~n10773;
  assign n10775 = n10325 & ~n10774;
  assign n10776 = n9396 & n10320;
  assign n10777 = P3_PHYADDRPOINTER_REG_20_ & n10316;
  assign n10778 = P3_REIP_REG_20_ & n10334;
  assign n10779 = n10332 & ~n10774;
  assign n10780 = n9420 & n10329;
  assign n10781 = ~n10777 & ~n10778;
  assign n10782 = ~n10779 & n10781;
  assign n10783 = ~n10780 & n10782;
  assign n10784 = n9367 & n10318;
  assign n10785 = ~n10770 & ~n10775;
  assign n10786 = ~n10776 & n10785;
  assign n10787 = n10783 & n10786;
  assign n1925 = n10784 | ~n10787;
  assign n10789 = P3_PHYADDRPOINTER_REG_20_ & n10766;
  assign n10790 = ~P3_PHYADDRPOINTER_REG_21_ & n10789;
  assign n10791 = P3_PHYADDRPOINTER_REG_21_ & ~n10789;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = n10323 & ~n10792;
  assign n10794 = P3_PHYADDRPOINTER_REG_20_ & n10771;
  assign n10795 = ~P3_PHYADDRPOINTER_REG_21_ & n10794;
  assign n10796 = P3_PHYADDRPOINTER_REG_21_ & ~n10794;
  assign n10797 = ~n10795 & ~n10796;
  assign n10798 = n10325 & ~n10797;
  assign n10799 = n9472 & n10320;
  assign n10800 = P3_PHYADDRPOINTER_REG_21_ & n10316;
  assign n10801 = P3_REIP_REG_21_ & n10334;
  assign n10802 = n10332 & ~n10797;
  assign n10803 = n9497 & n10329;
  assign n10804 = ~n10800 & ~n10801;
  assign n10805 = ~n10802 & n10804;
  assign n10806 = ~n10803 & n10805;
  assign n10807 = ~n9443 & n10318;
  assign n10808 = ~n10793 & ~n10798;
  assign n10809 = ~n10799 & n10808;
  assign n10810 = n10806 & n10809;
  assign n1930 = n10807 | ~n10810;
  assign n10812 = P3_PHYADDRPOINTER_REG_21_ & n10789;
  assign n10813 = ~P3_PHYADDRPOINTER_REG_22_ & n10812;
  assign n10814 = P3_PHYADDRPOINTER_REG_22_ & ~n10812;
  assign n10815 = ~n10813 & ~n10814;
  assign n10816 = n10323 & ~n10815;
  assign n10817 = P3_PHYADDRPOINTER_REG_21_ & n10794;
  assign n10818 = ~P3_PHYADDRPOINTER_REG_22_ & n10817;
  assign n10819 = P3_PHYADDRPOINTER_REG_22_ & ~n10817;
  assign n10820 = ~n10818 & ~n10819;
  assign n10821 = n10325 & ~n10820;
  assign n10822 = ~n9559 & n10318;
  assign n10823 = ~n9580 & n10320;
  assign n10824 = P3_PHYADDRPOINTER_REG_22_ & n10316;
  assign n10825 = P3_REIP_REG_22_ & n10334;
  assign n10826 = n10332 & ~n10820;
  assign n10827 = ~n9538 & n10329;
  assign n10828 = ~n10824 & ~n10825;
  assign n10829 = ~n10826 & n10828;
  assign n10830 = ~n10827 & n10829;
  assign n10831 = ~n10816 & ~n10821;
  assign n10832 = ~n10822 & n10831;
  assign n10833 = ~n10823 & n10832;
  assign n1935 = ~n10830 | ~n10833;
  assign n10835 = P3_PHYADDRPOINTER_REG_22_ & n10812;
  assign n10836 = ~P3_PHYADDRPOINTER_REG_23_ & n10835;
  assign n10837 = P3_PHYADDRPOINTER_REG_23_ & ~n10835;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = n10323 & ~n10838;
  assign n10840 = P3_PHYADDRPOINTER_REG_22_ & n10817;
  assign n10841 = ~P3_PHYADDRPOINTER_REG_23_ & n10840;
  assign n10842 = P3_PHYADDRPOINTER_REG_23_ & ~n10840;
  assign n10843 = ~n10841 & ~n10842;
  assign n10844 = n10325 & ~n10843;
  assign n10845 = ~n9639 & n10318;
  assign n10846 = n9662 & n10320;
  assign n10847 = P3_PHYADDRPOINTER_REG_23_ & n10316;
  assign n10848 = P3_REIP_REG_23_ & n10334;
  assign n10849 = n10332 & ~n10843;
  assign n10850 = n9621 & n10329;
  assign n10851 = ~n10847 & ~n10848;
  assign n10852 = ~n10849 & n10851;
  assign n10853 = ~n10850 & n10852;
  assign n10854 = ~n10839 & ~n10844;
  assign n10855 = ~n10845 & n10854;
  assign n10856 = ~n10846 & n10855;
  assign n1940 = ~n10853 | ~n10856;
  assign n10858 = P3_PHYADDRPOINTER_REG_23_ & n10835;
  assign n10859 = ~P3_PHYADDRPOINTER_REG_24_ & n10858;
  assign n10860 = P3_PHYADDRPOINTER_REG_24_ & ~n10858;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = n10323 & ~n10861;
  assign n10863 = ~n9719 & n10318;
  assign n10864 = P3_PHYADDRPOINTER_REG_23_ & n10840;
  assign n10865 = ~P3_PHYADDRPOINTER_REG_24_ & n10864;
  assign n10866 = P3_PHYADDRPOINTER_REG_24_ & ~n10864;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = n10325 & ~n10867;
  assign n10869 = ~n9727 & n10320;
  assign n10870 = P3_PHYADDRPOINTER_REG_24_ & n10316;
  assign n10871 = P3_REIP_REG_24_ & n10334;
  assign n10872 = n10332 & ~n10867;
  assign n10873 = ~n9692 & n10329;
  assign n10874 = ~n10870 & ~n10871;
  assign n10875 = ~n10872 & n10874;
  assign n10876 = ~n10873 & n10875;
  assign n10877 = ~n10862 & ~n10863;
  assign n10878 = ~n10868 & n10877;
  assign n10879 = ~n10869 & n10878;
  assign n1945 = ~n10876 | ~n10879;
  assign n10881 = P3_PHYADDRPOINTER_REG_24_ & n10858;
  assign n10882 = ~P3_PHYADDRPOINTER_REG_25_ & n10881;
  assign n10883 = P3_PHYADDRPOINTER_REG_25_ & ~n10881;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = n10323 & ~n10884;
  assign n10886 = ~n9802 & n10318;
  assign n10887 = P3_PHYADDRPOINTER_REG_24_ & n10864;
  assign n10888 = ~P3_PHYADDRPOINTER_REG_25_ & n10887;
  assign n10889 = P3_PHYADDRPOINTER_REG_25_ & ~n10887;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = n10325 & ~n10890;
  assign n10892 = n9808 & n10320;
  assign n10893 = P3_PHYADDRPOINTER_REG_25_ & n10316;
  assign n10894 = P3_REIP_REG_25_ & n10334;
  assign n10895 = n10332 & ~n10890;
  assign n10896 = n9772 & n10329;
  assign n10897 = ~n10893 & ~n10894;
  assign n10898 = ~n10895 & n10897;
  assign n10899 = ~n10896 & n10898;
  assign n10900 = ~n10885 & ~n10886;
  assign n10901 = ~n10891 & n10900;
  assign n10902 = ~n10892 & n10901;
  assign n1950 = ~n10899 | ~n10902;
  assign n10904 = P3_PHYADDRPOINTER_REG_25_ & n10881;
  assign n10905 = ~P3_PHYADDRPOINTER_REG_26_ & n10904;
  assign n10906 = P3_PHYADDRPOINTER_REG_26_ & ~n10904;
  assign n10907 = ~n10905 & ~n10906;
  assign n10908 = n10323 & ~n10907;
  assign n10909 = n9848 & n10318;
  assign n10910 = P3_PHYADDRPOINTER_REG_25_ & n10887;
  assign n10911 = ~P3_PHYADDRPOINTER_REG_26_ & n10910;
  assign n10912 = P3_PHYADDRPOINTER_REG_26_ & ~n10910;
  assign n10913 = ~n10911 & ~n10912;
  assign n10914 = n10325 & ~n10913;
  assign n10915 = n9852 & n10320;
  assign n10916 = P3_PHYADDRPOINTER_REG_26_ & n10316;
  assign n10917 = n9894 & n10329;
  assign n10918 = n10332 & ~n10913;
  assign n10919 = P3_REIP_REG_26_ & n10334;
  assign n10920 = ~n10916 & ~n10917;
  assign n10921 = ~n10918 & n10920;
  assign n10922 = ~n10919 & n10921;
  assign n10923 = ~n10908 & ~n10909;
  assign n10924 = ~n10914 & n10923;
  assign n10925 = ~n10915 & n10924;
  assign n1955 = ~n10922 | ~n10925;
  assign n10927 = P3_PHYADDRPOINTER_REG_26_ & n10904;
  assign n10928 = ~P3_PHYADDRPOINTER_REG_27_ & n10927;
  assign n10929 = P3_PHYADDRPOINTER_REG_27_ & ~n10927;
  assign n10930 = ~n10928 & ~n10929;
  assign n10931 = n10323 & ~n10930;
  assign n10932 = ~n9923 & n10318;
  assign n10933 = P3_PHYADDRPOINTER_REG_26_ & n10910;
  assign n10934 = ~P3_PHYADDRPOINTER_REG_27_ & n10933;
  assign n10935 = P3_PHYADDRPOINTER_REG_27_ & ~n10933;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = n10325 & ~n10936;
  assign n10938 = ~n9927 & n10320;
  assign n10939 = P3_PHYADDRPOINTER_REG_27_ & n10316;
  assign n10940 = ~n9969 & n10329;
  assign n10941 = n10332 & ~n10936;
  assign n10942 = P3_REIP_REG_27_ & n10334;
  assign n10943 = ~n10939 & ~n10940;
  assign n10944 = ~n10941 & n10943;
  assign n10945 = ~n10942 & n10944;
  assign n10946 = ~n10931 & ~n10932;
  assign n10947 = ~n10937 & n10946;
  assign n10948 = ~n10938 & n10947;
  assign n1960 = ~n10945 | ~n10948;
  assign n10950 = n10005 & n10318;
  assign n10951 = n10010 & n10320;
  assign n10952 = P3_PHYADDRPOINTER_REG_27_ & n10927;
  assign n10953 = ~P3_PHYADDRPOINTER_REG_28_ & n10952;
  assign n10954 = P3_PHYADDRPOINTER_REG_28_ & ~n10952;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = n10323 & ~n10955;
  assign n10957 = P3_PHYADDRPOINTER_REG_27_ & n10933;
  assign n10958 = ~P3_PHYADDRPOINTER_REG_28_ & n10957;
  assign n10959 = P3_PHYADDRPOINTER_REG_28_ & ~n10957;
  assign n10960 = ~n10958 & ~n10959;
  assign n10961 = n10325 & ~n10960;
  assign n10962 = P3_PHYADDRPOINTER_REG_28_ & n10316;
  assign n10963 = n10053 & n10329;
  assign n10964 = n10332 & ~n10960;
  assign n10965 = P3_REIP_REG_28_ & n10334;
  assign n10966 = ~n10962 & ~n10963;
  assign n10967 = ~n10964 & n10966;
  assign n10968 = ~n10965 & n10967;
  assign n10969 = ~n10950 & ~n10951;
  assign n10970 = ~n10956 & n10969;
  assign n10971 = ~n10961 & n10970;
  assign n1965 = ~n10968 | ~n10971;
  assign n10973 = ~n10082 & n10318;
  assign n10974 = n10086 & n10320;
  assign n10975 = P3_PHYADDRPOINTER_REG_28_ & n10952;
  assign n10976 = ~P3_PHYADDRPOINTER_REG_29_ & n10975;
  assign n10977 = P3_PHYADDRPOINTER_REG_29_ & ~n10975;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = n10323 & ~n10978;
  assign n10980 = P3_PHYADDRPOINTER_REG_28_ & n10957;
  assign n10981 = ~P3_PHYADDRPOINTER_REG_29_ & n10980;
  assign n10982 = P3_PHYADDRPOINTER_REG_29_ & ~n10980;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = n10325 & ~n10983;
  assign n10985 = P3_PHYADDRPOINTER_REG_29_ & n10316;
  assign n10986 = P3_REIP_REG_29_ & n10334;
  assign n10987 = n10128 & n10329;
  assign n10988 = n10332 & ~n10983;
  assign n10989 = ~n10985 & ~n10986;
  assign n10990 = ~n10987 & n10989;
  assign n10991 = ~n10988 & n10990;
  assign n10992 = ~n10973 & ~n10974;
  assign n10993 = ~n10979 & n10992;
  assign n10994 = ~n10984 & n10993;
  assign n1970 = ~n10991 | ~n10994;
  assign n10996 = ~n10159 & n10318;
  assign n10997 = ~n10163 & n10320;
  assign n10998 = P3_PHYADDRPOINTER_REG_29_ & n10975;
  assign n10999 = ~P3_PHYADDRPOINTER_REG_30_ & n10998;
  assign n11000 = P3_PHYADDRPOINTER_REG_30_ & ~n10998;
  assign n11001 = ~n10999 & ~n11000;
  assign n11002 = n10323 & ~n11001;
  assign n11003 = P3_PHYADDRPOINTER_REG_29_ & n10980;
  assign n11004 = ~P3_PHYADDRPOINTER_REG_30_ & n11003;
  assign n11005 = P3_PHYADDRPOINTER_REG_30_ & ~n11003;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = n10325 & ~n11006;
  assign n11008 = P3_PHYADDRPOINTER_REG_30_ & n10316;
  assign n11009 = P3_REIP_REG_30_ & n10334;
  assign n11010 = ~n10205 & n10329;
  assign n11011 = n10332 & ~n11006;
  assign n11012 = ~n11008 & ~n11009;
  assign n11013 = ~n11010 & n11012;
  assign n11014 = ~n11011 & n11013;
  assign n11015 = ~n10996 & ~n10997;
  assign n11016 = ~n11002 & n11015;
  assign n11017 = ~n11007 & n11016;
  assign n1975 = ~n11014 | ~n11017;
  assign n11019 = n10276 & n10318;
  assign n11020 = P3_PHYADDRPOINTER_REG_30_ & n10998;
  assign n11021 = ~P3_PHYADDRPOINTER_REG_31_ & n11020;
  assign n11022 = P3_PHYADDRPOINTER_REG_31_ & ~n11020;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = n10323 & ~n11023;
  assign n11025 = ~n10281 & n10320;
  assign n11026 = P3_PHYADDRPOINTER_REG_30_ & n11003;
  assign n11027 = ~P3_PHYADDRPOINTER_REG_31_ & n11026;
  assign n11028 = P3_PHYADDRPOINTER_REG_31_ & ~n11026;
  assign n11029 = ~n11027 & ~n11028;
  assign n11030 = n10325 & ~n11029;
  assign n11031 = P3_PHYADDRPOINTER_REG_31_ & n10316;
  assign n11032 = P3_REIP_REG_31_ & n10334;
  assign n11033 = ~n10229 & n10329;
  assign n11034 = n10332 & ~n11029;
  assign n11035 = ~n11031 & ~n11032;
  assign n11036 = ~n11033 & n11035;
  assign n11037 = ~n11034 & n11036;
  assign n11038 = ~n11019 & ~n11024;
  assign n11039 = ~n11025 & n11038;
  assign n11040 = ~n11030 & n11039;
  assign n1980 = ~n11037 | ~n11040;
  assign n11042 = ~n4986 & n5442;
  assign n11043 = n5411 & n11042;
  assign n11044 = ~n5598 & ~n11043;
  assign n11045 = n5713 & ~n11044;
  assign n11046 = ~n5327 & n11045;
  assign n11047 = BUF2_REG_15_ & n11046;
  assign n11048 = n5327 & n11045;
  assign n11049 = P3_EAX_REG_15_ & n11048;
  assign n11050 = P3_LWORD_REG_15_ & ~n11045;
  assign n11051 = ~n11047 & ~n11049;
  assign n1985 = n11050 | ~n11051;
  assign n11053 = BUF2_REG_14_ & n11046;
  assign n11054 = P3_EAX_REG_14_ & n11048;
  assign n11055 = P3_LWORD_REG_14_ & ~n11045;
  assign n11056 = ~n11053 & ~n11054;
  assign n1990 = n11055 | ~n11056;
  assign n11058 = BUF2_REG_13_ & n11046;
  assign n11059 = P3_EAX_REG_13_ & n11048;
  assign n11060 = P3_LWORD_REG_13_ & ~n11045;
  assign n11061 = ~n11058 & ~n11059;
  assign n1995 = n11060 | ~n11061;
  assign n11063 = BUF2_REG_12_ & n11046;
  assign n11064 = P3_EAX_REG_12_ & n11048;
  assign n11065 = P3_LWORD_REG_12_ & ~n11045;
  assign n11066 = ~n11063 & ~n11064;
  assign n2000 = n11065 | ~n11066;
  assign n11068 = BUF2_REG_11_ & n11046;
  assign n11069 = P3_EAX_REG_11_ & n11048;
  assign n11070 = P3_LWORD_REG_11_ & ~n11045;
  assign n11071 = ~n11068 & ~n11069;
  assign n2005 = n11070 | ~n11071;
  assign n11073 = BUF2_REG_10_ & n11046;
  assign n11074 = P3_EAX_REG_10_ & n11048;
  assign n11075 = P3_LWORD_REG_10_ & ~n11045;
  assign n11076 = ~n11073 & ~n11074;
  assign n2010 = n11075 | ~n11076;
  assign n11078 = BUF2_REG_9_ & n11046;
  assign n11079 = P3_EAX_REG_9_ & n11048;
  assign n11080 = P3_LWORD_REG_9_ & ~n11045;
  assign n11081 = ~n11078 & ~n11079;
  assign n2015 = n11080 | ~n11081;
  assign n11083 = BUF2_REG_8_ & n11046;
  assign n11084 = P3_EAX_REG_8_ & n11048;
  assign n11085 = P3_LWORD_REG_8_ & ~n11045;
  assign n11086 = ~n11083 & ~n11084;
  assign n2020 = n11085 | ~n11086;
  assign n11088 = BUF2_REG_7_ & n11046;
  assign n11089 = P3_EAX_REG_7_ & n11048;
  assign n11090 = P3_LWORD_REG_7_ & ~n11045;
  assign n11091 = ~n11088 & ~n11089;
  assign n2025 = n11090 | ~n11091;
  assign n11093 = BUF2_REG_6_ & n11046;
  assign n11094 = P3_EAX_REG_6_ & n11048;
  assign n11095 = P3_LWORD_REG_6_ & ~n11045;
  assign n11096 = ~n11093 & ~n11094;
  assign n2030 = n11095 | ~n11096;
  assign n11098 = BUF2_REG_5_ & n11046;
  assign n11099 = P3_EAX_REG_5_ & n11048;
  assign n11100 = P3_LWORD_REG_5_ & ~n11045;
  assign n11101 = ~n11098 & ~n11099;
  assign n2035 = n11100 | ~n11101;
  assign n11103 = BUF2_REG_4_ & n11046;
  assign n11104 = P3_EAX_REG_4_ & n11048;
  assign n11105 = P3_LWORD_REG_4_ & ~n11045;
  assign n11106 = ~n11103 & ~n11104;
  assign n2040 = n11105 | ~n11106;
  assign n11108 = BUF2_REG_3_ & n11046;
  assign n11109 = P3_EAX_REG_3_ & n11048;
  assign n11110 = P3_LWORD_REG_3_ & ~n11045;
  assign n11111 = ~n11108 & ~n11109;
  assign n2045 = n11110 | ~n11111;
  assign n11113 = BUF2_REG_2_ & n11046;
  assign n11114 = P3_EAX_REG_2_ & n11048;
  assign n11115 = P3_LWORD_REG_2_ & ~n11045;
  assign n11116 = ~n11113 & ~n11114;
  assign n2050 = n11115 | ~n11116;
  assign n11118 = BUF2_REG_1_ & n11046;
  assign n11119 = P3_EAX_REG_1_ & n11048;
  assign n11120 = P3_LWORD_REG_1_ & ~n11045;
  assign n11121 = ~n11118 & ~n11119;
  assign n2055 = n11120 | ~n11121;
  assign n11123 = BUF2_REG_0_ & n11046;
  assign n11124 = P3_EAX_REG_0_ & n11048;
  assign n11125 = P3_LWORD_REG_0_ & ~n11045;
  assign n11126 = ~n11123 & ~n11124;
  assign n2060 = n11125 | ~n11126;
  assign n11128 = P3_EAX_REG_30_ & n11048;
  assign n11129 = P3_UWORD_REG_14_ & ~n11045;
  assign n11130 = ~n11053 & ~n11128;
  assign n2065 = n11129 | ~n11130;
  assign n11132 = P3_EAX_REG_29_ & n11048;
  assign n11133 = P3_UWORD_REG_13_ & ~n11045;
  assign n11134 = ~n11058 & ~n11132;
  assign n2070 = n11133 | ~n11134;
  assign n11136 = P3_EAX_REG_28_ & n11048;
  assign n11137 = P3_UWORD_REG_12_ & ~n11045;
  assign n11138 = ~n11063 & ~n11136;
  assign n2075 = n11137 | ~n11138;
  assign n11140 = P3_EAX_REG_27_ & n11048;
  assign n11141 = P3_UWORD_REG_11_ & ~n11045;
  assign n11142 = ~n11068 & ~n11140;
  assign n2080 = n11141 | ~n11142;
  assign n11144 = P3_EAX_REG_26_ & n11048;
  assign n11145 = P3_UWORD_REG_10_ & ~n11045;
  assign n11146 = ~n11073 & ~n11144;
  assign n2085 = n11145 | ~n11146;
  assign n11148 = P3_EAX_REG_25_ & n11048;
  assign n11149 = P3_UWORD_REG_9_ & ~n11045;
  assign n11150 = ~n11078 & ~n11148;
  assign n2090 = n11149 | ~n11150;
  assign n11152 = P3_EAX_REG_24_ & n11048;
  assign n11153 = P3_UWORD_REG_8_ & ~n11045;
  assign n11154 = ~n11083 & ~n11152;
  assign n2095 = n11153 | ~n11154;
  assign n11156 = P3_EAX_REG_23_ & n11048;
  assign n11157 = P3_UWORD_REG_7_ & ~n11045;
  assign n11158 = ~n11088 & ~n11156;
  assign n2100 = n11157 | ~n11158;
  assign n11160 = P3_EAX_REG_22_ & n11048;
  assign n11161 = P3_UWORD_REG_6_ & ~n11045;
  assign n11162 = ~n11093 & ~n11160;
  assign n2105 = n11161 | ~n11162;
  assign n11164 = P3_EAX_REG_21_ & n11048;
  assign n11165 = P3_UWORD_REG_5_ & ~n11045;
  assign n11166 = ~n11098 & ~n11164;
  assign n2110 = n11165 | ~n11166;
  assign n11168 = P3_EAX_REG_20_ & n11048;
  assign n11169 = P3_UWORD_REG_4_ & ~n11045;
  assign n11170 = ~n11103 & ~n11168;
  assign n2115 = n11169 | ~n11170;
  assign n11172 = P3_EAX_REG_19_ & n11048;
  assign n11173 = P3_UWORD_REG_3_ & ~n11045;
  assign n11174 = ~n11108 & ~n11172;
  assign n2120 = n11173 | ~n11174;
  assign n11176 = P3_EAX_REG_18_ & n11048;
  assign n11177 = P3_UWORD_REG_2_ & ~n11045;
  assign n11178 = ~n11113 & ~n11176;
  assign n2125 = n11177 | ~n11178;
  assign n11180 = P3_EAX_REG_17_ & n11048;
  assign n11181 = P3_UWORD_REG_1_ & ~n11045;
  assign n11182 = ~n11118 & ~n11180;
  assign n2130 = n11181 | ~n11182;
  assign n11184 = P3_EAX_REG_16_ & n11048;
  assign n11185 = P3_UWORD_REG_0_ & ~n11045;
  assign n11186 = ~n11123 & ~n11184;
  assign n2135 = n11185 | ~n11186;
  assign n11188 = ~P3_STATE2_REG_0_ & n5071;
  assign n11189 = n5077 & n5713;
  assign n11190 = ~n5599_1 & n11189;
  assign n11191 = ~n11188 & ~n11190;
  assign n11192 = P3_STATE2_REG_0_ & ~n11191;
  assign n11193 = P3_EAX_REG_0_ & n11192;
  assign n11194 = ~P3_STATE2_REG_0_ & ~n11191;
  assign n11195 = P3_LWORD_REG_0_ & n11194;
  assign n11196 = P3_DATAO_REG_0_ & n11191;
  assign n11197 = ~n11193 & ~n11195;
  assign n2140 = n11196 | ~n11197;
  assign n11199 = P3_EAX_REG_1_ & n11192;
  assign n11200 = P3_LWORD_REG_1_ & n11194;
  assign n11201 = P3_DATAO_REG_1_ & n11191;
  assign n11202 = ~n11199 & ~n11200;
  assign n2144 = n11201 | ~n11202;
  assign n11204 = P3_EAX_REG_2_ & n11192;
  assign n11205 = P3_LWORD_REG_2_ & n11194;
  assign n11206 = P3_DATAO_REG_2_ & n11191;
  assign n11207 = ~n11204 & ~n11205;
  assign n2148 = n11206 | ~n11207;
  assign n11209 = P3_EAX_REG_3_ & n11192;
  assign n11210 = P3_LWORD_REG_3_ & n11194;
  assign n11211 = P3_DATAO_REG_3_ & n11191;
  assign n11212 = ~n11209 & ~n11210;
  assign n2152 = n11211 | ~n11212;
  assign n11214 = P3_EAX_REG_4_ & n11192;
  assign n11215 = P3_LWORD_REG_4_ & n11194;
  assign n11216 = P3_DATAO_REG_4_ & n11191;
  assign n11217 = ~n11214 & ~n11215;
  assign n2156 = n11216 | ~n11217;
  assign n11219 = P3_EAX_REG_5_ & n11192;
  assign n11220 = P3_LWORD_REG_5_ & n11194;
  assign n11221 = P3_DATAO_REG_5_ & n11191;
  assign n11222 = ~n11219 & ~n11220;
  assign n2160 = n11221 | ~n11222;
  assign n11224 = P3_EAX_REG_6_ & n11192;
  assign n11225 = P3_LWORD_REG_6_ & n11194;
  assign n11226 = P3_DATAO_REG_6_ & n11191;
  assign n11227 = ~n11224 & ~n11225;
  assign n2164 = n11226 | ~n11227;
  assign n11229 = P3_EAX_REG_7_ & n11192;
  assign n11230 = P3_LWORD_REG_7_ & n11194;
  assign n11231 = P3_DATAO_REG_7_ & n11191;
  assign n11232 = ~n11229 & ~n11230;
  assign n2168 = n11231 | ~n11232;
  assign n11234 = P3_EAX_REG_8_ & n11192;
  assign n11235 = P3_LWORD_REG_8_ & n11194;
  assign n11236 = P3_DATAO_REG_8_ & n11191;
  assign n11237 = ~n11234 & ~n11235;
  assign n2172 = n11236 | ~n11237;
  assign n11239 = P3_EAX_REG_9_ & n11192;
  assign n11240 = P3_LWORD_REG_9_ & n11194;
  assign n11241 = P3_DATAO_REG_9_ & n11191;
  assign n11242 = ~n11239 & ~n11240;
  assign n2176 = n11241 | ~n11242;
  assign n11244 = P3_EAX_REG_10_ & n11192;
  assign n11245 = P3_LWORD_REG_10_ & n11194;
  assign n11246 = P3_DATAO_REG_10_ & n11191;
  assign n11247 = ~n11244 & ~n11245;
  assign n2180 = n11246 | ~n11247;
  assign n11249 = P3_EAX_REG_11_ & n11192;
  assign n11250 = P3_LWORD_REG_11_ & n11194;
  assign n11251 = P3_DATAO_REG_11_ & n11191;
  assign n11252 = ~n11249 & ~n11250;
  assign n2184 = n11251 | ~n11252;
  assign n11254 = P3_EAX_REG_12_ & n11192;
  assign n11255 = P3_LWORD_REG_12_ & n11194;
  assign n11256 = P3_DATAO_REG_12_ & n11191;
  assign n11257 = ~n11254 & ~n11255;
  assign n2188 = n11256 | ~n11257;
  assign n11259 = P3_EAX_REG_13_ & n11192;
  assign n11260 = P3_LWORD_REG_13_ & n11194;
  assign n11261 = P3_DATAO_REG_13_ & n11191;
  assign n11262 = ~n11259 & ~n11260;
  assign n2192 = n11261 | ~n11262;
  assign n11264 = P3_EAX_REG_14_ & n11192;
  assign n11265 = P3_LWORD_REG_14_ & n11194;
  assign n11266 = P3_DATAO_REG_14_ & n11191;
  assign n11267 = ~n11264 & ~n11265;
  assign n2196 = n11266 | ~n11267;
  assign n11269 = P3_EAX_REG_15_ & n11192;
  assign n11270 = P3_LWORD_REG_15_ & n11194;
  assign n11271 = P3_DATAO_REG_15_ & n11191;
  assign n11272 = ~n11269 & ~n11270;
  assign n2200 = n11271 | ~n11272;
  assign n11274 = P3_UWORD_REG_0_ & n11194;
  assign n11275 = P3_DATAO_REG_16_ & n11191;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = ~n5358 & n11192;
  assign n11278 = P3_EAX_REG_16_ & n11277;
  assign n2204 = ~n11276 | n11278;
  assign n11280 = P3_UWORD_REG_1_ & n11194;
  assign n11281 = P3_DATAO_REG_17_ & n11191;
  assign n11282 = ~n11280 & ~n11281;
  assign n11283 = P3_EAX_REG_17_ & n11277;
  assign n2208 = ~n11282 | n11283;
  assign n11285 = P3_UWORD_REG_2_ & n11194;
  assign n11286 = P3_DATAO_REG_18_ & n11191;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = P3_EAX_REG_18_ & n11277;
  assign n2212 = ~n11287 | n11288;
  assign n11290 = P3_UWORD_REG_3_ & n11194;
  assign n11291 = P3_DATAO_REG_19_ & n11191;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = P3_EAX_REG_19_ & n11277;
  assign n2216 = ~n11292 | n11293;
  assign n11295 = P3_UWORD_REG_4_ & n11194;
  assign n11296 = P3_DATAO_REG_20_ & n11191;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = P3_EAX_REG_20_ & n11277;
  assign n2220 = ~n11297 | n11298;
  assign n11300 = P3_UWORD_REG_5_ & n11194;
  assign n11301 = P3_DATAO_REG_21_ & n11191;
  assign n11302 = ~n11300 & ~n11301;
  assign n11303 = P3_EAX_REG_21_ & n11277;
  assign n2224 = ~n11302 | n11303;
  assign n11305 = P3_UWORD_REG_6_ & n11194;
  assign n11306 = P3_DATAO_REG_22_ & n11191;
  assign n11307 = ~n11305 & ~n11306;
  assign n11308 = P3_EAX_REG_22_ & n11277;
  assign n2228 = ~n11307 | n11308;
  assign n11310 = P3_UWORD_REG_7_ & n11194;
  assign n11311 = P3_DATAO_REG_23_ & n11191;
  assign n11312 = ~n11310 & ~n11311;
  assign n11313 = P3_EAX_REG_23_ & n11277;
  assign n2232 = ~n11312 | n11313;
  assign n11315 = P3_UWORD_REG_8_ & n11194;
  assign n11316 = P3_DATAO_REG_24_ & n11191;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = P3_EAX_REG_24_ & n11277;
  assign n2236 = ~n11317 | n11318;
  assign n11320 = P3_UWORD_REG_9_ & n11194;
  assign n11321 = P3_DATAO_REG_25_ & n11191;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = P3_EAX_REG_25_ & n11277;
  assign n2240 = ~n11322 | n11323;
  assign n11325 = P3_UWORD_REG_10_ & n11194;
  assign n11326 = P3_DATAO_REG_26_ & n11191;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = P3_EAX_REG_26_ & n11277;
  assign n2244 = ~n11327 | n11328;
  assign n11330 = P3_UWORD_REG_11_ & n11194;
  assign n11331 = P3_DATAO_REG_27_ & n11191;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = P3_EAX_REG_27_ & n11277;
  assign n2248 = ~n11332 | n11333;
  assign n11335 = P3_UWORD_REG_12_ & n11194;
  assign n11336 = P3_DATAO_REG_28_ & n11191;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = P3_EAX_REG_28_ & n11277;
  assign n2252 = ~n11337 | n11338;
  assign n11340 = P3_UWORD_REG_13_ & n11194;
  assign n11341 = P3_DATAO_REG_29_ & n11191;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = P3_EAX_REG_29_ & n11277;
  assign n2256 = ~n11342 | n11343;
  assign n11345 = P3_UWORD_REG_14_ & n11194;
  assign n11346 = P3_DATAO_REG_30_ & n11191;
  assign n11347 = ~n11345 & ~n11346;
  assign n11348 = P3_EAX_REG_30_ & n11277;
  assign n2260 = ~n11347 | n11348;
  assign n2264 = P3_DATAO_REG_31_ & n11191;
  assign n11351 = n5593 & ~n5657;
  assign n11352 = n5713 & ~n11351;
  assign n11353 = n5447 & n11352;
  assign n11354 = ~n7423 & n11353;
  assign n11355 = ~n5230 & n11352;
  assign n11356 = ~n5447 & n11355;
  assign n11357 = BUF2_REG_0_ & n11356;
  assign n11358 = P3_EAX_REG_0_ & ~n11352;
  assign n11359 = n5230 & n11352;
  assign n11360 = ~P3_EAX_REG_0_ & n11359;
  assign n11361 = ~n11358 & ~n11360;
  assign n11362 = ~n11354 & ~n11357;
  assign n2268 = ~n11361 | ~n11362;
  assign n11364 = ~n7541 & n11353;
  assign n11365 = BUF2_REG_1_ & n11356;
  assign n11366 = P3_EAX_REG_1_ & ~n11352;
  assign n11367 = ~P3_EAX_REG_0_ & P3_EAX_REG_1_;
  assign n11368 = P3_EAX_REG_0_ & ~P3_EAX_REG_1_;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = n11359 & ~n11369;
  assign n11371 = ~n11366 & ~n11370;
  assign n11372 = ~n11364 & ~n11365;
  assign n2273 = ~n11371 | ~n11372;
  assign n11374 = ~n7652 & n11353;
  assign n11375 = BUF2_REG_2_ & n11356;
  assign n11376 = P3_EAX_REG_2_ & ~n11352;
  assign n11377 = P3_EAX_REG_0_ & P3_EAX_REG_1_;
  assign n11378 = ~P3_EAX_REG_2_ & n11377;
  assign n11379 = P3_EAX_REG_2_ & ~n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = n11359 & ~n11380;
  assign n11382 = ~n11376 & ~n11381;
  assign n11383 = ~n11374 & ~n11375;
  assign n2278 = ~n11382 | ~n11383;
  assign n11385 = ~n7782 & n11353;
  assign n11386 = BUF2_REG_3_ & n11356;
  assign n11387 = P3_EAX_REG_3_ & ~n11352;
  assign n11388 = P3_EAX_REG_0_ & P3_EAX_REG_2_;
  assign n11389 = P3_EAX_REG_1_ & n11388;
  assign n11390 = P3_EAX_REG_3_ & ~n11389;
  assign n11391 = ~P3_EAX_REG_3_ & n11389;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = n11359 & ~n11392;
  assign n11394 = ~n11387 & ~n11393;
  assign n11395 = ~n11385 & ~n11386;
  assign n2283 = ~n11394 | ~n11395;
  assign n11397 = ~n7913 & n11353;
  assign n11398 = BUF2_REG_4_ & n11356;
  assign n11399 = P3_EAX_REG_4_ & ~n11352;
  assign n11400 = P3_EAX_REG_3_ & n11389;
  assign n11401 = ~P3_EAX_REG_4_ & n11400;
  assign n11402 = P3_EAX_REG_4_ & ~n11400;
  assign n11403 = ~n11401 & ~n11402;
  assign n11404 = n11359 & ~n11403;
  assign n11405 = ~n11399 & ~n11404;
  assign n11406 = ~n11397 & ~n11398;
  assign n2288 = ~n11405 | ~n11406;
  assign n11408 = ~n8059 & n11353;
  assign n11409 = BUF2_REG_5_ & n11356;
  assign n11410 = P3_EAX_REG_5_ & ~n11352;
  assign n11411 = P3_EAX_REG_3_ & P3_EAX_REG_4_;
  assign n11412 = n11389 & n11411;
  assign n11413 = P3_EAX_REG_5_ & ~n11412;
  assign n11414 = ~P3_EAX_REG_5_ & n11412;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = n11359 & ~n11415;
  assign n11417 = ~n11410 & ~n11416;
  assign n11418 = ~n11408 & ~n11409;
  assign n2293 = ~n11417 | ~n11418;
  assign n11420 = ~n8195 & n11353;
  assign n11421 = BUF2_REG_6_ & n11356;
  assign n11422 = P3_EAX_REG_6_ & ~n11352;
  assign n11423 = P3_EAX_REG_5_ & n11412;
  assign n11424 = ~P3_EAX_REG_6_ & n11423;
  assign n11425 = P3_EAX_REG_6_ & ~n11423;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = n11359 & ~n11426;
  assign n11428 = ~n11422 & ~n11427;
  assign n11429 = ~n11420 & ~n11421;
  assign n2298 = ~n11428 | ~n11429;
  assign n11431 = ~n7457 & n11353;
  assign n11432 = BUF2_REG_7_ & n11356;
  assign n11433 = P3_EAX_REG_7_ & ~n11352;
  assign n11434 = P3_EAX_REG_5_ & P3_EAX_REG_6_;
  assign n11435 = n11412 & n11434;
  assign n11436 = P3_EAX_REG_7_ & ~n11435;
  assign n11437 = ~P3_EAX_REG_7_ & n11435;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = n11359 & ~n11438;
  assign n11440 = ~n11433 & ~n11439;
  assign n11441 = ~n11431 & ~n11432;
  assign n2303 = ~n11440 | ~n11441;
  assign n11443 = ~n5607 & ~n5614_1;
  assign n11444 = ~n5558 & ~n11443;
  assign n11445 = n5088_1 & n11444;
  assign n11446 = P3_INSTQUEUE_REG_15__0_ & n11445;
  assign n11447 = n5092_1 & n11444;
  assign n11448 = P3_INSTQUEUE_REG_14__0_ & n11447;
  assign n11449 = n5079_1 & n11444;
  assign n11450 = P3_INSTQUEUE_REG_13__0_ & n11449;
  assign n11451 = n5083 & n11444;
  assign n11452 = P3_INSTQUEUE_REG_12__0_ & n11451;
  assign n11453 = ~n11446 & ~n11448;
  assign n11454 = ~n11450 & n11453;
  assign n11455 = ~n11452 & n11454;
  assign n11456 = n5558 & ~n11443;
  assign n11457 = n5088_1 & n11456;
  assign n11458 = P3_INSTQUEUE_REG_11__0_ & n11457;
  assign n11459 = n5092_1 & n11456;
  assign n11460 = P3_INSTQUEUE_REG_10__0_ & n11459;
  assign n11461 = n5079_1 & n11456;
  assign n11462 = P3_INSTQUEUE_REG_9__0_ & n11461;
  assign n11463 = n5083 & n11456;
  assign n11464 = P3_INSTQUEUE_REG_8__0_ & n11463;
  assign n11465 = ~n11458 & ~n11460;
  assign n11466 = ~n11462 & n11465;
  assign n11467 = ~n11464 & n11466;
  assign n11468 = ~n5558 & n11443;
  assign n11469 = n5088_1 & n11468;
  assign n11470 = P3_INSTQUEUE_REG_7__0_ & n11469;
  assign n11471 = n5092_1 & n11468;
  assign n11472 = P3_INSTQUEUE_REG_6__0_ & n11471;
  assign n11473 = n5079_1 & n11468;
  assign n11474 = P3_INSTQUEUE_REG_5__0_ & n11473;
  assign n11475 = n5083 & n11468;
  assign n11476 = P3_INSTQUEUE_REG_4__0_ & n11475;
  assign n11477 = ~n11470 & ~n11472;
  assign n11478 = ~n11474 & n11477;
  assign n11479 = ~n11476 & n11478;
  assign n11480 = n5558 & n11443;
  assign n11481 = n5088_1 & n11480;
  assign n11482 = P3_INSTQUEUE_REG_3__0_ & n11481;
  assign n11483 = n5092_1 & n11480;
  assign n11484 = P3_INSTQUEUE_REG_2__0_ & n11483;
  assign n11485 = n5079_1 & n11480;
  assign n11486 = P3_INSTQUEUE_REG_1__0_ & n11485;
  assign n11487 = n5083 & n11480;
  assign n11488 = P3_INSTQUEUE_REG_0__0_ & n11487;
  assign n11489 = ~n11482 & ~n11484;
  assign n11490 = ~n11486 & n11489;
  assign n11491 = ~n11488 & n11490;
  assign n11492 = n11455 & n11467;
  assign n11493 = n11479 & n11492;
  assign n11494 = n11491 & n11493;
  assign n11495 = n11353 & ~n11494;
  assign n11496 = BUF2_REG_8_ & n11356;
  assign n11497 = P3_EAX_REG_8_ & ~n11352;
  assign n11498 = P3_EAX_REG_7_ & n11435;
  assign n11499 = ~P3_EAX_REG_8_ & n11498;
  assign n11500 = P3_EAX_REG_8_ & ~n11498;
  assign n11501 = ~n11499 & ~n11500;
  assign n11502 = n11359 & ~n11501;
  assign n11503 = ~n11497 & ~n11502;
  assign n11504 = ~n11495 & ~n11496;
  assign n2308 = ~n11503 | ~n11504;
  assign n11506 = P3_INSTQUEUE_REG_15__1_ & n11445;
  assign n11507 = P3_INSTQUEUE_REG_14__1_ & n11447;
  assign n11508 = P3_INSTQUEUE_REG_13__1_ & n11449;
  assign n11509 = P3_INSTQUEUE_REG_12__1_ & n11451;
  assign n11510 = ~n11506 & ~n11507;
  assign n11511 = ~n11508 & n11510;
  assign n11512 = ~n11509 & n11511;
  assign n11513 = P3_INSTQUEUE_REG_11__1_ & n11457;
  assign n11514 = P3_INSTQUEUE_REG_10__1_ & n11459;
  assign n11515 = P3_INSTQUEUE_REG_9__1_ & n11461;
  assign n11516 = P3_INSTQUEUE_REG_8__1_ & n11463;
  assign n11517 = ~n11513 & ~n11514;
  assign n11518 = ~n11515 & n11517;
  assign n11519 = ~n11516 & n11518;
  assign n11520 = P3_INSTQUEUE_REG_7__1_ & n11469;
  assign n11521 = P3_INSTQUEUE_REG_6__1_ & n11471;
  assign n11522 = P3_INSTQUEUE_REG_5__1_ & n11473;
  assign n11523 = P3_INSTQUEUE_REG_4__1_ & n11475;
  assign n11524 = ~n11520 & ~n11521;
  assign n11525 = ~n11522 & n11524;
  assign n11526 = ~n11523 & n11525;
  assign n11527 = P3_INSTQUEUE_REG_3__1_ & n11481;
  assign n11528 = P3_INSTQUEUE_REG_2__1_ & n11483;
  assign n11529 = P3_INSTQUEUE_REG_1__1_ & n11485;
  assign n11530 = P3_INSTQUEUE_REG_0__1_ & n11487;
  assign n11531 = ~n11527 & ~n11528;
  assign n11532 = ~n11529 & n11531;
  assign n11533 = ~n11530 & n11532;
  assign n11534 = n11512 & n11519;
  assign n11535 = n11526 & n11534;
  assign n11536 = n11533 & n11535;
  assign n11537 = n11353 & ~n11536;
  assign n11538 = BUF2_REG_9_ & n11356;
  assign n11539 = P3_EAX_REG_9_ & ~n11352;
  assign n11540 = P3_EAX_REG_7_ & P3_EAX_REG_8_;
  assign n11541 = n11435 & n11540;
  assign n11542 = P3_EAX_REG_9_ & ~n11541;
  assign n11543 = ~P3_EAX_REG_9_ & n11541;
  assign n11544 = ~n11542 & ~n11543;
  assign n11545 = n11359 & ~n11544;
  assign n11546 = ~n11539 & ~n11545;
  assign n11547 = ~n11537 & ~n11538;
  assign n2313 = ~n11546 | ~n11547;
  assign n11549 = P3_INSTQUEUE_REG_15__2_ & n11445;
  assign n11550 = P3_INSTQUEUE_REG_14__2_ & n11447;
  assign n11551 = P3_INSTQUEUE_REG_13__2_ & n11449;
  assign n11552 = P3_INSTQUEUE_REG_12__2_ & n11451;
  assign n11553 = ~n11549 & ~n11550;
  assign n11554 = ~n11551 & n11553;
  assign n11555 = ~n11552 & n11554;
  assign n11556 = P3_INSTQUEUE_REG_11__2_ & n11457;
  assign n11557 = P3_INSTQUEUE_REG_10__2_ & n11459;
  assign n11558 = P3_INSTQUEUE_REG_9__2_ & n11461;
  assign n11559 = P3_INSTQUEUE_REG_8__2_ & n11463;
  assign n11560 = ~n11556 & ~n11557;
  assign n11561 = ~n11558 & n11560;
  assign n11562 = ~n11559 & n11561;
  assign n11563 = P3_INSTQUEUE_REG_7__2_ & n11469;
  assign n11564 = P3_INSTQUEUE_REG_6__2_ & n11471;
  assign n11565 = P3_INSTQUEUE_REG_5__2_ & n11473;
  assign n11566 = P3_INSTQUEUE_REG_4__2_ & n11475;
  assign n11567 = ~n11563 & ~n11564;
  assign n11568 = ~n11565 & n11567;
  assign n11569 = ~n11566 & n11568;
  assign n11570 = P3_INSTQUEUE_REG_3__2_ & n11481;
  assign n11571 = P3_INSTQUEUE_REG_2__2_ & n11483;
  assign n11572 = P3_INSTQUEUE_REG_1__2_ & n11485;
  assign n11573 = P3_INSTQUEUE_REG_0__2_ & n11487;
  assign n11574 = ~n11570 & ~n11571;
  assign n11575 = ~n11572 & n11574;
  assign n11576 = ~n11573 & n11575;
  assign n11577 = n11555 & n11562;
  assign n11578 = n11569 & n11577;
  assign n11579 = n11576 & n11578;
  assign n11580 = n11353 & ~n11579;
  assign n11581 = BUF2_REG_10_ & n11356;
  assign n11582 = P3_EAX_REG_10_ & ~n11352;
  assign n11583 = P3_EAX_REG_9_ & n11541;
  assign n11584 = ~P3_EAX_REG_10_ & n11583;
  assign n11585 = P3_EAX_REG_10_ & ~n11583;
  assign n11586 = ~n11584 & ~n11585;
  assign n11587 = n11359 & ~n11586;
  assign n11588 = ~n11582 & ~n11587;
  assign n11589 = ~n11580 & ~n11581;
  assign n2318 = ~n11588 | ~n11589;
  assign n11591 = P3_INSTQUEUE_REG_15__3_ & n11445;
  assign n11592 = P3_INSTQUEUE_REG_14__3_ & n11447;
  assign n11593 = P3_INSTQUEUE_REG_13__3_ & n11449;
  assign n11594 = P3_INSTQUEUE_REG_12__3_ & n11451;
  assign n11595 = ~n11591 & ~n11592;
  assign n11596 = ~n11593 & n11595;
  assign n11597 = ~n11594 & n11596;
  assign n11598 = P3_INSTQUEUE_REG_11__3_ & n11457;
  assign n11599 = P3_INSTQUEUE_REG_10__3_ & n11459;
  assign n11600 = P3_INSTQUEUE_REG_9__3_ & n11461;
  assign n11601 = P3_INSTQUEUE_REG_8__3_ & n11463;
  assign n11602 = ~n11598 & ~n11599;
  assign n11603 = ~n11600 & n11602;
  assign n11604 = ~n11601 & n11603;
  assign n11605 = P3_INSTQUEUE_REG_7__3_ & n11469;
  assign n11606 = P3_INSTQUEUE_REG_6__3_ & n11471;
  assign n11607 = P3_INSTQUEUE_REG_5__3_ & n11473;
  assign n11608 = P3_INSTQUEUE_REG_4__3_ & n11475;
  assign n11609 = ~n11605 & ~n11606;
  assign n11610 = ~n11607 & n11609;
  assign n11611 = ~n11608 & n11610;
  assign n11612 = P3_INSTQUEUE_REG_3__3_ & n11481;
  assign n11613 = P3_INSTQUEUE_REG_2__3_ & n11483;
  assign n11614 = P3_INSTQUEUE_REG_1__3_ & n11485;
  assign n11615 = P3_INSTQUEUE_REG_0__3_ & n11487;
  assign n11616 = ~n11612 & ~n11613;
  assign n11617 = ~n11614 & n11616;
  assign n11618 = ~n11615 & n11617;
  assign n11619 = n11597 & n11604;
  assign n11620 = n11611 & n11619;
  assign n11621 = n11618 & n11620;
  assign n11622 = n11353 & ~n11621;
  assign n11623 = BUF2_REG_11_ & n11356;
  assign n11624 = P3_EAX_REG_11_ & ~n11352;
  assign n11625 = P3_EAX_REG_9_ & P3_EAX_REG_10_;
  assign n11626 = n11541 & n11625;
  assign n11627 = P3_EAX_REG_11_ & ~n11626;
  assign n11628 = ~P3_EAX_REG_11_ & n11626;
  assign n11629 = ~n11627 & ~n11628;
  assign n11630 = n11359 & ~n11629;
  assign n11631 = ~n11624 & ~n11630;
  assign n11632 = ~n11622 & ~n11623;
  assign n2323 = ~n11631 | ~n11632;
  assign n11634 = P3_INSTQUEUE_REG_15__4_ & n11445;
  assign n11635 = P3_INSTQUEUE_REG_14__4_ & n11447;
  assign n11636 = P3_INSTQUEUE_REG_13__4_ & n11449;
  assign n11637 = P3_INSTQUEUE_REG_12__4_ & n11451;
  assign n11638 = ~n11634 & ~n11635;
  assign n11639 = ~n11636 & n11638;
  assign n11640 = ~n11637 & n11639;
  assign n11641 = P3_INSTQUEUE_REG_11__4_ & n11457;
  assign n11642 = P3_INSTQUEUE_REG_10__4_ & n11459;
  assign n11643 = P3_INSTQUEUE_REG_9__4_ & n11461;
  assign n11644 = P3_INSTQUEUE_REG_8__4_ & n11463;
  assign n11645 = ~n11641 & ~n11642;
  assign n11646 = ~n11643 & n11645;
  assign n11647 = ~n11644 & n11646;
  assign n11648 = P3_INSTQUEUE_REG_7__4_ & n11469;
  assign n11649 = P3_INSTQUEUE_REG_6__4_ & n11471;
  assign n11650 = P3_INSTQUEUE_REG_5__4_ & n11473;
  assign n11651 = P3_INSTQUEUE_REG_4__4_ & n11475;
  assign n11652 = ~n11648 & ~n11649;
  assign n11653 = ~n11650 & n11652;
  assign n11654 = ~n11651 & n11653;
  assign n11655 = P3_INSTQUEUE_REG_3__4_ & n11481;
  assign n11656 = P3_INSTQUEUE_REG_2__4_ & n11483;
  assign n11657 = P3_INSTQUEUE_REG_1__4_ & n11485;
  assign n11658 = P3_INSTQUEUE_REG_0__4_ & n11487;
  assign n11659 = ~n11655 & ~n11656;
  assign n11660 = ~n11657 & n11659;
  assign n11661 = ~n11658 & n11660;
  assign n11662 = n11640 & n11647;
  assign n11663 = n11654 & n11662;
  assign n11664 = n11661 & n11663;
  assign n11665 = n11353 & ~n11664;
  assign n11666 = BUF2_REG_12_ & n11356;
  assign n11667 = P3_EAX_REG_12_ & ~n11352;
  assign n11668 = P3_EAX_REG_11_ & n11626;
  assign n11669 = ~P3_EAX_REG_12_ & n11668;
  assign n11670 = P3_EAX_REG_12_ & ~n11668;
  assign n11671 = ~n11669 & ~n11670;
  assign n11672 = n11359 & ~n11671;
  assign n11673 = ~n11667 & ~n11672;
  assign n11674 = ~n11665 & ~n11666;
  assign n2328 = ~n11673 | ~n11674;
  assign n11676 = BUF2_REG_13_ & n11356;
  assign n11677 = P3_INSTQUEUE_REG_15__5_ & n11445;
  assign n11678 = P3_INSTQUEUE_REG_14__5_ & n11447;
  assign n11679 = P3_INSTQUEUE_REG_13__5_ & n11449;
  assign n11680 = P3_INSTQUEUE_REG_12__5_ & n11451;
  assign n11681 = ~n11677 & ~n11678;
  assign n11682 = ~n11679 & n11681;
  assign n11683 = ~n11680 & n11682;
  assign n11684 = P3_INSTQUEUE_REG_11__5_ & n11457;
  assign n11685 = P3_INSTQUEUE_REG_10__5_ & n11459;
  assign n11686 = P3_INSTQUEUE_REG_9__5_ & n11461;
  assign n11687 = P3_INSTQUEUE_REG_8__5_ & n11463;
  assign n11688 = ~n11684 & ~n11685;
  assign n11689 = ~n11686 & n11688;
  assign n11690 = ~n11687 & n11689;
  assign n11691 = P3_INSTQUEUE_REG_7__5_ & n11469;
  assign n11692 = P3_INSTQUEUE_REG_6__5_ & n11471;
  assign n11693 = P3_INSTQUEUE_REG_5__5_ & n11473;
  assign n11694 = P3_INSTQUEUE_REG_4__5_ & n11475;
  assign n11695 = ~n11691 & ~n11692;
  assign n11696 = ~n11693 & n11695;
  assign n11697 = ~n11694 & n11696;
  assign n11698 = P3_INSTQUEUE_REG_3__5_ & n11481;
  assign n11699 = P3_INSTQUEUE_REG_2__5_ & n11483;
  assign n11700 = P3_INSTQUEUE_REG_1__5_ & n11485;
  assign n11701 = P3_INSTQUEUE_REG_0__5_ & n11487;
  assign n11702 = ~n11698 & ~n11699;
  assign n11703 = ~n11700 & n11702;
  assign n11704 = ~n11701 & n11703;
  assign n11705 = n11683 & n11690;
  assign n11706 = n11697 & n11705;
  assign n11707 = n11704 & n11706;
  assign n11708 = n11353 & ~n11707;
  assign n11709 = P3_EAX_REG_13_ & ~n11352;
  assign n11710 = ~n11708 & ~n11709;
  assign n11711 = P3_EAX_REG_11_ & P3_EAX_REG_12_;
  assign n11712 = n11626 & n11711;
  assign n11713 = P3_EAX_REG_13_ & ~n11712;
  assign n11714 = ~P3_EAX_REG_13_ & n11712;
  assign n11715 = ~n11713 & ~n11714;
  assign n11716 = n11359 & ~n11715;
  assign n11717 = ~n11676 & n11710;
  assign n2333 = n11716 | ~n11717;
  assign n11719 = BUF2_REG_14_ & n11356;
  assign n11720 = P3_INSTQUEUE_REG_15__6_ & n11445;
  assign n11721 = P3_INSTQUEUE_REG_14__6_ & n11447;
  assign n11722 = P3_INSTQUEUE_REG_13__6_ & n11449;
  assign n11723 = P3_INSTQUEUE_REG_12__6_ & n11451;
  assign n11724 = ~n11720 & ~n11721;
  assign n11725 = ~n11722 & n11724;
  assign n11726 = ~n11723 & n11725;
  assign n11727 = P3_INSTQUEUE_REG_11__6_ & n11457;
  assign n11728 = P3_INSTQUEUE_REG_10__6_ & n11459;
  assign n11729 = P3_INSTQUEUE_REG_9__6_ & n11461;
  assign n11730 = P3_INSTQUEUE_REG_8__6_ & n11463;
  assign n11731 = ~n11727 & ~n11728;
  assign n11732 = ~n11729 & n11731;
  assign n11733 = ~n11730 & n11732;
  assign n11734 = P3_INSTQUEUE_REG_7__6_ & n11469;
  assign n11735 = P3_INSTQUEUE_REG_6__6_ & n11471;
  assign n11736 = P3_INSTQUEUE_REG_5__6_ & n11473;
  assign n11737 = P3_INSTQUEUE_REG_4__6_ & n11475;
  assign n11738 = ~n11734 & ~n11735;
  assign n11739 = ~n11736 & n11738;
  assign n11740 = ~n11737 & n11739;
  assign n11741 = P3_INSTQUEUE_REG_3__6_ & n11481;
  assign n11742 = P3_INSTQUEUE_REG_2__6_ & n11483;
  assign n11743 = P3_INSTQUEUE_REG_1__6_ & n11485;
  assign n11744 = P3_INSTQUEUE_REG_0__6_ & n11487;
  assign n11745 = ~n11741 & ~n11742;
  assign n11746 = ~n11743 & n11745;
  assign n11747 = ~n11744 & n11746;
  assign n11748 = n11726 & n11733;
  assign n11749 = n11740 & n11748;
  assign n11750 = n11747 & n11749;
  assign n11751 = n11353 & ~n11750;
  assign n11752 = P3_EAX_REG_14_ & ~n11352;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = P3_EAX_REG_13_ & n11712;
  assign n11755 = ~P3_EAX_REG_14_ & n11754;
  assign n11756 = P3_EAX_REG_14_ & ~n11754;
  assign n11757 = ~n11755 & ~n11756;
  assign n11758 = n11359 & ~n11757;
  assign n11759 = ~n11719 & n11753;
  assign n2338 = n11758 | ~n11759;
  assign n11761 = BUF2_REG_15_ & n11356;
  assign n11762 = P3_INSTQUEUE_REG_15__7_ & n11445;
  assign n11763 = P3_INSTQUEUE_REG_14__7_ & n11447;
  assign n11764 = P3_INSTQUEUE_REG_13__7_ & n11449;
  assign n11765 = P3_INSTQUEUE_REG_12__7_ & n11451;
  assign n11766 = ~n11762 & ~n11763;
  assign n11767 = ~n11764 & n11766;
  assign n11768 = ~n11765 & n11767;
  assign n11769 = P3_INSTQUEUE_REG_11__7_ & n11457;
  assign n11770 = P3_INSTQUEUE_REG_10__7_ & n11459;
  assign n11771 = P3_INSTQUEUE_REG_9__7_ & n11461;
  assign n11772 = P3_INSTQUEUE_REG_8__7_ & n11463;
  assign n11773 = ~n11769 & ~n11770;
  assign n11774 = ~n11771 & n11773;
  assign n11775 = ~n11772 & n11774;
  assign n11776 = P3_INSTQUEUE_REG_7__7_ & n11469;
  assign n11777 = P3_INSTQUEUE_REG_6__7_ & n11471;
  assign n11778 = P3_INSTQUEUE_REG_5__7_ & n11473;
  assign n11779 = P3_INSTQUEUE_REG_4__7_ & n11475;
  assign n11780 = ~n11776 & ~n11777;
  assign n11781 = ~n11778 & n11780;
  assign n11782 = ~n11779 & n11781;
  assign n11783 = P3_INSTQUEUE_REG_3__7_ & n11481;
  assign n11784 = P3_INSTQUEUE_REG_2__7_ & n11483;
  assign n11785 = P3_INSTQUEUE_REG_1__7_ & n11485;
  assign n11786 = P3_INSTQUEUE_REG_0__7_ & n11487;
  assign n11787 = ~n11783 & ~n11784;
  assign n11788 = ~n11785 & n11787;
  assign n11789 = ~n11786 & n11788;
  assign n11790 = n11768 & n11775;
  assign n11791 = n11782 & n11790;
  assign n11792 = n11789 & n11791;
  assign n11793 = n11353 & ~n11792;
  assign n11794 = P3_EAX_REG_15_ & ~n11352;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = P3_EAX_REG_13_ & P3_EAX_REG_14_;
  assign n11797 = n11712 & n11796;
  assign n11798 = P3_EAX_REG_15_ & ~n11797;
  assign n11799 = ~P3_EAX_REG_15_ & n11797;
  assign n11800 = ~n11798 & ~n11799;
  assign n11801 = n11359 & ~n11800;
  assign n11802 = ~n11761 & n11795;
  assign n2343 = n11801 | ~n11802;
  assign n11804 = ~n5167 & n11355;
  assign n11805 = BUF2_REG_16_ & n11804;
  assign n11806 = n5136_1 & n11355;
  assign n11807 = BUF2_REG_0_ & n11806;
  assign n11808 = P3_EAX_REG_16_ & ~n11352;
  assign n11809 = P3_INSTQUEUERD_ADDR_REG_2_ & ~n5092_1;
  assign n11810 = ~P3_INSTQUEUERD_ADDR_REG_3_ & n11809;
  assign n11811 = P3_INSTQUEUERD_ADDR_REG_3_ & ~n11809;
  assign n11812 = ~n11810 & ~n11811;
  assign n11813 = ~n5093 & ~n11809;
  assign n11814 = n11812 & n11813;
  assign n11815 = n7373 & n11814;
  assign n11816 = P3_INSTQUEUE_REG_7__0_ & n11815;
  assign n11817 = n7370 & n11814;
  assign n11818 = P3_INSTQUEUE_REG_6__0_ & n11817;
  assign n11819 = n7379 & n11814;
  assign n11820 = P3_INSTQUEUE_REG_5__0_ & n11819;
  assign n11821 = n7376 & n11814;
  assign n11822 = P3_INSTQUEUE_REG_4__0_ & n11821;
  assign n11823 = ~n11816 & ~n11818;
  assign n11824 = ~n11820 & n11823;
  assign n11825 = ~n11822 & n11824;
  assign n11826 = n11812 & ~n11813;
  assign n11827 = n7373 & n11826;
  assign n11828 = P3_INSTQUEUE_REG_3__0_ & n11827;
  assign n11829 = n7370 & n11826;
  assign n11830 = P3_INSTQUEUE_REG_2__0_ & n11829;
  assign n11831 = n7379 & n11826;
  assign n11832 = P3_INSTQUEUE_REG_1__0_ & n11831;
  assign n11833 = n7376 & n11826;
  assign n11834 = P3_INSTQUEUE_REG_0__0_ & n11833;
  assign n11835 = ~n11828 & ~n11830;
  assign n11836 = ~n11832 & n11835;
  assign n11837 = ~n11834 & n11836;
  assign n11838 = ~n11812 & n11813;
  assign n11839 = n7373 & n11838;
  assign n11840 = P3_INSTQUEUE_REG_15__0_ & n11839;
  assign n11841 = n7370 & n11838;
  assign n11842 = P3_INSTQUEUE_REG_14__0_ & n11841;
  assign n11843 = n7379 & n11838;
  assign n11844 = P3_INSTQUEUE_REG_13__0_ & n11843;
  assign n11845 = n7376 & n11838;
  assign n11846 = P3_INSTQUEUE_REG_12__0_ & n11845;
  assign n11847 = ~n11840 & ~n11842;
  assign n11848 = ~n11844 & n11847;
  assign n11849 = ~n11846 & n11848;
  assign n11850 = ~n11812 & ~n11813;
  assign n11851 = n7373 & n11850;
  assign n11852 = P3_INSTQUEUE_REG_11__0_ & n11851;
  assign n11853 = n7370 & n11850;
  assign n11854 = P3_INSTQUEUE_REG_10__0_ & n11853;
  assign n11855 = n7379 & n11850;
  assign n11856 = P3_INSTQUEUE_REG_9__0_ & n11855;
  assign n11857 = n7376 & n11850;
  assign n11858 = P3_INSTQUEUE_REG_8__0_ & n11857;
  assign n11859 = ~n11852 & ~n11854;
  assign n11860 = ~n11856 & n11859;
  assign n11861 = ~n11858 & n11860;
  assign n11862 = n11825 & n11837;
  assign n11863 = n11849 & n11862;
  assign n11864 = n11861 & n11863;
  assign n11865 = n11353 & ~n11864;
  assign n11866 = ~n11808 & ~n11865;
  assign n11867 = P3_EAX_REG_15_ & n11797;
  assign n11868 = ~P3_EAX_REG_16_ & n11867;
  assign n11869 = P3_EAX_REG_16_ & ~n11867;
  assign n11870 = ~n11868 & ~n11869;
  assign n11871 = n11359 & ~n11870;
  assign n11872 = ~n11805 & ~n11807;
  assign n11873 = n11866 & n11872;
  assign n2348 = n11871 | ~n11873;
  assign n11875 = BUF2_REG_17_ & n11804;
  assign n11876 = BUF2_REG_1_ & n11806;
  assign n11877 = P3_EAX_REG_17_ & ~n11352;
  assign n11878 = P3_INSTQUEUE_REG_7__1_ & n11815;
  assign n11879 = P3_INSTQUEUE_REG_6__1_ & n11817;
  assign n11880 = P3_INSTQUEUE_REG_5__1_ & n11819;
  assign n11881 = P3_INSTQUEUE_REG_4__1_ & n11821;
  assign n11882 = ~n11878 & ~n11879;
  assign n11883 = ~n11880 & n11882;
  assign n11884 = ~n11881 & n11883;
  assign n11885 = P3_INSTQUEUE_REG_3__1_ & n11827;
  assign n11886 = P3_INSTQUEUE_REG_2__1_ & n11829;
  assign n11887 = P3_INSTQUEUE_REG_1__1_ & n11831;
  assign n11888 = P3_INSTQUEUE_REG_0__1_ & n11833;
  assign n11889 = ~n11885 & ~n11886;
  assign n11890 = ~n11887 & n11889;
  assign n11891 = ~n11888 & n11890;
  assign n11892 = P3_INSTQUEUE_REG_15__1_ & n11839;
  assign n11893 = P3_INSTQUEUE_REG_14__1_ & n11841;
  assign n11894 = P3_INSTQUEUE_REG_13__1_ & n11843;
  assign n11895 = P3_INSTQUEUE_REG_12__1_ & n11845;
  assign n11896 = ~n11892 & ~n11893;
  assign n11897 = ~n11894 & n11896;
  assign n11898 = ~n11895 & n11897;
  assign n11899 = P3_INSTQUEUE_REG_11__1_ & n11851;
  assign n11900 = P3_INSTQUEUE_REG_10__1_ & n11853;
  assign n11901 = P3_INSTQUEUE_REG_9__1_ & n11855;
  assign n11902 = P3_INSTQUEUE_REG_8__1_ & n11857;
  assign n11903 = ~n11899 & ~n11900;
  assign n11904 = ~n11901 & n11903;
  assign n11905 = ~n11902 & n11904;
  assign n11906 = n11884 & n11891;
  assign n11907 = n11898 & n11906;
  assign n11908 = n11905 & n11907;
  assign n11909 = n11353 & ~n11908;
  assign n11910 = ~n11877 & ~n11909;
  assign n11911 = P3_EAX_REG_15_ & P3_EAX_REG_16_;
  assign n11912 = n11797 & n11911;
  assign n11913 = P3_EAX_REG_17_ & ~n11912;
  assign n11914 = ~P3_EAX_REG_17_ & n11912;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 = n11359 & ~n11915;
  assign n11917 = ~n11875 & ~n11876;
  assign n11918 = n11910 & n11917;
  assign n2353 = n11916 | ~n11918;
  assign n11920 = BUF2_REG_18_ & n11804;
  assign n11921 = BUF2_REG_2_ & n11806;
  assign n11922 = P3_EAX_REG_18_ & ~n11352;
  assign n11923 = P3_INSTQUEUE_REG_7__2_ & n11815;
  assign n11924 = P3_INSTQUEUE_REG_6__2_ & n11817;
  assign n11925 = P3_INSTQUEUE_REG_5__2_ & n11819;
  assign n11926 = P3_INSTQUEUE_REG_4__2_ & n11821;
  assign n11927 = ~n11923 & ~n11924;
  assign n11928 = ~n11925 & n11927;
  assign n11929 = ~n11926 & n11928;
  assign n11930 = P3_INSTQUEUE_REG_3__2_ & n11827;
  assign n11931 = P3_INSTQUEUE_REG_2__2_ & n11829;
  assign n11932 = P3_INSTQUEUE_REG_1__2_ & n11831;
  assign n11933 = P3_INSTQUEUE_REG_0__2_ & n11833;
  assign n11934 = ~n11930 & ~n11931;
  assign n11935 = ~n11932 & n11934;
  assign n11936 = ~n11933 & n11935;
  assign n11937 = P3_INSTQUEUE_REG_15__2_ & n11839;
  assign n11938 = P3_INSTQUEUE_REG_14__2_ & n11841;
  assign n11939 = P3_INSTQUEUE_REG_13__2_ & n11843;
  assign n11940 = P3_INSTQUEUE_REG_12__2_ & n11845;
  assign n11941 = ~n11937 & ~n11938;
  assign n11942 = ~n11939 & n11941;
  assign n11943 = ~n11940 & n11942;
  assign n11944 = P3_INSTQUEUE_REG_11__2_ & n11851;
  assign n11945 = P3_INSTQUEUE_REG_10__2_ & n11853;
  assign n11946 = P3_INSTQUEUE_REG_9__2_ & n11855;
  assign n11947 = P3_INSTQUEUE_REG_8__2_ & n11857;
  assign n11948 = ~n11944 & ~n11945;
  assign n11949 = ~n11946 & n11948;
  assign n11950 = ~n11947 & n11949;
  assign n11951 = n11929 & n11936;
  assign n11952 = n11943 & n11951;
  assign n11953 = n11950 & n11952;
  assign n11954 = n11353 & ~n11953;
  assign n11955 = ~n11922 & ~n11954;
  assign n11956 = P3_EAX_REG_17_ & n11912;
  assign n11957 = ~P3_EAX_REG_18_ & n11956;
  assign n11958 = P3_EAX_REG_18_ & ~n11956;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = n11359 & ~n11959;
  assign n11961 = ~n11920 & ~n11921;
  assign n11962 = n11955 & n11961;
  assign n2358 = n11960 | ~n11962;
  assign n11964 = BUF2_REG_19_ & n11804;
  assign n11965 = BUF2_REG_3_ & n11806;
  assign n11966 = P3_EAX_REG_19_ & ~n11352;
  assign n11967 = P3_INSTQUEUE_REG_7__3_ & n11815;
  assign n11968 = P3_INSTQUEUE_REG_6__3_ & n11817;
  assign n11969 = P3_INSTQUEUE_REG_5__3_ & n11819;
  assign n11970 = P3_INSTQUEUE_REG_4__3_ & n11821;
  assign n11971 = ~n11967 & ~n11968;
  assign n11972 = ~n11969 & n11971;
  assign n11973 = ~n11970 & n11972;
  assign n11974 = P3_INSTQUEUE_REG_3__3_ & n11827;
  assign n11975 = P3_INSTQUEUE_REG_2__3_ & n11829;
  assign n11976 = P3_INSTQUEUE_REG_1__3_ & n11831;
  assign n11977 = P3_INSTQUEUE_REG_0__3_ & n11833;
  assign n11978 = ~n11974 & ~n11975;
  assign n11979 = ~n11976 & n11978;
  assign n11980 = ~n11977 & n11979;
  assign n11981 = P3_INSTQUEUE_REG_15__3_ & n11839;
  assign n11982 = P3_INSTQUEUE_REG_14__3_ & n11841;
  assign n11983 = P3_INSTQUEUE_REG_13__3_ & n11843;
  assign n11984 = P3_INSTQUEUE_REG_12__3_ & n11845;
  assign n11985 = ~n11981 & ~n11982;
  assign n11986 = ~n11983 & n11985;
  assign n11987 = ~n11984 & n11986;
  assign n11988 = P3_INSTQUEUE_REG_11__3_ & n11851;
  assign n11989 = P3_INSTQUEUE_REG_10__3_ & n11853;
  assign n11990 = P3_INSTQUEUE_REG_9__3_ & n11855;
  assign n11991 = P3_INSTQUEUE_REG_8__3_ & n11857;
  assign n11992 = ~n11988 & ~n11989;
  assign n11993 = ~n11990 & n11992;
  assign n11994 = ~n11991 & n11993;
  assign n11995 = n11973 & n11980;
  assign n11996 = n11987 & n11995;
  assign n11997 = n11994 & n11996;
  assign n11998 = n11353 & ~n11997;
  assign n11999 = ~n11966 & ~n11998;
  assign n12000 = P3_EAX_REG_17_ & P3_EAX_REG_18_;
  assign n12001 = n11912 & n12000;
  assign n12002 = P3_EAX_REG_19_ & ~n12001;
  assign n12003 = ~P3_EAX_REG_19_ & n12001;
  assign n12004 = ~n12002 & ~n12003;
  assign n12005 = n11359 & ~n12004;
  assign n12006 = ~n11964 & ~n11965;
  assign n12007 = n11999 & n12006;
  assign n2363 = n12005 | ~n12007;
  assign n12009 = BUF2_REG_20_ & n11804;
  assign n12010 = BUF2_REG_4_ & n11806;
  assign n12011 = P3_EAX_REG_20_ & ~n11352;
  assign n12012 = P3_INSTQUEUE_REG_7__4_ & n11815;
  assign n12013 = P3_INSTQUEUE_REG_6__4_ & n11817;
  assign n12014 = P3_INSTQUEUE_REG_5__4_ & n11819;
  assign n12015 = P3_INSTQUEUE_REG_4__4_ & n11821;
  assign n12016 = ~n12012 & ~n12013;
  assign n12017 = ~n12014 & n12016;
  assign n12018 = ~n12015 & n12017;
  assign n12019 = P3_INSTQUEUE_REG_3__4_ & n11827;
  assign n12020 = P3_INSTQUEUE_REG_2__4_ & n11829;
  assign n12021 = P3_INSTQUEUE_REG_1__4_ & n11831;
  assign n12022 = P3_INSTQUEUE_REG_0__4_ & n11833;
  assign n12023 = ~n12019 & ~n12020;
  assign n12024 = ~n12021 & n12023;
  assign n12025 = ~n12022 & n12024;
  assign n12026 = P3_INSTQUEUE_REG_15__4_ & n11839;
  assign n12027 = P3_INSTQUEUE_REG_14__4_ & n11841;
  assign n12028 = P3_INSTQUEUE_REG_13__4_ & n11843;
  assign n12029 = P3_INSTQUEUE_REG_12__4_ & n11845;
  assign n12030 = ~n12026 & ~n12027;
  assign n12031 = ~n12028 & n12030;
  assign n12032 = ~n12029 & n12031;
  assign n12033 = P3_INSTQUEUE_REG_11__4_ & n11851;
  assign n12034 = P3_INSTQUEUE_REG_10__4_ & n11853;
  assign n12035 = P3_INSTQUEUE_REG_9__4_ & n11855;
  assign n12036 = P3_INSTQUEUE_REG_8__4_ & n11857;
  assign n12037 = ~n12033 & ~n12034;
  assign n12038 = ~n12035 & n12037;
  assign n12039 = ~n12036 & n12038;
  assign n12040 = n12018 & n12025;
  assign n12041 = n12032 & n12040;
  assign n12042 = n12039 & n12041;
  assign n12043 = n11353 & ~n12042;
  assign n12044 = ~n12011 & ~n12043;
  assign n12045 = P3_EAX_REG_19_ & n12001;
  assign n12046 = ~P3_EAX_REG_20_ & n12045;
  assign n12047 = P3_EAX_REG_20_ & ~n12045;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = n11359 & ~n12048;
  assign n12050 = ~n12009 & ~n12010;
  assign n12051 = n12044 & n12050;
  assign n2368 = n12049 | ~n12051;
  assign n12053 = BUF2_REG_21_ & n11804;
  assign n12054 = BUF2_REG_5_ & n11806;
  assign n12055 = P3_EAX_REG_21_ & ~n11352;
  assign n12056 = P3_INSTQUEUE_REG_7__5_ & n11815;
  assign n12057 = P3_INSTQUEUE_REG_6__5_ & n11817;
  assign n12058 = P3_INSTQUEUE_REG_5__5_ & n11819;
  assign n12059 = P3_INSTQUEUE_REG_4__5_ & n11821;
  assign n12060 = ~n12056 & ~n12057;
  assign n12061 = ~n12058 & n12060;
  assign n12062 = ~n12059 & n12061;
  assign n12063 = P3_INSTQUEUE_REG_3__5_ & n11827;
  assign n12064 = P3_INSTQUEUE_REG_2__5_ & n11829;
  assign n12065 = P3_INSTQUEUE_REG_1__5_ & n11831;
  assign n12066 = P3_INSTQUEUE_REG_0__5_ & n11833;
  assign n12067 = ~n12063 & ~n12064;
  assign n12068 = ~n12065 & n12067;
  assign n12069 = ~n12066 & n12068;
  assign n12070 = P3_INSTQUEUE_REG_15__5_ & n11839;
  assign n12071 = P3_INSTQUEUE_REG_14__5_ & n11841;
  assign n12072 = P3_INSTQUEUE_REG_13__5_ & n11843;
  assign n12073 = P3_INSTQUEUE_REG_12__5_ & n11845;
  assign n12074 = ~n12070 & ~n12071;
  assign n12075 = ~n12072 & n12074;
  assign n12076 = ~n12073 & n12075;
  assign n12077 = P3_INSTQUEUE_REG_11__5_ & n11851;
  assign n12078 = P3_INSTQUEUE_REG_10__5_ & n11853;
  assign n12079 = P3_INSTQUEUE_REG_9__5_ & n11855;
  assign n12080 = P3_INSTQUEUE_REG_8__5_ & n11857;
  assign n12081 = ~n12077 & ~n12078;
  assign n12082 = ~n12079 & n12081;
  assign n12083 = ~n12080 & n12082;
  assign n12084 = n12062 & n12069;
  assign n12085 = n12076 & n12084;
  assign n12086 = n12083 & n12085;
  assign n12087 = n11353 & ~n12086;
  assign n12088 = ~n12055 & ~n12087;
  assign n12089 = P3_EAX_REG_19_ & P3_EAX_REG_20_;
  assign n12090 = n12001 & n12089;
  assign n12091 = P3_EAX_REG_21_ & ~n12090;
  assign n12092 = ~P3_EAX_REG_21_ & n12090;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = n11359 & ~n12093;
  assign n12095 = ~n12053 & ~n12054;
  assign n12096 = n12088 & n12095;
  assign n2373 = n12094 | ~n12096;
  assign n12098 = BUF2_REG_22_ & n11804;
  assign n12099 = BUF2_REG_6_ & n11806;
  assign n12100 = P3_EAX_REG_22_ & ~n11352;
  assign n12101 = P3_INSTQUEUE_REG_7__6_ & n11815;
  assign n12102 = P3_INSTQUEUE_REG_6__6_ & n11817;
  assign n12103 = P3_INSTQUEUE_REG_5__6_ & n11819;
  assign n12104 = P3_INSTQUEUE_REG_4__6_ & n11821;
  assign n12105 = ~n12101 & ~n12102;
  assign n12106 = ~n12103 & n12105;
  assign n12107 = ~n12104 & n12106;
  assign n12108 = P3_INSTQUEUE_REG_3__6_ & n11827;
  assign n12109 = P3_INSTQUEUE_REG_2__6_ & n11829;
  assign n12110 = P3_INSTQUEUE_REG_1__6_ & n11831;
  assign n12111 = P3_INSTQUEUE_REG_0__6_ & n11833;
  assign n12112 = ~n12108 & ~n12109;
  assign n12113 = ~n12110 & n12112;
  assign n12114 = ~n12111 & n12113;
  assign n12115 = P3_INSTQUEUE_REG_15__6_ & n11839;
  assign n12116 = P3_INSTQUEUE_REG_14__6_ & n11841;
  assign n12117 = P3_INSTQUEUE_REG_13__6_ & n11843;
  assign n12118 = P3_INSTQUEUE_REG_12__6_ & n11845;
  assign n12119 = ~n12115 & ~n12116;
  assign n12120 = ~n12117 & n12119;
  assign n12121 = ~n12118 & n12120;
  assign n12122 = P3_INSTQUEUE_REG_11__6_ & n11851;
  assign n12123 = P3_INSTQUEUE_REG_10__6_ & n11853;
  assign n12124 = P3_INSTQUEUE_REG_9__6_ & n11855;
  assign n12125 = P3_INSTQUEUE_REG_8__6_ & n11857;
  assign n12126 = ~n12122 & ~n12123;
  assign n12127 = ~n12124 & n12126;
  assign n12128 = ~n12125 & n12127;
  assign n12129 = n12107 & n12114;
  assign n12130 = n12121 & n12129;
  assign n12131 = n12128 & n12130;
  assign n12132 = n11353 & ~n12131;
  assign n12133 = ~n12100 & ~n12132;
  assign n12134 = P3_EAX_REG_21_ & n12090;
  assign n12135 = ~P3_EAX_REG_22_ & n12134;
  assign n12136 = P3_EAX_REG_22_ & ~n12134;
  assign n12137 = ~n12135 & ~n12136;
  assign n12138 = n11359 & ~n12137;
  assign n12139 = ~n12098 & ~n12099;
  assign n12140 = n12133 & n12139;
  assign n2378 = n12138 | ~n12140;
  assign n12142 = BUF2_REG_23_ & n11804;
  assign n12143 = BUF2_REG_7_ & n11806;
  assign n12144 = P3_EAX_REG_23_ & ~n11352;
  assign n12145 = P3_INSTQUEUERD_ADDR_REG_3_ & ~P3_INSTQUEUERD_ADDR_REG_2_;
  assign n12146 = ~n5109 & ~n12145;
  assign n12147 = n5080 & n12146;
  assign n12148 = P3_INSTQUEUE_REG_7__0_ & n12147;
  assign n12149 = n5084_1 & n12146;
  assign n12150 = P3_INSTQUEUE_REG_6__0_ & n12149;
  assign n12151 = n5089 & n12146;
  assign n12152 = P3_INSTQUEUE_REG_5__0_ & n12151;
  assign n12153 = n5093 & n12146;
  assign n12154 = P3_INSTQUEUE_REG_4__0_ & n12153;
  assign n12155 = ~n12148 & ~n12150;
  assign n12156 = ~n12152 & n12155;
  assign n12157 = ~n12154 & n12156;
  assign n12158 = P3_INSTQUEUERD_ADDR_REG_2_ & n12146;
  assign n12159 = n5079_1 & n12158;
  assign n12160 = P3_INSTQUEUE_REG_3__0_ & n12159;
  assign n12161 = n5083 & n12158;
  assign n12162 = P3_INSTQUEUE_REG_2__0_ & n12161;
  assign n12163 = n5088_1 & n12158;
  assign n12164 = P3_INSTQUEUE_REG_1__0_ & n12163;
  assign n12165 = n5092_1 & n12158;
  assign n12166 = P3_INSTQUEUE_REG_0__0_ & n12165;
  assign n12167 = ~n12160 & ~n12162;
  assign n12168 = ~n12164 & n12167;
  assign n12169 = ~n12166 & n12168;
  assign n12170 = n5080 & ~n12146;
  assign n12171 = P3_INSTQUEUE_REG_15__0_ & n12170;
  assign n12172 = n5084_1 & ~n12146;
  assign n12173 = P3_INSTQUEUE_REG_14__0_ & n12172;
  assign n12174 = n5089 & ~n12146;
  assign n12175 = P3_INSTQUEUE_REG_13__0_ & n12174;
  assign n12176 = n5093 & ~n12146;
  assign n12177 = P3_INSTQUEUE_REG_12__0_ & n12176;
  assign n12178 = ~n12171 & ~n12173;
  assign n12179 = ~n12175 & n12178;
  assign n12180 = ~n12177 & n12179;
  assign n12181 = P3_INSTQUEUERD_ADDR_REG_2_ & ~n12146;
  assign n12182 = n5079_1 & n12181;
  assign n12183 = P3_INSTQUEUE_REG_11__0_ & n12182;
  assign n12184 = n5083 & n12181;
  assign n12185 = P3_INSTQUEUE_REG_10__0_ & n12184;
  assign n12186 = n5088_1 & n12181;
  assign n12187 = P3_INSTQUEUE_REG_9__0_ & n12186;
  assign n12188 = n5092_1 & n12181;
  assign n12189 = P3_INSTQUEUE_REG_8__0_ & n12188;
  assign n12190 = ~n12183 & ~n12185;
  assign n12191 = ~n12187 & n12190;
  assign n12192 = ~n12189 & n12191;
  assign n12193 = n12157 & n12169;
  assign n12194 = n12180 & n12193;
  assign n12195 = n12192 & n12194;
  assign n12196 = P3_INSTQUEUE_REG_7__7_ & n11815;
  assign n12197 = P3_INSTQUEUE_REG_6__7_ & n11817;
  assign n12198 = P3_INSTQUEUE_REG_5__7_ & n11819;
  assign n12199 = P3_INSTQUEUE_REG_4__7_ & n11821;
  assign n12200 = ~n12196 & ~n12197;
  assign n12201 = ~n12198 & n12200;
  assign n12202 = ~n12199 & n12201;
  assign n12203 = P3_INSTQUEUE_REG_3__7_ & n11827;
  assign n12204 = P3_INSTQUEUE_REG_2__7_ & n11829;
  assign n12205 = P3_INSTQUEUE_REG_1__7_ & n11831;
  assign n12206 = P3_INSTQUEUE_REG_0__7_ & n11833;
  assign n12207 = ~n12203 & ~n12204;
  assign n12208 = ~n12205 & n12207;
  assign n12209 = ~n12206 & n12208;
  assign n12210 = P3_INSTQUEUE_REG_15__7_ & n11839;
  assign n12211 = P3_INSTQUEUE_REG_14__7_ & n11841;
  assign n12212 = P3_INSTQUEUE_REG_13__7_ & n11843;
  assign n12213 = P3_INSTQUEUE_REG_12__7_ & n11845;
  assign n12214 = ~n12210 & ~n12211;
  assign n12215 = ~n12212 & n12214;
  assign n12216 = ~n12213 & n12215;
  assign n12217 = P3_INSTQUEUE_REG_11__7_ & n11851;
  assign n12218 = P3_INSTQUEUE_REG_10__7_ & n11853;
  assign n12219 = P3_INSTQUEUE_REG_9__7_ & n11855;
  assign n12220 = P3_INSTQUEUE_REG_8__7_ & n11857;
  assign n12221 = ~n12217 & ~n12218;
  assign n12222 = ~n12219 & n12221;
  assign n12223 = ~n12220 & n12222;
  assign n12224 = n12202 & n12209;
  assign n12225 = n12216 & n12224;
  assign n12226 = n12223 & n12225;
  assign n12227 = ~n12195 & n12226;
  assign n12228 = n12195 & ~n12226;
  assign n12229 = ~n12227 & ~n12228;
  assign n12230 = n11353 & ~n12229;
  assign n12231 = ~n12144 & ~n12230;
  assign n12232 = P3_EAX_REG_21_ & P3_EAX_REG_22_;
  assign n12233 = n12090 & n12232;
  assign n12234 = P3_EAX_REG_23_ & ~n12233;
  assign n12235 = ~P3_EAX_REG_23_ & n12233;
  assign n12236 = ~n12234 & ~n12235;
  assign n12237 = n11359 & ~n12236;
  assign n12238 = ~n12142 & ~n12143;
  assign n12239 = n12231 & n12238;
  assign n2383 = n12237 | ~n12239;
  assign n12241 = BUF2_REG_24_ & n11804;
  assign n12242 = BUF2_REG_8_ & n11806;
  assign n12243 = P3_EAX_REG_24_ & ~n11352;
  assign n12244 = ~n12195 & ~n12226;
  assign n12245 = P3_INSTQUEUE_REG_7__1_ & n12147;
  assign n12246 = P3_INSTQUEUE_REG_6__1_ & n12149;
  assign n12247 = P3_INSTQUEUE_REG_5__1_ & n12151;
  assign n12248 = P3_INSTQUEUE_REG_4__1_ & n12153;
  assign n12249 = ~n12245 & ~n12246;
  assign n12250 = ~n12247 & n12249;
  assign n12251 = ~n12248 & n12250;
  assign n12252 = P3_INSTQUEUE_REG_3__1_ & n12159;
  assign n12253 = P3_INSTQUEUE_REG_2__1_ & n12161;
  assign n12254 = P3_INSTQUEUE_REG_1__1_ & n12163;
  assign n12255 = P3_INSTQUEUE_REG_0__1_ & n12165;
  assign n12256 = ~n12252 & ~n12253;
  assign n12257 = ~n12254 & n12256;
  assign n12258 = ~n12255 & n12257;
  assign n12259 = P3_INSTQUEUE_REG_15__1_ & n12170;
  assign n12260 = P3_INSTQUEUE_REG_14__1_ & n12172;
  assign n12261 = P3_INSTQUEUE_REG_13__1_ & n12174;
  assign n12262 = P3_INSTQUEUE_REG_12__1_ & n12176;
  assign n12263 = ~n12259 & ~n12260;
  assign n12264 = ~n12261 & n12263;
  assign n12265 = ~n12262 & n12264;
  assign n12266 = P3_INSTQUEUE_REG_11__1_ & n12182;
  assign n12267 = P3_INSTQUEUE_REG_10__1_ & n12184;
  assign n12268 = P3_INSTQUEUE_REG_9__1_ & n12186;
  assign n12269 = P3_INSTQUEUE_REG_8__1_ & n12188;
  assign n12270 = ~n12266 & ~n12267;
  assign n12271 = ~n12268 & n12270;
  assign n12272 = ~n12269 & n12271;
  assign n12273 = n12251 & n12258;
  assign n12274 = n12265 & n12273;
  assign n12275 = n12272 & n12274;
  assign n12276 = n12244 & n12275;
  assign n12277 = ~n12244 & ~n12275;
  assign n12278 = ~n12276 & ~n12277;
  assign n12279 = n11353 & ~n12278;
  assign n12280 = ~n12243 & ~n12279;
  assign n12281 = P3_EAX_REG_23_ & n12233;
  assign n12282 = ~P3_EAX_REG_24_ & n12281;
  assign n12283 = P3_EAX_REG_24_ & ~n12281;
  assign n12284 = ~n12282 & ~n12283;
  assign n12285 = n11359 & ~n12284;
  assign n12286 = ~n12241 & ~n12242;
  assign n12287 = n12280 & n12286;
  assign n2388 = n12285 | ~n12287;
  assign n12289 = BUF2_REG_25_ & n11804;
  assign n12290 = BUF2_REG_9_ & n11806;
  assign n12291 = P3_EAX_REG_25_ & ~n11352;
  assign n12292 = n12244 & ~n12275;
  assign n12293 = P3_INSTQUEUE_REG_7__2_ & n12147;
  assign n12294 = P3_INSTQUEUE_REG_6__2_ & n12149;
  assign n12295 = P3_INSTQUEUE_REG_5__2_ & n12151;
  assign n12296 = P3_INSTQUEUE_REG_4__2_ & n12153;
  assign n12297 = ~n12293 & ~n12294;
  assign n12298 = ~n12295 & n12297;
  assign n12299 = ~n12296 & n12298;
  assign n12300 = P3_INSTQUEUE_REG_3__2_ & n12159;
  assign n12301 = P3_INSTQUEUE_REG_2__2_ & n12161;
  assign n12302 = P3_INSTQUEUE_REG_1__2_ & n12163;
  assign n12303 = P3_INSTQUEUE_REG_0__2_ & n12165;
  assign n12304 = ~n12300 & ~n12301;
  assign n12305 = ~n12302 & n12304;
  assign n12306 = ~n12303 & n12305;
  assign n12307 = P3_INSTQUEUE_REG_15__2_ & n12170;
  assign n12308 = P3_INSTQUEUE_REG_14__2_ & n12172;
  assign n12309 = P3_INSTQUEUE_REG_13__2_ & n12174;
  assign n12310 = P3_INSTQUEUE_REG_12__2_ & n12176;
  assign n12311 = ~n12307 & ~n12308;
  assign n12312 = ~n12309 & n12311;
  assign n12313 = ~n12310 & n12312;
  assign n12314 = P3_INSTQUEUE_REG_11__2_ & n12182;
  assign n12315 = P3_INSTQUEUE_REG_10__2_ & n12184;
  assign n12316 = P3_INSTQUEUE_REG_9__2_ & n12186;
  assign n12317 = P3_INSTQUEUE_REG_8__2_ & n12188;
  assign n12318 = ~n12314 & ~n12315;
  assign n12319 = ~n12316 & n12318;
  assign n12320 = ~n12317 & n12319;
  assign n12321 = n12299 & n12306;
  assign n12322 = n12313 & n12321;
  assign n12323 = n12320 & n12322;
  assign n12324 = n12292 & n12323;
  assign n12325 = ~n12292 & ~n12323;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = n11353 & ~n12326;
  assign n12328 = ~n12291 & ~n12327;
  assign n12329 = P3_EAX_REG_23_ & P3_EAX_REG_24_;
  assign n12330 = n12233 & n12329;
  assign n12331 = P3_EAX_REG_25_ & ~n12330;
  assign n12332 = ~P3_EAX_REG_25_ & n12330;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = n11359 & ~n12333;
  assign n12335 = ~n12289 & ~n12290;
  assign n12336 = n12328 & n12335;
  assign n2393 = n12334 | ~n12336;
  assign n12338 = BUF2_REG_26_ & n11804;
  assign n12339 = BUF2_REG_10_ & n11806;
  assign n12340 = P3_EAX_REG_26_ & ~n11352;
  assign n12341 = n12292 & ~n12323;
  assign n12342 = P3_INSTQUEUE_REG_7__3_ & n12147;
  assign n12343 = P3_INSTQUEUE_REG_6__3_ & n12149;
  assign n12344 = P3_INSTQUEUE_REG_5__3_ & n12151;
  assign n12345 = P3_INSTQUEUE_REG_4__3_ & n12153;
  assign n12346 = ~n12342 & ~n12343;
  assign n12347 = ~n12344 & n12346;
  assign n12348 = ~n12345 & n12347;
  assign n12349 = P3_INSTQUEUE_REG_3__3_ & n12159;
  assign n12350 = P3_INSTQUEUE_REG_2__3_ & n12161;
  assign n12351 = P3_INSTQUEUE_REG_1__3_ & n12163;
  assign n12352 = P3_INSTQUEUE_REG_0__3_ & n12165;
  assign n12353 = ~n12349 & ~n12350;
  assign n12354 = ~n12351 & n12353;
  assign n12355 = ~n12352 & n12354;
  assign n12356 = P3_INSTQUEUE_REG_15__3_ & n12170;
  assign n12357 = P3_INSTQUEUE_REG_14__3_ & n12172;
  assign n12358 = P3_INSTQUEUE_REG_13__3_ & n12174;
  assign n12359 = P3_INSTQUEUE_REG_12__3_ & n12176;
  assign n12360 = ~n12356 & ~n12357;
  assign n12361 = ~n12358 & n12360;
  assign n12362 = ~n12359 & n12361;
  assign n12363 = P3_INSTQUEUE_REG_11__3_ & n12182;
  assign n12364 = P3_INSTQUEUE_REG_10__3_ & n12184;
  assign n12365 = P3_INSTQUEUE_REG_9__3_ & n12186;
  assign n12366 = P3_INSTQUEUE_REG_8__3_ & n12188;
  assign n12367 = ~n12363 & ~n12364;
  assign n12368 = ~n12365 & n12367;
  assign n12369 = ~n12366 & n12368;
  assign n12370 = n12348 & n12355;
  assign n12371 = n12362 & n12370;
  assign n12372 = n12369 & n12371;
  assign n12373 = n12341 & n12372;
  assign n12374 = ~n12341 & ~n12372;
  assign n12375 = ~n12373 & ~n12374;
  assign n12376 = n11353 & ~n12375;
  assign n12377 = ~n12340 & ~n12376;
  assign n12378 = P3_EAX_REG_25_ & n12330;
  assign n12379 = ~P3_EAX_REG_26_ & n12378;
  assign n12380 = P3_EAX_REG_26_ & ~n12378;
  assign n12381 = ~n12379 & ~n12380;
  assign n12382 = n11359 & ~n12381;
  assign n12383 = ~n12338 & ~n12339;
  assign n12384 = n12377 & n12383;
  assign n2398 = n12382 | ~n12384;
  assign n12386 = BUF2_REG_27_ & n11804;
  assign n12387 = BUF2_REG_11_ & n11806;
  assign n12388 = P3_EAX_REG_27_ & ~n11352;
  assign n12389 = n12341 & ~n12372;
  assign n12390 = P3_INSTQUEUE_REG_7__4_ & n12147;
  assign n12391 = P3_INSTQUEUE_REG_6__4_ & n12149;
  assign n12392 = P3_INSTQUEUE_REG_5__4_ & n12151;
  assign n12393 = P3_INSTQUEUE_REG_4__4_ & n12153;
  assign n12394 = ~n12390 & ~n12391;
  assign n12395 = ~n12392 & n12394;
  assign n12396 = ~n12393 & n12395;
  assign n12397 = P3_INSTQUEUE_REG_3__4_ & n12159;
  assign n12398 = P3_INSTQUEUE_REG_2__4_ & n12161;
  assign n12399 = P3_INSTQUEUE_REG_1__4_ & n12163;
  assign n12400 = P3_INSTQUEUE_REG_0__4_ & n12165;
  assign n12401 = ~n12397 & ~n12398;
  assign n12402 = ~n12399 & n12401;
  assign n12403 = ~n12400 & n12402;
  assign n12404 = P3_INSTQUEUE_REG_15__4_ & n12170;
  assign n12405 = P3_INSTQUEUE_REG_14__4_ & n12172;
  assign n12406 = P3_INSTQUEUE_REG_13__4_ & n12174;
  assign n12407 = P3_INSTQUEUE_REG_12__4_ & n12176;
  assign n12408 = ~n12404 & ~n12405;
  assign n12409 = ~n12406 & n12408;
  assign n12410 = ~n12407 & n12409;
  assign n12411 = P3_INSTQUEUE_REG_11__4_ & n12182;
  assign n12412 = P3_INSTQUEUE_REG_10__4_ & n12184;
  assign n12413 = P3_INSTQUEUE_REG_9__4_ & n12186;
  assign n12414 = P3_INSTQUEUE_REG_8__4_ & n12188;
  assign n12415 = ~n12411 & ~n12412;
  assign n12416 = ~n12413 & n12415;
  assign n12417 = ~n12414 & n12416;
  assign n12418 = n12396 & n12403;
  assign n12419 = n12410 & n12418;
  assign n12420 = n12417 & n12419;
  assign n12421 = n12389 & n12420;
  assign n12422 = ~n12389 & ~n12420;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = n11353 & ~n12423;
  assign n12425 = ~n12388 & ~n12424;
  assign n12426 = P3_EAX_REG_25_ & P3_EAX_REG_26_;
  assign n12427 = n12330 & n12426;
  assign n12428 = P3_EAX_REG_27_ & ~n12427;
  assign n12429 = ~P3_EAX_REG_27_ & n12427;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = n11359 & ~n12430;
  assign n12432 = ~n12386 & ~n12387;
  assign n12433 = n12425 & n12432;
  assign n2403 = n12431 | ~n12433;
  assign n12435 = BUF2_REG_28_ & n11804;
  assign n12436 = BUF2_REG_12_ & n11806;
  assign n12437 = P3_EAX_REG_28_ & ~n11352;
  assign n12438 = n12389 & ~n12420;
  assign n12439 = P3_INSTQUEUE_REG_7__5_ & n12147;
  assign n12440 = P3_INSTQUEUE_REG_6__5_ & n12149;
  assign n12441 = P3_INSTQUEUE_REG_5__5_ & n12151;
  assign n12442 = P3_INSTQUEUE_REG_4__5_ & n12153;
  assign n12443 = ~n12439 & ~n12440;
  assign n12444 = ~n12441 & n12443;
  assign n12445 = ~n12442 & n12444;
  assign n12446 = P3_INSTQUEUE_REG_3__5_ & n12159;
  assign n12447 = P3_INSTQUEUE_REG_2__5_ & n12161;
  assign n12448 = P3_INSTQUEUE_REG_1__5_ & n12163;
  assign n12449 = P3_INSTQUEUE_REG_0__5_ & n12165;
  assign n12450 = ~n12446 & ~n12447;
  assign n12451 = ~n12448 & n12450;
  assign n12452 = ~n12449 & n12451;
  assign n12453 = P3_INSTQUEUE_REG_15__5_ & n12170;
  assign n12454 = P3_INSTQUEUE_REG_14__5_ & n12172;
  assign n12455 = P3_INSTQUEUE_REG_13__5_ & n12174;
  assign n12456 = P3_INSTQUEUE_REG_12__5_ & n12176;
  assign n12457 = ~n12453 & ~n12454;
  assign n12458 = ~n12455 & n12457;
  assign n12459 = ~n12456 & n12458;
  assign n12460 = P3_INSTQUEUE_REG_11__5_ & n12182;
  assign n12461 = P3_INSTQUEUE_REG_10__5_ & n12184;
  assign n12462 = P3_INSTQUEUE_REG_9__5_ & n12186;
  assign n12463 = P3_INSTQUEUE_REG_8__5_ & n12188;
  assign n12464 = ~n12460 & ~n12461;
  assign n12465 = ~n12462 & n12464;
  assign n12466 = ~n12463 & n12465;
  assign n12467 = n12445 & n12452;
  assign n12468 = n12459 & n12467;
  assign n12469 = n12466 & n12468;
  assign n12470 = n12438 & n12469;
  assign n12471 = ~n12438 & ~n12469;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = n11353 & ~n12472;
  assign n12474 = P3_EAX_REG_27_ & n12427;
  assign n12475 = ~P3_EAX_REG_28_ & n12474;
  assign n12476 = P3_EAX_REG_28_ & ~n12474;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = n11359 & ~n12477;
  assign n12479 = ~n12435 & ~n12436;
  assign n12480 = ~n12437 & n12479;
  assign n12481 = ~n12473 & n12480;
  assign n2408 = n12478 | ~n12481;
  assign n12483 = BUF2_REG_29_ & n11804;
  assign n12484 = BUF2_REG_13_ & n11806;
  assign n12485 = P3_EAX_REG_29_ & ~n11352;
  assign n12486 = n12438 & ~n12469;
  assign n12487 = P3_INSTQUEUE_REG_7__6_ & n12147;
  assign n12488 = P3_INSTQUEUE_REG_6__6_ & n12149;
  assign n12489 = P3_INSTQUEUE_REG_5__6_ & n12151;
  assign n12490 = P3_INSTQUEUE_REG_4__6_ & n12153;
  assign n12491 = ~n12487 & ~n12488;
  assign n12492 = ~n12489 & n12491;
  assign n12493 = ~n12490 & n12492;
  assign n12494 = P3_INSTQUEUE_REG_3__6_ & n12159;
  assign n12495 = P3_INSTQUEUE_REG_2__6_ & n12161;
  assign n12496 = P3_INSTQUEUE_REG_1__6_ & n12163;
  assign n12497 = P3_INSTQUEUE_REG_0__6_ & n12165;
  assign n12498 = ~n12494 & ~n12495;
  assign n12499 = ~n12496 & n12498;
  assign n12500 = ~n12497 & n12499;
  assign n12501 = P3_INSTQUEUE_REG_15__6_ & n12170;
  assign n12502 = P3_INSTQUEUE_REG_14__6_ & n12172;
  assign n12503 = P3_INSTQUEUE_REG_13__6_ & n12174;
  assign n12504 = P3_INSTQUEUE_REG_12__6_ & n12176;
  assign n12505 = ~n12501 & ~n12502;
  assign n12506 = ~n12503 & n12505;
  assign n12507 = ~n12504 & n12506;
  assign n12508 = P3_INSTQUEUE_REG_11__6_ & n12182;
  assign n12509 = P3_INSTQUEUE_REG_10__6_ & n12184;
  assign n12510 = P3_INSTQUEUE_REG_9__6_ & n12186;
  assign n12511 = P3_INSTQUEUE_REG_8__6_ & n12188;
  assign n12512 = ~n12508 & ~n12509;
  assign n12513 = ~n12510 & n12512;
  assign n12514 = ~n12511 & n12513;
  assign n12515 = n12493 & n12500;
  assign n12516 = n12507 & n12515;
  assign n12517 = n12514 & n12516;
  assign n12518 = n12486 & n12517;
  assign n12519 = ~n12486 & ~n12517;
  assign n12520 = ~n12518 & ~n12519;
  assign n12521 = n11353 & ~n12520;
  assign n12522 = P3_EAX_REG_27_ & P3_EAX_REG_28_;
  assign n12523 = n12427 & n12522;
  assign n12524 = P3_EAX_REG_29_ & ~n12523;
  assign n12525 = ~P3_EAX_REG_29_ & n12523;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = n11359 & ~n12526;
  assign n12528 = ~n12483 & ~n12484;
  assign n12529 = ~n12485 & n12528;
  assign n12530 = ~n12521 & n12529;
  assign n2413 = n12527 | ~n12530;
  assign n12532 = BUF2_REG_30_ & n11804;
  assign n12533 = BUF2_REG_14_ & n11806;
  assign n12534 = P3_EAX_REG_30_ & ~n11352;
  assign n12535 = n12486 & ~n12517;
  assign n12536 = P3_INSTQUEUE_REG_7__7_ & n12147;
  assign n12537 = P3_INSTQUEUE_REG_6__7_ & n12149;
  assign n12538 = P3_INSTQUEUE_REG_5__7_ & n12151;
  assign n12539 = P3_INSTQUEUE_REG_4__7_ & n12153;
  assign n12540 = ~n12536 & ~n12537;
  assign n12541 = ~n12538 & n12540;
  assign n12542 = ~n12539 & n12541;
  assign n12543 = P3_INSTQUEUE_REG_3__7_ & n12159;
  assign n12544 = P3_INSTQUEUE_REG_2__7_ & n12161;
  assign n12545 = P3_INSTQUEUE_REG_1__7_ & n12163;
  assign n12546 = P3_INSTQUEUE_REG_0__7_ & n12165;
  assign n12547 = ~n12543 & ~n12544;
  assign n12548 = ~n12545 & n12547;
  assign n12549 = ~n12546 & n12548;
  assign n12550 = P3_INSTQUEUE_REG_15__7_ & n12170;
  assign n12551 = P3_INSTQUEUE_REG_14__7_ & n12172;
  assign n12552 = P3_INSTQUEUE_REG_13__7_ & n12174;
  assign n12553 = P3_INSTQUEUE_REG_12__7_ & n12176;
  assign n12554 = ~n12550 & ~n12551;
  assign n12555 = ~n12552 & n12554;
  assign n12556 = ~n12553 & n12555;
  assign n12557 = P3_INSTQUEUE_REG_11__7_ & n12182;
  assign n12558 = P3_INSTQUEUE_REG_10__7_ & n12184;
  assign n12559 = P3_INSTQUEUE_REG_9__7_ & n12186;
  assign n12560 = P3_INSTQUEUE_REG_8__7_ & n12188;
  assign n12561 = ~n12557 & ~n12558;
  assign n12562 = ~n12559 & n12561;
  assign n12563 = ~n12560 & n12562;
  assign n12564 = n12542 & n12549;
  assign n12565 = n12556 & n12564;
  assign n12566 = n12563 & n12565;
  assign n12567 = n12535 & n12566;
  assign n12568 = ~n12535 & ~n12566;
  assign n12569 = ~n12567 & ~n12568;
  assign n12570 = n11353 & ~n12569;
  assign n12571 = P3_EAX_REG_29_ & n12523;
  assign n12572 = ~P3_EAX_REG_30_ & n12571;
  assign n12573 = P3_EAX_REG_30_ & ~n12571;
  assign n12574 = ~n12572 & ~n12573;
  assign n12575 = n11359 & ~n12574;
  assign n12576 = ~n12532 & ~n12533;
  assign n12577 = ~n12534 & n12576;
  assign n12578 = ~n12570 & n12577;
  assign n2418 = n12575 | ~n12578;
  assign n12580 = P3_EAX_REG_31_ & ~n11352;
  assign n12581 = BUF2_REG_31_ & n11804;
  assign n12582 = P3_EAX_REG_30_ & n12571;
  assign n12583 = ~P3_EAX_REG_31_ & n12582;
  assign n12584 = P3_EAX_REG_31_ & ~n12582;
  assign n12585 = ~n12583 & ~n12584;
  assign n12586 = n11359 & ~n12585;
  assign n12587 = ~n12580 & ~n12581;
  assign n2423 = n12586 | ~n12587;
  assign n12589 = ~n5500 & ~n5594_1;
  assign n12590 = n5713 & ~n12589;
  assign n12591 = n5230 & n12590;
  assign n12592 = ~P3_EBX_REG_0_ & n12591;
  assign n12593 = ~n5230 & n12590;
  assign n12594 = P3_INSTQUEUE_REG_0__0_ & n12593;
  assign n12595 = P3_EBX_REG_0_ & ~n12590;
  assign n12596 = ~n12592 & ~n12594;
  assign n2428 = n12595 | ~n12596;
  assign n12598 = ~P3_EBX_REG_0_ & P3_EBX_REG_1_;
  assign n12599 = P3_EBX_REG_0_ & ~P3_EBX_REG_1_;
  assign n12600 = ~n12598 & ~n12599;
  assign n12601 = n12591 & ~n12600;
  assign n12602 = P3_INSTQUEUE_REG_0__1_ & n12593;
  assign n12603 = P3_EBX_REG_1_ & ~n12590;
  assign n12604 = ~n12601 & ~n12602;
  assign n2433 = n12603 | ~n12604;
  assign n12606 = P3_EBX_REG_0_ & P3_EBX_REG_1_;
  assign n12607 = ~P3_EBX_REG_2_ & n12606;
  assign n12608 = P3_EBX_REG_2_ & ~n12606;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = n12591 & ~n12609;
  assign n12611 = P3_INSTQUEUE_REG_0__2_ & n12593;
  assign n12612 = P3_EBX_REG_2_ & ~n12590;
  assign n12613 = ~n12610 & ~n12611;
  assign n2438 = n12612 | ~n12613;
  assign n12615 = P3_EBX_REG_0_ & P3_EBX_REG_2_;
  assign n12616 = P3_EBX_REG_1_ & n12615;
  assign n12617 = P3_EBX_REG_3_ & ~n12616;
  assign n12618 = ~P3_EBX_REG_3_ & n12616;
  assign n12619 = ~n12617 & ~n12618;
  assign n12620 = n12591 & ~n12619;
  assign n12621 = P3_INSTQUEUE_REG_0__3_ & n12593;
  assign n12622 = P3_EBX_REG_3_ & ~n12590;
  assign n12623 = ~n12620 & ~n12621;
  assign n2443 = n12622 | ~n12623;
  assign n12625 = P3_EBX_REG_3_ & n12616;
  assign n12626 = ~P3_EBX_REG_4_ & n12625;
  assign n12627 = P3_EBX_REG_4_ & ~n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = n12591 & ~n12628;
  assign n12630 = P3_INSTQUEUE_REG_0__4_ & n12593;
  assign n12631 = P3_EBX_REG_4_ & ~n12590;
  assign n12632 = ~n12629 & ~n12630;
  assign n2448 = n12631 | ~n12632;
  assign n12634 = P3_EBX_REG_3_ & P3_EBX_REG_4_;
  assign n12635 = n12616 & n12634;
  assign n12636 = P3_EBX_REG_5_ & ~n12635;
  assign n12637 = ~P3_EBX_REG_5_ & n12635;
  assign n12638 = ~n12636 & ~n12637;
  assign n12639 = n12591 & ~n12638;
  assign n12640 = P3_INSTQUEUE_REG_0__5_ & n12593;
  assign n12641 = P3_EBX_REG_5_ & ~n12590;
  assign n12642 = ~n12639 & ~n12640;
  assign n2453 = n12641 | ~n12642;
  assign n12644 = P3_EBX_REG_5_ & n12635;
  assign n12645 = ~P3_EBX_REG_6_ & n12644;
  assign n12646 = P3_EBX_REG_6_ & ~n12644;
  assign n12647 = ~n12645 & ~n12646;
  assign n12648 = n12591 & ~n12647;
  assign n12649 = P3_INSTQUEUE_REG_0__6_ & n12593;
  assign n12650 = P3_EBX_REG_6_ & ~n12590;
  assign n12651 = ~n12648 & ~n12649;
  assign n2458 = n12650 | ~n12651;
  assign n12653 = P3_EBX_REG_5_ & P3_EBX_REG_6_;
  assign n12654 = n12635 & n12653;
  assign n12655 = P3_EBX_REG_7_ & ~n12654;
  assign n12656 = ~P3_EBX_REG_7_ & n12654;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = n12591 & ~n12657;
  assign n12659 = P3_INSTQUEUE_REG_0__7_ & n12593;
  assign n12660 = P3_EBX_REG_7_ & ~n12590;
  assign n12661 = ~n12658 & ~n12659;
  assign n2463 = n12660 | ~n12661;
  assign n12663 = P3_EBX_REG_7_ & n12654;
  assign n12664 = ~P3_EBX_REG_8_ & n12663;
  assign n12665 = P3_EBX_REG_8_ & ~n12663;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = n12591 & ~n12666;
  assign n12668 = ~n11494 & n12593;
  assign n12669 = P3_EBX_REG_8_ & ~n12590;
  assign n12670 = ~n12667 & ~n12668;
  assign n2468 = n12669 | ~n12670;
  assign n12672 = P3_EBX_REG_7_ & P3_EBX_REG_8_;
  assign n12673 = n12654 & n12672;
  assign n12674 = P3_EBX_REG_9_ & ~n12673;
  assign n12675 = ~P3_EBX_REG_9_ & n12673;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = n12591 & ~n12676;
  assign n12678 = ~n11536 & n12593;
  assign n12679 = P3_EBX_REG_9_ & ~n12590;
  assign n12680 = ~n12677 & ~n12678;
  assign n2473 = n12679 | ~n12680;
  assign n12682 = P3_EBX_REG_10_ & ~n12590;
  assign n12683 = ~n11579 & n12593;
  assign n12684 = P3_EBX_REG_9_ & n12673;
  assign n12685 = ~P3_EBX_REG_10_ & n12684;
  assign n12686 = P3_EBX_REG_10_ & ~n12684;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = n12591 & ~n12687;
  assign n12689 = ~n12682 & ~n12683;
  assign n2478 = n12688 | ~n12689;
  assign n12691 = P3_EBX_REG_11_ & ~n12590;
  assign n12692 = ~n11621 & n12593;
  assign n12693 = P3_EBX_REG_9_ & P3_EBX_REG_10_;
  assign n12694 = n12673 & n12693;
  assign n12695 = P3_EBX_REG_11_ & ~n12694;
  assign n12696 = ~P3_EBX_REG_11_ & n12694;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = n12591 & ~n12697;
  assign n12699 = ~n12691 & ~n12692;
  assign n2483 = n12698 | ~n12699;
  assign n12701 = P3_EBX_REG_12_ & ~n12590;
  assign n12702 = ~n11664 & n12593;
  assign n12703 = P3_EBX_REG_11_ & n12694;
  assign n12704 = ~P3_EBX_REG_12_ & n12703;
  assign n12705 = P3_EBX_REG_12_ & ~n12703;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = n12591 & ~n12706;
  assign n12708 = ~n12701 & ~n12702;
  assign n2488 = n12707 | ~n12708;
  assign n12710 = P3_EBX_REG_13_ & ~n12590;
  assign n12711 = ~n11707 & n12593;
  assign n12712 = P3_EBX_REG_11_ & P3_EBX_REG_12_;
  assign n12713 = n12694 & n12712;
  assign n12714 = P3_EBX_REG_13_ & ~n12713;
  assign n12715 = ~P3_EBX_REG_13_ & n12713;
  assign n12716 = ~n12714 & ~n12715;
  assign n12717 = n12591 & ~n12716;
  assign n12718 = ~n12710 & ~n12711;
  assign n2493 = n12717 | ~n12718;
  assign n12720 = P3_EBX_REG_14_ & ~n12590;
  assign n12721 = ~n11750 & n12593;
  assign n12722 = P3_EBX_REG_13_ & n12713;
  assign n12723 = ~P3_EBX_REG_14_ & n12722;
  assign n12724 = P3_EBX_REG_14_ & ~n12722;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = n12591 & ~n12725;
  assign n12727 = ~n12720 & ~n12721;
  assign n2498 = n12726 | ~n12727;
  assign n12729 = P3_EBX_REG_15_ & ~n12590;
  assign n12730 = ~n11792 & n12593;
  assign n12731 = P3_EBX_REG_13_ & P3_EBX_REG_14_;
  assign n12732 = n12713 & n12731;
  assign n12733 = P3_EBX_REG_15_ & ~n12732;
  assign n12734 = ~P3_EBX_REG_15_ & n12732;
  assign n12735 = ~n12733 & ~n12734;
  assign n12736 = n12591 & ~n12735;
  assign n12737 = ~n12729 & ~n12730;
  assign n2503 = n12736 | ~n12737;
  assign n12739 = P3_EBX_REG_16_ & ~n12590;
  assign n12740 = ~n11864 & n12593;
  assign n12741 = P3_EBX_REG_15_ & n12732;
  assign n12742 = ~P3_EBX_REG_16_ & n12741;
  assign n12743 = P3_EBX_REG_16_ & ~n12741;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = n12591 & ~n12744;
  assign n12746 = ~n12739 & ~n12740;
  assign n2508 = n12745 | ~n12746;
  assign n12748 = P3_EBX_REG_17_ & ~n12590;
  assign n12749 = ~n11908 & n12593;
  assign n12750 = P3_EBX_REG_15_ & P3_EBX_REG_16_;
  assign n12751 = n12732 & n12750;
  assign n12752 = P3_EBX_REG_17_ & ~n12751;
  assign n12753 = ~P3_EBX_REG_17_ & n12751;
  assign n12754 = ~n12752 & ~n12753;
  assign n12755 = n12591 & ~n12754;
  assign n12756 = ~n12748 & ~n12749;
  assign n2513 = n12755 | ~n12756;
  assign n12758 = P3_EBX_REG_18_ & ~n12590;
  assign n12759 = ~n11953 & n12593;
  assign n12760 = P3_EBX_REG_17_ & n12751;
  assign n12761 = ~P3_EBX_REG_18_ & n12760;
  assign n12762 = P3_EBX_REG_18_ & ~n12760;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = n12591 & ~n12763;
  assign n12765 = ~n12758 & ~n12759;
  assign n2518 = n12764 | ~n12765;
  assign n12767 = P3_EBX_REG_19_ & ~n12590;
  assign n12768 = ~n11997 & n12593;
  assign n12769 = P3_EBX_REG_17_ & P3_EBX_REG_18_;
  assign n12770 = n12751 & n12769;
  assign n12771 = P3_EBX_REG_19_ & ~n12770;
  assign n12772 = ~P3_EBX_REG_19_ & n12770;
  assign n12773 = ~n12771 & ~n12772;
  assign n12774 = n12591 & ~n12773;
  assign n12775 = ~n12767 & ~n12768;
  assign n2523 = n12774 | ~n12775;
  assign n12777 = P3_EBX_REG_20_ & ~n12590;
  assign n12778 = ~n12042 & n12593;
  assign n12779 = P3_EBX_REG_19_ & n12770;
  assign n12780 = ~P3_EBX_REG_20_ & n12779;
  assign n12781 = P3_EBX_REG_20_ & ~n12779;
  assign n12782 = ~n12780 & ~n12781;
  assign n12783 = n12591 & ~n12782;
  assign n12784 = ~n12777 & ~n12778;
  assign n2528 = n12783 | ~n12784;
  assign n12786 = P3_EBX_REG_21_ & ~n12590;
  assign n12787 = ~n12086 & n12593;
  assign n12788 = P3_EBX_REG_19_ & P3_EBX_REG_20_;
  assign n12789 = n12770 & n12788;
  assign n12790 = P3_EBX_REG_21_ & ~n12789;
  assign n12791 = ~P3_EBX_REG_21_ & n12789;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = n12591 & ~n12792;
  assign n12794 = ~n12786 & ~n12787;
  assign n2533 = n12793 | ~n12794;
  assign n12796 = P3_EBX_REG_22_ & ~n12590;
  assign n12797 = ~n12131 & n12593;
  assign n12798 = P3_EBX_REG_21_ & n12789;
  assign n12799 = ~P3_EBX_REG_22_ & n12798;
  assign n12800 = P3_EBX_REG_22_ & ~n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = n12591 & ~n12801;
  assign n12803 = ~n12796 & ~n12797;
  assign n2538 = n12802 | ~n12803;
  assign n12805 = P3_EBX_REG_23_ & ~n12590;
  assign n12806 = ~n12229 & n12593;
  assign n12807 = P3_EBX_REG_21_ & P3_EBX_REG_22_;
  assign n12808 = n12789 & n12807;
  assign n12809 = P3_EBX_REG_23_ & ~n12808;
  assign n12810 = ~P3_EBX_REG_23_ & n12808;
  assign n12811 = ~n12809 & ~n12810;
  assign n12812 = n12591 & ~n12811;
  assign n12813 = ~n12805 & ~n12806;
  assign n2543 = n12812 | ~n12813;
  assign n12815 = P3_EBX_REG_24_ & ~n12590;
  assign n12816 = ~n12278 & n12593;
  assign n12817 = P3_EBX_REG_23_ & n12808;
  assign n12818 = ~P3_EBX_REG_24_ & n12817;
  assign n12819 = P3_EBX_REG_24_ & ~n12817;
  assign n12820 = ~n12818 & ~n12819;
  assign n12821 = n12591 & ~n12820;
  assign n12822 = ~n12815 & ~n12816;
  assign n2548 = n12821 | ~n12822;
  assign n12824 = P3_EBX_REG_25_ & ~n12590;
  assign n12825 = ~n12326 & n12593;
  assign n12826 = P3_EBX_REG_23_ & P3_EBX_REG_24_;
  assign n12827 = n12808 & n12826;
  assign n12828 = P3_EBX_REG_25_ & ~n12827;
  assign n12829 = ~P3_EBX_REG_25_ & n12827;
  assign n12830 = ~n12828 & ~n12829;
  assign n12831 = n12591 & ~n12830;
  assign n12832 = ~n12824 & ~n12825;
  assign n2553 = n12831 | ~n12832;
  assign n12834 = P3_EBX_REG_26_ & ~n12590;
  assign n12835 = ~n12375 & n12593;
  assign n12836 = P3_EBX_REG_25_ & n12827;
  assign n12837 = ~P3_EBX_REG_26_ & n12836;
  assign n12838 = P3_EBX_REG_26_ & ~n12836;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = n12591 & ~n12839;
  assign n12841 = ~n12834 & ~n12835;
  assign n2558 = n12840 | ~n12841;
  assign n12843 = P3_EBX_REG_27_ & ~n12590;
  assign n12844 = ~n12423 & n12593;
  assign n12845 = P3_EBX_REG_25_ & P3_EBX_REG_26_;
  assign n12846 = n12827 & n12845;
  assign n12847 = P3_EBX_REG_27_ & ~n12846;
  assign n12848 = ~P3_EBX_REG_27_ & n12846;
  assign n12849 = ~n12847 & ~n12848;
  assign n12850 = n12591 & ~n12849;
  assign n12851 = ~n12843 & ~n12844;
  assign n2563 = n12850 | ~n12851;
  assign n12853 = P3_EBX_REG_28_ & ~n12590;
  assign n12854 = ~n12472 & n12593;
  assign n12855 = P3_EBX_REG_27_ & n12846;
  assign n12856 = ~P3_EBX_REG_28_ & n12855;
  assign n12857 = P3_EBX_REG_28_ & ~n12855;
  assign n12858 = ~n12856 & ~n12857;
  assign n12859 = n12591 & ~n12858;
  assign n12860 = ~n12853 & ~n12854;
  assign n2568 = n12859 | ~n12860;
  assign n12862 = P3_EBX_REG_29_ & ~n12590;
  assign n12863 = ~n12520 & n12593;
  assign n12864 = P3_EBX_REG_27_ & P3_EBX_REG_28_;
  assign n12865 = n12846 & n12864;
  assign n12866 = P3_EBX_REG_29_ & ~n12865;
  assign n12867 = ~P3_EBX_REG_29_ & n12865;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = n12591 & ~n12868;
  assign n12870 = ~n12862 & ~n12863;
  assign n2573 = n12869 | ~n12870;
  assign n12872 = P3_EBX_REG_30_ & ~n12590;
  assign n12873 = ~n12569 & n12593;
  assign n12874 = P3_EBX_REG_29_ & n12865;
  assign n12875 = ~P3_EBX_REG_30_ & n12874;
  assign n12876 = P3_EBX_REG_30_ & ~n12874;
  assign n12877 = ~n12875 & ~n12876;
  assign n12878 = n12591 & ~n12877;
  assign n12879 = ~n12872 & ~n12873;
  assign n2578 = n12878 | ~n12879;
  assign n12881 = P3_EBX_REG_31_ & ~n12590;
  assign n12882 = P3_EBX_REG_30_ & n12874;
  assign n12883 = ~P3_EBX_REG_31_ & n12882;
  assign n12884 = P3_EBX_REG_31_ & ~n12882;
  assign n12885 = ~n12883 & ~n12884;
  assign n12886 = n12591 & ~n12885;
  assign n2583 = n12881 | n12886;
  assign n12888 = ~n5724_1 & ~n5763;
  assign n12889 = ~n7327 & n12888;
  assign n12890 = n5591 & n5599_1;
  assign n12891 = n5713 & ~n12890;
  assign n12892 = n12889 & ~n12891;
  assign n12893 = P3_STATE2_REG_2_ & ~n12892;
  assign n12894 = n5441 & n12893;
  assign n12895 = ~n5074_1 & n12894;
  assign n12896 = ~P3_EBX_REG_31_ & n12895;
  assign n12897 = n5359_1 & n12893;
  assign n12898 = ~n5077 & n12897;
  assign n12899 = n5077 & n12897;
  assign n12900 = ~n5074_1 & n12899;
  assign n12901 = ~n12896 & ~n12898;
  assign n12902 = ~n12900 & n12901;
  assign n12903 = P3_EBX_REG_0_ & ~n12902;
  assign n12904 = n5074_1 & n12899;
  assign n12905 = P3_REIP_REG_0_ & n12904;
  assign n12906 = P3_EBX_REG_31_ & n12895;
  assign n12907 = P3_EBX_REG_0_ & n12906;
  assign n12908 = n5436 & n12893;
  assign n12909 = ~P3_INSTQUEUERD_ADDR_REG_0_ & n12908;
  assign n12910 = n5432 & n12893;
  assign n12911 = ~P3_INSTQUEUERD_ADDR_REG_0_ & n12910;
  assign n12912 = ~n12909 & ~n12911;
  assign n12913 = ~n12905 & ~n12907;
  assign n12914 = n12912 & n12913;
  assign n12915 = n5074_1 & n12894;
  assign n12916 = P3_REIP_REG_0_ & n12915;
  assign n12917 = P3_STATE2_REG_1_ & ~n12892;
  assign n12918 = n11029 & n12917;
  assign n12919 = P3_PHYADDRPOINTER_REG_0_ & n12918;
  assign n12920 = P3_REIP_REG_0_ & n12892;
  assign n12921 = P3_STATE2_REG_3_ & ~n12892;
  assign n12922 = P3_PHYADDRPOINTER_REG_0_ & n12921;
  assign n12923 = ~n12920 & ~n12922;
  assign n12924 = ~n11029 & n12917;
  assign n12925 = P3_PHYADDRPOINTER_REG_0_ & n12924;
  assign n12926 = n12923 & ~n12925;
  assign n12927 = ~n12903 & n12914;
  assign n12928 = ~n12916 & n12927;
  assign n12929 = ~n12919 & n12928;
  assign n2588 = ~n12926 | ~n12929;
  assign n12931 = P3_EBX_REG_1_ & ~n12902;
  assign n12932 = ~P3_REIP_REG_1_ & n12904;
  assign n12933 = ~n12600 & n12906;
  assign n12934 = ~n5083 & ~n5088_1;
  assign n12935 = n12908 & ~n12934;
  assign n12936 = n12910 & ~n12934;
  assign n12937 = ~n12935 & ~n12936;
  assign n12938 = ~n12932 & ~n12933;
  assign n12939 = n12937 & n12938;
  assign n12940 = ~P3_REIP_REG_1_ & n12915;
  assign n12941 = ~P3_PHYADDRPOINTER_REG_1_ & n12918;
  assign n12942 = P3_REIP_REG_1_ & n12892;
  assign n12943 = P3_PHYADDRPOINTER_REG_1_ & n12921;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = P3_PHYADDRPOINTER_REG_0_ & P3_PHYADDRPOINTER_REG_1_;
  assign n12946 = ~P3_PHYADDRPOINTER_REG_0_ & ~P3_PHYADDRPOINTER_REG_1_;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = n12924 & ~n12947;
  assign n12949 = n12944 & ~n12948;
  assign n12950 = ~n12931 & n12939;
  assign n12951 = ~n12940 & n12950;
  assign n12952 = ~n12941 & n12951;
  assign n2593 = ~n12949 | ~n12952;
  assign n12954 = P3_EBX_REG_2_ & ~n12902;
  assign n12955 = P3_REIP_REG_1_ & ~P3_REIP_REG_2_;
  assign n12956 = ~P3_REIP_REG_1_ & P3_REIP_REG_2_;
  assign n12957 = ~n12955 & ~n12956;
  assign n12958 = n12904 & ~n12957;
  assign n12959 = ~P3_EBX_REG_0_ & ~P3_EBX_REG_1_;
  assign n12960 = P3_EBX_REG_2_ & ~n12959;
  assign n12961 = ~P3_EBX_REG_2_ & n12959;
  assign n12962 = ~n12960 & ~n12961;
  assign n12963 = n12906 & n12962;
  assign n12964 = ~n5561 & n12908;
  assign n12965 = ~n5561 & n12910;
  assign n12966 = ~n12964 & ~n12965;
  assign n12967 = ~n12958 & ~n12963;
  assign n12968 = n12966 & n12967;
  assign n12969 = n12915 & ~n12957;
  assign n12970 = ~n10363 & n12918;
  assign n12971 = P3_REIP_REG_2_ & n12892;
  assign n12972 = P3_PHYADDRPOINTER_REG_2_ & n12921;
  assign n12973 = ~n12971 & ~n12972;
  assign n12974 = ~P3_PHYADDRPOINTER_REG_0_ & P3_PHYADDRPOINTER_REG_1_;
  assign n12975 = ~n10363 & ~n12974;
  assign n12976 = n10363 & n12974;
  assign n12977 = ~n12975 & ~n12976;
  assign n12978 = n12924 & n12977;
  assign n12979 = n12973 & ~n12978;
  assign n12980 = ~n12954 & n12968;
  assign n12981 = ~n12969 & n12980;
  assign n12982 = ~n12970 & n12981;
  assign n2598 = ~n12979 | ~n12982;
  assign n12984 = P3_EBX_REG_3_ & ~n12902;
  assign n12985 = P3_REIP_REG_1_ & P3_REIP_REG_2_;
  assign n12986 = ~P3_REIP_REG_3_ & n12985;
  assign n12987 = P3_REIP_REG_3_ & ~n12985;
  assign n12988 = ~n12986 & ~n12987;
  assign n12989 = n12904 & ~n12988;
  assign n12990 = ~P3_EBX_REG_3_ & n12961;
  assign n12991 = P3_EBX_REG_3_ & ~n12961;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = n12906 & n12992;
  assign n12994 = ~P3_INSTQUEUERD_ADDR_REG_3_ & n5609_1;
  assign n12995 = ~n5610 & ~n12994;
  assign n12996 = n12908 & ~n12995;
  assign n12997 = n12910 & ~n12995;
  assign n12998 = ~n12996 & ~n12997;
  assign n12999 = ~n12989 & ~n12993;
  assign n13000 = n12998 & n12999;
  assign n13001 = n12915 & ~n12988;
  assign n13002 = ~n10385 & n12918;
  assign n13003 = P3_REIP_REG_3_ & n12892;
  assign n13004 = P3_PHYADDRPOINTER_REG_3_ & n12921;
  assign n13005 = ~n13003 & ~n13004;
  assign n13006 = n10385 & n12976;
  assign n13007 = ~n10385 & ~n12976;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = n12924 & n13008;
  assign n13010 = n13005 & ~n13009;
  assign n13011 = ~n12984 & n13000;
  assign n13012 = ~n13001 & n13011;
  assign n13013 = ~n13002 & n13012;
  assign n2603 = ~n13010 | ~n13013;
  assign n13015 = P3_INSTQUEUERD_ADDR_REG_3_ & n5609_1;
  assign n13016 = ~P3_INSTQUEUERD_ADDR_REG_4_ & n13015;
  assign n13017 = P3_INSTQUEUERD_ADDR_REG_4_ & ~n13015;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = n12910 & ~n13018;
  assign n13020 = n12908 & ~n13018;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = P3_EBX_REG_4_ & ~n12902;
  assign n13023 = P3_EBX_REG_4_ & ~n12990;
  assign n13024 = ~P3_EBX_REG_3_ & ~P3_EBX_REG_4_;
  assign n13025 = n12961 & n13024;
  assign n13026 = ~n13023 & ~n13025;
  assign n13027 = n12906 & n13026;
  assign n13028 = n7326 & ~n12892;
  assign n13029 = P3_REIP_REG_3_ & n12985;
  assign n13030 = ~P3_REIP_REG_4_ & n13029;
  assign n13031 = P3_REIP_REG_4_ & ~n13029;
  assign n13032 = ~n13030 & ~n13031;
  assign n13033 = n12904 & ~n13032;
  assign n13034 = ~n13027 & ~n13028;
  assign n13035 = ~n13033 & n13034;
  assign n13036 = n12915 & ~n13032;
  assign n13037 = ~n10406 & n12918;
  assign n13038 = n13021 & ~n13022;
  assign n13039 = n13035 & n13038;
  assign n13040 = ~n13036 & n13039;
  assign n13041 = ~n13037 & n13040;
  assign n13042 = P3_REIP_REG_4_ & n12892;
  assign n13043 = P3_PHYADDRPOINTER_REG_4_ & n12921;
  assign n13044 = ~n13042 & ~n13043;
  assign n13045 = ~n10406 & ~n13006;
  assign n13046 = n10385 & n10406;
  assign n13047 = n12976 & n13046;
  assign n13048 = ~n13045 & ~n13047;
  assign n13049 = n12924 & n13048;
  assign n13050 = n13044 & ~n13049;
  assign n2608 = ~n13041 | ~n13050;
  assign n13052 = P3_INSTQUEUERD_ADDR_REG_4_ & n13015;
  assign n13053 = n12910 & n13052;
  assign n13054 = n12908 & n13052;
  assign n13055 = ~n13053 & ~n13054;
  assign n13056 = P3_EBX_REG_5_ & ~n12902;
  assign n13057 = ~P3_EBX_REG_5_ & n13025;
  assign n13058 = P3_EBX_REG_5_ & ~n13025;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = n12906 & n13059;
  assign n13061 = P3_REIP_REG_4_ & n13029;
  assign n13062 = ~P3_REIP_REG_5_ & n13061;
  assign n13063 = P3_REIP_REG_5_ & ~n13061;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = n12904 & ~n13064;
  assign n13066 = ~n13028 & ~n13060;
  assign n13067 = ~n13065 & n13066;
  assign n13068 = n12915 & ~n13064;
  assign n13069 = ~n10429 & n12918;
  assign n13070 = n13055 & ~n13056;
  assign n13071 = n13067 & n13070;
  assign n13072 = ~n13068 & n13071;
  assign n13073 = ~n13069 & n13072;
  assign n13074 = P3_REIP_REG_5_ & n12892;
  assign n13075 = P3_PHYADDRPOINTER_REG_5_ & n12921;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = n10429 & n13047;
  assign n13078 = ~n10429 & ~n13047;
  assign n13079 = ~n13077 & ~n13078;
  assign n13080 = n12924 & n13079;
  assign n13081 = n13076 & ~n13080;
  assign n2613 = ~n13073 | ~n13081;
  assign n13083 = P3_REIP_REG_5_ & n13061;
  assign n13084 = ~P3_REIP_REG_6_ & n13083;
  assign n13085 = P3_REIP_REG_6_ & ~n13083;
  assign n13086 = ~n13084 & ~n13085;
  assign n13087 = n12915 & ~n13086;
  assign n13088 = P3_EBX_REG_6_ & ~n12902;
  assign n13089 = P3_EBX_REG_6_ & ~n13057;
  assign n13090 = ~P3_EBX_REG_5_ & ~P3_EBX_REG_6_;
  assign n13091 = n13025 & n13090;
  assign n13092 = ~n13089 & ~n13091;
  assign n13093 = n12906 & n13092;
  assign n13094 = n12904 & ~n13086;
  assign n13095 = ~n13028 & ~n13093;
  assign n13096 = ~n13094 & n13095;
  assign n13097 = ~n10452 & ~n13077;
  assign n13098 = n10429 & n10452;
  assign n13099 = n13047 & n13098;
  assign n13100 = ~n13097 & ~n13099;
  assign n13101 = n12924 & n13100;
  assign n13102 = P3_REIP_REG_6_ & n12892;
  assign n13103 = P3_PHYADDRPOINTER_REG_6_ & n12921;
  assign n13104 = ~n13102 & ~n13103;
  assign n13105 = ~n10452 & n12918;
  assign n13106 = n13104 & ~n13105;
  assign n13107 = ~n13087 & ~n13088;
  assign n13108 = n13096 & n13107;
  assign n13109 = ~n13101 & n13108;
  assign n2618 = ~n13106 | ~n13109;
  assign n13111 = P3_REIP_REG_6_ & n13083;
  assign n13112 = ~P3_REIP_REG_7_ & n13111;
  assign n13113 = P3_REIP_REG_7_ & ~n13111;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = n12915 & ~n13114;
  assign n13116 = P3_EBX_REG_7_ & ~n12902;
  assign n13117 = ~P3_EBX_REG_7_ & n13091;
  assign n13118 = P3_EBX_REG_7_ & ~n13091;
  assign n13119 = ~n13117 & ~n13118;
  assign n13120 = n12906 & n13119;
  assign n13121 = n12904 & ~n13114;
  assign n13122 = ~n13028 & ~n13120;
  assign n13123 = ~n13121 & n13122;
  assign n13124 = n10475 & n13099;
  assign n13125 = ~n10475 & ~n13099;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = n12924 & n13126;
  assign n13128 = P3_REIP_REG_7_ & n12892;
  assign n13129 = P3_PHYADDRPOINTER_REG_7_ & n12921;
  assign n13130 = ~n13128 & ~n13129;
  assign n13131 = ~n10475 & n12918;
  assign n13132 = n13130 & ~n13131;
  assign n13133 = ~n13115 & ~n13116;
  assign n13134 = n13123 & n13133;
  assign n13135 = ~n13127 & n13134;
  assign n2623 = ~n13132 | ~n13135;
  assign n13137 = P3_REIP_REG_7_ & n13111;
  assign n13138 = ~P3_REIP_REG_8_ & n13137;
  assign n13139 = P3_REIP_REG_8_ & ~n13137;
  assign n13140 = ~n13138 & ~n13139;
  assign n13141 = n12915 & ~n13140;
  assign n13142 = P3_EBX_REG_8_ & ~n12902;
  assign n13143 = P3_EBX_REG_8_ & ~n13117;
  assign n13144 = ~P3_EBX_REG_7_ & ~P3_EBX_REG_8_;
  assign n13145 = n13091 & n13144;
  assign n13146 = ~n13143 & ~n13145;
  assign n13147 = n12906 & n13146;
  assign n13148 = n12904 & ~n13140;
  assign n13149 = ~n13028 & ~n13147;
  assign n13150 = ~n13148 & n13149;
  assign n13151 = ~n10498 & ~n13124;
  assign n13152 = n10475 & n10498;
  assign n13153 = n13099 & n13152;
  assign n13154 = ~n13151 & ~n13153;
  assign n13155 = n12924 & n13154;
  assign n13156 = P3_REIP_REG_8_ & n12892;
  assign n13157 = P3_PHYADDRPOINTER_REG_8_ & n12921;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = ~n10498 & n12918;
  assign n13160 = n13158 & ~n13159;
  assign n13161 = ~n13141 & ~n13142;
  assign n13162 = n13150 & n13161;
  assign n13163 = ~n13155 & n13162;
  assign n2628 = ~n13160 | ~n13163;
  assign n13165 = P3_REIP_REG_8_ & n13137;
  assign n13166 = ~P3_REIP_REG_9_ & n13165;
  assign n13167 = P3_REIP_REG_9_ & ~n13165;
  assign n13168 = ~n13166 & ~n13167;
  assign n13169 = n12915 & ~n13168;
  assign n13170 = P3_EBX_REG_9_ & ~n12902;
  assign n13171 = ~P3_EBX_REG_9_ & n13145;
  assign n13172 = P3_EBX_REG_9_ & ~n13145;
  assign n13173 = ~n13171 & ~n13172;
  assign n13174 = n12906 & n13173;
  assign n13175 = n12904 & ~n13168;
  assign n13176 = ~n13028 & ~n13174;
  assign n13177 = ~n13175 & n13176;
  assign n13178 = n10521 & n13153;
  assign n13179 = ~n10521 & ~n13153;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = n12924 & n13180;
  assign n13182 = P3_REIP_REG_9_ & n12892;
  assign n13183 = P3_PHYADDRPOINTER_REG_9_ & n12921;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = ~n10521 & n12918;
  assign n13186 = n13184 & ~n13185;
  assign n13187 = ~n13169 & ~n13170;
  assign n13188 = n13177 & n13187;
  assign n13189 = ~n13181 & n13188;
  assign n2633 = ~n13186 | ~n13189;
  assign n13191 = P3_REIP_REG_9_ & n13165;
  assign n13192 = ~P3_REIP_REG_10_ & n13191;
  assign n13193 = P3_REIP_REG_10_ & ~n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = n12915 & ~n13194;
  assign n13196 = P3_EBX_REG_10_ & ~n12902;
  assign n13197 = P3_EBX_REG_10_ & ~n13171;
  assign n13198 = ~P3_EBX_REG_9_ & ~P3_EBX_REG_10_;
  assign n13199 = n13145 & n13198;
  assign n13200 = ~n13197 & ~n13199;
  assign n13201 = n12906 & n13200;
  assign n13202 = n12904 & ~n13194;
  assign n13203 = ~n13028 & ~n13201;
  assign n13204 = ~n13202 & n13203;
  assign n13205 = ~n10544 & ~n13178;
  assign n13206 = n10521 & n10544;
  assign n13207 = n13153 & n13206;
  assign n13208 = ~n13205 & ~n13207;
  assign n13209 = n12924 & n13208;
  assign n13210 = P3_REIP_REG_10_ & n12892;
  assign n13211 = P3_PHYADDRPOINTER_REG_10_ & n12921;
  assign n13212 = ~n13210 & ~n13211;
  assign n13213 = ~n10544 & n12918;
  assign n13214 = n13212 & ~n13213;
  assign n13215 = ~n13195 & ~n13196;
  assign n13216 = n13204 & n13215;
  assign n13217 = ~n13209 & n13216;
  assign n2638 = ~n13214 | ~n13217;
  assign n13219 = P3_REIP_REG_10_ & n13191;
  assign n13220 = ~P3_REIP_REG_11_ & n13219;
  assign n13221 = P3_REIP_REG_11_ & ~n13219;
  assign n13222 = ~n13220 & ~n13221;
  assign n13223 = n12915 & ~n13222;
  assign n13224 = P3_EBX_REG_11_ & ~n12902;
  assign n13225 = ~P3_EBX_REG_11_ & n13199;
  assign n13226 = P3_EBX_REG_11_ & ~n13199;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = n12906 & n13227;
  assign n13229 = n12904 & ~n13222;
  assign n13230 = ~n13028 & ~n13228;
  assign n13231 = ~n13229 & n13230;
  assign n13232 = n10567 & n13207;
  assign n13233 = ~n10567 & ~n13207;
  assign n13234 = ~n13232 & ~n13233;
  assign n13235 = n12924 & n13234;
  assign n13236 = P3_REIP_REG_11_ & n12892;
  assign n13237 = P3_PHYADDRPOINTER_REG_11_ & n12921;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = ~n10567 & n12918;
  assign n13240 = n13238 & ~n13239;
  assign n13241 = ~n13223 & ~n13224;
  assign n13242 = n13231 & n13241;
  assign n13243 = ~n13235 & n13242;
  assign n2643 = ~n13240 | ~n13243;
  assign n13245 = P3_REIP_REG_11_ & n13219;
  assign n13246 = ~P3_REIP_REG_12_ & n13245;
  assign n13247 = P3_REIP_REG_12_ & ~n13245;
  assign n13248 = ~n13246 & ~n13247;
  assign n13249 = n12915 & ~n13248;
  assign n13250 = P3_EBX_REG_12_ & ~n12902;
  assign n13251 = P3_EBX_REG_12_ & ~n13225;
  assign n13252 = ~P3_EBX_REG_11_ & ~P3_EBX_REG_12_;
  assign n13253 = n13199 & n13252;
  assign n13254 = ~n13251 & ~n13253;
  assign n13255 = n12906 & n13254;
  assign n13256 = n12904 & ~n13248;
  assign n13257 = ~n13028 & ~n13255;
  assign n13258 = ~n13256 & n13257;
  assign n13259 = ~n10590 & ~n13232;
  assign n13260 = n10567 & n10590;
  assign n13261 = n13207 & n13260;
  assign n13262 = ~n13259 & ~n13261;
  assign n13263 = n12924 & n13262;
  assign n13264 = P3_REIP_REG_12_ & n12892;
  assign n13265 = P3_PHYADDRPOINTER_REG_12_ & n12921;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = ~n10590 & n12918;
  assign n13268 = n13266 & ~n13267;
  assign n13269 = ~n13249 & ~n13250;
  assign n13270 = n13258 & n13269;
  assign n13271 = ~n13263 & n13270;
  assign n2648 = ~n13268 | ~n13271;
  assign n13273 = P3_REIP_REG_12_ & n13245;
  assign n13274 = ~P3_REIP_REG_13_ & n13273;
  assign n13275 = P3_REIP_REG_13_ & ~n13273;
  assign n13276 = ~n13274 & ~n13275;
  assign n13277 = n12915 & ~n13276;
  assign n13278 = P3_EBX_REG_13_ & ~n12902;
  assign n13279 = ~P3_EBX_REG_13_ & n13253;
  assign n13280 = P3_EBX_REG_13_ & ~n13253;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = n12906 & n13281;
  assign n13283 = n12904 & ~n13276;
  assign n13284 = ~n13028 & ~n13282;
  assign n13285 = ~n13283 & n13284;
  assign n13286 = n10613 & n13261;
  assign n13287 = ~n10613 & ~n13261;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = n12924 & n13288;
  assign n13290 = P3_REIP_REG_13_ & n12892;
  assign n13291 = P3_PHYADDRPOINTER_REG_13_ & n12921;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = ~n10613 & n12918;
  assign n13294 = n13292 & ~n13293;
  assign n13295 = ~n13277 & ~n13278;
  assign n13296 = n13285 & n13295;
  assign n13297 = ~n13289 & n13296;
  assign n2653 = ~n13294 | ~n13297;
  assign n13299 = P3_REIP_REG_13_ & n13273;
  assign n13300 = ~P3_REIP_REG_14_ & n13299;
  assign n13301 = P3_REIP_REG_14_ & ~n13299;
  assign n13302 = ~n13300 & ~n13301;
  assign n13303 = n12915 & ~n13302;
  assign n13304 = P3_EBX_REG_14_ & ~n12902;
  assign n13305 = P3_EBX_REG_14_ & ~n13279;
  assign n13306 = ~P3_EBX_REG_13_ & ~P3_EBX_REG_14_;
  assign n13307 = n13253 & n13306;
  assign n13308 = ~n13305 & ~n13307;
  assign n13309 = n12906 & n13308;
  assign n13310 = n12904 & ~n13302;
  assign n13311 = ~n13028 & ~n13309;
  assign n13312 = ~n13310 & n13311;
  assign n13313 = ~n10636 & ~n13286;
  assign n13314 = n10613 & n10636;
  assign n13315 = n13261 & n13314;
  assign n13316 = ~n13313 & ~n13315;
  assign n13317 = n12924 & n13316;
  assign n13318 = P3_REIP_REG_14_ & n12892;
  assign n13319 = P3_PHYADDRPOINTER_REG_14_ & n12921;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n10636 & n12918;
  assign n13322 = n13320 & ~n13321;
  assign n13323 = ~n13303 & ~n13304;
  assign n13324 = n13312 & n13323;
  assign n13325 = ~n13317 & n13324;
  assign n2658 = ~n13322 | ~n13325;
  assign n13327 = P3_REIP_REG_14_ & n13299;
  assign n13328 = ~P3_REIP_REG_15_ & n13327;
  assign n13329 = P3_REIP_REG_15_ & ~n13327;
  assign n13330 = ~n13328 & ~n13329;
  assign n13331 = n12915 & ~n13330;
  assign n13332 = P3_EBX_REG_15_ & ~n12902;
  assign n13333 = ~P3_EBX_REG_15_ & n13307;
  assign n13334 = P3_EBX_REG_15_ & ~n13307;
  assign n13335 = ~n13333 & ~n13334;
  assign n13336 = n12906 & n13335;
  assign n13337 = n12904 & ~n13330;
  assign n13338 = ~n13028 & ~n13336;
  assign n13339 = ~n13337 & n13338;
  assign n13340 = n10659 & n13315;
  assign n13341 = ~n10659 & ~n13315;
  assign n13342 = ~n13340 & ~n13341;
  assign n13343 = n12924 & n13342;
  assign n13344 = P3_REIP_REG_15_ & n12892;
  assign n13345 = P3_PHYADDRPOINTER_REG_15_ & n12921;
  assign n13346 = ~n13344 & ~n13345;
  assign n13347 = ~n10659 & n12918;
  assign n13348 = n13346 & ~n13347;
  assign n13349 = ~n13331 & ~n13332;
  assign n13350 = n13339 & n13349;
  assign n13351 = ~n13343 & n13350;
  assign n2663 = ~n13348 | ~n13351;
  assign n13353 = P3_REIP_REG_15_ & n13327;
  assign n13354 = ~P3_REIP_REG_16_ & n13353;
  assign n13355 = P3_REIP_REG_16_ & ~n13353;
  assign n13356 = ~n13354 & ~n13355;
  assign n13357 = n12915 & ~n13356;
  assign n13358 = P3_EBX_REG_16_ & ~n12902;
  assign n13359 = P3_EBX_REG_16_ & ~n13333;
  assign n13360 = ~P3_EBX_REG_15_ & ~P3_EBX_REG_16_;
  assign n13361 = n13307 & n13360;
  assign n13362 = ~n13359 & ~n13361;
  assign n13363 = n12906 & n13362;
  assign n13364 = n12904 & ~n13356;
  assign n13365 = ~n13028 & ~n13363;
  assign n13366 = ~n13364 & n13365;
  assign n13367 = ~n10682 & ~n13340;
  assign n13368 = n10659 & n10682;
  assign n13369 = n13315 & n13368;
  assign n13370 = ~n13367 & ~n13369;
  assign n13371 = n12924 & n13370;
  assign n13372 = P3_REIP_REG_16_ & n12892;
  assign n13373 = P3_PHYADDRPOINTER_REG_16_ & n12921;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = ~n10682 & n12918;
  assign n13376 = n13374 & ~n13375;
  assign n13377 = ~n13357 & ~n13358;
  assign n13378 = n13366 & n13377;
  assign n13379 = ~n13371 & n13378;
  assign n2668 = ~n13376 | ~n13379;
  assign n13381 = P3_REIP_REG_16_ & n13353;
  assign n13382 = ~P3_REIP_REG_17_ & n13381;
  assign n13383 = P3_REIP_REG_17_ & ~n13381;
  assign n13384 = ~n13382 & ~n13383;
  assign n13385 = n12915 & ~n13384;
  assign n13386 = P3_EBX_REG_17_ & ~n12902;
  assign n13387 = ~P3_EBX_REG_17_ & n13361;
  assign n13388 = P3_EBX_REG_17_ & ~n13361;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = n12906 & n13389;
  assign n13391 = n12904 & ~n13384;
  assign n13392 = ~n13028 & ~n13390;
  assign n13393 = ~n13391 & n13392;
  assign n13394 = n10705 & n13369;
  assign n13395 = ~n10705 & ~n13369;
  assign n13396 = ~n13394 & ~n13395;
  assign n13397 = n12924 & n13396;
  assign n13398 = P3_REIP_REG_17_ & n12892;
  assign n13399 = P3_PHYADDRPOINTER_REG_17_ & n12921;
  assign n13400 = ~n13398 & ~n13399;
  assign n13401 = ~n10705 & n12918;
  assign n13402 = n13400 & ~n13401;
  assign n13403 = ~n13385 & ~n13386;
  assign n13404 = n13393 & n13403;
  assign n13405 = ~n13397 & n13404;
  assign n2673 = ~n13402 | ~n13405;
  assign n13407 = P3_REIP_REG_17_ & n13381;
  assign n13408 = ~P3_REIP_REG_18_ & n13407;
  assign n13409 = P3_REIP_REG_18_ & ~n13407;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = n12915 & ~n13410;
  assign n13412 = P3_EBX_REG_18_ & ~n12902;
  assign n13413 = P3_EBX_REG_18_ & ~n13387;
  assign n13414 = ~P3_EBX_REG_17_ & ~P3_EBX_REG_18_;
  assign n13415 = n13361 & n13414;
  assign n13416 = ~n13413 & ~n13415;
  assign n13417 = n12906 & n13416;
  assign n13418 = n12904 & ~n13410;
  assign n13419 = ~n13028 & ~n13417;
  assign n13420 = ~n13418 & n13419;
  assign n13421 = ~n10728 & ~n13394;
  assign n13422 = n10705 & n10728;
  assign n13423 = n13369 & n13422;
  assign n13424 = ~n13421 & ~n13423;
  assign n13425 = n12924 & n13424;
  assign n13426 = P3_REIP_REG_18_ & n12892;
  assign n13427 = P3_PHYADDRPOINTER_REG_18_ & n12921;
  assign n13428 = ~n13426 & ~n13427;
  assign n13429 = ~n10728 & n12918;
  assign n13430 = n13428 & ~n13429;
  assign n13431 = ~n13411 & ~n13412;
  assign n13432 = n13420 & n13431;
  assign n13433 = ~n13425 & n13432;
  assign n2678 = ~n13430 | ~n13433;
  assign n13435 = P3_REIP_REG_18_ & n13407;
  assign n13436 = ~P3_REIP_REG_19_ & n13435;
  assign n13437 = P3_REIP_REG_19_ & ~n13435;
  assign n13438 = ~n13436 & ~n13437;
  assign n13439 = n12915 & ~n13438;
  assign n13440 = P3_EBX_REG_19_ & ~n12902;
  assign n13441 = ~P3_EBX_REG_19_ & n13415;
  assign n13442 = P3_EBX_REG_19_ & ~n13415;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = n12906 & n13443;
  assign n13445 = n12904 & ~n13438;
  assign n13446 = ~n13028 & ~n13444;
  assign n13447 = ~n13445 & n13446;
  assign n13448 = n10751 & n13423;
  assign n13449 = ~n10751 & ~n13423;
  assign n13450 = ~n13448 & ~n13449;
  assign n13451 = n12924 & n13450;
  assign n13452 = P3_REIP_REG_19_ & n12892;
  assign n13453 = P3_PHYADDRPOINTER_REG_19_ & n12921;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = ~n10751 & n12918;
  assign n13456 = n13454 & ~n13455;
  assign n13457 = ~n13439 & ~n13440;
  assign n13458 = n13447 & n13457;
  assign n13459 = ~n13451 & n13458;
  assign n2683 = ~n13456 | ~n13459;
  assign n13461 = P3_REIP_REG_19_ & n13435;
  assign n13462 = ~P3_REIP_REG_20_ & n13461;
  assign n13463 = P3_REIP_REG_20_ & ~n13461;
  assign n13464 = ~n13462 & ~n13463;
  assign n13465 = n12915 & ~n13464;
  assign n13466 = P3_EBX_REG_20_ & ~n12902;
  assign n13467 = n12904 & ~n13464;
  assign n13468 = P3_EBX_REG_20_ & ~n13441;
  assign n13469 = ~P3_EBX_REG_19_ & ~P3_EBX_REG_20_;
  assign n13470 = n13415 & n13469;
  assign n13471 = ~n13468 & ~n13470;
  assign n13472 = n12906 & n13471;
  assign n13473 = ~n13467 & ~n13472;
  assign n13474 = ~n10774 & ~n13448;
  assign n13475 = n10751 & n10774;
  assign n13476 = n13423 & n13475;
  assign n13477 = ~n13474 & ~n13476;
  assign n13478 = n12924 & n13477;
  assign n13479 = P3_REIP_REG_20_ & n12892;
  assign n13480 = P3_PHYADDRPOINTER_REG_20_ & n12921;
  assign n13481 = ~n13479 & ~n13480;
  assign n13482 = ~n10774 & n12918;
  assign n13483 = n13481 & ~n13482;
  assign n13484 = ~n13465 & ~n13466;
  assign n13485 = n13473 & n13484;
  assign n13486 = ~n13478 & n13485;
  assign n2688 = ~n13483 | ~n13486;
  assign n13488 = P3_REIP_REG_20_ & n13461;
  assign n13489 = ~P3_REIP_REG_21_ & n13488;
  assign n13490 = P3_REIP_REG_21_ & ~n13488;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = n12915 & ~n13491;
  assign n13493 = P3_EBX_REG_21_ & ~n12902;
  assign n13494 = n12904 & ~n13491;
  assign n13495 = ~P3_EBX_REG_21_ & n13470;
  assign n13496 = P3_EBX_REG_21_ & ~n13470;
  assign n13497 = ~n13495 & ~n13496;
  assign n13498 = n12906 & n13497;
  assign n13499 = ~n13494 & ~n13498;
  assign n13500 = n10797 & n13476;
  assign n13501 = ~n10797 & ~n13476;
  assign n13502 = ~n13500 & ~n13501;
  assign n13503 = n12924 & n13502;
  assign n13504 = P3_REIP_REG_21_ & n12892;
  assign n13505 = P3_PHYADDRPOINTER_REG_21_ & n12921;
  assign n13506 = ~n13504 & ~n13505;
  assign n13507 = ~n10797 & n12918;
  assign n13508 = n13506 & ~n13507;
  assign n13509 = ~n13492 & ~n13493;
  assign n13510 = n13499 & n13509;
  assign n13511 = ~n13503 & n13510;
  assign n2693 = ~n13508 | ~n13511;
  assign n13513 = P3_REIP_REG_21_ & n13488;
  assign n13514 = ~P3_REIP_REG_22_ & n13513;
  assign n13515 = P3_REIP_REG_22_ & ~n13513;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = n12915 & ~n13516;
  assign n13518 = P3_EBX_REG_22_ & ~n12902;
  assign n13519 = n12904 & ~n13516;
  assign n13520 = P3_EBX_REG_22_ & ~n13495;
  assign n13521 = ~P3_EBX_REG_21_ & ~P3_EBX_REG_22_;
  assign n13522 = n13470 & n13521;
  assign n13523 = ~n13520 & ~n13522;
  assign n13524 = n12906 & n13523;
  assign n13525 = ~n13519 & ~n13524;
  assign n13526 = ~n10820 & ~n13500;
  assign n13527 = n10797 & n10820;
  assign n13528 = n13476 & n13527;
  assign n13529 = ~n13526 & ~n13528;
  assign n13530 = n12924 & n13529;
  assign n13531 = P3_REIP_REG_22_ & n12892;
  assign n13532 = P3_PHYADDRPOINTER_REG_22_ & n12921;
  assign n13533 = ~n13531 & ~n13532;
  assign n13534 = ~n10820 & n12918;
  assign n13535 = n13533 & ~n13534;
  assign n13536 = ~n13517 & ~n13518;
  assign n13537 = n13525 & n13536;
  assign n13538 = ~n13530 & n13537;
  assign n2698 = ~n13535 | ~n13538;
  assign n13540 = P3_REIP_REG_22_ & n13513;
  assign n13541 = ~P3_REIP_REG_23_ & n13540;
  assign n13542 = P3_REIP_REG_23_ & ~n13540;
  assign n13543 = ~n13541 & ~n13542;
  assign n13544 = n12915 & ~n13543;
  assign n13545 = P3_EBX_REG_23_ & ~n12902;
  assign n13546 = n12904 & ~n13543;
  assign n13547 = ~P3_EBX_REG_23_ & n13522;
  assign n13548 = P3_EBX_REG_23_ & ~n13522;
  assign n13549 = ~n13547 & ~n13548;
  assign n13550 = n12906 & n13549;
  assign n13551 = ~n13546 & ~n13550;
  assign n13552 = n10843 & n13528;
  assign n13553 = ~n10843 & ~n13528;
  assign n13554 = ~n13552 & ~n13553;
  assign n13555 = n12924 & n13554;
  assign n13556 = P3_REIP_REG_23_ & n12892;
  assign n13557 = P3_PHYADDRPOINTER_REG_23_ & n12921;
  assign n13558 = ~n13556 & ~n13557;
  assign n13559 = ~n10843 & n12918;
  assign n13560 = n13558 & ~n13559;
  assign n13561 = ~n13544 & ~n13545;
  assign n13562 = n13551 & n13561;
  assign n13563 = ~n13555 & n13562;
  assign n2703 = ~n13560 | ~n13563;
  assign n13565 = P3_REIP_REG_23_ & n13540;
  assign n13566 = ~P3_REIP_REG_24_ & n13565;
  assign n13567 = P3_REIP_REG_24_ & ~n13565;
  assign n13568 = ~n13566 & ~n13567;
  assign n13569 = n12915 & ~n13568;
  assign n13570 = P3_EBX_REG_24_ & ~n12902;
  assign n13571 = n12904 & ~n13568;
  assign n13572 = P3_EBX_REG_24_ & ~n13547;
  assign n13573 = ~P3_EBX_REG_23_ & ~P3_EBX_REG_24_;
  assign n13574 = n13522 & n13573;
  assign n13575 = ~n13572 & ~n13574;
  assign n13576 = n12906 & n13575;
  assign n13577 = ~n13571 & ~n13576;
  assign n13578 = ~n10867 & ~n13552;
  assign n13579 = n10843 & n10867;
  assign n13580 = n13528 & n13579;
  assign n13581 = ~n13578 & ~n13580;
  assign n13582 = n12924 & n13581;
  assign n13583 = P3_REIP_REG_24_ & n12892;
  assign n13584 = P3_PHYADDRPOINTER_REG_24_ & n12921;
  assign n13585 = ~n13583 & ~n13584;
  assign n13586 = ~n10867 & n12918;
  assign n13587 = n13585 & ~n13586;
  assign n13588 = ~n13569 & ~n13570;
  assign n13589 = n13577 & n13588;
  assign n13590 = ~n13582 & n13589;
  assign n2708 = ~n13587 | ~n13590;
  assign n13592 = P3_REIP_REG_24_ & n13565;
  assign n13593 = ~P3_REIP_REG_25_ & n13592;
  assign n13594 = P3_REIP_REG_25_ & ~n13592;
  assign n13595 = ~n13593 & ~n13594;
  assign n13596 = n12915 & ~n13595;
  assign n13597 = P3_EBX_REG_25_ & ~n12902;
  assign n13598 = n12904 & ~n13595;
  assign n13599 = ~P3_EBX_REG_25_ & n13574;
  assign n13600 = P3_EBX_REG_25_ & ~n13574;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = n12906 & n13601;
  assign n13603 = ~n13598 & ~n13602;
  assign n13604 = n10890 & n13580;
  assign n13605 = ~n10890 & ~n13580;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = n12924 & n13606;
  assign n13608 = P3_REIP_REG_25_ & n12892;
  assign n13609 = P3_PHYADDRPOINTER_REG_25_ & n12921;
  assign n13610 = ~n13608 & ~n13609;
  assign n13611 = ~n10890 & n12918;
  assign n13612 = n13610 & ~n13611;
  assign n13613 = ~n13596 & ~n13597;
  assign n13614 = n13603 & n13613;
  assign n13615 = ~n13607 & n13614;
  assign n2713 = ~n13612 | ~n13615;
  assign n13617 = P3_REIP_REG_25_ & n13592;
  assign n13618 = ~P3_REIP_REG_26_ & n13617;
  assign n13619 = P3_REIP_REG_26_ & ~n13617;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = n12915 & ~n13620;
  assign n13622 = P3_EBX_REG_26_ & ~n12902;
  assign n13623 = n12904 & ~n13620;
  assign n13624 = P3_EBX_REG_26_ & ~n13599;
  assign n13625 = ~P3_EBX_REG_25_ & ~P3_EBX_REG_26_;
  assign n13626 = n13574 & n13625;
  assign n13627 = ~n13624 & ~n13626;
  assign n13628 = n12906 & n13627;
  assign n13629 = ~n13623 & ~n13628;
  assign n13630 = ~n10913 & ~n13604;
  assign n13631 = n10890 & n10913;
  assign n13632 = n13580 & n13631;
  assign n13633 = ~n13630 & ~n13632;
  assign n13634 = n12924 & n13633;
  assign n13635 = P3_REIP_REG_26_ & n12892;
  assign n13636 = P3_PHYADDRPOINTER_REG_26_ & n12921;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = ~n10913 & n12918;
  assign n13639 = n13637 & ~n13638;
  assign n13640 = ~n13621 & ~n13622;
  assign n13641 = n13629 & n13640;
  assign n13642 = ~n13634 & n13641;
  assign n2718 = ~n13639 | ~n13642;
  assign n13644 = P3_REIP_REG_26_ & n13617;
  assign n13645 = ~P3_REIP_REG_27_ & n13644;
  assign n13646 = P3_REIP_REG_27_ & ~n13644;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = n12915 & ~n13647;
  assign n13649 = P3_EBX_REG_27_ & ~n12902;
  assign n13650 = n12904 & ~n13647;
  assign n13651 = ~P3_EBX_REG_27_ & n13626;
  assign n13652 = P3_EBX_REG_27_ & ~n13626;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = n12906 & n13653;
  assign n13655 = ~n13650 & ~n13654;
  assign n13656 = n10936 & n13632;
  assign n13657 = ~n10936 & ~n13632;
  assign n13658 = ~n13656 & ~n13657;
  assign n13659 = n12924 & n13658;
  assign n13660 = P3_REIP_REG_27_ & n12892;
  assign n13661 = P3_PHYADDRPOINTER_REG_27_ & n12921;
  assign n13662 = ~n13660 & ~n13661;
  assign n13663 = ~n10936 & n12918;
  assign n13664 = n13662 & ~n13663;
  assign n13665 = ~n13648 & ~n13649;
  assign n13666 = n13655 & n13665;
  assign n13667 = ~n13659 & n13666;
  assign n2723 = ~n13664 | ~n13667;
  assign n13669 = P3_REIP_REG_27_ & n13644;
  assign n13670 = ~P3_REIP_REG_28_ & n13669;
  assign n13671 = P3_REIP_REG_28_ & ~n13669;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = n12915 & ~n13672;
  assign n13674 = P3_EBX_REG_28_ & ~n12902;
  assign n13675 = n12904 & ~n13672;
  assign n13676 = P3_EBX_REG_28_ & ~n13651;
  assign n13677 = ~P3_EBX_REG_27_ & ~P3_EBX_REG_28_;
  assign n13678 = n13626 & n13677;
  assign n13679 = ~n13676 & ~n13678;
  assign n13680 = n12906 & n13679;
  assign n13681 = ~n13675 & ~n13680;
  assign n13682 = ~n10960 & ~n13656;
  assign n13683 = n10936 & n10960;
  assign n13684 = n13632 & n13683;
  assign n13685 = ~n13682 & ~n13684;
  assign n13686 = n12924 & n13685;
  assign n13687 = P3_REIP_REG_28_ & n12892;
  assign n13688 = P3_PHYADDRPOINTER_REG_28_ & n12921;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = ~n10960 & n12918;
  assign n13691 = n13689 & ~n13690;
  assign n13692 = ~n13673 & ~n13674;
  assign n13693 = n13681 & n13692;
  assign n13694 = ~n13686 & n13693;
  assign n2728 = ~n13691 | ~n13694;
  assign n13696 = P3_REIP_REG_28_ & n13669;
  assign n13697 = ~P3_REIP_REG_29_ & n13696;
  assign n13698 = P3_REIP_REG_29_ & ~n13696;
  assign n13699 = ~n13697 & ~n13698;
  assign n13700 = n12915 & ~n13699;
  assign n13701 = P3_EBX_REG_29_ & ~n12902;
  assign n13702 = n12904 & ~n13699;
  assign n13703 = P3_EBX_REG_29_ & ~n13678;
  assign n13704 = ~P3_EBX_REG_29_ & n13678;
  assign n13705 = ~n13703 & ~n13704;
  assign n13706 = n12906 & n13705;
  assign n13707 = ~n13702 & ~n13706;
  assign n13708 = ~n10983 & ~n13684;
  assign n13709 = n10983 & n13684;
  assign n13710 = ~n13708 & ~n13709;
  assign n13711 = n12924 & n13710;
  assign n13712 = P3_REIP_REG_29_ & n12892;
  assign n13713 = P3_PHYADDRPOINTER_REG_29_ & n12921;
  assign n13714 = ~n13712 & ~n13713;
  assign n13715 = ~n10983 & n12918;
  assign n13716 = n13714 & ~n13715;
  assign n13717 = ~n13700 & ~n13701;
  assign n13718 = n13707 & n13717;
  assign n13719 = ~n13711 & n13718;
  assign n2733 = ~n13716 | ~n13719;
  assign n13721 = P3_REIP_REG_29_ & n13696;
  assign n13722 = ~P3_REIP_REG_30_ & n13721;
  assign n13723 = P3_REIP_REG_30_ & ~n13721;
  assign n13724 = ~n13722 & ~n13723;
  assign n13725 = n12915 & ~n13724;
  assign n13726 = P3_EBX_REG_30_ & ~n12902;
  assign n13727 = n12904 & ~n13724;
  assign n13728 = ~P3_EBX_REG_30_ & n13704;
  assign n13729 = P3_EBX_REG_30_ & ~n13704;
  assign n13730 = ~n13728 & ~n13729;
  assign n13731 = n12906 & n13730;
  assign n13732 = ~n13727 & ~n13731;
  assign n13733 = n11006 & n13709;
  assign n13734 = ~n11006 & ~n13709;
  assign n13735 = ~n13733 & ~n13734;
  assign n13736 = n12924 & n13735;
  assign n13737 = P3_REIP_REG_30_ & n12892;
  assign n13738 = P3_PHYADDRPOINTER_REG_30_ & n12921;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = ~n11006 & n12918;
  assign n13741 = n13739 & ~n13740;
  assign n13742 = ~n13725 & ~n13726;
  assign n13743 = n13732 & n13742;
  assign n13744 = ~n13736 & n13743;
  assign n2738 = ~n13741 | ~n13744;
  assign n13746 = ~n11029 & n13733;
  assign n13747 = n11029 & ~n13733;
  assign n13748 = ~n13746 & ~n13747;
  assign n13749 = ~n11029 & n12918;
  assign n13750 = n13748 & ~n13749;
  assign n13751 = P3_EBX_REG_31_ & ~n12902;
  assign n13752 = P3_EBX_REG_31_ & n13728;
  assign n13753 = ~P3_EBX_REG_31_ & ~n13728;
  assign n13754 = ~n13752 & ~n13753;
  assign n13755 = n12906 & ~n13754;
  assign n13756 = P3_REIP_REG_30_ & n13721;
  assign n13757 = ~P3_REIP_REG_31_ & n13756;
  assign n13758 = P3_REIP_REG_31_ & ~n13756;
  assign n13759 = ~n13757 & ~n13758;
  assign n13760 = n12904 & ~n13759;
  assign n13761 = P3_PHYADDRPOINTER_REG_31_ & n12921;
  assign n13762 = P3_REIP_REG_31_ & n12892;
  assign n13763 = ~n13761 & ~n13762;
  assign n13764 = n12915 & ~n13759;
  assign n13765 = n13763 & ~n13764;
  assign n13766 = ~n13751 & ~n13755;
  assign n13767 = ~n13760 & n13766;
  assign n13768 = n13765 & n13767;
  assign n13769 = n13750 & n13768;
  assign n13770 = ~n12924 & ~n13749;
  assign n13771 = n13768 & n13770;
  assign n2743 = ~n13769 & ~n13771;
  assign n13773 = ~P3_DATAWIDTH_REG_1_ & ~P3_REIP_REG_1_;
  assign n13774 = ~P3_DATAWIDTH_REG_30_ & ~P3_DATAWIDTH_REG_31_;
  assign n13775 = P3_DATAWIDTH_REG_0_ & P3_DATAWIDTH_REG_1_;
  assign n13776 = ~P3_DATAWIDTH_REG_28_ & ~P3_DATAWIDTH_REG_29_;
  assign n13777 = ~P3_DATAWIDTH_REG_26_ & ~P3_DATAWIDTH_REG_27_;
  assign n13778 = n13774 & ~n13775;
  assign n13779 = n13776 & n13778;
  assign n13780 = n13777 & n13779;
  assign n13781 = ~P3_DATAWIDTH_REG_22_ & ~P3_DATAWIDTH_REG_23_;
  assign n13782 = ~P3_DATAWIDTH_REG_24_ & n13781;
  assign n13783 = ~P3_DATAWIDTH_REG_25_ & n13782;
  assign n13784 = ~P3_DATAWIDTH_REG_18_ & ~P3_DATAWIDTH_REG_19_;
  assign n13785 = ~P3_DATAWIDTH_REG_20_ & n13784;
  assign n13786 = ~P3_DATAWIDTH_REG_21_ & n13785;
  assign n13787 = n13783 & n13786;
  assign n13788 = ~P3_DATAWIDTH_REG_14_ & ~P3_DATAWIDTH_REG_15_;
  assign n13789 = ~P3_DATAWIDTH_REG_16_ & n13788;
  assign n13790 = ~P3_DATAWIDTH_REG_17_ & n13789;
  assign n13791 = ~P3_DATAWIDTH_REG_10_ & ~P3_DATAWIDTH_REG_11_;
  assign n13792 = ~P3_DATAWIDTH_REG_12_ & n13791;
  assign n13793 = ~P3_DATAWIDTH_REG_13_ & n13792;
  assign n13794 = n13790 & n13793;
  assign n13795 = ~P3_DATAWIDTH_REG_6_ & ~P3_DATAWIDTH_REG_7_;
  assign n13796 = ~P3_DATAWIDTH_REG_8_ & n13795;
  assign n13797 = ~P3_DATAWIDTH_REG_9_ & n13796;
  assign n13798 = ~P3_DATAWIDTH_REG_2_ & ~P3_DATAWIDTH_REG_3_;
  assign n13799 = ~P3_DATAWIDTH_REG_4_ & n13798;
  assign n13800 = ~P3_DATAWIDTH_REG_5_ & n13799;
  assign n13801 = n13797 & n13800;
  assign n13802 = n13780 & n13787;
  assign n13803 = n13794 & n13802;
  assign n13804 = n13801 & n13803;
  assign n13805 = n13773 & n13804;
  assign n13806 = P3_BYTEENABLE_REG_3_ & ~n13804;
  assign n13807 = ~P3_DATAWIDTH_REG_0_ & ~P3_REIP_REG_0_;
  assign n13808 = ~P3_DATAWIDTH_REG_1_ & n13807;
  assign n13809 = n13804 & n13808;
  assign n13810 = ~n13805 & ~n13806;
  assign n2748 = n13809 | ~n13810;
  assign n13812 = P3_REIP_REG_0_ & P3_REIP_REG_1_;
  assign n13813 = P3_DATAWIDTH_REG_0_ & ~P3_REIP_REG_0_;
  assign n13814 = ~P3_DATAWIDTH_REG_0_ & ~P3_DATAWIDTH_REG_1_;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816 = ~P3_REIP_REG_1_ & ~n13815;
  assign n13817 = ~n13812 & ~n13816;
  assign n13818 = n13804 & ~n13817;
  assign n13819 = P3_BYTEENABLE_REG_2_ & ~n13804;
  assign n2753 = n13818 | n13819;
  assign n13821 = P3_REIP_REG_1_ & n13804;
  assign n13822 = P3_BYTEENABLE_REG_1_ & ~n13804;
  assign n13823 = ~n13821 & ~n13822;
  assign n2758 = n13809 | ~n13823;
  assign n13825 = ~P3_REIP_REG_0_ & ~P3_REIP_REG_1_;
  assign n13826 = n13804 & ~n13825;
  assign n13827 = P3_BYTEENABLE_REG_0_ & ~n13804;
  assign n2763 = n13826 | n13827;
  assign n13829 = P3_W_R_N_REG & ~n4817;
  assign n13830 = ~P3_READREQUEST_REG & n4817;
  assign n2768 = n13829 | n13830;
  assign n13832 = n5481 & n5713;
  assign n13833 = ~n5429_1 & n5713;
  assign n13834 = P3_FLUSH_REG & ~n13833;
  assign n2772 = n13832 | n13834;
  assign n13836 = P3_MORE_REG & ~n13833;
  assign n13837 = ~n5475 & n13833;
  assign n2777 = n13836 | n13837;
  assign n13839 = BS16 & ~n5034_1;
  assign n13840 = P3_STATEBS16_REG & n5034_1;
  assign n13841 = ~P3_STATE_REG_0_ & n4989_1;
  assign n13842 = ~n13839 & ~n13840;
  assign n2782 = n13841 | ~n13842;
  assign n13844 = ~n5359_1 & ~n5432;
  assign n13845 = ~n5077 & ~n13844;
  assign n13846 = ~P3_STATEBS16_REG & n5359_1;
  assign n13847 = ~n4986 & ~n13846;
  assign n13848 = P3_STATE2_REG_2_ & ~n13845;
  assign n13849 = n13847 & n13848;
  assign n13850 = P3_STATE2_REG_0_ & ~n13849;
  assign n13851 = ~n5729_1 & ~n13850;
  assign n13852 = ~n4986 & n5071;
  assign n13853 = ~n5719_1 & ~n13852;
  assign n13854 = ~P3_STATE2_REG_0_ & ~n13853;
  assign n13855 = ~n5791 & ~n13854;
  assign n13856 = ~n12891 & n13855;
  assign n13857 = ~n13851 & ~n13856;
  assign n13858 = P3_REQUESTPENDING_REG & n13856;
  assign n2787 = n13857 | n13858;
  assign n13860 = P3_D_C_N_REG & ~n4817;
  assign n13861 = ~P3_CODEFETCH_REG & n4817;
  assign n13862 = ~n13860 & ~n13861;
  assign n2792 = n13841 | ~n13862;
  assign n13864 = P3_MEMORYFETCH_REG & n4817;
  assign n13865 = P3_M_IO_N_REG & ~n4817;
  assign n2796 = n13864 | n13865;
  assign n13867 = P3_STATE2_REG_0_ & n7326;
  assign n13868 = n5428 & n5713;
  assign n13869 = P3_CODEFETCH_REG & ~n13868;
  assign n2800 = n13867 | n13869;
  assign n13871 = P3_STATE_REG_0_ & P3_ADS_N_REG;
  assign n2805 = ~n5034_1 | n13871;
  assign n13873 = P3_STATE2_REG_2_ & ~n5441;
  assign n13874 = ~n5436 & n13873;
  assign n13875 = ~n7326 & ~n12891;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = P3_READREQUEST_REG & n13875;
  assign n2809 = n13876 | n13877;
  assign n13879 = P3_STATE2_REG_2_ & n5358;
  assign n13880 = ~n13875 & ~n13879;
  assign n13881 = P3_MEMORYFETCH_REG & n13875;
  assign n2814 = n13880 | n13881;
  assign n13883 = P2_STATE_REG_1_ & ~P2_STATE_REG_0_;
  assign n13884 = P2_BYTEENABLE_REG_3_ & n13883;
  assign n13885 = P2_BE_N_REG_3_ & ~n13883;
  assign n2819 = n13884 | n13885;
  assign n13887 = P2_BYTEENABLE_REG_2_ & n13883;
  assign n13888 = P2_BE_N_REG_2_ & ~n13883;
  assign n2824 = n13887 | n13888;
  assign n13890 = P2_BYTEENABLE_REG_1_ & n13883;
  assign n13891 = P2_BE_N_REG_1_ & ~n13883;
  assign n2829 = n13890 | n13891;
  assign n13893 = P2_BYTEENABLE_REG_0_ & n13883;
  assign n13894 = P2_BE_N_REG_0_ & ~n13883;
  assign n2834 = n13893 | n13894;
  assign n13896 = P2_STATE_REG_2_ & n13883;
  assign n13897 = P2_REIP_REG_30_ & n13896;
  assign n13898 = ~P2_STATE_REG_2_ & n13883;
  assign n13899 = P2_REIP_REG_31_ & n13898;
  assign n13900 = P2_ADDRESS_REG_29_ & ~n13883;
  assign n13901 = ~n13897 & ~n13899;
  assign n2839 = n13900 | ~n13901;
  assign n13903 = P2_REIP_REG_29_ & n13896;
  assign n13904 = P2_REIP_REG_30_ & n13898;
  assign n13905 = P2_ADDRESS_REG_28_ & ~n13883;
  assign n13906 = ~n13903 & ~n13904;
  assign n2844 = n13905 | ~n13906;
  assign n13908 = P2_REIP_REG_28_ & n13896;
  assign n13909 = P2_REIP_REG_29_ & n13898;
  assign n13910 = P2_ADDRESS_REG_27_ & ~n13883;
  assign n13911 = ~n13908 & ~n13909;
  assign n2849 = n13910 | ~n13911;
  assign n13913 = P2_REIP_REG_27_ & n13896;
  assign n13914 = P2_REIP_REG_28_ & n13898;
  assign n13915 = P2_ADDRESS_REG_26_ & ~n13883;
  assign n13916 = ~n13913 & ~n13914;
  assign n2854 = n13915 | ~n13916;
  assign n13918 = P2_REIP_REG_26_ & n13896;
  assign n13919 = P2_REIP_REG_27_ & n13898;
  assign n13920 = P2_ADDRESS_REG_25_ & ~n13883;
  assign n13921 = ~n13918 & ~n13919;
  assign n2859 = n13920 | ~n13921;
  assign n13923 = P2_REIP_REG_25_ & n13896;
  assign n13924 = P2_REIP_REG_26_ & n13898;
  assign n13925 = P2_ADDRESS_REG_24_ & ~n13883;
  assign n13926 = ~n13923 & ~n13924;
  assign n2864 = n13925 | ~n13926;
  assign n13928 = P2_REIP_REG_24_ & n13896;
  assign n13929 = P2_REIP_REG_25_ & n13898;
  assign n13930 = P2_ADDRESS_REG_23_ & ~n13883;
  assign n13931 = ~n13928 & ~n13929;
  assign n2869 = n13930 | ~n13931;
  assign n13933 = P2_REIP_REG_23_ & n13896;
  assign n13934 = P2_REIP_REG_24_ & n13898;
  assign n13935 = P2_ADDRESS_REG_22_ & ~n13883;
  assign n13936 = ~n13933 & ~n13934;
  assign n2874 = n13935 | ~n13936;
  assign n13938 = P2_REIP_REG_22_ & n13896;
  assign n13939 = P2_REIP_REG_23_ & n13898;
  assign n13940 = P2_ADDRESS_REG_21_ & ~n13883;
  assign n13941 = ~n13938 & ~n13939;
  assign n2879 = n13940 | ~n13941;
  assign n13943 = P2_REIP_REG_21_ & n13896;
  assign n13944 = P2_REIP_REG_22_ & n13898;
  assign n13945 = P2_ADDRESS_REG_20_ & ~n13883;
  assign n13946 = ~n13943 & ~n13944;
  assign n2884 = n13945 | ~n13946;
  assign n13948 = P2_REIP_REG_20_ & n13896;
  assign n13949 = P2_REIP_REG_21_ & n13898;
  assign n13950 = P2_ADDRESS_REG_19_ & ~n13883;
  assign n13951 = ~n13948 & ~n13949;
  assign n2889 = n13950 | ~n13951;
  assign n13953 = P2_REIP_REG_19_ & n13896;
  assign n13954 = P2_REIP_REG_20_ & n13898;
  assign n13955 = P2_ADDRESS_REG_18_ & ~n13883;
  assign n13956 = ~n13953 & ~n13954;
  assign n2894 = n13955 | ~n13956;
  assign n13958 = P2_REIP_REG_18_ & n13896;
  assign n13959 = P2_REIP_REG_19_ & n13898;
  assign n13960 = P2_ADDRESS_REG_17_ & ~n13883;
  assign n13961 = ~n13958 & ~n13959;
  assign n2899 = n13960 | ~n13961;
  assign n13963 = P2_REIP_REG_17_ & n13896;
  assign n13964 = P2_REIP_REG_18_ & n13898;
  assign n13965 = P2_ADDRESS_REG_16_ & ~n13883;
  assign n13966 = ~n13963 & ~n13964;
  assign n2904 = n13965 | ~n13966;
  assign n13968 = P2_REIP_REG_16_ & n13896;
  assign n13969 = P2_REIP_REG_17_ & n13898;
  assign n13970 = P2_ADDRESS_REG_15_ & ~n13883;
  assign n13971 = ~n13968 & ~n13969;
  assign n2909 = n13970 | ~n13971;
  assign n13973 = P2_REIP_REG_15_ & n13896;
  assign n13974 = P2_REIP_REG_16_ & n13898;
  assign n13975 = P2_ADDRESS_REG_14_ & ~n13883;
  assign n13976 = ~n13973 & ~n13974;
  assign n2914 = n13975 | ~n13976;
  assign n13978 = P2_REIP_REG_14_ & n13896;
  assign n13979 = P2_REIP_REG_15_ & n13898;
  assign n13980 = P2_ADDRESS_REG_13_ & ~n13883;
  assign n13981 = ~n13978 & ~n13979;
  assign n2919 = n13980 | ~n13981;
  assign n13983 = P2_REIP_REG_13_ & n13896;
  assign n13984 = P2_REIP_REG_14_ & n13898;
  assign n13985 = P2_ADDRESS_REG_12_ & ~n13883;
  assign n13986 = ~n13983 & ~n13984;
  assign n2924 = n13985 | ~n13986;
  assign n13988 = P2_REIP_REG_12_ & n13896;
  assign n13989 = P2_REIP_REG_13_ & n13898;
  assign n13990 = P2_ADDRESS_REG_11_ & ~n13883;
  assign n13991 = ~n13988 & ~n13989;
  assign n2929 = n13990 | ~n13991;
  assign n13993 = P2_REIP_REG_11_ & n13896;
  assign n13994 = P2_REIP_REG_12_ & n13898;
  assign n13995 = P2_ADDRESS_REG_10_ & ~n13883;
  assign n13996 = ~n13993 & ~n13994;
  assign n2934 = n13995 | ~n13996;
  assign n13998 = P2_REIP_REG_10_ & n13896;
  assign n13999 = P2_REIP_REG_11_ & n13898;
  assign n14000 = P2_ADDRESS_REG_9_ & ~n13883;
  assign n14001 = ~n13998 & ~n13999;
  assign n2939 = n14000 | ~n14001;
  assign n14003 = P2_REIP_REG_9_ & n13896;
  assign n14004 = P2_REIP_REG_10_ & n13898;
  assign n14005 = P2_ADDRESS_REG_8_ & ~n13883;
  assign n14006 = ~n14003 & ~n14004;
  assign n2944 = n14005 | ~n14006;
  assign n14008 = P2_REIP_REG_8_ & n13896;
  assign n14009 = P2_REIP_REG_9_ & n13898;
  assign n14010 = P2_ADDRESS_REG_7_ & ~n13883;
  assign n14011 = ~n14008 & ~n14009;
  assign n2949 = n14010 | ~n14011;
  assign n14013 = P2_REIP_REG_7_ & n13896;
  assign n14014 = P2_REIP_REG_8_ & n13898;
  assign n14015 = P2_ADDRESS_REG_6_ & ~n13883;
  assign n14016 = ~n14013 & ~n14014;
  assign n2954 = n14015 | ~n14016;
  assign n14018 = P2_REIP_REG_6_ & n13896;
  assign n14019 = P2_REIP_REG_7_ & n13898;
  assign n14020 = P2_ADDRESS_REG_5_ & ~n13883;
  assign n14021 = ~n14018 & ~n14019;
  assign n2959 = n14020 | ~n14021;
  assign n14023 = P2_REIP_REG_5_ & n13896;
  assign n14024 = P2_REIP_REG_6_ & n13898;
  assign n14025 = P2_ADDRESS_REG_4_ & ~n13883;
  assign n14026 = ~n14023 & ~n14024;
  assign n2964 = n14025 | ~n14026;
  assign n14028 = P2_REIP_REG_4_ & n13896;
  assign n14029 = P2_REIP_REG_5_ & n13898;
  assign n14030 = P2_ADDRESS_REG_3_ & ~n13883;
  assign n14031 = ~n14028 & ~n14029;
  assign n2969 = n14030 | ~n14031;
  assign n14033 = P2_REIP_REG_3_ & n13896;
  assign n14034 = P2_REIP_REG_4_ & n13898;
  assign n14035 = P2_ADDRESS_REG_2_ & ~n13883;
  assign n14036 = ~n14033 & ~n14034;
  assign n2974 = n14035 | ~n14036;
  assign n14038 = P2_REIP_REG_2_ & n13896;
  assign n14039 = P2_REIP_REG_3_ & n13898;
  assign n14040 = P2_ADDRESS_REG_1_ & ~n13883;
  assign n14041 = ~n14038 & ~n14039;
  assign n2979 = n14040 | ~n14041;
  assign n14043 = P2_REIP_REG_1_ & n13896;
  assign n14044 = P2_REIP_REG_2_ & n13898;
  assign n14045 = P2_ADDRESS_REG_0_ & ~n13883;
  assign n14046 = ~n14043 & ~n14044;
  assign n2984 = n14045 | ~n14046;
  assign n14048 = ~P2_STATE_REG_2_ & P2_STATE_REG_1_;
  assign n14049 = NA & n14048;
  assign n14050 = ~HOLD & ~P2_REQUESTPENDING_REG;
  assign n14051 = READY12_REG & READY21_REG;
  assign n14052 = P2_STATE_REG_1_ & ~n14050;
  assign n14053 = n14051 & n14052;
  assign n14054 = ~P2_STATE_REG_2_ & ~P2_STATE_REG_1_;
  assign n14055 = HOLD & ~P2_REQUESTPENDING_REG;
  assign n14056 = n14054 & n14055;
  assign n14057 = ~n14053 & ~n14056;
  assign n14058 = P2_STATE_REG_0_ & ~n14049;
  assign n14059 = ~n14057 & n14058;
  assign n14060 = ~n13896 & ~n14059;
  assign n14061 = ~NA & ~P2_STATE_REG_0_;
  assign n14062 = ~HOLD & P2_REQUESTPENDING_REG;
  assign n14063 = ~n14050 & ~n14062;
  assign n14064 = P2_STATE_REG_0_ & n14063;
  assign n14065 = ~n14061 & ~n14064;
  assign n14066 = n14050 & ~n14051;
  assign n14067 = ~n14051 & n14062;
  assign n14068 = P2_STATE_REG_1_ & ~n14066;
  assign n14069 = ~n14067 & n14068;
  assign n14070 = n14065 & ~n14069;
  assign n14071 = P2_STATE_REG_2_ & ~n14070;
  assign n2989 = ~n14060 | n14071;
  assign n14073 = P2_STATE_REG_0_ & n14062;
  assign n14074 = P2_STATE_REG_2_ & ~P2_STATE_REG_0_;
  assign n14075 = ~P2_STATE_REG_2_ & P2_REQUESTPENDING_REG;
  assign n14076 = P2_STATE_REG_0_ & n14075;
  assign n14077 = ~n14073 & ~n14074;
  assign n14078 = ~n14076 & n14077;
  assign n14079 = ~P2_STATE_REG_1_ & ~n14078;
  assign n14080 = HOLD & ~n14051;
  assign n14081 = P2_STATE_REG_0_ & ~n14080;
  assign n14082 = P2_STATE_REG_2_ & ~n14081;
  assign n14083 = ~n14066 & ~n14082;
  assign n14084 = P2_STATE_REG_1_ & n14083;
  assign n14085 = n13883 & n14051;
  assign n14086 = ~n13898 & ~n14085;
  assign n14087 = ~n14079 & ~n14084;
  assign n2994 = ~n14086 | ~n14087;
  assign n14089 = P2_STATE_REG_0_ & P2_REQUESTPENDING_REG;
  assign n14090 = P2_STATE_REG_1_ & ~n14067;
  assign n14091 = n14089 & ~n14090;
  assign n14092 = ~P2_STATE_REG_2_ & ~n14091;
  assign n14093 = P2_STATE_REG_0_ & ~n14062;
  assign n14094 = P2_STATE_REG_2_ & n14093;
  assign n14095 = NA & ~P2_STATE_REG_0_;
  assign n14096 = P2_STATE_REG_2_ & ~n14062;
  assign n14097 = ~n14095 & ~n14096;
  assign n14098 = ~P2_STATE_REG_1_ & ~n14097;
  assign n14099 = ~n14092 & ~n14094;
  assign n2999 = n14098 | ~n14099;
  assign n14101 = ~BS16 & ~n14054;
  assign n14102 = P2_STATE_REG_0_ & n14048;
  assign n14103 = ~P2_STATE_REG_1_ & ~P2_STATE_REG_0_;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = n14101 & ~n14104;
  assign n14106 = P2_DATAWIDTH_REG_0_ & n14104;
  assign n3004 = n14105 | n14106;
  assign n14108 = P2_DATAWIDTH_REG_1_ & n14104;
  assign n14109 = ~n14101 & ~n14104;
  assign n3009 = n14108 | n14109;
  assign n3014 = P2_DATAWIDTH_REG_2_ & n14104;
  assign n3019 = P2_DATAWIDTH_REG_3_ & n14104;
  assign n3024 = P2_DATAWIDTH_REG_4_ & n14104;
  assign n3029 = P2_DATAWIDTH_REG_5_ & n14104;
  assign n3034 = P2_DATAWIDTH_REG_6_ & n14104;
  assign n3039 = P2_DATAWIDTH_REG_7_ & n14104;
  assign n3044 = P2_DATAWIDTH_REG_8_ & n14104;
  assign n3049 = P2_DATAWIDTH_REG_9_ & n14104;
  assign n3054 = P2_DATAWIDTH_REG_10_ & n14104;
  assign n3059 = P2_DATAWIDTH_REG_11_ & n14104;
  assign n3064 = P2_DATAWIDTH_REG_12_ & n14104;
  assign n3069 = P2_DATAWIDTH_REG_13_ & n14104;
  assign n3074 = P2_DATAWIDTH_REG_14_ & n14104;
  assign n3079 = P2_DATAWIDTH_REG_15_ & n14104;
  assign n3084 = P2_DATAWIDTH_REG_16_ & n14104;
  assign n3089 = P2_DATAWIDTH_REG_17_ & n14104;
  assign n3094 = P2_DATAWIDTH_REG_18_ & n14104;
  assign n3099 = P2_DATAWIDTH_REG_19_ & n14104;
  assign n3104 = P2_DATAWIDTH_REG_20_ & n14104;
  assign n3109 = P2_DATAWIDTH_REG_21_ & n14104;
  assign n3114 = P2_DATAWIDTH_REG_22_ & n14104;
  assign n3119 = P2_DATAWIDTH_REG_23_ & n14104;
  assign n3124 = P2_DATAWIDTH_REG_24_ & n14104;
  assign n3129 = P2_DATAWIDTH_REG_25_ & n14104;
  assign n3134 = P2_DATAWIDTH_REG_26_ & n14104;
  assign n3139 = P2_DATAWIDTH_REG_27_ & n14104;
  assign n3144 = P2_DATAWIDTH_REG_28_ & n14104;
  assign n3149 = P2_DATAWIDTH_REG_29_ & n14104;
  assign n3154 = P2_DATAWIDTH_REG_30_ & n14104;
  assign n3159 = P2_DATAWIDTH_REG_31_ & n14104;
  assign n14141 = P2_STATE2_REG_2_ & P2_STATE2_REG_1_;
  assign n14142 = P2_STATE_REG_2_ & ~P2_STATE_REG_1_;
  assign n14143 = ~n14048 & ~n14142;
  assign n14144 = ~P2_STATE_REG_0_ & ~n14143;
  assign n14145 = ~n14051 & n14144;
  assign n14146 = ~P2_INSTQUEUE_REG_2__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14147 = ~P2_INSTQUEUE_REG_10__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14148 = ~P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14149 = P2_INSTQUEUERD_ADDR_REG_1_ & n14148;
  assign n14150 = ~n14146 & ~n14147;
  assign n14151 = n14149 & n14150;
  assign n14152 = ~P2_INSTQUEUE_REG_6__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14153 = ~P2_INSTQUEUE_REG_14__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14154 = P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14155 = P2_INSTQUEUERD_ADDR_REG_2_ & n14154;
  assign n14156 = ~n14152 & ~n14153;
  assign n14157 = n14155 & n14156;
  assign n14158 = ~P2_INSTQUEUE_REG_5__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14159 = ~P2_INSTQUEUE_REG_13__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14160 = ~P2_INSTQUEUERD_ADDR_REG_1_ & P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14161 = P2_INSTQUEUERD_ADDR_REG_2_ & n14160;
  assign n14162 = ~n14158 & ~n14159;
  assign n14163 = n14161 & n14162;
  assign n14164 = ~P2_INSTQUEUE_REG_7__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14165 = ~P2_INSTQUEUE_REG_15__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14166 = P2_INSTQUEUERD_ADDR_REG_1_ & P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14167 = P2_INSTQUEUERD_ADDR_REG_2_ & n14166;
  assign n14168 = ~n14164 & ~n14165;
  assign n14169 = n14167 & n14168;
  assign n14170 = ~n14151 & ~n14157;
  assign n14171 = ~n14163 & n14170;
  assign n14172 = ~n14169 & n14171;
  assign n14173 = ~P2_INSTQUEUE_REG_4__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14174 = ~P2_INSTQUEUE_REG_12__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14175 = ~P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14176 = P2_INSTQUEUERD_ADDR_REG_2_ & n14175;
  assign n14177 = ~n14173 & ~n14174;
  assign n14178 = n14176 & n14177;
  assign n14179 = ~P2_INSTQUEUE_REG_9__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14180 = ~P2_INSTQUEUE_REG_1__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14181 = ~P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign n14182 = P2_INSTQUEUERD_ADDR_REG_0_ & n14181;
  assign n14183 = ~n14179 & ~n14180;
  assign n14184 = n14182 & n14183;
  assign n14185 = ~P2_INSTQUEUE_REG_8__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14186 = ~P2_INSTQUEUE_REG_0__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14187 = ~P2_INSTQUEUERD_ADDR_REG_2_ & n14175;
  assign n14188 = ~n14185 & ~n14186;
  assign n14189 = n14187 & n14188;
  assign n14190 = ~P2_INSTQUEUE_REG_3__0_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14191 = ~P2_INSTQUEUE_REG_11__0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14192 = ~P2_INSTQUEUERD_ADDR_REG_2_ & P2_INSTQUEUERD_ADDR_REG_1_;
  assign n14193 = P2_INSTQUEUERD_ADDR_REG_0_ & n14192;
  assign n14194 = ~n14190 & ~n14191;
  assign n14195 = n14193 & n14194;
  assign n14196 = ~n14178 & ~n14184;
  assign n14197 = ~n14189 & n14196;
  assign n14198 = ~n14195 & n14197;
  assign n14199 = n14172 & n14198;
  assign n14200 = ~P2_INSTQUEUE_REG_2__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14201 = ~P2_INSTQUEUE_REG_10__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = n14149 & n14202;
  assign n14204 = ~P2_INSTQUEUE_REG_6__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14205 = ~P2_INSTQUEUE_REG_14__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14206 = ~n14204 & ~n14205;
  assign n14207 = n14155 & n14206;
  assign n14208 = ~P2_INSTQUEUE_REG_5__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14209 = ~P2_INSTQUEUE_REG_13__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14210 = ~n14208 & ~n14209;
  assign n14211 = n14161 & n14210;
  assign n14212 = ~P2_INSTQUEUE_REG_7__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14213 = ~P2_INSTQUEUE_REG_15__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = n14167 & n14214;
  assign n14216 = ~n14203 & ~n14207;
  assign n14217 = ~n14211 & n14216;
  assign n14218 = ~n14215 & n14217;
  assign n14219 = ~P2_INSTQUEUE_REG_4__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14220 = ~P2_INSTQUEUE_REG_12__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14221 = ~n14219 & ~n14220;
  assign n14222 = n14176 & n14221;
  assign n14223 = ~P2_INSTQUEUE_REG_9__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14224 = ~P2_INSTQUEUE_REG_1__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14225 = ~n14223 & ~n14224;
  assign n14226 = n14182 & n14225;
  assign n14227 = ~P2_INSTQUEUE_REG_8__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14228 = ~P2_INSTQUEUE_REG_0__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14229 = ~n14227 & ~n14228;
  assign n14230 = n14187 & n14229;
  assign n14231 = ~P2_INSTQUEUE_REG_3__1_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14232 = ~P2_INSTQUEUE_REG_11__1_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14233 = ~n14231 & ~n14232;
  assign n14234 = n14193 & n14233;
  assign n14235 = ~n14222 & ~n14226;
  assign n14236 = ~n14230 & n14235;
  assign n14237 = ~n14234 & n14236;
  assign n14238 = n14218 & n14237;
  assign n14239 = ~n14199 & n14238;
  assign n14240 = n14199 & ~n14238;
  assign n14241 = ~n14239 & ~n14240;
  assign n14242 = n14145 & ~n14241;
  assign n14243 = n14199 & n14238;
  assign n14244 = ~n14199 & ~n14238;
  assign n14245 = ~n14243 & ~n14244;
  assign n14246 = ~n14051 & ~n14245;
  assign n14247 = ~n14242 & ~n14246;
  assign n14248 = ~P2_INSTQUEUE_REG_2__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14249 = ~P2_INSTQUEUE_REG_10__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14250 = ~n14248 & ~n14249;
  assign n14251 = n14149 & n14250;
  assign n14252 = ~P2_INSTQUEUE_REG_6__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14253 = ~P2_INSTQUEUE_REG_14__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = n14155 & n14254;
  assign n14256 = ~P2_INSTQUEUE_REG_5__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14257 = ~P2_INSTQUEUE_REG_13__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14258 = ~n14256 & ~n14257;
  assign n14259 = n14161 & n14258;
  assign n14260 = ~P2_INSTQUEUE_REG_7__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14261 = ~P2_INSTQUEUE_REG_15__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14262 = ~n14260 & ~n14261;
  assign n14263 = n14167 & n14262;
  assign n14264 = ~n14251 & ~n14255;
  assign n14265 = ~n14259 & n14264;
  assign n14266 = ~n14263 & n14265;
  assign n14267 = ~P2_INSTQUEUE_REG_4__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14268 = ~P2_INSTQUEUE_REG_12__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14269 = ~n14267 & ~n14268;
  assign n14270 = n14176 & n14269;
  assign n14271 = ~P2_INSTQUEUE_REG_9__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14272 = ~P2_INSTQUEUE_REG_1__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14273 = ~n14271 & ~n14272;
  assign n14274 = n14182 & n14273;
  assign n14275 = ~P2_INSTQUEUE_REG_8__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14276 = ~P2_INSTQUEUE_REG_0__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = n14187 & n14277;
  assign n14279 = ~P2_INSTQUEUE_REG_3__7_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14280 = ~P2_INSTQUEUE_REG_11__7_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = n14193 & n14281;
  assign n14283 = ~n14270 & ~n14274;
  assign n14284 = ~n14278 & n14283;
  assign n14285 = ~n14282 & n14284;
  assign n14286 = n14266 & n14285;
  assign n14287 = ~P2_INSTQUEUE_REG_2__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14288 = ~P2_INSTQUEUE_REG_10__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = n14149 & n14289;
  assign n14291 = ~P2_INSTQUEUE_REG_6__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14292 = ~P2_INSTQUEUE_REG_14__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14293 = ~n14291 & ~n14292;
  assign n14294 = n14155 & n14293;
  assign n14295 = ~P2_INSTQUEUE_REG_5__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14296 = ~P2_INSTQUEUE_REG_13__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = n14161 & n14297;
  assign n14299 = ~P2_INSTQUEUE_REG_7__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14300 = ~P2_INSTQUEUE_REG_15__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = n14167 & n14301;
  assign n14303 = ~n14290 & ~n14294;
  assign n14304 = ~n14298 & n14303;
  assign n14305 = ~n14302 & n14304;
  assign n14306 = ~P2_INSTQUEUE_REG_4__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14307 = ~P2_INSTQUEUE_REG_12__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14308 = ~n14306 & ~n14307;
  assign n14309 = n14176 & n14308;
  assign n14310 = ~P2_INSTQUEUE_REG_9__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14311 = ~P2_INSTQUEUE_REG_1__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14312 = ~n14310 & ~n14311;
  assign n14313 = n14182 & n14312;
  assign n14314 = ~P2_INSTQUEUE_REG_8__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14315 = ~P2_INSTQUEUE_REG_0__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = n14187 & n14316;
  assign n14318 = ~P2_INSTQUEUE_REG_3__3_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14319 = ~P2_INSTQUEUE_REG_11__3_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14320 = ~n14318 & ~n14319;
  assign n14321 = n14193 & n14320;
  assign n14322 = ~n14309 & ~n14313;
  assign n14323 = ~n14317 & n14322;
  assign n14324 = ~n14321 & n14323;
  assign n14325 = n14305 & n14324;
  assign n14326 = ~n14286 & ~n14325;
  assign n14327 = ~P2_INSTQUEUE_REG_2__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14328 = ~P2_INSTQUEUE_REG_10__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14329 = ~n14327 & ~n14328;
  assign n14330 = n14149 & n14329;
  assign n14331 = ~P2_INSTQUEUE_REG_6__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14332 = ~P2_INSTQUEUE_REG_14__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14333 = ~n14331 & ~n14332;
  assign n14334 = n14155 & n14333;
  assign n14335 = ~P2_INSTQUEUE_REG_5__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14336 = ~P2_INSTQUEUE_REG_13__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14337 = ~n14335 & ~n14336;
  assign n14338 = n14161 & n14337;
  assign n14339 = ~P2_INSTQUEUE_REG_7__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14340 = ~P2_INSTQUEUE_REG_15__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14341 = ~n14339 & ~n14340;
  assign n14342 = n14167 & n14341;
  assign n14343 = ~n14330 & ~n14334;
  assign n14344 = ~n14338 & n14343;
  assign n14345 = ~n14342 & n14344;
  assign n14346 = ~P2_INSTQUEUE_REG_4__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14347 = ~P2_INSTQUEUE_REG_12__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14348 = ~n14346 & ~n14347;
  assign n14349 = n14176 & n14348;
  assign n14350 = ~P2_INSTQUEUE_REG_9__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14351 = ~P2_INSTQUEUE_REG_1__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = n14182 & n14352;
  assign n14354 = ~P2_INSTQUEUE_REG_8__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14355 = ~P2_INSTQUEUE_REG_0__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14356 = ~n14354 & ~n14355;
  assign n14357 = n14187 & n14356;
  assign n14358 = ~P2_INSTQUEUE_REG_3__5_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14359 = ~P2_INSTQUEUE_REG_11__5_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14360 = ~n14358 & ~n14359;
  assign n14361 = n14193 & n14360;
  assign n14362 = ~n14349 & ~n14353;
  assign n14363 = ~n14357 & n14362;
  assign n14364 = ~n14361 & n14363;
  assign n14365 = n14345 & n14364;
  assign n14366 = ~P2_INSTQUEUE_REG_2__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14367 = ~P2_INSTQUEUE_REG_10__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14368 = ~n14366 & ~n14367;
  assign n14369 = n14149 & n14368;
  assign n14370 = ~P2_INSTQUEUE_REG_6__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14371 = ~P2_INSTQUEUE_REG_14__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14372 = ~n14370 & ~n14371;
  assign n14373 = n14155 & n14372;
  assign n14374 = ~P2_INSTQUEUE_REG_5__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14375 = ~P2_INSTQUEUE_REG_13__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14376 = ~n14374 & ~n14375;
  assign n14377 = n14161 & n14376;
  assign n14378 = ~P2_INSTQUEUE_REG_7__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14379 = ~P2_INSTQUEUE_REG_15__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14380 = ~n14378 & ~n14379;
  assign n14381 = n14167 & n14380;
  assign n14382 = ~n14369 & ~n14373;
  assign n14383 = ~n14377 & n14382;
  assign n14384 = ~n14381 & n14383;
  assign n14385 = ~P2_INSTQUEUE_REG_4__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14386 = ~P2_INSTQUEUE_REG_12__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = n14176 & n14387;
  assign n14389 = ~P2_INSTQUEUE_REG_9__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14390 = ~P2_INSTQUEUE_REG_1__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14391 = ~n14389 & ~n14390;
  assign n14392 = n14182 & n14391;
  assign n14393 = ~P2_INSTQUEUE_REG_8__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14394 = ~P2_INSTQUEUE_REG_0__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14395 = ~n14393 & ~n14394;
  assign n14396 = n14187 & n14395;
  assign n14397 = ~P2_INSTQUEUE_REG_3__6_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14398 = ~P2_INSTQUEUE_REG_11__6_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14399 = ~n14397 & ~n14398;
  assign n14400 = n14193 & n14399;
  assign n14401 = ~n14388 & ~n14392;
  assign n14402 = ~n14396 & n14401;
  assign n14403 = ~n14400 & n14402;
  assign n14404 = n14384 & n14403;
  assign n14405 = ~P2_INSTQUEUE_REG_2__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14406 = ~P2_INSTQUEUE_REG_10__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14407 = ~n14405 & ~n14406;
  assign n14408 = n14149 & n14407;
  assign n14409 = ~P2_INSTQUEUE_REG_6__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14410 = ~P2_INSTQUEUE_REG_14__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14411 = ~n14409 & ~n14410;
  assign n14412 = n14155 & n14411;
  assign n14413 = ~P2_INSTQUEUE_REG_5__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14414 = ~P2_INSTQUEUE_REG_13__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14415 = ~n14413 & ~n14414;
  assign n14416 = n14161 & n14415;
  assign n14417 = ~P2_INSTQUEUE_REG_7__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14418 = ~P2_INSTQUEUE_REG_15__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14419 = ~n14417 & ~n14418;
  assign n14420 = n14167 & n14419;
  assign n14421 = ~n14408 & ~n14412;
  assign n14422 = ~n14416 & n14421;
  assign n14423 = ~n14420 & n14422;
  assign n14424 = ~P2_INSTQUEUE_REG_4__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14425 = ~P2_INSTQUEUE_REG_12__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14426 = ~n14424 & ~n14425;
  assign n14427 = n14176 & n14426;
  assign n14428 = ~P2_INSTQUEUE_REG_9__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14429 = ~P2_INSTQUEUE_REG_1__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14430 = ~n14428 & ~n14429;
  assign n14431 = n14182 & n14430;
  assign n14432 = ~P2_INSTQUEUE_REG_8__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14433 = ~P2_INSTQUEUE_REG_0__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14434 = ~n14432 & ~n14433;
  assign n14435 = n14187 & n14434;
  assign n14436 = ~P2_INSTQUEUE_REG_3__4_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14437 = ~P2_INSTQUEUE_REG_11__4_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14438 = ~n14436 & ~n14437;
  assign n14439 = n14193 & n14438;
  assign n14440 = ~n14427 & ~n14431;
  assign n14441 = ~n14435 & n14440;
  assign n14442 = ~n14439 & n14441;
  assign n14443 = n14423 & n14442;
  assign n14444 = ~P2_INSTQUEUE_REG_2__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14445 = ~P2_INSTQUEUE_REG_10__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14446 = ~n14444 & ~n14445;
  assign n14447 = n14149 & n14446;
  assign n14448 = ~P2_INSTQUEUE_REG_6__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14449 = ~P2_INSTQUEUE_REG_14__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14450 = ~n14448 & ~n14449;
  assign n14451 = n14155 & n14450;
  assign n14452 = ~P2_INSTQUEUE_REG_5__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14453 = ~P2_INSTQUEUE_REG_13__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14454 = ~n14452 & ~n14453;
  assign n14455 = n14161 & n14454;
  assign n14456 = ~P2_INSTQUEUE_REG_7__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14457 = ~P2_INSTQUEUE_REG_15__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14458 = ~n14456 & ~n14457;
  assign n14459 = n14167 & n14458;
  assign n14460 = ~n14447 & ~n14451;
  assign n14461 = ~n14455 & n14460;
  assign n14462 = ~n14459 & n14461;
  assign n14463 = ~P2_INSTQUEUE_REG_4__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14464 = ~P2_INSTQUEUE_REG_12__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14465 = ~n14463 & ~n14464;
  assign n14466 = n14176 & n14465;
  assign n14467 = ~P2_INSTQUEUE_REG_9__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14468 = ~P2_INSTQUEUE_REG_1__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = n14182 & n14469;
  assign n14471 = ~P2_INSTQUEUE_REG_8__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14472 = ~P2_INSTQUEUE_REG_0__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14473 = ~n14471 & ~n14472;
  assign n14474 = n14187 & n14473;
  assign n14475 = ~P2_INSTQUEUE_REG_3__2_ & ~P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14476 = ~P2_INSTQUEUE_REG_11__2_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14477 = ~n14475 & ~n14476;
  assign n14478 = n14193 & n14477;
  assign n14479 = ~n14466 & ~n14470;
  assign n14480 = ~n14474 & n14479;
  assign n14481 = ~n14478 & n14480;
  assign n14482 = n14462 & n14481;
  assign n14483 = n14404 & n14443;
  assign n14484 = n14482 & n14483;
  assign n14485 = n14326 & n14365;
  assign n14486 = n14484 & n14485;
  assign n14487 = ~n14199 & ~n14486;
  assign n14488 = ~n14286 & n14325;
  assign n14489 = ~n14365 & ~n14404;
  assign n14490 = n14443 & n14489;
  assign n14491 = n14488 & n14490;
  assign n14492 = ~n14482 & n14491;
  assign n14493 = n14199 & ~n14492;
  assign n14494 = P2_INSTQUEUERD_ADDR_REG_4_ & ~P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n14495 = ~P2_INSTQUEUERD_ADDR_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n14496 = P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n14497 = ~P2_INSTQUEUERD_ADDR_REG_2_ & P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n14498 = P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n14499 = P2_INSTQUEUERD_ADDR_REG_0_ & ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n14500 = P2_INSTQUEUEWR_ADDR_REG_1_ & ~n14499;
  assign n14501 = ~P2_INSTQUEUEWR_ADDR_REG_1_ & n14499;
  assign n14502 = ~P2_INSTQUEUERD_ADDR_REG_1_ & ~n14501;
  assign n14503 = ~n14500 & ~n14502;
  assign n14504 = ~n14498 & ~n14503;
  assign n14505 = ~n14497 & ~n14504;
  assign n14506 = ~n14496 & ~n14505;
  assign n14507 = ~n14495 & ~n14506;
  assign n14508 = ~P2_INSTQUEUERD_ADDR_REG_4_ & P2_INSTQUEUEWR_ADDR_REG_4_;
  assign n14509 = n14507 & ~n14508;
  assign n14510 = ~n14494 & ~n14509;
  assign n14511 = n14239 & ~n14510;
  assign n14512 = ~n14239 & ~n14510;
  assign n14513 = ~n14511 & ~n14512;
  assign n14514 = ~n14494 & ~n14508;
  assign n14515 = ~n14507 & ~n14514;
  assign n14516 = n14507 & n14514;
  assign n14517 = ~n14515 & ~n14516;
  assign n14518 = n14239 & ~n14517;
  assign n14519 = ~n14239 & ~n14517;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521 = ~n14495 & ~n14496;
  assign n14522 = ~n14505 & ~n14521;
  assign n14523 = n14505 & n14521;
  assign n14524 = ~n14522 & ~n14523;
  assign n14525 = n14239 & ~n14524;
  assign n14526 = ~n14239 & ~n14524;
  assign n14527 = ~n14525 & ~n14526;
  assign n14528 = ~P2_INSTQUEUERD_ADDR_REG_1_ & P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n14529 = P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n14530 = ~n14528 & ~n14529;
  assign n14531 = ~n14499 & ~n14530;
  assign n14532 = n14499 & n14530;
  assign n14533 = ~n14531 & ~n14532;
  assign n14534 = n14239 & ~n14533;
  assign n14535 = ~n14239 & ~n14533;
  assign n14536 = ~n14534 & ~n14535;
  assign n14537 = ~n14497 & ~n14498;
  assign n14538 = ~n14503 & ~n14537;
  assign n14539 = n14503 & n14537;
  assign n14540 = ~n14538 & ~n14539;
  assign n14541 = n14239 & ~n14540;
  assign n14542 = ~n14239 & ~n14540;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = n14513 & n14520;
  assign n14545 = n14527 & n14544;
  assign n14546 = n14536 & n14545;
  assign n14547 = n14543 & n14546;
  assign n14548 = n14513 & ~n14547;
  assign n14549 = ~n14240 & ~n14548;
  assign n14550 = P2_STATE2_REG_0_ & ~n14199;
  assign n14551 = ~n14510 & n14550;
  assign n14552 = ~P2_INSTQUEUERD_ADDR_REG_3_ & n14167;
  assign n14553 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n14167;
  assign n14554 = ~n14552 & ~n14553;
  assign n14555 = ~n14154 & ~n14160;
  assign n14556 = n14554 & n14555;
  assign n14557 = P2_INSTQUEUERD_ADDR_REG_2_ & ~n14166;
  assign n14558 = ~n14193 & ~n14557;
  assign n14559 = P2_INSTQUEUERD_ADDR_REG_0_ & n14558;
  assign n14560 = n14556 & n14559;
  assign n14561 = P2_INSTQUEUE_REG_0__6_ & n14560;
  assign n14562 = ~P2_INSTQUEUERD_ADDR_REG_0_ & n14558;
  assign n14563 = n14556 & n14562;
  assign n14564 = P2_INSTQUEUE_REG_1__6_ & n14563;
  assign n14565 = n14554 & ~n14555;
  assign n14566 = n14559 & n14565;
  assign n14567 = P2_INSTQUEUE_REG_2__6_ & n14566;
  assign n14568 = n14562 & n14565;
  assign n14569 = P2_INSTQUEUE_REG_3__6_ & n14568;
  assign n14570 = ~n14561 & ~n14564;
  assign n14571 = ~n14567 & n14570;
  assign n14572 = ~n14569 & n14571;
  assign n14573 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n14558;
  assign n14574 = n14556 & n14573;
  assign n14575 = P2_INSTQUEUE_REG_4__6_ & n14574;
  assign n14576 = ~P2_INSTQUEUERD_ADDR_REG_0_ & ~n14558;
  assign n14577 = n14556 & n14576;
  assign n14578 = P2_INSTQUEUE_REG_5__6_ & n14577;
  assign n14579 = n14565 & n14573;
  assign n14580 = P2_INSTQUEUE_REG_6__6_ & n14579;
  assign n14581 = n14565 & n14576;
  assign n14582 = P2_INSTQUEUE_REG_7__6_ & n14581;
  assign n14583 = ~n14575 & ~n14578;
  assign n14584 = ~n14580 & n14583;
  assign n14585 = ~n14582 & n14584;
  assign n14586 = ~n14554 & ~n14555;
  assign n14587 = n14576 & n14586;
  assign n14588 = P2_INSTQUEUE_REG_15__6_ & n14587;
  assign n14589 = n14573 & n14586;
  assign n14590 = P2_INSTQUEUE_REG_14__6_ & n14589;
  assign n14591 = ~n14554 & n14555;
  assign n14592 = n14576 & n14591;
  assign n14593 = P2_INSTQUEUE_REG_13__6_ & n14592;
  assign n14594 = n14573 & n14591;
  assign n14595 = P2_INSTQUEUE_REG_12__6_ & n14594;
  assign n14596 = ~n14588 & ~n14590;
  assign n14597 = ~n14593 & n14596;
  assign n14598 = ~n14595 & n14597;
  assign n14599 = n14562 & n14586;
  assign n14600 = P2_INSTQUEUE_REG_11__6_ & n14599;
  assign n14601 = n14559 & n14586;
  assign n14602 = P2_INSTQUEUE_REG_10__6_ & n14601;
  assign n14603 = n14562 & n14591;
  assign n14604 = P2_INSTQUEUE_REG_9__6_ & n14603;
  assign n14605 = n14559 & n14591;
  assign n14606 = P2_INSTQUEUE_REG_8__6_ & n14605;
  assign n14607 = ~n14600 & ~n14602;
  assign n14608 = ~n14604 & n14607;
  assign n14609 = ~n14606 & n14608;
  assign n14610 = n14572 & n14585;
  assign n14611 = n14598 & n14610;
  assign n14612 = n14609 & n14611;
  assign n14613 = n14244 & ~n14612;
  assign n14614 = n14244 & ~n14613;
  assign n14615 = ~n14244 & n14613;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = P2_INSTQUEUE_REG_0__5_ & n14560;
  assign n14618 = P2_INSTQUEUE_REG_1__5_ & n14563;
  assign n14619 = P2_INSTQUEUE_REG_2__5_ & n14566;
  assign n14620 = P2_INSTQUEUE_REG_3__5_ & n14568;
  assign n14621 = ~n14617 & ~n14618;
  assign n14622 = ~n14619 & n14621;
  assign n14623 = ~n14620 & n14622;
  assign n14624 = P2_INSTQUEUE_REG_4__5_ & n14574;
  assign n14625 = P2_INSTQUEUE_REG_5__5_ & n14577;
  assign n14626 = P2_INSTQUEUE_REG_6__5_ & n14579;
  assign n14627 = P2_INSTQUEUE_REG_7__5_ & n14581;
  assign n14628 = ~n14624 & ~n14625;
  assign n14629 = ~n14626 & n14628;
  assign n14630 = ~n14627 & n14629;
  assign n14631 = P2_INSTQUEUE_REG_15__5_ & n14587;
  assign n14632 = P2_INSTQUEUE_REG_14__5_ & n14589;
  assign n14633 = P2_INSTQUEUE_REG_13__5_ & n14592;
  assign n14634 = P2_INSTQUEUE_REG_12__5_ & n14594;
  assign n14635 = ~n14631 & ~n14632;
  assign n14636 = ~n14633 & n14635;
  assign n14637 = ~n14634 & n14636;
  assign n14638 = P2_INSTQUEUE_REG_11__5_ & n14599;
  assign n14639 = P2_INSTQUEUE_REG_10__5_ & n14601;
  assign n14640 = P2_INSTQUEUE_REG_9__5_ & n14603;
  assign n14641 = P2_INSTQUEUE_REG_8__5_ & n14605;
  assign n14642 = ~n14638 & ~n14639;
  assign n14643 = ~n14640 & n14642;
  assign n14644 = ~n14641 & n14643;
  assign n14645 = n14623 & n14630;
  assign n14646 = n14637 & n14645;
  assign n14647 = n14644 & n14646;
  assign n14648 = n14244 & ~n14647;
  assign n14649 = n14244 & ~n14648;
  assign n14650 = ~n14244 & n14648;
  assign n14651 = n14241 & ~n14243;
  assign n14652 = P2_INSTQUEUEWR_ADDR_REG_3_ & ~n14651;
  assign n14653 = ~n14244 & ~n14652;
  assign n14654 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n14651;
  assign n14655 = P2_INSTQUEUE_REG_0__3_ & n14560;
  assign n14656 = P2_INSTQUEUE_REG_1__3_ & n14563;
  assign n14657 = P2_INSTQUEUE_REG_2__3_ & n14566;
  assign n14658 = P2_INSTQUEUE_REG_3__3_ & n14568;
  assign n14659 = ~n14655 & ~n14656;
  assign n14660 = ~n14657 & n14659;
  assign n14661 = ~n14658 & n14660;
  assign n14662 = P2_INSTQUEUE_REG_4__3_ & n14574;
  assign n14663 = P2_INSTQUEUE_REG_5__3_ & n14577;
  assign n14664 = P2_INSTQUEUE_REG_6__3_ & n14579;
  assign n14665 = P2_INSTQUEUE_REG_7__3_ & n14581;
  assign n14666 = ~n14662 & ~n14663;
  assign n14667 = ~n14664 & n14666;
  assign n14668 = ~n14665 & n14667;
  assign n14669 = P2_INSTQUEUE_REG_15__3_ & n14587;
  assign n14670 = P2_INSTQUEUE_REG_14__3_ & n14589;
  assign n14671 = P2_INSTQUEUE_REG_13__3_ & n14592;
  assign n14672 = P2_INSTQUEUE_REG_12__3_ & n14594;
  assign n14673 = ~n14669 & ~n14670;
  assign n14674 = ~n14671 & n14673;
  assign n14675 = ~n14672 & n14674;
  assign n14676 = P2_INSTQUEUE_REG_11__3_ & n14599;
  assign n14677 = P2_INSTQUEUE_REG_10__3_ & n14601;
  assign n14678 = P2_INSTQUEUE_REG_9__3_ & n14603;
  assign n14679 = P2_INSTQUEUE_REG_8__3_ & n14605;
  assign n14680 = ~n14676 & ~n14677;
  assign n14681 = ~n14678 & n14680;
  assign n14682 = ~n14679 & n14681;
  assign n14683 = n14661 & n14668;
  assign n14684 = n14675 & n14683;
  assign n14685 = n14682 & n14684;
  assign n14686 = n14244 & ~n14685;
  assign n14687 = ~n14654 & ~n14686;
  assign n14688 = ~n14653 & n14687;
  assign n14689 = P2_INSTQUEUEWR_ADDR_REG_2_ & ~n14651;
  assign n14690 = ~n14244 & ~n14689;
  assign n14691 = P2_INSTQUEUERD_ADDR_REG_2_ & ~n14651;
  assign n14692 = P2_INSTQUEUE_REG_0__2_ & n14560;
  assign n14693 = P2_INSTQUEUE_REG_1__2_ & n14563;
  assign n14694 = P2_INSTQUEUE_REG_2__2_ & n14566;
  assign n14695 = P2_INSTQUEUE_REG_3__2_ & n14568;
  assign n14696 = ~n14692 & ~n14693;
  assign n14697 = ~n14694 & n14696;
  assign n14698 = ~n14695 & n14697;
  assign n14699 = P2_INSTQUEUE_REG_4__2_ & n14574;
  assign n14700 = P2_INSTQUEUE_REG_5__2_ & n14577;
  assign n14701 = P2_INSTQUEUE_REG_6__2_ & n14579;
  assign n14702 = P2_INSTQUEUE_REG_7__2_ & n14581;
  assign n14703 = ~n14699 & ~n14700;
  assign n14704 = ~n14701 & n14703;
  assign n14705 = ~n14702 & n14704;
  assign n14706 = P2_INSTQUEUE_REG_15__2_ & n14587;
  assign n14707 = P2_INSTQUEUE_REG_14__2_ & n14589;
  assign n14708 = P2_INSTQUEUE_REG_13__2_ & n14592;
  assign n14709 = P2_INSTQUEUE_REG_12__2_ & n14594;
  assign n14710 = ~n14706 & ~n14707;
  assign n14711 = ~n14708 & n14710;
  assign n14712 = ~n14709 & n14711;
  assign n14713 = P2_INSTQUEUE_REG_11__2_ & n14599;
  assign n14714 = P2_INSTQUEUE_REG_10__2_ & n14601;
  assign n14715 = P2_INSTQUEUE_REG_9__2_ & n14603;
  assign n14716 = P2_INSTQUEUE_REG_8__2_ & n14605;
  assign n14717 = ~n14713 & ~n14714;
  assign n14718 = ~n14715 & n14717;
  assign n14719 = ~n14716 & n14718;
  assign n14720 = n14698 & n14705;
  assign n14721 = n14712 & n14720;
  assign n14722 = n14719 & n14721;
  assign n14723 = n14244 & ~n14722;
  assign n14724 = ~n14691 & ~n14723;
  assign n14725 = ~n14690 & n14724;
  assign n14726 = ~n14688 & ~n14725;
  assign n14727 = n14653 & ~n14687;
  assign n14728 = ~n14726 & ~n14727;
  assign n14729 = P2_INSTQUEUERD_ADDR_REG_4_ & ~n14651;
  assign n14730 = P2_INSTQUEUE_REG_0__4_ & n14560;
  assign n14731 = P2_INSTQUEUE_REG_1__4_ & n14563;
  assign n14732 = P2_INSTQUEUE_REG_2__4_ & n14566;
  assign n14733 = P2_INSTQUEUE_REG_3__4_ & n14568;
  assign n14734 = ~n14730 & ~n14731;
  assign n14735 = ~n14732 & n14734;
  assign n14736 = ~n14733 & n14735;
  assign n14737 = P2_INSTQUEUE_REG_4__4_ & n14574;
  assign n14738 = P2_INSTQUEUE_REG_5__4_ & n14577;
  assign n14739 = P2_INSTQUEUE_REG_6__4_ & n14579;
  assign n14740 = P2_INSTQUEUE_REG_7__4_ & n14581;
  assign n14741 = ~n14737 & ~n14738;
  assign n14742 = ~n14739 & n14741;
  assign n14743 = ~n14740 & n14742;
  assign n14744 = P2_INSTQUEUE_REG_15__4_ & n14587;
  assign n14745 = P2_INSTQUEUE_REG_14__4_ & n14589;
  assign n14746 = P2_INSTQUEUE_REG_13__4_ & n14592;
  assign n14747 = P2_INSTQUEUE_REG_12__4_ & n14594;
  assign n14748 = ~n14744 & ~n14745;
  assign n14749 = ~n14746 & n14748;
  assign n14750 = ~n14747 & n14749;
  assign n14751 = P2_INSTQUEUE_REG_11__4_ & n14599;
  assign n14752 = P2_INSTQUEUE_REG_10__4_ & n14601;
  assign n14753 = P2_INSTQUEUE_REG_9__4_ & n14603;
  assign n14754 = P2_INSTQUEUE_REG_8__4_ & n14605;
  assign n14755 = ~n14751 & ~n14752;
  assign n14756 = ~n14753 & n14755;
  assign n14757 = ~n14754 & n14756;
  assign n14758 = n14736 & n14743;
  assign n14759 = n14750 & n14758;
  assign n14760 = n14757 & n14759;
  assign n14761 = n14244 & ~n14760;
  assign n14762 = ~n14729 & ~n14761;
  assign n14763 = P2_INSTQUEUEWR_ADDR_REG_4_ & ~n14651;
  assign n14764 = ~n14244 & ~n14763;
  assign n14765 = ~n14762 & n14764;
  assign n14766 = n14728 & ~n14765;
  assign n14767 = n14762 & ~n14764;
  assign n14768 = n14690 & ~n14724;
  assign n14769 = ~n14727 & ~n14768;
  assign n14770 = ~n14765 & n14769;
  assign n14771 = P2_INSTQUEUERD_ADDR_REG_1_ & ~n14651;
  assign n14772 = P2_INSTQUEUE_REG_0__1_ & n14560;
  assign n14773 = P2_INSTQUEUE_REG_1__1_ & n14563;
  assign n14774 = P2_INSTQUEUE_REG_2__1_ & n14566;
  assign n14775 = P2_INSTQUEUE_REG_3__1_ & n14568;
  assign n14776 = ~n14772 & ~n14773;
  assign n14777 = ~n14774 & n14776;
  assign n14778 = ~n14775 & n14777;
  assign n14779 = P2_INSTQUEUE_REG_4__1_ & n14574;
  assign n14780 = P2_INSTQUEUE_REG_5__1_ & n14577;
  assign n14781 = P2_INSTQUEUE_REG_6__1_ & n14579;
  assign n14782 = P2_INSTQUEUE_REG_7__1_ & n14581;
  assign n14783 = ~n14779 & ~n14780;
  assign n14784 = ~n14781 & n14783;
  assign n14785 = ~n14782 & n14784;
  assign n14786 = P2_INSTQUEUE_REG_15__1_ & n14587;
  assign n14787 = P2_INSTQUEUE_REG_14__1_ & n14589;
  assign n14788 = P2_INSTQUEUE_REG_13__1_ & n14592;
  assign n14789 = P2_INSTQUEUE_REG_12__1_ & n14594;
  assign n14790 = ~n14786 & ~n14787;
  assign n14791 = ~n14788 & n14790;
  assign n14792 = ~n14789 & n14791;
  assign n14793 = P2_INSTQUEUE_REG_11__1_ & n14599;
  assign n14794 = P2_INSTQUEUE_REG_10__1_ & n14601;
  assign n14795 = P2_INSTQUEUE_REG_9__1_ & n14603;
  assign n14796 = P2_INSTQUEUE_REG_8__1_ & n14605;
  assign n14797 = ~n14793 & ~n14794;
  assign n14798 = ~n14795 & n14797;
  assign n14799 = ~n14796 & n14798;
  assign n14800 = n14778 & n14785;
  assign n14801 = n14792 & n14800;
  assign n14802 = n14799 & n14801;
  assign n14803 = n14244 & ~n14802;
  assign n14804 = ~n14771 & ~n14803;
  assign n14805 = P2_INSTQUEUEWR_ADDR_REG_1_ & ~n14651;
  assign n14806 = ~n14244 & ~n14805;
  assign n14807 = ~n14804 & n14806;
  assign n14808 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n14651;
  assign n14809 = P2_INSTQUEUE_REG_0__0_ & n14560;
  assign n14810 = P2_INSTQUEUE_REG_1__0_ & n14563;
  assign n14811 = P2_INSTQUEUE_REG_2__0_ & n14566;
  assign n14812 = P2_INSTQUEUE_REG_3__0_ & n14568;
  assign n14813 = ~n14809 & ~n14810;
  assign n14814 = ~n14811 & n14813;
  assign n14815 = ~n14812 & n14814;
  assign n14816 = P2_INSTQUEUE_REG_4__0_ & n14574;
  assign n14817 = P2_INSTQUEUE_REG_5__0_ & n14577;
  assign n14818 = P2_INSTQUEUE_REG_6__0_ & n14579;
  assign n14819 = P2_INSTQUEUE_REG_7__0_ & n14581;
  assign n14820 = ~n14816 & ~n14817;
  assign n14821 = ~n14818 & n14820;
  assign n14822 = ~n14819 & n14821;
  assign n14823 = P2_INSTQUEUE_REG_15__0_ & n14587;
  assign n14824 = P2_INSTQUEUE_REG_14__0_ & n14589;
  assign n14825 = P2_INSTQUEUE_REG_13__0_ & n14592;
  assign n14826 = P2_INSTQUEUE_REG_12__0_ & n14594;
  assign n14827 = ~n14823 & ~n14824;
  assign n14828 = ~n14825 & n14827;
  assign n14829 = ~n14826 & n14828;
  assign n14830 = P2_INSTQUEUE_REG_11__0_ & n14599;
  assign n14831 = P2_INSTQUEUE_REG_10__0_ & n14601;
  assign n14832 = P2_INSTQUEUE_REG_9__0_ & n14603;
  assign n14833 = P2_INSTQUEUE_REG_8__0_ & n14605;
  assign n14834 = ~n14830 & ~n14831;
  assign n14835 = ~n14832 & n14834;
  assign n14836 = ~n14833 & n14835;
  assign n14837 = n14815 & n14822;
  assign n14838 = n14829 & n14837;
  assign n14839 = n14836 & n14838;
  assign n14840 = n14244 & ~n14839;
  assign n14841 = ~n14808 & ~n14840;
  assign n14842 = P2_INSTQUEUEWR_ADDR_REG_0_ & ~n14651;
  assign n14843 = ~n14244 & ~n14842;
  assign n14844 = ~n14841 & n14843;
  assign n14845 = ~n14807 & ~n14844;
  assign n14846 = n14804 & ~n14806;
  assign n14847 = ~n14845 & ~n14846;
  assign n14848 = n14770 & ~n14847;
  assign n14849 = ~n14766 & ~n14767;
  assign n14850 = ~n14848 & n14849;
  assign n14851 = ~n14650 & ~n14850;
  assign n14852 = ~n14649 & ~n14851;
  assign n14853 = ~n14616 & ~n14852;
  assign n14854 = n14616 & n14852;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = P2_STATE2_REG_0_ & n14240;
  assign n14857 = P2_STATE2_REG_0_ & n14238;
  assign n14858 = ~n14856 & ~n14857;
  assign n14859 = ~n14855 & ~n14858;
  assign n14860 = ~P2_STATE2_REG_0_ & ~n14551;
  assign n14861 = n14859 & n14860;
  assign n14862 = P2_STATE2_REG_0_ & n14551;
  assign n14863 = ~n14859 & n14862;
  assign n14864 = ~n14551 & n14859;
  assign n14865 = n14551 & ~n14859;
  assign n14866 = ~n14649 & ~n14650;
  assign n14867 = ~n14850 & ~n14866;
  assign n14868 = n14850 & n14866;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = ~n14858 & ~n14869;
  assign n14871 = ~n14551 & n14870;
  assign n14872 = ~P2_STATE2_REG_0_ & P2_INSTQUEUERD_ADDR_REG_4_;
  assign n14873 = ~n14517 & n14550;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = ~n14765 & ~n14767;
  assign n14876 = n14769 & ~n14847;
  assign n14877 = ~n14728 & ~n14876;
  assign n14878 = ~n14875 & ~n14877;
  assign n14879 = n14875 & n14877;
  assign n14880 = ~n14878 & ~n14879;
  assign n14881 = ~n14858 & ~n14880;
  assign n14882 = ~n14874 & ~n14881;
  assign n14883 = ~n14688 & ~n14727;
  assign n14884 = ~n14768 & ~n14847;
  assign n14885 = ~n14725 & ~n14884;
  assign n14886 = ~n14883 & ~n14885;
  assign n14887 = n14883 & n14885;
  assign n14888 = ~n14886 & ~n14887;
  assign n14889 = ~n14858 & ~n14888;
  assign n14890 = P2_STATE2_REG_0_ & ~n14889;
  assign n14891 = ~P2_STATE2_REG_0_ & P2_INSTQUEUERD_ADDR_REG_3_;
  assign n14892 = ~n14524 & n14550;
  assign n14893 = ~n14891 & ~n14892;
  assign n14894 = ~n14890 & n14893;
  assign n14895 = ~P2_STATE2_REG_0_ & P2_INSTQUEUERD_ADDR_REG_2_;
  assign n14896 = ~n14857 & ~n14895;
  assign n14897 = ~n14540 & n14550;
  assign n14898 = n14896 & ~n14897;
  assign n14899 = ~n14725 & ~n14768;
  assign n14900 = ~n14847 & ~n14899;
  assign n14901 = n14847 & n14899;
  assign n14902 = ~n14900 & ~n14901;
  assign n14903 = P2_STATE2_REG_0_ & n14199;
  assign n14904 = n14902 & n14903;
  assign n14905 = ~n14898 & n14904;
  assign n14906 = n14890 & ~n14893;
  assign n14907 = ~n14807 & ~n14846;
  assign n14908 = ~n14844 & ~n14907;
  assign n14909 = n14844 & n14907;
  assign n14910 = ~n14908 & ~n14909;
  assign n14911 = ~n14858 & ~n14910;
  assign n14912 = P2_STATE2_REG_0_ & ~n14911;
  assign n14913 = ~n14533 & n14550;
  assign n14914 = ~P2_STATE2_REG_0_ & P2_INSTQUEUERD_ADDR_REG_1_;
  assign n14915 = ~n14913 & ~n14914;
  assign n14916 = ~n14856 & n14915;
  assign n14917 = ~n14912 & n14916;
  assign n14918 = n14898 & ~n14904;
  assign n14919 = n14841 & ~n14843;
  assign n14920 = ~n14844 & ~n14919;
  assign n14921 = n14903 & n14920;
  assign n14922 = ~n14238 & n14550;
  assign n14923 = n14921 & n14922;
  assign n14924 = ~P2_STATE2_REG_0_ & P2_INSTQUEUERD_ADDR_REG_0_;
  assign n14925 = ~n14857 & ~n14924;
  assign n14926 = ~P2_INSTQUEUERD_ADDR_REG_0_ & P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n14927 = ~n14499 & ~n14926;
  assign n14928 = n14550 & ~n14927;
  assign n14929 = n14925 & ~n14928;
  assign n14930 = ~n14921 & ~n14922;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = n14912 & ~n14916;
  assign n14933 = ~n14923 & ~n14931;
  assign n14934 = ~n14932 & n14933;
  assign n14935 = ~n14917 & ~n14918;
  assign n14936 = ~n14934 & n14935;
  assign n14937 = ~n14905 & ~n14906;
  assign n14938 = ~n14936 & n14937;
  assign n14939 = n14874 & n14881;
  assign n14940 = ~n14894 & ~n14938;
  assign n14941 = ~n14939 & n14940;
  assign n14942 = n14551 & ~n14870;
  assign n14943 = ~n14882 & ~n14941;
  assign n14944 = ~n14942 & n14943;
  assign n14945 = ~n14871 & ~n14944;
  assign n14946 = ~n14864 & ~n14865;
  assign n14947 = ~n14945 & n14946;
  assign n14948 = ~n14861 & ~n14863;
  assign n14949 = ~n14947 & n14948;
  assign n14950 = n14240 & n14949;
  assign n14951 = ~n14549 & ~n14950;
  assign n14952 = ~n14487 & ~n14493;
  assign n14953 = n14951 & n14952;
  assign n14954 = n14247 & n14953;
  assign n14955 = ~P2_FLUSH_REG & ~P2_MORE_REG;
  assign n14956 = n14954 & ~n14955;
  assign n14957 = n14286 & n14443;
  assign n14958 = ~n14404 & n14957;
  assign n14959 = n14365 & n14958;
  assign n14960 = n14325 & n14482;
  assign n14961 = n14959 & n14960;
  assign n14962 = n14244 & n14961;
  assign n14963 = n14404 & ~n14443;
  assign n14964 = n14243 & n14963;
  assign n14965 = ~n14286 & n14365;
  assign n14966 = n14960 & n14965;
  assign n14967 = n14964 & n14966;
  assign n14968 = ~n14962 & ~n14967;
  assign n14969 = ~n14554 & ~n14968;
  assign n14970 = ~P2_INSTQUEUERD_ADDR_REG_2_ & ~n14166;
  assign n14971 = ~P2_INSTQUEUERD_ADDR_REG_3_ & n14970;
  assign n14972 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n14970;
  assign n14973 = ~n14971 & ~n14972;
  assign n14974 = ~n14365 & n14404;
  assign n14975 = ~n14443 & n14482;
  assign n14976 = n14326 & n14974;
  assign n14977 = n14975 & n14976;
  assign n14978 = n14244 & n14977;
  assign n14979 = n14243 & n14977;
  assign n14980 = ~n14978 & ~n14979;
  assign n14981 = n14973 & ~n14980;
  assign n14982 = ~n14969 & ~n14981;
  assign n14983 = P2_INSTQUEUERD_ADDR_REG_2_ & P2_INSTQUEUERD_ADDR_REG_1_;
  assign n14984 = ~P2_INSTQUEUERD_ADDR_REG_3_ & n14983;
  assign n14985 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n14983;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = n14199 & n14492;
  assign n14988 = ~n14199 & n14486;
  assign n14989 = n14243 & ~n14404;
  assign n14990 = n14966 & n14989;
  assign n14991 = ~n14987 & ~n14988;
  assign n14992 = ~n14990 & n14991;
  assign n14993 = ~n14986 & ~n14992;
  assign n14994 = n14982 & ~n14993;
  assign n14995 = P2_STATE2_REG_0_ & n14962;
  assign n14996 = P2_EBX_REG_2_ & n14995;
  assign n14997 = n14486 & n14922;
  assign n14998 = P2_REIP_REG_2_ & n14997;
  assign n14999 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_2_;
  assign n15000 = ~n14404 & n14857;
  assign n15001 = n14199 & n14966;
  assign n15002 = n15000 & n15001;
  assign n15003 = P2_STATE2_REG_0_ & ~n14143;
  assign n15004 = n14239 & n15003;
  assign n15005 = n14486 & n15004;
  assign n15006 = n14238 & n14404;
  assign n15007 = P2_STATE2_REG_0_ & n15006;
  assign n15008 = n14199 & n15007;
  assign n15009 = ~n14443 & n14966;
  assign n15010 = n15008 & n15009;
  assign n15011 = P2_STATE2_REG_0_ & ~n14482;
  assign n15012 = n14199 & n15011;
  assign n15013 = n14491 & n15012;
  assign n15014 = ~n15002 & ~n15005;
  assign n15015 = ~n15010 & n15014;
  assign n15016 = ~n15013 & n15015;
  assign n15017 = P2_INSTADDRPOINTER_REG_2_ & ~n15016;
  assign n15018 = ~n14996 & ~n14998;
  assign n15019 = ~n14999 & n15018;
  assign n15020 = ~n15017 & n15019;
  assign n15021 = ~P2_STATE2_REG_0_ & P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n15022 = ~P2_STATE2_REG_1_ & ~n15021;
  assign n15023 = n14199 & n14857;
  assign n15024 = n14482 & n14489;
  assign n15025 = ~n14286 & n14443;
  assign n15026 = ~n14365 & ~n14974;
  assign n15027 = n15025 & n15026;
  assign n15028 = ~n14482 & ~n15027;
  assign n15029 = ~n14325 & ~n14974;
  assign n15030 = n14286 & ~n14443;
  assign n15031 = ~n15029 & ~n15030;
  assign n15032 = ~n14484 & n15031;
  assign n15033 = ~n15024 & ~n15028;
  assign n15034 = n15032 & n15033;
  assign n15035 = n15023 & ~n15034;
  assign n15036 = n14238 & n14550;
  assign n15037 = ~n14325 & n14443;
  assign n15038 = n14365 & ~n14404;
  assign n15039 = ~n14974 & ~n15038;
  assign n15040 = ~n14286 & n15039;
  assign n15041 = n15037 & n15040;
  assign n15042 = n15036 & ~n15041;
  assign n15043 = n14922 & ~n14959;
  assign n15044 = n14325 & n15043;
  assign n15045 = ~n14482 & n14550;
  assign n15046 = n14326 & n14482;
  assign n15047 = n14490 & n15046;
  assign n15048 = n14550 & n15047;
  assign n15049 = ~n14856 & ~n15044;
  assign n15050 = ~n15045 & n15049;
  assign n15051 = ~n15048 & n15050;
  assign n15052 = ~n14365 & n15008;
  assign n15053 = ~n14325 & n14922;
  assign n15054 = ~n14443 & ~n14974;
  assign n15055 = ~n14365 & n14443;
  assign n15056 = n14404 & n15055;
  assign n15057 = ~n14286 & ~n15054;
  assign n15058 = ~n15056 & n15057;
  assign n15059 = ~n15038 & n15058;
  assign n15060 = n15053 & ~n15059;
  assign n15061 = n14243 & n14961;
  assign n15062 = P2_STATE2_REG_0_ & n15061;
  assign n15063 = ~n15052 & ~n15060;
  assign n15064 = ~n15062 & n15063;
  assign n15065 = ~n15035 & ~n15042;
  assign n15066 = n15051 & n15065;
  assign n15067 = n15064 & n15066;
  assign n15068 = P2_INSTQUEUERD_ADDR_REG_2_ & ~n15067;
  assign n15069 = n15022 & ~n15068;
  assign n15070 = ~n15020 & ~n15069;
  assign n15071 = n15020 & n15069;
  assign n15072 = P2_EBX_REG_1_ & n14995;
  assign n15073 = P2_REIP_REG_1_ & n14997;
  assign n15074 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_1_;
  assign n15075 = P2_INSTADDRPOINTER_REG_1_ & ~n15016;
  assign n15076 = ~n15072 & ~n15073;
  assign n15077 = ~n15074 & n15076;
  assign n15078 = ~n15075 & n15077;
  assign n15079 = P2_REIP_REG_0_ & n14997;
  assign n15080 = ~n15023 & ~n15079;
  assign n15081 = ~n15034 & ~n15080;
  assign n15082 = P2_EBX_REG_0_ & n14995;
  assign n15083 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_0_;
  assign n15084 = P2_INSTADDRPOINTER_REG_0_ & ~n15016;
  assign n15085 = ~n15083 & ~n15084;
  assign n15086 = ~P2_STATE2_REG_1_ & ~P2_STATE2_REG_0_;
  assign n15087 = ~n15042 & ~n15086;
  assign n15088 = ~n15045 & n15087;
  assign n15089 = ~n15048 & n15088;
  assign n15090 = n14238 & ~n14974;
  assign n15091 = ~n14959 & n15090;
  assign n15092 = P2_STATE2_REG_0_ & ~n15091;
  assign n15093 = n14325 & ~n14959;
  assign n15094 = ~n14325 & ~n15059;
  assign n15095 = ~n15093 & ~n15094;
  assign n15096 = ~n14199 & n15095;
  assign n15097 = n15092 & ~n15096;
  assign n15098 = ~n15081 & ~n15082;
  assign n15099 = n15085 & n15098;
  assign n15100 = n15089 & n15099;
  assign n15101 = ~n15097 & n15100;
  assign n15102 = P2_INSTQUEUEWR_ADDR_REG_0_ & n15086;
  assign n15103 = n14922 & n14961;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = ~n15042 & ~n15060;
  assign n15106 = ~n15010 & ~n15052;
  assign n15107 = ~n15062 & n15106;
  assign n15108 = ~n15035 & n15104;
  assign n15109 = n15051 & n15108;
  assign n15110 = n15105 & n15109;
  assign n15111 = n15107 & n15110;
  assign n15112 = ~n15010 & n15104;
  assign n15113 = ~P2_INSTQUEUERD_ADDR_REG_0_ & n15112;
  assign n15114 = ~n15111 & ~n15113;
  assign n15115 = ~n15078 & ~n15101;
  assign n15116 = n15114 & n15115;
  assign n15117 = P2_INSTQUEUEWR_ADDR_REG_1_ & n15086;
  assign n15118 = ~n14143 & n14550;
  assign n15119 = n14486 & n15118;
  assign n15120 = ~n14997 & ~n15013;
  assign n15121 = ~n15002 & n15120;
  assign n15122 = ~n15117 & n15121;
  assign n15123 = ~n15119 & n15122;
  assign n15124 = P2_INSTQUEUERD_ADDR_REG_1_ & ~n15067;
  assign n15125 = n15123 & ~n15124;
  assign n15126 = ~n15101 & n15114;
  assign n15127 = n15078 & ~n15126;
  assign n15128 = ~n15125 & ~n15127;
  assign n15129 = ~n15116 & ~n15128;
  assign n15130 = ~n15071 & ~n15129;
  assign n15131 = ~n15070 & ~n15130;
  assign n15132 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n15067;
  assign n15133 = P2_INSTQUEUEWR_ADDR_REG_3_ & n15086;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = P2_EBX_REG_3_ & n14995;
  assign n15136 = P2_REIP_REG_3_ & n14997;
  assign n15137 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_3_;
  assign n15138 = P2_INSTADDRPOINTER_REG_3_ & ~n15016;
  assign n15139 = ~n15135 & ~n15136;
  assign n15140 = ~n15137 & n15139;
  assign n15141 = ~n15138 & n15140;
  assign n15142 = ~n15134 & n15141;
  assign n15143 = n15134 & ~n15141;
  assign n15144 = ~n15142 & ~n15143;
  assign n15145 = n15131 & ~n15144;
  assign n15146 = ~n15131 & n15144;
  assign n15147 = ~n15145 & ~n15146;
  assign n15148 = ~n14959 & ~n15090;
  assign n15149 = n14241 & ~n15148;
  assign n15150 = n14960 & ~n15149;
  assign n15151 = n14199 & ~n14404;
  assign n15152 = ~n14482 & ~n15151;
  assign n15153 = ~n14286 & ~n14365;
  assign n15154 = n14240 & ~n15153;
  assign n15155 = ~n15061 & ~n15154;
  assign n15156 = ~n15150 & ~n15152;
  assign n15157 = n15155 & n15156;
  assign n15158 = n14239 & ~n15040;
  assign n15159 = n14482 & ~n15158;
  assign n15160 = ~n14238 & ~n15059;
  assign n15161 = n15159 & ~n15160;
  assign n15162 = ~n14325 & ~n15161;
  assign n15163 = n14243 & ~n15034;
  assign n15164 = ~n14241 & ~n14443;
  assign n15165 = ~n15163 & ~n15164;
  assign n15166 = n15157 & ~n15162;
  assign n15167 = n15165 & n15166;
  assign n15168 = ~n15047 & n15167;
  assign n15169 = ~n15147 & ~n15168;
  assign n15170 = n14994 & ~n15169;
  assign n15171 = ~n14949 & n14979;
  assign n15172 = n14243 & n14492;
  assign n15173 = n14244 & n14486;
  assign n15174 = ~n15172 & ~n15173;
  assign n15175 = ~n14051 & ~n15174;
  assign n15176 = n14548 & n15175;
  assign n15177 = ~n15171 & ~n15176;
  assign n15178 = n14240 & n14492;
  assign n15179 = n14145 & n15178;
  assign n15180 = ~n14949 & n15179;
  assign n15181 = n14949 & n14978;
  assign n15182 = ~n14974 & n14975;
  assign n15183 = n14486 & n14548;
  assign n15184 = n14145 & n15183;
  assign n15185 = ~n15182 & ~n15184;
  assign n15186 = n14199 & n14491;
  assign n15187 = ~n14482 & ~n15186;
  assign n15188 = n14199 & n14443;
  assign n15189 = ~n14286 & ~n15188;
  assign n15190 = ~n14325 & n15189;
  assign n15191 = ~n14240 & n15190;
  assign n15192 = n14482 & ~n15191;
  assign n15193 = ~n15038 & ~n15056;
  assign n15194 = ~n15158 & n15193;
  assign n15195 = ~n15187 & ~n15192;
  assign n15196 = n15194 & n15195;
  assign n15197 = ~n15180 & ~n15181;
  assign n15198 = n15185 & n15197;
  assign n15199 = n15196 & n15198;
  assign n15200 = n15177 & n15199;
  assign n15201 = ~n15170 & ~n15200;
  assign n15202 = P2_INSTQUEUERD_ADDR_REG_3_ & n15200;
  assign n15203 = ~n15201 & ~n15202;
  assign n15204 = ~n14558 & ~n14968;
  assign n15205 = n14558 & ~n14980;
  assign n15206 = ~n15204 & ~n15205;
  assign n15207 = P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_INSTQUEUERD_ADDR_REG_1_;
  assign n15208 = ~n14192 & ~n15207;
  assign n15209 = ~n14992 & ~n15208;
  assign n15210 = n15206 & ~n15209;
  assign n15211 = n15020 & ~n15069;
  assign n15212 = ~n15020 & n15069;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = n15129 & ~n15213;
  assign n15215 = ~n15129 & n15213;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = ~n15168 & ~n15216;
  assign n15218 = n15210 & ~n15217;
  assign n15219 = ~n15200 & ~n15218;
  assign n15220 = P2_INSTQUEUERD_ADDR_REG_2_ & n15200;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = ~n15203 & ~n15221;
  assign n15223 = P2_INSTQUEUERD_ADDR_REG_4_ & n15200;
  assign n15224 = P2_INSTQUEUERD_ADDR_REG_3_ & P2_INSTQUEUERD_ADDR_REG_1_;
  assign n15225 = P2_INSTQUEUERD_ADDR_REG_2_ & n15224;
  assign n15226 = P2_INSTQUEUERD_ADDR_REG_4_ & ~n14482;
  assign n15227 = n14238 & n15226;
  assign n15228 = n15225 & ~n15227;
  assign n15229 = ~n15225 & n15227;
  assign n15230 = ~n15228 & ~n15229;
  assign n15231 = n15172 & ~n15230;
  assign n15232 = ~n15200 & n15231;
  assign n15233 = ~n15223 & ~n15232;
  assign n15234 = ~n15222 & n15233;
  assign n15235 = ~P2_INSTQUEUEWR_ADDR_REG_4_ & ~n15233;
  assign n15236 = P2_INSTQUEUEWR_ADDR_REG_3_ & n15203;
  assign n15237 = P2_INSTQUEUEWR_ADDR_REG_4_ & n15233;
  assign n15238 = ~P2_INSTQUEUEWR_ADDR_REG_2_ & ~n15221;
  assign n15239 = ~P2_INSTQUEUEWR_ADDR_REG_3_ & ~n15203;
  assign n15240 = ~P2_INSTQUEUERD_ADDR_REG_1_ & ~n14992;
  assign n15241 = n14482 & ~n14555;
  assign n15242 = n14244 & n14959;
  assign n15243 = ~n14286 & ~n14443;
  assign n15244 = n14404 & n15243;
  assign n15245 = n14243 & n15244;
  assign n15246 = ~n15242 & ~n15245;
  assign n15247 = n14365 & ~n15246;
  assign n15248 = n14325 & n15247;
  assign n15249 = n14974 & n15243;
  assign n15250 = ~n14245 & n15249;
  assign n15251 = ~n14325 & n15250;
  assign n15252 = ~n15248 & ~n15251;
  assign n15253 = n15241 & ~n15252;
  assign n15254 = ~n15240 & ~n15253;
  assign n15255 = n15116 & ~n15125;
  assign n15256 = ~n15078 & ~n15126;
  assign n15257 = n15125 & n15256;
  assign n15258 = ~n15255 & ~n15257;
  assign n15259 = n15125 & n15126;
  assign n15260 = ~n15125 & ~n15126;
  assign n15261 = ~n15259 & ~n15260;
  assign n15262 = n15078 & ~n15261;
  assign n15263 = n15258 & ~n15262;
  assign n15264 = ~n15168 & ~n15263;
  assign n15265 = n15254 & ~n15264;
  assign n15266 = ~n15200 & ~n15265;
  assign n15267 = P2_INSTQUEUERD_ADDR_REG_1_ & n15200;
  assign n15268 = ~n15266 & ~n15267;
  assign n15269 = P2_INSTQUEUEWR_ADDR_REG_1_ & n15268;
  assign n15270 = P2_INSTQUEUEWR_ADDR_REG_2_ & n15221;
  assign n15271 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n14992;
  assign n15272 = ~P2_INSTQUEUERD_ADDR_REG_0_ & n14482;
  assign n15273 = ~n15252 & n15272;
  assign n15274 = ~n15271 & ~n15273;
  assign n15275 = ~n15101 & ~n15114;
  assign n15276 = n15101 & n15114;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = ~n15168 & ~n15277;
  assign n15279 = n15274 & ~n15278;
  assign n15280 = ~n15200 & ~n15279;
  assign n15281 = P2_INSTQUEUERD_ADDR_REG_0_ & n15200;
  assign n15282 = ~n15280 & ~n15281;
  assign n15283 = ~P2_INSTQUEUEWR_ADDR_REG_1_ & ~n15268;
  assign n15284 = P2_INSTQUEUEWR_ADDR_REG_0_ & n15282;
  assign n15285 = ~n15283 & n15284;
  assign n15286 = ~n15269 & ~n15270;
  assign n15287 = ~n15285 & n15286;
  assign n15288 = ~n15238 & ~n15239;
  assign n15289 = ~n15287 & n15288;
  assign n15290 = ~n15236 & ~n15237;
  assign n15291 = ~n15289 & n15290;
  assign n15292 = ~n15235 & ~n15291;
  assign n15293 = n14910 & n14920;
  assign n15294 = ~n14902 & ~n15293;
  assign n15295 = n14869 & n14880;
  assign n15296 = n14888 & n15295;
  assign n15297 = ~n15294 & n15296;
  assign n15298 = n14855 & ~n15297;
  assign n15299 = n14239 & n15298;
  assign n15300 = P2_INSTQUEUERD_ADDR_REG_4_ & ~P2_FLUSH_REG;
  assign n15301 = P2_STATE2_REG_1_ & n15300;
  assign n15302 = ~P2_STATE2_REG_1_ & ~n14510;
  assign n15303 = ~n15301 & ~n15302;
  assign n15304 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_31_;
  assign n15305 = P2_PHYADDRPOINTER_REG_1_ & P2_PHYADDRPOINTER_REG_3_;
  assign n15306 = P2_PHYADDRPOINTER_REG_2_ & n15305;
  assign n15307 = P2_PHYADDRPOINTER_REG_4_ & n15306;
  assign n15308 = P2_PHYADDRPOINTER_REG_5_ & n15307;
  assign n15309 = P2_PHYADDRPOINTER_REG_6_ & n15308;
  assign n15310 = P2_PHYADDRPOINTER_REG_7_ & n15309;
  assign n15311 = P2_PHYADDRPOINTER_REG_8_ & n15310;
  assign n15312 = P2_PHYADDRPOINTER_REG_9_ & n15311;
  assign n15313 = P2_PHYADDRPOINTER_REG_10_ & n15312;
  assign n15314 = P2_PHYADDRPOINTER_REG_11_ & n15313;
  assign n15315 = P2_PHYADDRPOINTER_REG_12_ & n15314;
  assign n15316 = P2_PHYADDRPOINTER_REG_13_ & n15315;
  assign n15317 = P2_PHYADDRPOINTER_REG_14_ & n15316;
  assign n15318 = P2_PHYADDRPOINTER_REG_15_ & n15317;
  assign n15319 = P2_PHYADDRPOINTER_REG_16_ & n15318;
  assign n15320 = P2_PHYADDRPOINTER_REG_17_ & n15319;
  assign n15321 = P2_PHYADDRPOINTER_REG_18_ & n15320;
  assign n15322 = P2_PHYADDRPOINTER_REG_19_ & n15321;
  assign n15323 = P2_PHYADDRPOINTER_REG_20_ & n15322;
  assign n15324 = P2_PHYADDRPOINTER_REG_21_ & n15323;
  assign n15325 = P2_PHYADDRPOINTER_REG_22_ & n15324;
  assign n15326 = P2_PHYADDRPOINTER_REG_23_ & n15325;
  assign n15327 = P2_PHYADDRPOINTER_REG_24_ & n15326;
  assign n15328 = P2_PHYADDRPOINTER_REG_25_ & n15327;
  assign n15329 = P2_PHYADDRPOINTER_REG_26_ & n15328;
  assign n15330 = P2_PHYADDRPOINTER_REG_27_ & n15329;
  assign n15331 = P2_PHYADDRPOINTER_REG_28_ & n15330;
  assign n15332 = P2_PHYADDRPOINTER_REG_29_ & n15331;
  assign n15333 = P2_PHYADDRPOINTER_REG_30_ & n15332;
  assign n15334 = ~P2_PHYADDRPOINTER_REG_31_ & n15333;
  assign n15335 = P2_PHYADDRPOINTER_REG_31_ & ~n15333;
  assign n15336 = ~n15334 & ~n15335;
  assign n15337 = ~P2_STATE2_REG_0_ & ~n15336;
  assign n15338 = ~n15304 & ~n15337;
  assign n15339 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_0_;
  assign n15340 = ~P2_STATE2_REG_0_ & P2_PHYADDRPOINTER_REG_0_;
  assign n15341 = ~n15339 & ~n15340;
  assign n15342 = ~n15338 & ~n15341;
  assign n15343 = P2_INSTADDRPOINTER_REG_0_ & n15338;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = P2_FLUSH_REG & n15344;
  assign n15346 = P2_INSTQUEUERD_ADDR_REG_0_ & ~P2_FLUSH_REG;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = P2_STATE2_REG_1_ & n15347;
  assign n15349 = ~P2_STATE2_REG_1_ & ~n14927;
  assign n15350 = ~n15348 & ~n15349;
  assign n15351 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_1_;
  assign n15352 = ~P2_STATE2_REG_0_ & ~P2_PHYADDRPOINTER_REG_1_;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = ~n15341 & n15353;
  assign n15355 = n15341 & ~n15353;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = ~n15338 & ~n15356;
  assign n15358 = P2_INSTADDRPOINTER_REG_1_ & n15338;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = ~n15344 & ~n15359;
  assign n15361 = P2_FLUSH_REG & n15360;
  assign n15362 = P2_INSTQUEUERD_ADDR_REG_2_ & ~P2_FLUSH_REG;
  assign n15363 = ~n15361 & ~n15362;
  assign n15364 = P2_STATE2_REG_1_ & n15363;
  assign n15365 = ~P2_STATE2_REG_1_ & ~n14540;
  assign n15366 = ~n15364 & ~n15365;
  assign n15367 = P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_FLUSH_REG;
  assign n15368 = P2_STATE2_REG_1_ & ~n15367;
  assign n15369 = ~P2_STATE2_REG_1_ & ~n14524;
  assign n15370 = ~n15368 & ~n15369;
  assign n15371 = ~P2_STATE2_REG_1_ & ~n14517;
  assign n15372 = ~n15301 & ~n15371;
  assign n15373 = n15350 & n15366;
  assign n15374 = n15303 & n15373;
  assign n15375 = n15370 & n15374;
  assign n15376 = n15372 & n15375;
  assign n15377 = n15303 & ~n15376;
  assign n15378 = n15370 & n15372;
  assign n15379 = n15303 & n15378;
  assign n15380 = n15366 & n15379;
  assign n15381 = ~n15344 & n15359;
  assign n15382 = P2_FLUSH_REG & n15381;
  assign n15383 = P2_INSTQUEUERD_ADDR_REG_1_ & ~P2_FLUSH_REG;
  assign n15384 = ~n15382 & ~n15383;
  assign n15385 = P2_STATE2_REG_1_ & n15384;
  assign n15386 = ~P2_STATE2_REG_1_ & ~n14533;
  assign n15387 = ~n15385 & ~n15386;
  assign n15388 = n15380 & n15387;
  assign n15389 = n15377 & ~n15388;
  assign n15390 = n14244 & n15389;
  assign n15391 = ~n15299 & ~n15390;
  assign n15392 = n15047 & ~n15391;
  assign n15393 = ~n14979 & ~n15178;
  assign n15394 = n14949 & ~n15393;
  assign n15395 = ~n14949 & n14978;
  assign n15396 = ~n14988 & ~n15172;
  assign n15397 = ~n14548 & ~n15396;
  assign n15398 = n14239 & ~n15298;
  assign n15399 = n14244 & ~n15389;
  assign n15400 = ~n15398 & ~n15399;
  assign n15401 = n15047 & ~n15400;
  assign n15402 = ~n15394 & ~n15395;
  assign n15403 = ~n15397 & n15402;
  assign n15404 = ~n15401 & n15403;
  assign n15405 = ~n14956 & n15234;
  assign n15406 = n15292 & n15405;
  assign n15407 = ~n15392 & n15406;
  assign n15408 = n15404 & n15407;
  assign n15409 = ~P2_STATE2_REG_1_ & n15408;
  assign n15410 = P2_STATE2_REG_0_ & ~n15409;
  assign n15411 = ~P2_STATE2_REG_0_ & ~n14051;
  assign n15412 = P2_STATE2_REG_2_ & ~n15086;
  assign n15413 = ~P2_STATEBS16_REG & ~n14051;
  assign n15414 = ~P2_STATE_REG_0_ & n15413;
  assign n15415 = n15005 & n15414;
  assign n15416 = n15412 & ~n15415;
  assign n15417 = ~n15410 & ~n15411;
  assign n15418 = n15416 & n15417;
  assign n15419 = P2_STATE2_REG_0_ & ~n15418;
  assign n15420 = n14141 & n15419;
  assign n15421 = P2_STATE2_REG_3_ & ~n15419;
  assign n3164 = n15420 | n15421;
  assign n15423 = ~P2_STATE2_REG_0_ & P2_STATEBS16_REG;
  assign n15424 = ~P2_STATE2_REG_2_ & P2_STATE2_REG_0_;
  assign n15425 = ~n14051 & n15424;
  assign n15426 = ~n15423 & ~n15425;
  assign n15427 = P2_STATE2_REG_1_ & ~n15426;
  assign n15428 = P2_STATE2_REG_2_ & ~P2_STATE2_REG_1_;
  assign n15429 = ~n15427 & ~n15428;
  assign n15430 = P2_STATE2_REG_2_ & ~n15419;
  assign n3169 = ~n15429 | n15430;
  assign n15432 = P2_STATE2_REG_0_ & n15428;
  assign n15433 = ~n15418 & n15432;
  assign n15434 = n14051 & n15424;
  assign n15435 = ~n15418 & ~n15434;
  assign n15436 = P2_STATE2_REG_1_ & ~n15435;
  assign n15437 = ~P2_STATE2_REG_3_ & ~P2_STATE2_REG_1_;
  assign n15438 = ~n14051 & n15437;
  assign n15439 = n15419 & n15438;
  assign n15440 = P2_STATE2_REG_1_ & ~P2_STATEBS16_REG;
  assign n15441 = ~P2_STATE2_REG_2_ & n15440;
  assign n15442 = ~P2_STATE2_REG_0_ & n15441;
  assign n15443 = ~n15433 & ~n15436;
  assign n15444 = ~n15439 & n15443;
  assign n3174 = n15442 | ~n15444;
  assign n15446 = ~P2_STATE2_REG_2_ & ~P2_STATE2_REG_1_;
  assign n15447 = P2_STATE2_REG_3_ & ~n14949;
  assign n15448 = n15446 & n15447;
  assign n15449 = ~n15418 & ~n15448;
  assign n15450 = ~P2_STATE2_REG_0_ & n15449;
  assign n15451 = n14141 & n15389;
  assign n15452 = ~n15418 & ~n15451;
  assign n15453 = P2_STATE2_REG_0_ & ~n15452;
  assign n15454 = P2_STATE2_REG_3_ & ~P2_STATE2_REG_1_;
  assign n15455 = n15424 & n15454;
  assign n15456 = ~n15434 & ~n15455;
  assign n15457 = ~n15408 & n15432;
  assign n15458 = n15456 & ~n15457;
  assign n15459 = ~n15450 & ~n15453;
  assign n3179 = ~n15458 | ~n15459;
  assign n15461 = P2_INSTQUEUEWR_ADDR_REG_1_ & P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n15462 = P2_INSTQUEUEWR_ADDR_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n15463 = n15461 & n15462;
  assign n15464 = ~P2_INSTQUEUEWR_ADDR_REG_2_ & n15461;
  assign n15465 = P2_INSTQUEUEWR_ADDR_REG_2_ & ~n15461;
  assign n15466 = ~n15464 & ~n15465;
  assign n15467 = P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n15468 = P2_INSTQUEUEWR_ADDR_REG_3_ & ~n15461;
  assign n15469 = ~P2_INSTQUEUEWR_ADDR_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n15470 = n15461 & n15469;
  assign n15471 = ~n15467 & ~n15468;
  assign n15472 = ~n15470 & n15471;
  assign n15473 = ~n15466 & ~n15472;
  assign n15474 = ~P2_INSTQUEUEWR_ADDR_REG_1_ & P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n15475 = P2_INSTQUEUEWR_ADDR_REG_1_ & ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~P2_INSTQUEUEWR_ADDR_REG_0_ & ~n15476;
  assign n15478 = n15473 & n15477;
  assign n15479 = ~n15463 & ~n15478;
  assign n15480 = ~P2_STATE2_REG_3_ & ~P2_STATE2_REG_2_;
  assign n15481 = ~P2_STATEBS16_REG & n15480;
  assign n15482 = P2_STATE2_REG_0_ & ~n14238;
  assign n15483 = n14404 & n15482;
  assign n15484 = P2_INSTQUEUE_REG_0__1_ & n15483;
  assign n15485 = P2_INSTQUEUE_REG_0__0_ & n15483;
  assign n15486 = ~P2_STATE2_REG_3_ & P2_STATE2_REG_2_;
  assign n15487 = P2_STATE2_REG_0_ & n15486;
  assign n15488 = n14404 & n15487;
  assign n15489 = ~n15485 & n15488;
  assign n15490 = ~n14404 & n15482;
  assign n15491 = ~n15000 & ~n15490;
  assign n15492 = ~P2_STATE2_REG_3_ & n15491;
  assign n15493 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n15492;
  assign n15494 = ~P2_INSTQUEUEWR_ADDR_REG_0_ & n15480;
  assign n15495 = P2_STATE2_REG_2_ & ~P2_STATE2_REG_0_;
  assign n15496 = ~n15277 & n15495;
  assign n15497 = ~n15493 & ~n15494;
  assign n15498 = ~n15496 & n15497;
  assign n15499 = ~n15489 & ~n15498;
  assign n15500 = n15484 & ~n15499;
  assign n15501 = ~n15484 & n15499;
  assign n15502 = ~n15500 & ~n15501;
  assign n15503 = P2_INSTQUEUERD_ADDR_REG_1_ & ~n15492;
  assign n15504 = ~n15476 & n15480;
  assign n15505 = ~n15263 & n15495;
  assign n15506 = ~n15503 & ~n15504;
  assign n15507 = ~n15505 & n15506;
  assign n15508 = ~n15502 & n15507;
  assign n15509 = n15502 & ~n15507;
  assign n15510 = ~n15508 & ~n15509;
  assign n15511 = n15489 & ~n15498;
  assign n15512 = ~n15489 & n15498;
  assign n15513 = ~n15511 & ~n15512;
  assign n15514 = ~n15510 & n15513;
  assign n15515 = n15510 & ~n15513;
  assign n15516 = ~n15514 & ~n15515;
  assign n15517 = n15513 & ~n15516;
  assign n15518 = ~n15510 & ~n15513;
  assign n15519 = P2_INSTQUEUE_REG_0__2_ & n15483;
  assign n15520 = P2_INSTQUEUERD_ADDR_REG_2_ & ~n15492;
  assign n15521 = ~n15466 & n15480;
  assign n15522 = ~n15216 & n15495;
  assign n15523 = ~n15520 & ~n15521;
  assign n15524 = ~n15522 & n15523;
  assign n15525 = ~n15519 & n15524;
  assign n15526 = n15484 & n15499;
  assign n15527 = n15507 & ~n15526;
  assign n15528 = n15519 & ~n15524;
  assign n15529 = ~n15484 & ~n15499;
  assign n15530 = ~n15528 & ~n15529;
  assign n15531 = ~n15525 & ~n15527;
  assign n15532 = n15530 & n15531;
  assign n15533 = ~n15519 & ~n15524;
  assign n15534 = n15519 & n15524;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = ~n15526 & n15535;
  assign n15537 = ~n15507 & ~n15529;
  assign n15538 = n15536 & ~n15537;
  assign n15539 = ~n15532 & ~n15538;
  assign n15540 = n15518 & ~n15539;
  assign n15541 = ~n15518 & n15539;
  assign n15542 = ~n15540 & ~n15541;
  assign n15543 = ~n15527 & ~n15529;
  assign n15544 = ~n15525 & n15543;
  assign n15545 = ~n15528 & ~n15544;
  assign n15546 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n15492;
  assign n15547 = ~n15472 & n15480;
  assign n15548 = ~n15147 & n15495;
  assign n15549 = ~n15546 & ~n15547;
  assign n15550 = ~n15548 & n15549;
  assign n15551 = P2_INSTQUEUE_REG_0__3_ & n15483;
  assign n15552 = ~n15550 & ~n15551;
  assign n15553 = n15550 & n15551;
  assign n15554 = ~n15552 & ~n15553;
  assign n15555 = n15545 & ~n15554;
  assign n15556 = ~n15545 & n15554;
  assign n15557 = ~n15555 & ~n15556;
  assign n15558 = ~n15539 & ~n15557;
  assign n15559 = ~n15518 & ~n15557;
  assign n15560 = n15539 & n15557;
  assign n15561 = n15518 & n15560;
  assign n15562 = ~n15558 & ~n15559;
  assign n15563 = ~n15561 & n15562;
  assign n15564 = ~n15542 & ~n15563;
  assign n15565 = n15517 & n15564;
  assign n15566 = n15539 & ~n15557;
  assign n15567 = n15518 & n15566;
  assign n15568 = ~n15565 & ~n15567;
  assign n15569 = P2_STATEBS16_REG & n15480;
  assign n15570 = ~P2_STATE2_REG_2_ & P2_STATE2_REG_1_;
  assign n15571 = ~n15428 & ~n15570;
  assign n15572 = ~n15447 & n15571;
  assign n15573 = ~P2_STATE2_REG_0_ & ~n15572;
  assign n15574 = n15569 & n15573;
  assign n15575 = n15568 & n15574;
  assign n15576 = ~n15481 & ~n15575;
  assign n15577 = n15479 & ~n15576;
  assign n15578 = ~n15147 & ~n15216;
  assign n15579 = ~n15263 & ~n15277;
  assign n15580 = n15578 & n15579;
  assign n15581 = ~n15463 & ~n15580;
  assign n15582 = P2_STATE2_REG_2_ & n15581;
  assign n15583 = P2_STATE2_REG_3_ & ~n15463;
  assign n15584 = ~n15582 & ~n15583;
  assign n15585 = n15573 & n15584;
  assign n15586 = ~n15577 & n15585;
  assign n15587 = P2_INSTQUEUE_REG_15__7_ & ~n15586;
  assign n15588 = BUF1_REG_7_ & n4541;
  assign n15589 = BUF2_REG_7_ & ~n4541;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = n15573 & ~n15590;
  assign n15592 = P2_STATE2_REG_2_ & ~n15581;
  assign n15593 = n15568 & n15569;
  assign n15594 = ~n15481 & ~n15593;
  assign n15595 = ~n15479 & ~n15594;
  assign n15596 = ~n15592 & ~n15595;
  assign n15597 = n15591 & ~n15596;
  assign n15598 = BUF1_REG_23_ & n4541;
  assign n15599 = BUF2_REG_23_ & ~n4541;
  assign n15600 = ~n15598 & ~n15599;
  assign n15601 = n15574 & ~n15600;
  assign n15602 = n15567 & n15601;
  assign n15603 = P2_STATE2_REG_3_ & n15573;
  assign n15604 = ~n14286 & n15603;
  assign n15605 = n15463 & n15604;
  assign n15606 = BUF1_REG_31_ & n4541;
  assign n15607 = BUF2_REG_31_ & ~n4541;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = n15574 & ~n15608;
  assign n15610 = n15565 & n15609;
  assign n15611 = ~n15602 & ~n15605;
  assign n15612 = ~n15610 & n15611;
  assign n15613 = ~n15587 & ~n15597;
  assign n3184 = ~n15612 | ~n15613;
  assign n15615 = P2_INSTQUEUE_REG_15__6_ & ~n15586;
  assign n15616 = BUF1_REG_6_ & n4541;
  assign n15617 = BUF2_REG_6_ & ~n4541;
  assign n15618 = ~n15616 & ~n15617;
  assign n15619 = n15573 & ~n15618;
  assign n15620 = ~n15596 & n15619;
  assign n15621 = BUF1_REG_22_ & n4541;
  assign n15622 = BUF2_REG_22_ & ~n4541;
  assign n15623 = ~n15621 & ~n15622;
  assign n15624 = n15574 & ~n15623;
  assign n15625 = n15567 & n15624;
  assign n15626 = ~n14404 & n15603;
  assign n15627 = n15463 & n15626;
  assign n15628 = BUF1_REG_30_ & n4541;
  assign n15629 = BUF2_REG_30_ & ~n4541;
  assign n15630 = ~n15628 & ~n15629;
  assign n15631 = n15574 & ~n15630;
  assign n15632 = n15565 & n15631;
  assign n15633 = ~n15625 & ~n15627;
  assign n15634 = ~n15632 & n15633;
  assign n15635 = ~n15615 & ~n15620;
  assign n3189 = ~n15634 | ~n15635;
  assign n15637 = P2_INSTQUEUE_REG_15__5_ & ~n15586;
  assign n15638 = BUF1_REG_5_ & n4541;
  assign n15639 = BUF2_REG_5_ & ~n4541;
  assign n15640 = ~n15638 & ~n15639;
  assign n15641 = n15573 & ~n15640;
  assign n15642 = ~n15596 & n15641;
  assign n15643 = BUF1_REG_21_ & n4541;
  assign n15644 = BUF2_REG_21_ & ~n4541;
  assign n15645 = ~n15643 & ~n15644;
  assign n15646 = n15574 & ~n15645;
  assign n15647 = n15567 & n15646;
  assign n15648 = ~n14365 & n15603;
  assign n15649 = n15463 & n15648;
  assign n15650 = BUF1_REG_29_ & n4541;
  assign n15651 = BUF2_REG_29_ & ~n4541;
  assign n15652 = ~n15650 & ~n15651;
  assign n15653 = n15574 & ~n15652;
  assign n15654 = n15565 & n15653;
  assign n15655 = ~n15647 & ~n15649;
  assign n15656 = ~n15654 & n15655;
  assign n15657 = ~n15637 & ~n15642;
  assign n3194 = ~n15656 | ~n15657;
  assign n15659 = P2_INSTQUEUE_REG_15__4_ & ~n15586;
  assign n15660 = BUF1_REG_4_ & n4541;
  assign n15661 = BUF2_REG_4_ & ~n4541;
  assign n15662 = ~n15660 & ~n15661;
  assign n15663 = n15573 & ~n15662;
  assign n15664 = ~n15596 & n15663;
  assign n15665 = BUF1_REG_20_ & n4541;
  assign n15666 = BUF2_REG_20_ & ~n4541;
  assign n15667 = ~n15665 & ~n15666;
  assign n15668 = n15574 & ~n15667;
  assign n15669 = n15567 & n15668;
  assign n15670 = ~n14443 & n15603;
  assign n15671 = n15463 & n15670;
  assign n15672 = BUF1_REG_28_ & n4541;
  assign n15673 = BUF2_REG_28_ & ~n4541;
  assign n15674 = ~n15672 & ~n15673;
  assign n15675 = n15574 & ~n15674;
  assign n15676 = n15565 & n15675;
  assign n15677 = ~n15669 & ~n15671;
  assign n15678 = ~n15676 & n15677;
  assign n15679 = ~n15659 & ~n15664;
  assign n3199 = ~n15678 | ~n15679;
  assign n15681 = P2_INSTQUEUE_REG_15__3_ & ~n15586;
  assign n15682 = BUF1_REG_3_ & n4541;
  assign n15683 = BUF2_REG_3_ & ~n4541;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = n15573 & ~n15684;
  assign n15686 = ~n15596 & n15685;
  assign n15687 = BUF1_REG_19_ & n4541;
  assign n15688 = BUF2_REG_19_ & ~n4541;
  assign n15689 = ~n15687 & ~n15688;
  assign n15690 = n15574 & ~n15689;
  assign n15691 = n15567 & n15690;
  assign n15692 = ~n14325 & n15603;
  assign n15693 = n15463 & n15692;
  assign n15694 = BUF1_REG_27_ & n4541;
  assign n15695 = BUF2_REG_27_ & ~n4541;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = n15574 & ~n15696;
  assign n15698 = n15565 & n15697;
  assign n15699 = ~n15691 & ~n15693;
  assign n15700 = ~n15698 & n15699;
  assign n15701 = ~n15681 & ~n15686;
  assign n3204 = ~n15700 | ~n15701;
  assign n15703 = P2_INSTQUEUE_REG_15__2_ & ~n15586;
  assign n15704 = BUF1_REG_2_ & n4541;
  assign n15705 = BUF2_REG_2_ & ~n4541;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = n15573 & ~n15706;
  assign n15708 = ~n15596 & n15707;
  assign n15709 = BUF1_REG_18_ & n4541;
  assign n15710 = BUF2_REG_18_ & ~n4541;
  assign n15711 = ~n15709 & ~n15710;
  assign n15712 = n15574 & ~n15711;
  assign n15713 = n15567 & n15712;
  assign n15714 = ~n14482 & n15603;
  assign n15715 = n15463 & n15714;
  assign n15716 = BUF1_REG_26_ & n4541;
  assign n15717 = BUF2_REG_26_ & ~n4541;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = n15574 & ~n15718;
  assign n15720 = n15565 & n15719;
  assign n15721 = ~n15713 & ~n15715;
  assign n15722 = ~n15720 & n15721;
  assign n15723 = ~n15703 & ~n15708;
  assign n3209 = ~n15722 | ~n15723;
  assign n15725 = P2_INSTQUEUE_REG_15__1_ & ~n15586;
  assign n15726 = BUF1_REG_1_ & n4541;
  assign n15727 = BUF2_REG_1_ & ~n4541;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = n15573 & ~n15728;
  assign n15730 = ~n15596 & n15729;
  assign n15731 = BUF1_REG_17_ & n4541;
  assign n15732 = BUF2_REG_17_ & ~n4541;
  assign n15733 = ~n15731 & ~n15732;
  assign n15734 = n15574 & ~n15733;
  assign n15735 = n15567 & n15734;
  assign n15736 = ~n14238 & n15603;
  assign n15737 = n15463 & n15736;
  assign n15738 = BUF1_REG_25_ & n4541;
  assign n15739 = BUF2_REG_25_ & ~n4541;
  assign n15740 = ~n15738 & ~n15739;
  assign n15741 = n15574 & ~n15740;
  assign n15742 = n15565 & n15741;
  assign n15743 = ~n15735 & ~n15737;
  assign n15744 = ~n15742 & n15743;
  assign n15745 = ~n15725 & ~n15730;
  assign n3214 = ~n15744 | ~n15745;
  assign n15747 = P2_INSTQUEUE_REG_15__0_ & ~n15586;
  assign n15748 = BUF1_REG_0_ & n4541;
  assign n15749 = BUF2_REG_0_ & ~n4541;
  assign n15750 = ~n15748 & ~n15749;
  assign n15751 = n15573 & ~n15750;
  assign n15752 = ~n15596 & n15751;
  assign n15753 = BUF1_REG_16_ & n4541;
  assign n15754 = BUF2_REG_16_ & ~n4541;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = n15574 & ~n15755;
  assign n15757 = n15567 & n15756;
  assign n15758 = ~n14199 & n15603;
  assign n15759 = n15463 & n15758;
  assign n15760 = BUF1_REG_24_ & n4541;
  assign n15761 = BUF2_REG_24_ & ~n4541;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = n15574 & ~n15762;
  assign n15764 = n15565 & n15763;
  assign n15765 = ~n15757 & ~n15759;
  assign n15766 = ~n15764 & n15765;
  assign n15767 = ~n15747 & ~n15752;
  assign n3219 = ~n15766 | ~n15767;
  assign n15769 = ~n15513 & ~n15516;
  assign n15770 = n15564 & n15769;
  assign n15771 = n15514 & n15566;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = n15574 & n15772;
  assign n15774 = ~n15481 & ~n15773;
  assign n15775 = n15473 & ~n15476;
  assign n15776 = ~n15774 & ~n15775;
  assign n15777 = ~n15263 & n15277;
  assign n15778 = n15578 & n15777;
  assign n15779 = n15462 & n15475;
  assign n15780 = ~n15778 & ~n15779;
  assign n15781 = P2_STATE2_REG_2_ & n15780;
  assign n15782 = P2_STATE2_REG_3_ & ~n15779;
  assign n15783 = ~n15781 & ~n15782;
  assign n15784 = n15573 & n15783;
  assign n15785 = ~n15776 & n15784;
  assign n15786 = P2_INSTQUEUE_REG_14__7_ & ~n15785;
  assign n15787 = P2_STATE2_REG_2_ & ~n15780;
  assign n15788 = n15569 & n15772;
  assign n15789 = ~n15481 & ~n15788;
  assign n15790 = n15775 & ~n15789;
  assign n15791 = ~n15787 & ~n15790;
  assign n15792 = n15591 & ~n15791;
  assign n15793 = n15601 & n15771;
  assign n15794 = n15604 & n15779;
  assign n15795 = n15609 & n15770;
  assign n15796 = ~n15793 & ~n15794;
  assign n15797 = ~n15795 & n15796;
  assign n15798 = ~n15786 & ~n15792;
  assign n3224 = ~n15797 | ~n15798;
  assign n15800 = P2_INSTQUEUE_REG_14__6_ & ~n15785;
  assign n15801 = n15619 & ~n15791;
  assign n15802 = n15624 & n15771;
  assign n15803 = n15626 & n15779;
  assign n15804 = n15631 & n15770;
  assign n15805 = ~n15802 & ~n15803;
  assign n15806 = ~n15804 & n15805;
  assign n15807 = ~n15800 & ~n15801;
  assign n3229 = ~n15806 | ~n15807;
  assign n15809 = P2_INSTQUEUE_REG_14__5_ & ~n15785;
  assign n15810 = n15641 & ~n15791;
  assign n15811 = n15646 & n15771;
  assign n15812 = n15648 & n15779;
  assign n15813 = n15653 & n15770;
  assign n15814 = ~n15811 & ~n15812;
  assign n15815 = ~n15813 & n15814;
  assign n15816 = ~n15809 & ~n15810;
  assign n3234 = ~n15815 | ~n15816;
  assign n15818 = P2_INSTQUEUE_REG_14__4_ & ~n15785;
  assign n15819 = n15663 & ~n15791;
  assign n15820 = n15668 & n15771;
  assign n15821 = n15670 & n15779;
  assign n15822 = n15675 & n15770;
  assign n15823 = ~n15820 & ~n15821;
  assign n15824 = ~n15822 & n15823;
  assign n15825 = ~n15818 & ~n15819;
  assign n3239 = ~n15824 | ~n15825;
  assign n15827 = P2_INSTQUEUE_REG_14__3_ & ~n15785;
  assign n15828 = n15685 & ~n15791;
  assign n15829 = n15690 & n15771;
  assign n15830 = n15692 & n15779;
  assign n15831 = n15697 & n15770;
  assign n15832 = ~n15829 & ~n15830;
  assign n15833 = ~n15831 & n15832;
  assign n15834 = ~n15827 & ~n15828;
  assign n3244 = ~n15833 | ~n15834;
  assign n15836 = P2_INSTQUEUE_REG_14__2_ & ~n15785;
  assign n15837 = n15707 & ~n15791;
  assign n15838 = n15712 & n15771;
  assign n15839 = n15714 & n15779;
  assign n15840 = n15719 & n15770;
  assign n15841 = ~n15838 & ~n15839;
  assign n15842 = ~n15840 & n15841;
  assign n15843 = ~n15836 & ~n15837;
  assign n3249 = ~n15842 | ~n15843;
  assign n15845 = P2_INSTQUEUE_REG_14__1_ & ~n15785;
  assign n15846 = n15729 & ~n15791;
  assign n15847 = n15734 & n15771;
  assign n15848 = n15736 & n15779;
  assign n15849 = n15741 & n15770;
  assign n15850 = ~n15847 & ~n15848;
  assign n15851 = ~n15849 & n15850;
  assign n15852 = ~n15845 & ~n15846;
  assign n3254 = ~n15851 | ~n15852;
  assign n15854 = P2_INSTQUEUE_REG_14__0_ & ~n15785;
  assign n15855 = n15751 & ~n15791;
  assign n15856 = n15756 & n15771;
  assign n15857 = n15758 & n15779;
  assign n15858 = n15763 & n15770;
  assign n15859 = ~n15856 & ~n15857;
  assign n15860 = ~n15858 & n15859;
  assign n15861 = ~n15854 & ~n15855;
  assign n3259 = ~n15860 | ~n15861;
  assign n15863 = n15462 & n15474;
  assign n15864 = ~P2_INSTQUEUEWR_ADDR_REG_0_ & n15476;
  assign n15865 = n15473 & n15864;
  assign n15866 = ~n15863 & ~n15865;
  assign n15867 = n15513 & n15516;
  assign n15868 = n15564 & n15867;
  assign n15869 = n15515 & n15566;
  assign n15870 = ~n15868 & ~n15869;
  assign n15871 = n15574 & n15870;
  assign n15872 = ~n15481 & ~n15871;
  assign n15873 = n15866 & ~n15872;
  assign n15874 = n15263 & ~n15277;
  assign n15875 = n15578 & n15874;
  assign n15876 = ~n15863 & ~n15875;
  assign n15877 = P2_STATE2_REG_2_ & n15876;
  assign n15878 = P2_STATE2_REG_3_ & ~n15863;
  assign n15879 = ~n15877 & ~n15878;
  assign n15880 = n15573 & n15879;
  assign n15881 = ~n15873 & n15880;
  assign n15882 = P2_INSTQUEUE_REG_13__7_ & ~n15881;
  assign n15883 = P2_STATE2_REG_2_ & ~n15876;
  assign n15884 = n15569 & n15870;
  assign n15885 = ~n15481 & ~n15884;
  assign n15886 = ~n15866 & ~n15885;
  assign n15887 = ~n15883 & ~n15886;
  assign n15888 = n15591 & ~n15887;
  assign n15889 = n15601 & n15869;
  assign n15890 = n15604 & n15863;
  assign n15891 = n15609 & n15868;
  assign n15892 = ~n15889 & ~n15890;
  assign n15893 = ~n15891 & n15892;
  assign n15894 = ~n15882 & ~n15888;
  assign n3264 = ~n15893 | ~n15894;
  assign n15896 = P2_INSTQUEUE_REG_13__6_ & ~n15881;
  assign n15897 = n15619 & ~n15887;
  assign n15898 = n15624 & n15869;
  assign n15899 = n15626 & n15863;
  assign n15900 = n15631 & n15868;
  assign n15901 = ~n15898 & ~n15899;
  assign n15902 = ~n15900 & n15901;
  assign n15903 = ~n15896 & ~n15897;
  assign n3269 = ~n15902 | ~n15903;
  assign n15905 = P2_INSTQUEUE_REG_13__5_ & ~n15881;
  assign n15906 = n15641 & ~n15887;
  assign n15907 = n15646 & n15869;
  assign n15908 = n15648 & n15863;
  assign n15909 = n15653 & n15868;
  assign n15910 = ~n15907 & ~n15908;
  assign n15911 = ~n15909 & n15910;
  assign n15912 = ~n15905 & ~n15906;
  assign n3274 = ~n15911 | ~n15912;
  assign n15914 = P2_INSTQUEUE_REG_13__4_ & ~n15881;
  assign n15915 = n15663 & ~n15887;
  assign n15916 = n15668 & n15869;
  assign n15917 = n15670 & n15863;
  assign n15918 = n15675 & n15868;
  assign n15919 = ~n15916 & ~n15917;
  assign n15920 = ~n15918 & n15919;
  assign n15921 = ~n15914 & ~n15915;
  assign n3279 = ~n15920 | ~n15921;
  assign n15923 = P2_INSTQUEUE_REG_13__3_ & ~n15881;
  assign n15924 = n15685 & ~n15887;
  assign n15925 = n15690 & n15869;
  assign n15926 = n15692 & n15863;
  assign n15927 = n15697 & n15868;
  assign n15928 = ~n15925 & ~n15926;
  assign n15929 = ~n15927 & n15928;
  assign n15930 = ~n15923 & ~n15924;
  assign n3284 = ~n15929 | ~n15930;
  assign n15932 = P2_INSTQUEUE_REG_13__2_ & ~n15881;
  assign n15933 = n15707 & ~n15887;
  assign n15934 = n15712 & n15869;
  assign n15935 = n15714 & n15863;
  assign n15936 = n15719 & n15868;
  assign n15937 = ~n15934 & ~n15935;
  assign n15938 = ~n15936 & n15937;
  assign n15939 = ~n15932 & ~n15933;
  assign n3289 = ~n15938 | ~n15939;
  assign n15941 = P2_INSTQUEUE_REG_13__1_ & ~n15881;
  assign n15942 = n15729 & ~n15887;
  assign n15943 = n15734 & n15869;
  assign n15944 = n15736 & n15863;
  assign n15945 = n15741 & n15868;
  assign n15946 = ~n15943 & ~n15944;
  assign n15947 = ~n15945 & n15946;
  assign n15948 = ~n15941 & ~n15942;
  assign n3294 = ~n15947 | ~n15948;
  assign n15950 = P2_INSTQUEUE_REG_13__0_ & ~n15881;
  assign n15951 = n15751 & ~n15887;
  assign n15952 = n15756 & n15869;
  assign n15953 = n15758 & n15863;
  assign n15954 = n15763 & n15868;
  assign n15955 = ~n15952 & ~n15953;
  assign n15956 = ~n15954 & n15955;
  assign n15957 = ~n15950 & ~n15951;
  assign n3299 = ~n15956 | ~n15957;
  assign n15959 = ~n15513 & n15516;
  assign n15960 = n15564 & n15959;
  assign n15961 = n15510 & n15513;
  assign n15962 = n15566 & n15961;
  assign n15963 = ~n15960 & ~n15962;
  assign n15964 = n15574 & n15963;
  assign n15965 = ~n15481 & ~n15964;
  assign n15966 = n15473 & n15476;
  assign n15967 = ~n15965 & ~n15966;
  assign n15968 = n15263 & n15277;
  assign n15969 = n15578 & n15968;
  assign n15970 = ~P2_INSTQUEUEWR_ADDR_REG_1_ & ~P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n15971 = n15462 & n15970;
  assign n15972 = ~n15969 & ~n15971;
  assign n15973 = P2_STATE2_REG_2_ & n15972;
  assign n15974 = P2_STATE2_REG_3_ & ~n15971;
  assign n15975 = ~n15973 & ~n15974;
  assign n15976 = n15573 & n15975;
  assign n15977 = ~n15967 & n15976;
  assign n15978 = P2_INSTQUEUE_REG_12__7_ & ~n15977;
  assign n15979 = P2_STATE2_REG_2_ & ~n15972;
  assign n15980 = n15569 & n15963;
  assign n15981 = ~n15481 & ~n15980;
  assign n15982 = n15966 & ~n15981;
  assign n15983 = ~n15979 & ~n15982;
  assign n15984 = n15591 & ~n15983;
  assign n15985 = n15601 & n15962;
  assign n15986 = n15604 & n15971;
  assign n15987 = n15609 & n15960;
  assign n15988 = ~n15985 & ~n15986;
  assign n15989 = ~n15987 & n15988;
  assign n15990 = ~n15978 & ~n15984;
  assign n3304 = ~n15989 | ~n15990;
  assign n15992 = P2_INSTQUEUE_REG_12__6_ & ~n15977;
  assign n15993 = n15619 & ~n15983;
  assign n15994 = n15624 & n15962;
  assign n15995 = n15626 & n15971;
  assign n15996 = n15631 & n15960;
  assign n15997 = ~n15994 & ~n15995;
  assign n15998 = ~n15996 & n15997;
  assign n15999 = ~n15992 & ~n15993;
  assign n3309 = ~n15998 | ~n15999;
  assign n16001 = P2_INSTQUEUE_REG_12__5_ & ~n15977;
  assign n16002 = n15641 & ~n15983;
  assign n16003 = n15646 & n15962;
  assign n16004 = n15648 & n15971;
  assign n16005 = n15653 & n15960;
  assign n16006 = ~n16003 & ~n16004;
  assign n16007 = ~n16005 & n16006;
  assign n16008 = ~n16001 & ~n16002;
  assign n3314 = ~n16007 | ~n16008;
  assign n16010 = P2_INSTQUEUE_REG_12__4_ & ~n15977;
  assign n16011 = n15663 & ~n15983;
  assign n16012 = n15668 & n15962;
  assign n16013 = n15670 & n15971;
  assign n16014 = n15675 & n15960;
  assign n16015 = ~n16012 & ~n16013;
  assign n16016 = ~n16014 & n16015;
  assign n16017 = ~n16010 & ~n16011;
  assign n3319 = ~n16016 | ~n16017;
  assign n16019 = P2_INSTQUEUE_REG_12__3_ & ~n15977;
  assign n16020 = n15685 & ~n15983;
  assign n16021 = n15690 & n15962;
  assign n16022 = n15692 & n15971;
  assign n16023 = n15697 & n15960;
  assign n16024 = ~n16021 & ~n16022;
  assign n16025 = ~n16023 & n16024;
  assign n16026 = ~n16019 & ~n16020;
  assign n3324 = ~n16025 | ~n16026;
  assign n16028 = P2_INSTQUEUE_REG_12__2_ & ~n15977;
  assign n16029 = n15707 & ~n15983;
  assign n16030 = n15712 & n15962;
  assign n16031 = n15714 & n15971;
  assign n16032 = n15719 & n15960;
  assign n16033 = ~n16030 & ~n16031;
  assign n16034 = ~n16032 & n16033;
  assign n16035 = ~n16028 & ~n16029;
  assign n3329 = ~n16034 | ~n16035;
  assign n16037 = P2_INSTQUEUE_REG_12__1_ & ~n15977;
  assign n16038 = n15729 & ~n15983;
  assign n16039 = n15734 & n15962;
  assign n16040 = n15736 & n15971;
  assign n16041 = n15741 & n15960;
  assign n16042 = ~n16039 & ~n16040;
  assign n16043 = ~n16041 & n16042;
  assign n16044 = ~n16037 & ~n16038;
  assign n3334 = ~n16043 | ~n16044;
  assign n16046 = P2_INSTQUEUE_REG_12__0_ & ~n15977;
  assign n16047 = n15751 & ~n15983;
  assign n16048 = n15756 & n15962;
  assign n16049 = n15758 & n15971;
  assign n16050 = n15763 & n15960;
  assign n16051 = ~n16048 & ~n16049;
  assign n16052 = ~n16050 & n16051;
  assign n16053 = ~n16046 & ~n16047;
  assign n3339 = ~n16052 | ~n16053;
  assign n16055 = n15461 & n15467;
  assign n16056 = n15466 & ~n15472;
  assign n16057 = n15477 & n16056;
  assign n16058 = ~n16055 & ~n16057;
  assign n16059 = n15542 & ~n15563;
  assign n16060 = n15517 & n16059;
  assign n16061 = n15518 & n15558;
  assign n16062 = ~n16060 & ~n16061;
  assign n16063 = n15574 & n16062;
  assign n16064 = ~n15481 & ~n16063;
  assign n16065 = n16058 & ~n16064;
  assign n16066 = ~n15147 & n15216;
  assign n16067 = n15579 & n16066;
  assign n16068 = ~n16055 & ~n16067;
  assign n16069 = P2_STATE2_REG_2_ & n16068;
  assign n16070 = P2_STATE2_REG_3_ & ~n16055;
  assign n16071 = ~n16069 & ~n16070;
  assign n16072 = n15573 & n16071;
  assign n16073 = ~n16065 & n16072;
  assign n16074 = P2_INSTQUEUE_REG_11__7_ & ~n16073;
  assign n16075 = P2_STATE2_REG_2_ & ~n16068;
  assign n16076 = n15569 & n16062;
  assign n16077 = ~n15481 & ~n16076;
  assign n16078 = ~n16058 & ~n16077;
  assign n16079 = ~n16075 & ~n16078;
  assign n16080 = n15591 & ~n16079;
  assign n16081 = n15601 & n16061;
  assign n16082 = n15604 & n16055;
  assign n16083 = n15609 & n16060;
  assign n16084 = ~n16081 & ~n16082;
  assign n16085 = ~n16083 & n16084;
  assign n16086 = ~n16074 & ~n16080;
  assign n3344 = ~n16085 | ~n16086;
  assign n16088 = P2_INSTQUEUE_REG_11__6_ & ~n16073;
  assign n16089 = n15619 & ~n16079;
  assign n16090 = n15624 & n16061;
  assign n16091 = n15626 & n16055;
  assign n16092 = n15631 & n16060;
  assign n16093 = ~n16090 & ~n16091;
  assign n16094 = ~n16092 & n16093;
  assign n16095 = ~n16088 & ~n16089;
  assign n3349 = ~n16094 | ~n16095;
  assign n16097 = P2_INSTQUEUE_REG_11__5_ & ~n16073;
  assign n16098 = n15641 & ~n16079;
  assign n16099 = n15646 & n16061;
  assign n16100 = n15648 & n16055;
  assign n16101 = n15653 & n16060;
  assign n16102 = ~n16099 & ~n16100;
  assign n16103 = ~n16101 & n16102;
  assign n16104 = ~n16097 & ~n16098;
  assign n3354 = ~n16103 | ~n16104;
  assign n16106 = P2_INSTQUEUE_REG_11__4_ & ~n16073;
  assign n16107 = n15663 & ~n16079;
  assign n16108 = n15668 & n16061;
  assign n16109 = n15670 & n16055;
  assign n16110 = n15675 & n16060;
  assign n16111 = ~n16108 & ~n16109;
  assign n16112 = ~n16110 & n16111;
  assign n16113 = ~n16106 & ~n16107;
  assign n3359 = ~n16112 | ~n16113;
  assign n16115 = P2_INSTQUEUE_REG_11__3_ & ~n16073;
  assign n16116 = n15685 & ~n16079;
  assign n16117 = n15690 & n16061;
  assign n16118 = n15692 & n16055;
  assign n16119 = n15697 & n16060;
  assign n16120 = ~n16117 & ~n16118;
  assign n16121 = ~n16119 & n16120;
  assign n16122 = ~n16115 & ~n16116;
  assign n3364 = ~n16121 | ~n16122;
  assign n16124 = P2_INSTQUEUE_REG_11__2_ & ~n16073;
  assign n16125 = n15707 & ~n16079;
  assign n16126 = n15712 & n16061;
  assign n16127 = n15714 & n16055;
  assign n16128 = n15719 & n16060;
  assign n16129 = ~n16126 & ~n16127;
  assign n16130 = ~n16128 & n16129;
  assign n16131 = ~n16124 & ~n16125;
  assign n3369 = ~n16130 | ~n16131;
  assign n16133 = P2_INSTQUEUE_REG_11__1_ & ~n16073;
  assign n16134 = n15729 & ~n16079;
  assign n16135 = n15734 & n16061;
  assign n16136 = n15736 & n16055;
  assign n16137 = n15741 & n16060;
  assign n16138 = ~n16135 & ~n16136;
  assign n16139 = ~n16137 & n16138;
  assign n16140 = ~n16133 & ~n16134;
  assign n3374 = ~n16139 | ~n16140;
  assign n16142 = P2_INSTQUEUE_REG_11__0_ & ~n16073;
  assign n16143 = n15751 & ~n16079;
  assign n16144 = n15756 & n16061;
  assign n16145 = n15758 & n16055;
  assign n16146 = n15763 & n16060;
  assign n16147 = ~n16144 & ~n16145;
  assign n16148 = ~n16146 & n16147;
  assign n16149 = ~n16142 & ~n16143;
  assign n3379 = ~n16148 | ~n16149;
  assign n16151 = n15769 & n16059;
  assign n16152 = n15514 & n15558;
  assign n16153 = ~n16151 & ~n16152;
  assign n16154 = n15574 & n16153;
  assign n16155 = ~n15481 & ~n16154;
  assign n16156 = ~n15476 & n16056;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = n15777 & n16066;
  assign n16159 = n15467 & n15475;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = P2_STATE2_REG_2_ & n16160;
  assign n16162 = P2_STATE2_REG_3_ & ~n16159;
  assign n16163 = ~n16161 & ~n16162;
  assign n16164 = n15573 & n16163;
  assign n16165 = ~n16157 & n16164;
  assign n16166 = P2_INSTQUEUE_REG_10__7_ & ~n16165;
  assign n16167 = P2_STATE2_REG_2_ & ~n16160;
  assign n16168 = n15569 & n16153;
  assign n16169 = ~n15481 & ~n16168;
  assign n16170 = n16156 & ~n16169;
  assign n16171 = ~n16167 & ~n16170;
  assign n16172 = n15591 & ~n16171;
  assign n16173 = n15601 & n16152;
  assign n16174 = n15604 & n16159;
  assign n16175 = n15609 & n16151;
  assign n16176 = ~n16173 & ~n16174;
  assign n16177 = ~n16175 & n16176;
  assign n16178 = ~n16166 & ~n16172;
  assign n3384 = ~n16177 | ~n16178;
  assign n16180 = P2_INSTQUEUE_REG_10__6_ & ~n16165;
  assign n16181 = n15619 & ~n16171;
  assign n16182 = n15624 & n16152;
  assign n16183 = n15626 & n16159;
  assign n16184 = n15631 & n16151;
  assign n16185 = ~n16182 & ~n16183;
  assign n16186 = ~n16184 & n16185;
  assign n16187 = ~n16180 & ~n16181;
  assign n3389 = ~n16186 | ~n16187;
  assign n16189 = P2_INSTQUEUE_REG_10__5_ & ~n16165;
  assign n16190 = n15641 & ~n16171;
  assign n16191 = n15646 & n16152;
  assign n16192 = n15648 & n16159;
  assign n16193 = n15653 & n16151;
  assign n16194 = ~n16191 & ~n16192;
  assign n16195 = ~n16193 & n16194;
  assign n16196 = ~n16189 & ~n16190;
  assign n3394 = ~n16195 | ~n16196;
  assign n16198 = P2_INSTQUEUE_REG_10__4_ & ~n16165;
  assign n16199 = n15663 & ~n16171;
  assign n16200 = n15668 & n16152;
  assign n16201 = n15670 & n16159;
  assign n16202 = n15675 & n16151;
  assign n16203 = ~n16200 & ~n16201;
  assign n16204 = ~n16202 & n16203;
  assign n16205 = ~n16198 & ~n16199;
  assign n3399 = ~n16204 | ~n16205;
  assign n16207 = P2_INSTQUEUE_REG_10__3_ & ~n16165;
  assign n16208 = n15685 & ~n16171;
  assign n16209 = n15690 & n16152;
  assign n16210 = n15692 & n16159;
  assign n16211 = n15697 & n16151;
  assign n16212 = ~n16209 & ~n16210;
  assign n16213 = ~n16211 & n16212;
  assign n16214 = ~n16207 & ~n16208;
  assign n3404 = ~n16213 | ~n16214;
  assign n16216 = P2_INSTQUEUE_REG_10__2_ & ~n16165;
  assign n16217 = n15707 & ~n16171;
  assign n16218 = n15712 & n16152;
  assign n16219 = n15714 & n16159;
  assign n16220 = n15719 & n16151;
  assign n16221 = ~n16218 & ~n16219;
  assign n16222 = ~n16220 & n16221;
  assign n16223 = ~n16216 & ~n16217;
  assign n3409 = ~n16222 | ~n16223;
  assign n16225 = P2_INSTQUEUE_REG_10__1_ & ~n16165;
  assign n16226 = n15729 & ~n16171;
  assign n16227 = n15734 & n16152;
  assign n16228 = n15736 & n16159;
  assign n16229 = n15741 & n16151;
  assign n16230 = ~n16227 & ~n16228;
  assign n16231 = ~n16229 & n16230;
  assign n16232 = ~n16225 & ~n16226;
  assign n3414 = ~n16231 | ~n16232;
  assign n16234 = P2_INSTQUEUE_REG_10__0_ & ~n16165;
  assign n16235 = n15751 & ~n16171;
  assign n16236 = n15756 & n16152;
  assign n16237 = n15758 & n16159;
  assign n16238 = n15763 & n16151;
  assign n16239 = ~n16236 & ~n16237;
  assign n16240 = ~n16238 & n16239;
  assign n16241 = ~n16234 & ~n16235;
  assign n3419 = ~n16240 | ~n16241;
  assign n16243 = n15467 & n15474;
  assign n16244 = n15864 & n16056;
  assign n16245 = ~n16243 & ~n16244;
  assign n16246 = n15867 & n16059;
  assign n16247 = n15515 & n15558;
  assign n16248 = ~n16246 & ~n16247;
  assign n16249 = n15574 & n16248;
  assign n16250 = ~n15481 & ~n16249;
  assign n16251 = n16245 & ~n16250;
  assign n16252 = n15874 & n16066;
  assign n16253 = ~n16243 & ~n16252;
  assign n16254 = P2_STATE2_REG_2_ & n16253;
  assign n16255 = P2_STATE2_REG_3_ & ~n16243;
  assign n16256 = ~n16254 & ~n16255;
  assign n16257 = n15573 & n16256;
  assign n16258 = ~n16251 & n16257;
  assign n16259 = P2_INSTQUEUE_REG_9__7_ & ~n16258;
  assign n16260 = P2_STATE2_REG_2_ & ~n16253;
  assign n16261 = n15569 & n16248;
  assign n16262 = ~n15481 & ~n16261;
  assign n16263 = ~n16245 & ~n16262;
  assign n16264 = ~n16260 & ~n16263;
  assign n16265 = n15591 & ~n16264;
  assign n16266 = n15601 & n16247;
  assign n16267 = n15604 & n16243;
  assign n16268 = n15609 & n16246;
  assign n16269 = ~n16266 & ~n16267;
  assign n16270 = ~n16268 & n16269;
  assign n16271 = ~n16259 & ~n16265;
  assign n3424 = ~n16270 | ~n16271;
  assign n16273 = P2_INSTQUEUE_REG_9__6_ & ~n16258;
  assign n16274 = n15619 & ~n16264;
  assign n16275 = n15624 & n16247;
  assign n16276 = n15626 & n16243;
  assign n16277 = n15631 & n16246;
  assign n16278 = ~n16275 & ~n16276;
  assign n16279 = ~n16277 & n16278;
  assign n16280 = ~n16273 & ~n16274;
  assign n3429 = ~n16279 | ~n16280;
  assign n16282 = P2_INSTQUEUE_REG_9__5_ & ~n16258;
  assign n16283 = n15641 & ~n16264;
  assign n16284 = n15646 & n16247;
  assign n16285 = n15648 & n16243;
  assign n16286 = n15653 & n16246;
  assign n16287 = ~n16284 & ~n16285;
  assign n16288 = ~n16286 & n16287;
  assign n16289 = ~n16282 & ~n16283;
  assign n3434 = ~n16288 | ~n16289;
  assign n16291 = P2_INSTQUEUE_REG_9__4_ & ~n16258;
  assign n16292 = n15663 & ~n16264;
  assign n16293 = n15668 & n16247;
  assign n16294 = n15670 & n16243;
  assign n16295 = n15675 & n16246;
  assign n16296 = ~n16293 & ~n16294;
  assign n16297 = ~n16295 & n16296;
  assign n16298 = ~n16291 & ~n16292;
  assign n3439 = ~n16297 | ~n16298;
  assign n16300 = P2_INSTQUEUE_REG_9__3_ & ~n16258;
  assign n16301 = n15685 & ~n16264;
  assign n16302 = n15690 & n16247;
  assign n16303 = n15692 & n16243;
  assign n16304 = n15697 & n16246;
  assign n16305 = ~n16302 & ~n16303;
  assign n16306 = ~n16304 & n16305;
  assign n16307 = ~n16300 & ~n16301;
  assign n3444 = ~n16306 | ~n16307;
  assign n16309 = P2_INSTQUEUE_REG_9__2_ & ~n16258;
  assign n16310 = n15707 & ~n16264;
  assign n16311 = n15712 & n16247;
  assign n16312 = n15714 & n16243;
  assign n16313 = n15719 & n16246;
  assign n16314 = ~n16311 & ~n16312;
  assign n16315 = ~n16313 & n16314;
  assign n16316 = ~n16309 & ~n16310;
  assign n3449 = ~n16315 | ~n16316;
  assign n16318 = P2_INSTQUEUE_REG_9__1_ & ~n16258;
  assign n16319 = n15729 & ~n16264;
  assign n16320 = n15734 & n16247;
  assign n16321 = n15736 & n16243;
  assign n16322 = n15741 & n16246;
  assign n16323 = ~n16320 & ~n16321;
  assign n16324 = ~n16322 & n16323;
  assign n16325 = ~n16318 & ~n16319;
  assign n3454 = ~n16324 | ~n16325;
  assign n16327 = P2_INSTQUEUE_REG_9__0_ & ~n16258;
  assign n16328 = n15751 & ~n16264;
  assign n16329 = n15756 & n16247;
  assign n16330 = n15758 & n16243;
  assign n16331 = n15763 & n16246;
  assign n16332 = ~n16329 & ~n16330;
  assign n16333 = ~n16331 & n16332;
  assign n16334 = ~n16327 & ~n16328;
  assign n3459 = ~n16333 | ~n16334;
  assign n16336 = n15959 & n16059;
  assign n16337 = n15558 & n15961;
  assign n16338 = ~n16336 & ~n16337;
  assign n16339 = n15574 & n16338;
  assign n16340 = ~n15481 & ~n16339;
  assign n16341 = n15476 & n16056;
  assign n16342 = ~n16340 & ~n16341;
  assign n16343 = n15968 & n16066;
  assign n16344 = n15467 & n15970;
  assign n16345 = ~n16343 & ~n16344;
  assign n16346 = P2_STATE2_REG_2_ & n16345;
  assign n16347 = P2_STATE2_REG_3_ & ~n16344;
  assign n16348 = ~n16346 & ~n16347;
  assign n16349 = n15573 & n16348;
  assign n16350 = ~n16342 & n16349;
  assign n16351 = P2_INSTQUEUE_REG_8__7_ & ~n16350;
  assign n16352 = P2_STATE2_REG_2_ & ~n16345;
  assign n16353 = n15569 & n16338;
  assign n16354 = ~n15481 & ~n16353;
  assign n16355 = n16341 & ~n16354;
  assign n16356 = ~n16352 & ~n16355;
  assign n16357 = n15591 & ~n16356;
  assign n16358 = n15601 & n16337;
  assign n16359 = n15604 & n16344;
  assign n16360 = n15609 & n16336;
  assign n16361 = ~n16358 & ~n16359;
  assign n16362 = ~n16360 & n16361;
  assign n16363 = ~n16351 & ~n16357;
  assign n3464 = ~n16362 | ~n16363;
  assign n16365 = P2_INSTQUEUE_REG_8__6_ & ~n16350;
  assign n16366 = n15619 & ~n16356;
  assign n16367 = n15624 & n16337;
  assign n16368 = n15626 & n16344;
  assign n16369 = n15631 & n16336;
  assign n16370 = ~n16367 & ~n16368;
  assign n16371 = ~n16369 & n16370;
  assign n16372 = ~n16365 & ~n16366;
  assign n3469 = ~n16371 | ~n16372;
  assign n16374 = P2_INSTQUEUE_REG_8__5_ & ~n16350;
  assign n16375 = n15641 & ~n16356;
  assign n16376 = n15646 & n16337;
  assign n16377 = n15648 & n16344;
  assign n16378 = n15653 & n16336;
  assign n16379 = ~n16376 & ~n16377;
  assign n16380 = ~n16378 & n16379;
  assign n16381 = ~n16374 & ~n16375;
  assign n3474 = ~n16380 | ~n16381;
  assign n16383 = P2_INSTQUEUE_REG_8__4_ & ~n16350;
  assign n16384 = n15663 & ~n16356;
  assign n16385 = n15668 & n16337;
  assign n16386 = n15670 & n16344;
  assign n16387 = n15675 & n16336;
  assign n16388 = ~n16385 & ~n16386;
  assign n16389 = ~n16387 & n16388;
  assign n16390 = ~n16383 & ~n16384;
  assign n3479 = ~n16389 | ~n16390;
  assign n16392 = P2_INSTQUEUE_REG_8__3_ & ~n16350;
  assign n16393 = n15685 & ~n16356;
  assign n16394 = n15690 & n16337;
  assign n16395 = n15692 & n16344;
  assign n16396 = n15697 & n16336;
  assign n16397 = ~n16394 & ~n16395;
  assign n16398 = ~n16396 & n16397;
  assign n16399 = ~n16392 & ~n16393;
  assign n3484 = ~n16398 | ~n16399;
  assign n16401 = P2_INSTQUEUE_REG_8__2_ & ~n16350;
  assign n16402 = n15707 & ~n16356;
  assign n16403 = n15712 & n16337;
  assign n16404 = n15714 & n16344;
  assign n16405 = n15719 & n16336;
  assign n16406 = ~n16403 & ~n16404;
  assign n16407 = ~n16405 & n16406;
  assign n16408 = ~n16401 & ~n16402;
  assign n3489 = ~n16407 | ~n16408;
  assign n16410 = P2_INSTQUEUE_REG_8__1_ & ~n16350;
  assign n16411 = n15729 & ~n16356;
  assign n16412 = n15734 & n16337;
  assign n16413 = n15736 & n16344;
  assign n16414 = n15741 & n16336;
  assign n16415 = ~n16412 & ~n16413;
  assign n16416 = ~n16414 & n16415;
  assign n16417 = ~n16410 & ~n16411;
  assign n3494 = ~n16416 | ~n16417;
  assign n16419 = P2_INSTQUEUE_REG_8__0_ & ~n16350;
  assign n16420 = n15751 & ~n16356;
  assign n16421 = n15756 & n16337;
  assign n16422 = n15758 & n16344;
  assign n16423 = n15763 & n16336;
  assign n16424 = ~n16421 & ~n16422;
  assign n16425 = ~n16423 & n16424;
  assign n16426 = ~n16419 & ~n16420;
  assign n3499 = ~n16425 | ~n16426;
  assign n16428 = ~n15466 & n15472;
  assign n16429 = n15477 & n16428;
  assign n16430 = ~n15470 & ~n16429;
  assign n16431 = ~n15542 & n15563;
  assign n16432 = n15517 & n16431;
  assign n16433 = ~n15561 & ~n16432;
  assign n16434 = n15574 & n16433;
  assign n16435 = ~n15481 & ~n16434;
  assign n16436 = n16430 & ~n16435;
  assign n16437 = n15147 & ~n15216;
  assign n16438 = n15579 & n16437;
  assign n16439 = ~n15470 & ~n16438;
  assign n16440 = P2_STATE2_REG_2_ & n16439;
  assign n16441 = P2_STATE2_REG_3_ & ~n15470;
  assign n16442 = ~n16440 & ~n16441;
  assign n16443 = n15573 & n16442;
  assign n16444 = ~n16436 & n16443;
  assign n16445 = P2_INSTQUEUE_REG_7__7_ & ~n16444;
  assign n16446 = P2_STATE2_REG_2_ & ~n16439;
  assign n16447 = n15569 & n16433;
  assign n16448 = ~n15481 & ~n16447;
  assign n16449 = ~n16430 & ~n16448;
  assign n16450 = ~n16446 & ~n16449;
  assign n16451 = n15591 & ~n16450;
  assign n16452 = n15561 & n15601;
  assign n16453 = n15470 & n15604;
  assign n16454 = n15609 & n16432;
  assign n16455 = ~n16452 & ~n16453;
  assign n16456 = ~n16454 & n16455;
  assign n16457 = ~n16445 & ~n16451;
  assign n3504 = ~n16456 | ~n16457;
  assign n16459 = P2_INSTQUEUE_REG_7__6_ & ~n16444;
  assign n16460 = n15619 & ~n16450;
  assign n16461 = n15561 & n15624;
  assign n16462 = n15470 & n15626;
  assign n16463 = n15631 & n16432;
  assign n16464 = ~n16461 & ~n16462;
  assign n16465 = ~n16463 & n16464;
  assign n16466 = ~n16459 & ~n16460;
  assign n3509 = ~n16465 | ~n16466;
  assign n16468 = P2_INSTQUEUE_REG_7__5_ & ~n16444;
  assign n16469 = n15641 & ~n16450;
  assign n16470 = n15561 & n15646;
  assign n16471 = n15470 & n15648;
  assign n16472 = n15653 & n16432;
  assign n16473 = ~n16470 & ~n16471;
  assign n16474 = ~n16472 & n16473;
  assign n16475 = ~n16468 & ~n16469;
  assign n3514 = ~n16474 | ~n16475;
  assign n16477 = P2_INSTQUEUE_REG_7__4_ & ~n16444;
  assign n16478 = n15663 & ~n16450;
  assign n16479 = n15561 & n15668;
  assign n16480 = n15470 & n15670;
  assign n16481 = n15675 & n16432;
  assign n16482 = ~n16479 & ~n16480;
  assign n16483 = ~n16481 & n16482;
  assign n16484 = ~n16477 & ~n16478;
  assign n3519 = ~n16483 | ~n16484;
  assign n16486 = P2_INSTQUEUE_REG_7__3_ & ~n16444;
  assign n16487 = n15685 & ~n16450;
  assign n16488 = n15561 & n15690;
  assign n16489 = n15470 & n15692;
  assign n16490 = n15697 & n16432;
  assign n16491 = ~n16488 & ~n16489;
  assign n16492 = ~n16490 & n16491;
  assign n16493 = ~n16486 & ~n16487;
  assign n3524 = ~n16492 | ~n16493;
  assign n16495 = P2_INSTQUEUE_REG_7__2_ & ~n16444;
  assign n16496 = n15707 & ~n16450;
  assign n16497 = n15561 & n15712;
  assign n16498 = n15470 & n15714;
  assign n16499 = n15719 & n16432;
  assign n16500 = ~n16497 & ~n16498;
  assign n16501 = ~n16499 & n16500;
  assign n16502 = ~n16495 & ~n16496;
  assign n3529 = ~n16501 | ~n16502;
  assign n16504 = P2_INSTQUEUE_REG_7__1_ & ~n16444;
  assign n16505 = n15729 & ~n16450;
  assign n16506 = n15561 & n15734;
  assign n16507 = n15470 & n15736;
  assign n16508 = n15741 & n16432;
  assign n16509 = ~n16506 & ~n16507;
  assign n16510 = ~n16508 & n16509;
  assign n16511 = ~n16504 & ~n16505;
  assign n3534 = ~n16510 | ~n16511;
  assign n16513 = P2_INSTQUEUE_REG_7__0_ & ~n16444;
  assign n16514 = n15751 & ~n16450;
  assign n16515 = n15561 & n15756;
  assign n16516 = n15470 & n15758;
  assign n16517 = n15763 & n16432;
  assign n16518 = ~n16515 & ~n16516;
  assign n16519 = ~n16517 & n16518;
  assign n16520 = ~n16513 & ~n16514;
  assign n3539 = ~n16519 | ~n16520;
  assign n16522 = n15769 & n16431;
  assign n16523 = n15514 & n15560;
  assign n16524 = ~n16522 & ~n16523;
  assign n16525 = n15574 & n16524;
  assign n16526 = ~n15481 & ~n16525;
  assign n16527 = ~n15476 & n16428;
  assign n16528 = ~n16526 & ~n16527;
  assign n16529 = n15777 & n16437;
  assign n16530 = n15469 & n15475;
  assign n16531 = ~n16529 & ~n16530;
  assign n16532 = P2_STATE2_REG_2_ & n16531;
  assign n16533 = P2_STATE2_REG_3_ & ~n16530;
  assign n16534 = ~n16532 & ~n16533;
  assign n16535 = n15573 & n16534;
  assign n16536 = ~n16528 & n16535;
  assign n16537 = P2_INSTQUEUE_REG_6__7_ & ~n16536;
  assign n16538 = P2_STATE2_REG_2_ & ~n16531;
  assign n16539 = n15569 & n16524;
  assign n16540 = ~n15481 & ~n16539;
  assign n16541 = n16527 & ~n16540;
  assign n16542 = ~n16538 & ~n16541;
  assign n16543 = n15591 & ~n16542;
  assign n16544 = n15601 & n16523;
  assign n16545 = n15604 & n16530;
  assign n16546 = n15609 & n16522;
  assign n16547 = ~n16544 & ~n16545;
  assign n16548 = ~n16546 & n16547;
  assign n16549 = ~n16537 & ~n16543;
  assign n3544 = ~n16548 | ~n16549;
  assign n16551 = P2_INSTQUEUE_REG_6__6_ & ~n16536;
  assign n16552 = n15619 & ~n16542;
  assign n16553 = n15624 & n16523;
  assign n16554 = n15626 & n16530;
  assign n16555 = n15631 & n16522;
  assign n16556 = ~n16553 & ~n16554;
  assign n16557 = ~n16555 & n16556;
  assign n16558 = ~n16551 & ~n16552;
  assign n3549 = ~n16557 | ~n16558;
  assign n16560 = P2_INSTQUEUE_REG_6__5_ & ~n16536;
  assign n16561 = n15641 & ~n16542;
  assign n16562 = n15646 & n16523;
  assign n16563 = n15648 & n16530;
  assign n16564 = n15653 & n16522;
  assign n16565 = ~n16562 & ~n16563;
  assign n16566 = ~n16564 & n16565;
  assign n16567 = ~n16560 & ~n16561;
  assign n3554 = ~n16566 | ~n16567;
  assign n16569 = P2_INSTQUEUE_REG_6__4_ & ~n16536;
  assign n16570 = n15663 & ~n16542;
  assign n16571 = n15668 & n16523;
  assign n16572 = n15670 & n16530;
  assign n16573 = n15675 & n16522;
  assign n16574 = ~n16571 & ~n16572;
  assign n16575 = ~n16573 & n16574;
  assign n16576 = ~n16569 & ~n16570;
  assign n3559 = ~n16575 | ~n16576;
  assign n16578 = P2_INSTQUEUE_REG_6__3_ & ~n16536;
  assign n16579 = n15685 & ~n16542;
  assign n16580 = n15690 & n16523;
  assign n16581 = n15692 & n16530;
  assign n16582 = n15697 & n16522;
  assign n16583 = ~n16580 & ~n16581;
  assign n16584 = ~n16582 & n16583;
  assign n16585 = ~n16578 & ~n16579;
  assign n3564 = ~n16584 | ~n16585;
  assign n16587 = P2_INSTQUEUE_REG_6__2_ & ~n16536;
  assign n16588 = n15707 & ~n16542;
  assign n16589 = n15712 & n16523;
  assign n16590 = n15714 & n16530;
  assign n16591 = n15719 & n16522;
  assign n16592 = ~n16589 & ~n16590;
  assign n16593 = ~n16591 & n16592;
  assign n16594 = ~n16587 & ~n16588;
  assign n3569 = ~n16593 | ~n16594;
  assign n16596 = P2_INSTQUEUE_REG_6__1_ & ~n16536;
  assign n16597 = n15729 & ~n16542;
  assign n16598 = n15734 & n16523;
  assign n16599 = n15736 & n16530;
  assign n16600 = n15741 & n16522;
  assign n16601 = ~n16598 & ~n16599;
  assign n16602 = ~n16600 & n16601;
  assign n16603 = ~n16596 & ~n16597;
  assign n3574 = ~n16602 | ~n16603;
  assign n16605 = P2_INSTQUEUE_REG_6__0_ & ~n16536;
  assign n16606 = n15751 & ~n16542;
  assign n16607 = n15756 & n16523;
  assign n16608 = n15758 & n16530;
  assign n16609 = n15763 & n16522;
  assign n16610 = ~n16607 & ~n16608;
  assign n16611 = ~n16609 & n16610;
  assign n16612 = ~n16605 & ~n16606;
  assign n3579 = ~n16611 | ~n16612;
  assign n16614 = n15469 & n15474;
  assign n16615 = n15864 & n16428;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = n15867 & n16431;
  assign n16618 = n15515 & n15560;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = n15574 & n16619;
  assign n16621 = ~n15481 & ~n16620;
  assign n16622 = n16616 & ~n16621;
  assign n16623 = n15874 & n16437;
  assign n16624 = ~n16614 & ~n16623;
  assign n16625 = P2_STATE2_REG_2_ & n16624;
  assign n16626 = P2_STATE2_REG_3_ & ~n16614;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = n15573 & n16627;
  assign n16629 = ~n16622 & n16628;
  assign n16630 = P2_INSTQUEUE_REG_5__7_ & ~n16629;
  assign n16631 = P2_STATE2_REG_2_ & ~n16624;
  assign n16632 = n15569 & n16619;
  assign n16633 = ~n15481 & ~n16632;
  assign n16634 = ~n16616 & ~n16633;
  assign n16635 = ~n16631 & ~n16634;
  assign n16636 = n15591 & ~n16635;
  assign n16637 = n15601 & n16618;
  assign n16638 = n15604 & n16614;
  assign n16639 = n15609 & n16617;
  assign n16640 = ~n16637 & ~n16638;
  assign n16641 = ~n16639 & n16640;
  assign n16642 = ~n16630 & ~n16636;
  assign n3584 = ~n16641 | ~n16642;
  assign n16644 = P2_INSTQUEUE_REG_5__6_ & ~n16629;
  assign n16645 = n15619 & ~n16635;
  assign n16646 = n15624 & n16618;
  assign n16647 = n15626 & n16614;
  assign n16648 = n15631 & n16617;
  assign n16649 = ~n16646 & ~n16647;
  assign n16650 = ~n16648 & n16649;
  assign n16651 = ~n16644 & ~n16645;
  assign n3589 = ~n16650 | ~n16651;
  assign n16653 = P2_INSTQUEUE_REG_5__5_ & ~n16629;
  assign n16654 = n15641 & ~n16635;
  assign n16655 = n15646 & n16618;
  assign n16656 = n15648 & n16614;
  assign n16657 = n15653 & n16617;
  assign n16658 = ~n16655 & ~n16656;
  assign n16659 = ~n16657 & n16658;
  assign n16660 = ~n16653 & ~n16654;
  assign n3594 = ~n16659 | ~n16660;
  assign n16662 = P2_INSTQUEUE_REG_5__4_ & ~n16629;
  assign n16663 = n15663 & ~n16635;
  assign n16664 = n15668 & n16618;
  assign n16665 = n15670 & n16614;
  assign n16666 = n15675 & n16617;
  assign n16667 = ~n16664 & ~n16665;
  assign n16668 = ~n16666 & n16667;
  assign n16669 = ~n16662 & ~n16663;
  assign n3599 = ~n16668 | ~n16669;
  assign n16671 = P2_INSTQUEUE_REG_5__3_ & ~n16629;
  assign n16672 = n15685 & ~n16635;
  assign n16673 = n15690 & n16618;
  assign n16674 = n15692 & n16614;
  assign n16675 = n15697 & n16617;
  assign n16676 = ~n16673 & ~n16674;
  assign n16677 = ~n16675 & n16676;
  assign n16678 = ~n16671 & ~n16672;
  assign n3604 = ~n16677 | ~n16678;
  assign n16680 = P2_INSTQUEUE_REG_5__2_ & ~n16629;
  assign n16681 = n15707 & ~n16635;
  assign n16682 = n15712 & n16618;
  assign n16683 = n15714 & n16614;
  assign n16684 = n15719 & n16617;
  assign n16685 = ~n16682 & ~n16683;
  assign n16686 = ~n16684 & n16685;
  assign n16687 = ~n16680 & ~n16681;
  assign n3609 = ~n16686 | ~n16687;
  assign n16689 = P2_INSTQUEUE_REG_5__1_ & ~n16629;
  assign n16690 = n15729 & ~n16635;
  assign n16691 = n15734 & n16618;
  assign n16692 = n15736 & n16614;
  assign n16693 = n15741 & n16617;
  assign n16694 = ~n16691 & ~n16692;
  assign n16695 = ~n16693 & n16694;
  assign n16696 = ~n16689 & ~n16690;
  assign n3614 = ~n16695 | ~n16696;
  assign n16698 = P2_INSTQUEUE_REG_5__0_ & ~n16629;
  assign n16699 = n15751 & ~n16635;
  assign n16700 = n15756 & n16618;
  assign n16701 = n15758 & n16614;
  assign n16702 = n15763 & n16617;
  assign n16703 = ~n16700 & ~n16701;
  assign n16704 = ~n16702 & n16703;
  assign n16705 = ~n16698 & ~n16699;
  assign n3619 = ~n16704 | ~n16705;
  assign n16707 = n15959 & n16431;
  assign n16708 = n15560 & n15961;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = n15574 & n16709;
  assign n16711 = ~n15481 & ~n16710;
  assign n16712 = n15476 & n16428;
  assign n16713 = ~n16711 & ~n16712;
  assign n16714 = n15968 & n16437;
  assign n16715 = n15469 & n15970;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = P2_STATE2_REG_2_ & n16716;
  assign n16718 = P2_STATE2_REG_3_ & ~n16715;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = n15573 & n16719;
  assign n16721 = ~n16713 & n16720;
  assign n16722 = P2_INSTQUEUE_REG_4__7_ & ~n16721;
  assign n16723 = P2_STATE2_REG_2_ & ~n16716;
  assign n16724 = n15569 & n16709;
  assign n16725 = ~n15481 & ~n16724;
  assign n16726 = n16712 & ~n16725;
  assign n16727 = ~n16723 & ~n16726;
  assign n16728 = n15591 & ~n16727;
  assign n16729 = n15601 & n16708;
  assign n16730 = n15604 & n16715;
  assign n16731 = n15609 & n16707;
  assign n16732 = ~n16729 & ~n16730;
  assign n16733 = ~n16731 & n16732;
  assign n16734 = ~n16722 & ~n16728;
  assign n3624 = ~n16733 | ~n16734;
  assign n16736 = P2_INSTQUEUE_REG_4__6_ & ~n16721;
  assign n16737 = n15619 & ~n16727;
  assign n16738 = n15624 & n16708;
  assign n16739 = n15626 & n16715;
  assign n16740 = n15631 & n16707;
  assign n16741 = ~n16738 & ~n16739;
  assign n16742 = ~n16740 & n16741;
  assign n16743 = ~n16736 & ~n16737;
  assign n3629 = ~n16742 | ~n16743;
  assign n16745 = P2_INSTQUEUE_REG_4__5_ & ~n16721;
  assign n16746 = n15641 & ~n16727;
  assign n16747 = n15646 & n16708;
  assign n16748 = n15648 & n16715;
  assign n16749 = n15653 & n16707;
  assign n16750 = ~n16747 & ~n16748;
  assign n16751 = ~n16749 & n16750;
  assign n16752 = ~n16745 & ~n16746;
  assign n3634 = ~n16751 | ~n16752;
  assign n16754 = P2_INSTQUEUE_REG_4__4_ & ~n16721;
  assign n16755 = n15663 & ~n16727;
  assign n16756 = n15668 & n16708;
  assign n16757 = n15670 & n16715;
  assign n16758 = n15675 & n16707;
  assign n16759 = ~n16756 & ~n16757;
  assign n16760 = ~n16758 & n16759;
  assign n16761 = ~n16754 & ~n16755;
  assign n3639 = ~n16760 | ~n16761;
  assign n16763 = P2_INSTQUEUE_REG_4__3_ & ~n16721;
  assign n16764 = n15685 & ~n16727;
  assign n16765 = n15690 & n16708;
  assign n16766 = n15692 & n16715;
  assign n16767 = n15697 & n16707;
  assign n16768 = ~n16765 & ~n16766;
  assign n16769 = ~n16767 & n16768;
  assign n16770 = ~n16763 & ~n16764;
  assign n3644 = ~n16769 | ~n16770;
  assign n16772 = P2_INSTQUEUE_REG_4__2_ & ~n16721;
  assign n16773 = n15707 & ~n16727;
  assign n16774 = n15712 & n16708;
  assign n16775 = n15714 & n16715;
  assign n16776 = n15719 & n16707;
  assign n16777 = ~n16774 & ~n16775;
  assign n16778 = ~n16776 & n16777;
  assign n16779 = ~n16772 & ~n16773;
  assign n3649 = ~n16778 | ~n16779;
  assign n16781 = P2_INSTQUEUE_REG_4__1_ & ~n16721;
  assign n16782 = n15729 & ~n16727;
  assign n16783 = n15734 & n16708;
  assign n16784 = n15736 & n16715;
  assign n16785 = n15741 & n16707;
  assign n16786 = ~n16783 & ~n16784;
  assign n16787 = ~n16785 & n16786;
  assign n16788 = ~n16781 & ~n16782;
  assign n3654 = ~n16787 | ~n16788;
  assign n16790 = P2_INSTQUEUE_REG_4__0_ & ~n16721;
  assign n16791 = n15751 & ~n16727;
  assign n16792 = n15756 & n16708;
  assign n16793 = n15758 & n16715;
  assign n16794 = n15763 & n16707;
  assign n16795 = ~n16792 & ~n16793;
  assign n16796 = ~n16794 & n16795;
  assign n16797 = ~n16790 & ~n16791;
  assign n3659 = ~n16796 | ~n16797;
  assign n16799 = ~P2_INSTQUEUEWR_ADDR_REG_3_ & ~P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n16800 = n15461 & n16799;
  assign n16801 = n15466 & n15472;
  assign n16802 = n15477 & n16801;
  assign n16803 = ~n16800 & ~n16802;
  assign n16804 = n15542 & n15563;
  assign n16805 = n15517 & n16804;
  assign n16806 = ~n15539 & n15557;
  assign n16807 = n15518 & n16806;
  assign n16808 = ~n16805 & ~n16807;
  assign n16809 = n15574 & n16808;
  assign n16810 = ~n15481 & ~n16809;
  assign n16811 = n16803 & ~n16810;
  assign n16812 = n15147 & n15216;
  assign n16813 = n15579 & n16812;
  assign n16814 = ~n16800 & ~n16813;
  assign n16815 = P2_STATE2_REG_2_ & n16814;
  assign n16816 = P2_STATE2_REG_3_ & ~n16800;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = n15573 & n16817;
  assign n16819 = ~n16811 & n16818;
  assign n16820 = P2_INSTQUEUE_REG_3__7_ & ~n16819;
  assign n16821 = P2_STATE2_REG_2_ & ~n16814;
  assign n16822 = n15569 & n16808;
  assign n16823 = ~n15481 & ~n16822;
  assign n16824 = ~n16803 & ~n16823;
  assign n16825 = ~n16821 & ~n16824;
  assign n16826 = n15591 & ~n16825;
  assign n16827 = n15601 & n16807;
  assign n16828 = n15604 & n16800;
  assign n16829 = n15609 & n16805;
  assign n16830 = ~n16827 & ~n16828;
  assign n16831 = ~n16829 & n16830;
  assign n16832 = ~n16820 & ~n16826;
  assign n3664 = ~n16831 | ~n16832;
  assign n16834 = P2_INSTQUEUE_REG_3__6_ & ~n16819;
  assign n16835 = n15619 & ~n16825;
  assign n16836 = n15624 & n16807;
  assign n16837 = n15626 & n16800;
  assign n16838 = n15631 & n16805;
  assign n16839 = ~n16836 & ~n16837;
  assign n16840 = ~n16838 & n16839;
  assign n16841 = ~n16834 & ~n16835;
  assign n3669 = ~n16840 | ~n16841;
  assign n16843 = P2_INSTQUEUE_REG_3__5_ & ~n16819;
  assign n16844 = n15641 & ~n16825;
  assign n16845 = n15646 & n16807;
  assign n16846 = n15648 & n16800;
  assign n16847 = n15653 & n16805;
  assign n16848 = ~n16845 & ~n16846;
  assign n16849 = ~n16847 & n16848;
  assign n16850 = ~n16843 & ~n16844;
  assign n3674 = ~n16849 | ~n16850;
  assign n16852 = P2_INSTQUEUE_REG_3__4_ & ~n16819;
  assign n16853 = n15663 & ~n16825;
  assign n16854 = n15668 & n16807;
  assign n16855 = n15670 & n16800;
  assign n16856 = n15675 & n16805;
  assign n16857 = ~n16854 & ~n16855;
  assign n16858 = ~n16856 & n16857;
  assign n16859 = ~n16852 & ~n16853;
  assign n3679 = ~n16858 | ~n16859;
  assign n16861 = P2_INSTQUEUE_REG_3__3_ & ~n16819;
  assign n16862 = n15685 & ~n16825;
  assign n16863 = n15690 & n16807;
  assign n16864 = n15692 & n16800;
  assign n16865 = n15697 & n16805;
  assign n16866 = ~n16863 & ~n16864;
  assign n16867 = ~n16865 & n16866;
  assign n16868 = ~n16861 & ~n16862;
  assign n3684 = ~n16867 | ~n16868;
  assign n16870 = P2_INSTQUEUE_REG_3__2_ & ~n16819;
  assign n16871 = n15707 & ~n16825;
  assign n16872 = n15712 & n16807;
  assign n16873 = n15714 & n16800;
  assign n16874 = n15719 & n16805;
  assign n16875 = ~n16872 & ~n16873;
  assign n16876 = ~n16874 & n16875;
  assign n16877 = ~n16870 & ~n16871;
  assign n3689 = ~n16876 | ~n16877;
  assign n16879 = P2_INSTQUEUE_REG_3__1_ & ~n16819;
  assign n16880 = n15729 & ~n16825;
  assign n16881 = n15734 & n16807;
  assign n16882 = n15736 & n16800;
  assign n16883 = n15741 & n16805;
  assign n16884 = ~n16881 & ~n16882;
  assign n16885 = ~n16883 & n16884;
  assign n16886 = ~n16879 & ~n16880;
  assign n3694 = ~n16885 | ~n16886;
  assign n16888 = P2_INSTQUEUE_REG_3__0_ & ~n16819;
  assign n16889 = n15751 & ~n16825;
  assign n16890 = n15756 & n16807;
  assign n16891 = n15758 & n16800;
  assign n16892 = n15763 & n16805;
  assign n16893 = ~n16890 & ~n16891;
  assign n16894 = ~n16892 & n16893;
  assign n16895 = ~n16888 & ~n16889;
  assign n3699 = ~n16894 | ~n16895;
  assign n16897 = n15769 & n16804;
  assign n16898 = n15514 & n16806;
  assign n16899 = ~n16897 & ~n16898;
  assign n16900 = n15574 & n16899;
  assign n16901 = ~n15481 & ~n16900;
  assign n16902 = ~n15476 & n16801;
  assign n16903 = ~n16901 & ~n16902;
  assign n16904 = n15777 & n16812;
  assign n16905 = n15475 & n16799;
  assign n16906 = ~n16904 & ~n16905;
  assign n16907 = P2_STATE2_REG_2_ & n16906;
  assign n16908 = P2_STATE2_REG_3_ & ~n16905;
  assign n16909 = ~n16907 & ~n16908;
  assign n16910 = n15573 & n16909;
  assign n16911 = ~n16903 & n16910;
  assign n16912 = P2_INSTQUEUE_REG_2__7_ & ~n16911;
  assign n16913 = P2_STATE2_REG_2_ & ~n16906;
  assign n16914 = n15569 & n16899;
  assign n16915 = ~n15481 & ~n16914;
  assign n16916 = n16902 & ~n16915;
  assign n16917 = ~n16913 & ~n16916;
  assign n16918 = n15591 & ~n16917;
  assign n16919 = n15601 & n16898;
  assign n16920 = n15604 & n16905;
  assign n16921 = n15609 & n16897;
  assign n16922 = ~n16919 & ~n16920;
  assign n16923 = ~n16921 & n16922;
  assign n16924 = ~n16912 & ~n16918;
  assign n3704 = ~n16923 | ~n16924;
  assign n16926 = P2_INSTQUEUE_REG_2__6_ & ~n16911;
  assign n16927 = n15619 & ~n16917;
  assign n16928 = n15624 & n16898;
  assign n16929 = n15626 & n16905;
  assign n16930 = n15631 & n16897;
  assign n16931 = ~n16928 & ~n16929;
  assign n16932 = ~n16930 & n16931;
  assign n16933 = ~n16926 & ~n16927;
  assign n3709 = ~n16932 | ~n16933;
  assign n16935 = P2_INSTQUEUE_REG_2__5_ & ~n16911;
  assign n16936 = n15641 & ~n16917;
  assign n16937 = n15646 & n16898;
  assign n16938 = n15648 & n16905;
  assign n16939 = n15653 & n16897;
  assign n16940 = ~n16937 & ~n16938;
  assign n16941 = ~n16939 & n16940;
  assign n16942 = ~n16935 & ~n16936;
  assign n3714 = ~n16941 | ~n16942;
  assign n16944 = P2_INSTQUEUE_REG_2__4_ & ~n16911;
  assign n16945 = n15663 & ~n16917;
  assign n16946 = n15668 & n16898;
  assign n16947 = n15670 & n16905;
  assign n16948 = n15675 & n16897;
  assign n16949 = ~n16946 & ~n16947;
  assign n16950 = ~n16948 & n16949;
  assign n16951 = ~n16944 & ~n16945;
  assign n3719 = ~n16950 | ~n16951;
  assign n16953 = P2_INSTQUEUE_REG_2__3_ & ~n16911;
  assign n16954 = n15685 & ~n16917;
  assign n16955 = n15690 & n16898;
  assign n16956 = n15692 & n16905;
  assign n16957 = n15697 & n16897;
  assign n16958 = ~n16955 & ~n16956;
  assign n16959 = ~n16957 & n16958;
  assign n16960 = ~n16953 & ~n16954;
  assign n3724 = ~n16959 | ~n16960;
  assign n16962 = P2_INSTQUEUE_REG_2__2_ & ~n16911;
  assign n16963 = n15707 & ~n16917;
  assign n16964 = n15712 & n16898;
  assign n16965 = n15714 & n16905;
  assign n16966 = n15719 & n16897;
  assign n16967 = ~n16964 & ~n16965;
  assign n16968 = ~n16966 & n16967;
  assign n16969 = ~n16962 & ~n16963;
  assign n3729 = ~n16968 | ~n16969;
  assign n16971 = P2_INSTQUEUE_REG_2__1_ & ~n16911;
  assign n16972 = n15729 & ~n16917;
  assign n16973 = n15734 & n16898;
  assign n16974 = n15736 & n16905;
  assign n16975 = n15741 & n16897;
  assign n16976 = ~n16973 & ~n16974;
  assign n16977 = ~n16975 & n16976;
  assign n16978 = ~n16971 & ~n16972;
  assign n3734 = ~n16977 | ~n16978;
  assign n16980 = P2_INSTQUEUE_REG_2__0_ & ~n16911;
  assign n16981 = n15751 & ~n16917;
  assign n16982 = n15756 & n16898;
  assign n16983 = n15758 & n16905;
  assign n16984 = n15763 & n16897;
  assign n16985 = ~n16982 & ~n16983;
  assign n16986 = ~n16984 & n16985;
  assign n16987 = ~n16980 & ~n16981;
  assign n3739 = ~n16986 | ~n16987;
  assign n16989 = n15474 & n16799;
  assign n16990 = n15864 & n16801;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = n15867 & n16804;
  assign n16993 = n15515 & n16806;
  assign n16994 = ~n16992 & ~n16993;
  assign n16995 = n15574 & n16994;
  assign n16996 = ~n15481 & ~n16995;
  assign n16997 = n16991 & ~n16996;
  assign n16998 = n15874 & n16812;
  assign n16999 = ~n16989 & ~n16998;
  assign n17000 = P2_STATE2_REG_2_ & n16999;
  assign n17001 = P2_STATE2_REG_3_ & ~n16989;
  assign n17002 = ~n17000 & ~n17001;
  assign n17003 = n15573 & n17002;
  assign n17004 = ~n16997 & n17003;
  assign n17005 = P2_INSTQUEUE_REG_1__7_ & ~n17004;
  assign n17006 = P2_STATE2_REG_2_ & ~n16999;
  assign n17007 = n15569 & n16994;
  assign n17008 = ~n15481 & ~n17007;
  assign n17009 = ~n16991 & ~n17008;
  assign n17010 = ~n17006 & ~n17009;
  assign n17011 = n15591 & ~n17010;
  assign n17012 = n15601 & n16993;
  assign n17013 = n15604 & n16989;
  assign n17014 = n15609 & n16992;
  assign n17015 = ~n17012 & ~n17013;
  assign n17016 = ~n17014 & n17015;
  assign n17017 = ~n17005 & ~n17011;
  assign n3744 = ~n17016 | ~n17017;
  assign n17019 = P2_INSTQUEUE_REG_1__6_ & ~n17004;
  assign n17020 = n15619 & ~n17010;
  assign n17021 = n15624 & n16993;
  assign n17022 = n15626 & n16989;
  assign n17023 = n15631 & n16992;
  assign n17024 = ~n17021 & ~n17022;
  assign n17025 = ~n17023 & n17024;
  assign n17026 = ~n17019 & ~n17020;
  assign n3749 = ~n17025 | ~n17026;
  assign n17028 = P2_INSTQUEUE_REG_1__5_ & ~n17004;
  assign n17029 = n15641 & ~n17010;
  assign n17030 = n15646 & n16993;
  assign n17031 = n15648 & n16989;
  assign n17032 = n15653 & n16992;
  assign n17033 = ~n17030 & ~n17031;
  assign n17034 = ~n17032 & n17033;
  assign n17035 = ~n17028 & ~n17029;
  assign n3754 = ~n17034 | ~n17035;
  assign n17037 = P2_INSTQUEUE_REG_1__4_ & ~n17004;
  assign n17038 = n15663 & ~n17010;
  assign n17039 = n15668 & n16993;
  assign n17040 = n15670 & n16989;
  assign n17041 = n15675 & n16992;
  assign n17042 = ~n17039 & ~n17040;
  assign n17043 = ~n17041 & n17042;
  assign n17044 = ~n17037 & ~n17038;
  assign n3759 = ~n17043 | ~n17044;
  assign n17046 = P2_INSTQUEUE_REG_1__3_ & ~n17004;
  assign n17047 = n15685 & ~n17010;
  assign n17048 = n15690 & n16993;
  assign n17049 = n15692 & n16989;
  assign n17050 = n15697 & n16992;
  assign n17051 = ~n17048 & ~n17049;
  assign n17052 = ~n17050 & n17051;
  assign n17053 = ~n17046 & ~n17047;
  assign n3764 = ~n17052 | ~n17053;
  assign n17055 = P2_INSTQUEUE_REG_1__2_ & ~n17004;
  assign n17056 = n15707 & ~n17010;
  assign n17057 = n15712 & n16993;
  assign n17058 = n15714 & n16989;
  assign n17059 = n15719 & n16992;
  assign n17060 = ~n17057 & ~n17058;
  assign n17061 = ~n17059 & n17060;
  assign n17062 = ~n17055 & ~n17056;
  assign n3769 = ~n17061 | ~n17062;
  assign n17064 = P2_INSTQUEUE_REG_1__1_ & ~n17004;
  assign n17065 = n15729 & ~n17010;
  assign n17066 = n15734 & n16993;
  assign n17067 = n15736 & n16989;
  assign n17068 = n15741 & n16992;
  assign n17069 = ~n17066 & ~n17067;
  assign n17070 = ~n17068 & n17069;
  assign n17071 = ~n17064 & ~n17065;
  assign n3774 = ~n17070 | ~n17071;
  assign n17073 = P2_INSTQUEUE_REG_1__0_ & ~n17004;
  assign n17074 = n15751 & ~n17010;
  assign n17075 = n15756 & n16993;
  assign n17076 = n15758 & n16989;
  assign n17077 = n15763 & n16992;
  assign n17078 = ~n17075 & ~n17076;
  assign n17079 = ~n17077 & n17078;
  assign n17080 = ~n17073 & ~n17074;
  assign n3779 = ~n17079 | ~n17080;
  assign n17082 = n15959 & n16804;
  assign n17083 = n15961 & n16806;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = n15574 & n17084;
  assign n17086 = ~n15481 & ~n17085;
  assign n17087 = n15476 & n16801;
  assign n17088 = ~n17086 & ~n17087;
  assign n17089 = n15968 & n16812;
  assign n17090 = n15970 & n16799;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = P2_STATE2_REG_2_ & n17091;
  assign n17093 = P2_STATE2_REG_3_ & ~n17090;
  assign n17094 = ~n17092 & ~n17093;
  assign n17095 = n15573 & n17094;
  assign n17096 = ~n17088 & n17095;
  assign n17097 = P2_INSTQUEUE_REG_0__7_ & ~n17096;
  assign n17098 = P2_STATE2_REG_2_ & ~n17091;
  assign n17099 = n15569 & n17084;
  assign n17100 = ~n15481 & ~n17099;
  assign n17101 = n17087 & ~n17100;
  assign n17102 = ~n17098 & ~n17101;
  assign n17103 = n15591 & ~n17102;
  assign n17104 = n15601 & n17083;
  assign n17105 = n15604 & n17090;
  assign n17106 = n15609 & n17082;
  assign n17107 = ~n17104 & ~n17105;
  assign n17108 = ~n17106 & n17107;
  assign n17109 = ~n17097 & ~n17103;
  assign n3784 = ~n17108 | ~n17109;
  assign n17111 = P2_INSTQUEUE_REG_0__6_ & ~n17096;
  assign n17112 = n15619 & ~n17102;
  assign n17113 = n15624 & n17083;
  assign n17114 = n15626 & n17090;
  assign n17115 = n15631 & n17082;
  assign n17116 = ~n17113 & ~n17114;
  assign n17117 = ~n17115 & n17116;
  assign n17118 = ~n17111 & ~n17112;
  assign n3789 = ~n17117 | ~n17118;
  assign n17120 = P2_INSTQUEUE_REG_0__5_ & ~n17096;
  assign n17121 = n15641 & ~n17102;
  assign n17122 = n15646 & n17083;
  assign n17123 = n15648 & n17090;
  assign n17124 = n15653 & n17082;
  assign n17125 = ~n17122 & ~n17123;
  assign n17126 = ~n17124 & n17125;
  assign n17127 = ~n17120 & ~n17121;
  assign n3794 = ~n17126 | ~n17127;
  assign n17129 = P2_INSTQUEUE_REG_0__4_ & ~n17096;
  assign n17130 = n15663 & ~n17102;
  assign n17131 = n15668 & n17083;
  assign n17132 = n15670 & n17090;
  assign n17133 = n15675 & n17082;
  assign n17134 = ~n17131 & ~n17132;
  assign n17135 = ~n17133 & n17134;
  assign n17136 = ~n17129 & ~n17130;
  assign n3799 = ~n17135 | ~n17136;
  assign n17138 = P2_INSTQUEUE_REG_0__3_ & ~n17096;
  assign n17139 = n15685 & ~n17102;
  assign n17140 = n15690 & n17083;
  assign n17141 = n15692 & n17090;
  assign n17142 = n15697 & n17082;
  assign n17143 = ~n17140 & ~n17141;
  assign n17144 = ~n17142 & n17143;
  assign n17145 = ~n17138 & ~n17139;
  assign n3804 = ~n17144 | ~n17145;
  assign n17147 = P2_INSTQUEUE_REG_0__2_ & ~n17096;
  assign n17148 = n15707 & ~n17102;
  assign n17149 = n15712 & n17083;
  assign n17150 = n15714 & n17090;
  assign n17151 = n15719 & n17082;
  assign n17152 = ~n17149 & ~n17150;
  assign n17153 = ~n17151 & n17152;
  assign n17154 = ~n17147 & ~n17148;
  assign n3809 = ~n17153 | ~n17154;
  assign n17156 = P2_INSTQUEUE_REG_0__1_ & ~n17096;
  assign n17157 = n15729 & ~n17102;
  assign n17158 = n15734 & n17083;
  assign n17159 = n15736 & n17090;
  assign n17160 = n15741 & n17082;
  assign n17161 = ~n17158 & ~n17159;
  assign n17162 = ~n17160 & n17161;
  assign n17163 = ~n17156 & ~n17157;
  assign n3814 = ~n17162 | ~n17163;
  assign n17165 = P2_INSTQUEUE_REG_0__0_ & ~n17096;
  assign n17166 = n15751 & ~n17102;
  assign n17167 = n15756 & n17083;
  assign n17168 = n15758 & n17090;
  assign n17169 = n15763 & n17082;
  assign n17170 = ~n17167 & ~n17168;
  assign n17171 = ~n17169 & n17170;
  assign n17172 = ~n17165 & ~n17166;
  assign n3819 = ~n17171 | ~n17172;
  assign n17174 = P2_STATE2_REG_3_ & ~P2_STATE2_REG_0_;
  assign n17175 = P2_STATE2_REG_0_ & P2_FLUSH_REG;
  assign n17176 = n14141 & n17175;
  assign n17177 = ~n17174 & ~n17176;
  assign n17178 = ~n15200 & n15432;
  assign n17179 = n17177 & ~n17178;
  assign n17180 = P2_INSTQUEUERD_ADDR_REG_4_ & n17179;
  assign n17181 = ~n15230 & n15437;
  assign n17182 = n15172 & n17181;
  assign n17183 = ~n17179 & n17182;
  assign n3824 = n17180 | n17183;
  assign n17185 = ~n15170 & n15437;
  assign n17186 = n15447 & ~n15557;
  assign n17187 = ~n17185 & ~n17186;
  assign n17188 = ~n17179 & ~n17187;
  assign n17189 = P2_INSTQUEUERD_ADDR_REG_3_ & n17179;
  assign n3829 = n17188 | n17189;
  assign n17191 = n15447 & n15539;
  assign n17192 = ~n15218 & n15437;
  assign n17193 = P2_STATE2_REG_1_ & n15360;
  assign n17194 = ~n17191 & ~n17192;
  assign n17195 = ~n17193 & n17194;
  assign n17196 = ~n17179 & ~n17195;
  assign n17197 = P2_INSTQUEUERD_ADDR_REG_2_ & n17179;
  assign n3834 = n17196 | n17197;
  assign n17199 = n15447 & ~n15510;
  assign n17200 = ~n15265 & n15437;
  assign n17201 = P2_STATE2_REG_1_ & n15359;
  assign n17202 = ~n15344 & n17201;
  assign n17203 = ~n17199 & ~n17200;
  assign n17204 = ~n17202 & n17203;
  assign n17205 = ~n17179 & ~n17204;
  assign n17206 = P2_INSTQUEUERD_ADDR_REG_1_ & n17179;
  assign n3839 = n17205 | n17206;
  assign n17208 = ~n15279 & n15437;
  assign n17209 = n15447 & ~n15513;
  assign n17210 = P2_STATE2_REG_1_ & n15344;
  assign n17211 = ~n17208 & ~n17209;
  assign n17212 = ~n17210 & n17211;
  assign n17213 = ~n17179 & ~n17212;
  assign n17214 = P2_INSTQUEUERD_ADDR_REG_0_ & n17179;
  assign n3844 = n17213 | n17214;
  assign n17216 = P2_STATE2_REG_0_ & n14141;
  assign n17217 = ~n15389 & n17216;
  assign n17218 = ~n15573 & ~n17176;
  assign n17219 = ~n17217 & n17218;
  assign n3849 = P2_INSTQUEUEWR_ADDR_REG_4_ & n17219;
  assign n17221 = ~n15437 & ~n15481;
  assign n17222 = ~n15557 & ~n17221;
  assign n17223 = n14238 & n14365;
  assign n17224 = ~P2_STATE2_REG_3_ & ~n14143;
  assign n17225 = ~n14286 & n17224;
  assign n17226 = n17223 & n17225;
  assign n17227 = P2_REIP_REG_2_ & n17226;
  assign n17228 = ~P2_STATE2_REG_3_ & n14286;
  assign n17229 = P2_EAX_REG_2_ & n17228;
  assign n17230 = ~n17227 & ~n17229;
  assign n17231 = ~P2_STATE2_REG_3_ & ~n14238;
  assign n17232 = n14365 & n17231;
  assign n17233 = ~n14404 & n17225;
  assign n17234 = n14974 & n17231;
  assign n17235 = ~n17232 & ~n17233;
  assign n17236 = ~n17234 & n17235;
  assign n17237 = P2_INSTADDRPOINTER_REG_2_ & ~n17236;
  assign n17238 = n17230 & ~n17237;
  assign n17239 = P2_STATE2_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_2_;
  assign n17240 = ~n17234 & ~n17239;
  assign n17241 = ~P2_STATE2_REG_3_ & ~n14365;
  assign n17242 = n14238 & n17241;
  assign n17243 = ~n14722 & n17242;
  assign n17244 = n17240 & ~n17243;
  assign n17245 = ~n17238 & ~n17244;
  assign n17246 = n17238 & n17244;
  assign n17247 = P2_INSTADDRPOINTER_REG_0_ & ~n17236;
  assign n17248 = P2_EAX_REG_0_ & n17228;
  assign n17249 = P2_REIP_REG_0_ & n17226;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = ~P2_STATE2_REG_3_ & ~n17247;
  assign n17252 = n17250 & n17251;
  assign n17253 = P2_STATE2_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_0_;
  assign n17254 = ~n17228 & ~n17253;
  assign n17255 = ~n17234 & n17254;
  assign n17256 = ~n14839 & n17242;
  assign n17257 = n17255 & ~n17256;
  assign n17258 = ~n14974 & n17225;
  assign n17259 = P2_STATE2_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_1_;
  assign n17260 = ~n17232 & ~n17258;
  assign n17261 = ~n17259 & n17260;
  assign n17262 = ~n14802 & n17242;
  assign n17263 = n17261 & ~n17262;
  assign n17264 = ~n17252 & ~n17257;
  assign n17265 = ~n17263 & n17264;
  assign n17266 = P2_REIP_REG_1_ & n17226;
  assign n17267 = P2_EAX_REG_1_ & n17228;
  assign n17268 = ~n17266 & ~n17267;
  assign n17269 = P2_INSTADDRPOINTER_REG_1_ & ~n17236;
  assign n17270 = n17268 & ~n17269;
  assign n17271 = n17263 & ~n17264;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = ~n17265 & ~n17272;
  assign n17274 = ~n17246 & ~n17273;
  assign n17275 = ~n17245 & ~n17274;
  assign n17276 = P2_STATE2_REG_3_ & P2_INSTQUEUEWR_ADDR_REG_3_;
  assign n17277 = ~n14685 & n17242;
  assign n17278 = ~n17276 & ~n17277;
  assign n17279 = P2_REIP_REG_3_ & n17226;
  assign n17280 = P2_EAX_REG_3_ & n17228;
  assign n17281 = ~n17279 & ~n17280;
  assign n17282 = P2_INSTADDRPOINTER_REG_3_ & ~n17236;
  assign n17283 = n17281 & ~n17282;
  assign n17284 = ~n17278 & n17283;
  assign n17285 = n17278 & ~n17283;
  assign n17286 = ~n17284 & ~n17285;
  assign n17287 = n17275 & ~n17286;
  assign n17288 = ~n17275 & n17286;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = P2_STATE2_REG_3_ & ~n17289;
  assign n17291 = ~n17222 & ~n17290;
  assign n17292 = n15517 & ~n15542;
  assign n17293 = ~n15563 & ~n17292;
  assign n17294 = ~n16432 & ~n17293;
  assign n17295 = n15569 & ~n17294;
  assign n17296 = n17291 & ~n17295;
  assign n17297 = ~n17219 & ~n17296;
  assign n17298 = P2_INSTQUEUEWR_ADDR_REG_3_ & n17219;
  assign n3854 = n17297 | n17298;
  assign n17300 = n15539 & ~n17221;
  assign n17301 = n17238 & ~n17244;
  assign n17302 = ~n17238 & n17244;
  assign n17303 = ~n17301 & ~n17302;
  assign n17304 = n17273 & ~n17303;
  assign n17305 = ~n17273 & n17303;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = P2_STATE2_REG_3_ & ~n17306;
  assign n17308 = ~n17300 & ~n17307;
  assign n17309 = ~n15517 & ~n15542;
  assign n17310 = n15517 & n15542;
  assign n17311 = ~n17309 & ~n17310;
  assign n17312 = n15569 & ~n17311;
  assign n17313 = n17308 & ~n17312;
  assign n17314 = ~n17219 & ~n17313;
  assign n17315 = P2_INSTQUEUEWR_ADDR_REG_2_ & n17219;
  assign n3859 = n17314 | n17315;
  assign n17317 = ~n15510 & ~n17221;
  assign n17318 = n17265 & ~n17270;
  assign n17319 = ~n17263 & ~n17264;
  assign n17320 = n17270 & n17319;
  assign n17321 = ~n17318 & ~n17320;
  assign n17322 = n17264 & n17270;
  assign n17323 = ~n17264 & ~n17270;
  assign n17324 = ~n17322 & ~n17323;
  assign n17325 = n17263 & ~n17324;
  assign n17326 = n17321 & ~n17325;
  assign n17327 = P2_STATE2_REG_3_ & ~n17326;
  assign n17328 = ~n17317 & ~n17327;
  assign n17329 = ~n15769 & ~n15867;
  assign n17330 = n15569 & ~n17329;
  assign n17331 = n17328 & ~n17330;
  assign n17332 = ~n17219 & ~n17331;
  assign n17333 = P2_INSTQUEUEWR_ADDR_REG_1_ & n17219;
  assign n3864 = n17332 | n17333;
  assign n17335 = ~n15437 & ~n15480;
  assign n17336 = ~n15513 & ~n17335;
  assign n17337 = n17252 & ~n17257;
  assign n17338 = ~n17252 & n17257;
  assign n17339 = ~n17337 & ~n17338;
  assign n17340 = P2_STATE2_REG_3_ & ~n17339;
  assign n17341 = ~n17336 & ~n17340;
  assign n17342 = ~n15451 & n17341;
  assign n17343 = ~n17219 & ~n17342;
  assign n17344 = P2_INSTQUEUEWR_ADDR_REG_0_ & n17219;
  assign n3869 = n17343 | n17344;
  assign n17346 = P2_INSTQUEUE_REG_15__0_ & n15580;
  assign n17347 = P2_INSTQUEUE_REG_14__0_ & n15778;
  assign n17348 = P2_INSTQUEUE_REG_13__0_ & n15875;
  assign n17349 = P2_INSTQUEUE_REG_12__0_ & n15969;
  assign n17350 = ~n17346 & ~n17347;
  assign n17351 = ~n17348 & n17350;
  assign n17352 = ~n17349 & n17351;
  assign n17353 = P2_INSTQUEUE_REG_11__0_ & n16067;
  assign n17354 = P2_INSTQUEUE_REG_10__0_ & n16158;
  assign n17355 = P2_INSTQUEUE_REG_9__0_ & n16252;
  assign n17356 = P2_INSTQUEUE_REG_8__0_ & n16343;
  assign n17357 = ~n17353 & ~n17354;
  assign n17358 = ~n17355 & n17357;
  assign n17359 = ~n17356 & n17358;
  assign n17360 = P2_INSTQUEUE_REG_7__0_ & n16438;
  assign n17361 = P2_INSTQUEUE_REG_6__0_ & n16529;
  assign n17362 = P2_INSTQUEUE_REG_5__0_ & n16623;
  assign n17363 = P2_INSTQUEUE_REG_4__0_ & n16714;
  assign n17364 = ~n17360 & ~n17361;
  assign n17365 = ~n17362 & n17364;
  assign n17366 = ~n17363 & n17365;
  assign n17367 = P2_INSTQUEUE_REG_3__0_ & n16813;
  assign n17368 = P2_INSTQUEUE_REG_2__0_ & n16904;
  assign n17369 = P2_INSTQUEUE_REG_1__0_ & n16998;
  assign n17370 = P2_INSTQUEUE_REG_0__0_ & n17089;
  assign n17371 = ~n17367 & ~n17368;
  assign n17372 = ~n17369 & n17371;
  assign n17373 = ~n17370 & n17372;
  assign n17374 = n17352 & n17359;
  assign n17375 = n17366 & n17374;
  assign n17376 = n17373 & n17375;
  assign n17377 = ~n14238 & ~n17376;
  assign n17378 = n14238 & ~n14839;
  assign n17379 = ~n17377 & ~n17378;
  assign n17380 = ~n14238 & ~n17379;
  assign n17381 = n14238 & n17379;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = ~P2_INSTADDRPOINTER_REG_0_ & ~n17382;
  assign n17384 = P2_INSTADDRPOINTER_REG_0_ & n17382;
  assign n17385 = ~n17383 & ~n17384;
  assign n17386 = ~P2_STATE2_REG_1_ & n15480;
  assign n17387 = ~P2_STATE2_REG_0_ & n17386;
  assign n17388 = ~n14238 & ~n14486;
  assign n17389 = n14238 & n14482;
  assign n17390 = ~n17388 & ~n17389;
  assign n17391 = ~n14051 & n17390;
  assign n17392 = n14548 & n17391;
  assign n17393 = ~n15182 & ~n17392;
  assign n17394 = ~n15184 & n17393;
  assign n17395 = n14238 & n14975;
  assign n17396 = n14145 & ~n14482;
  assign n17397 = ~n14238 & n17396;
  assign n17398 = ~n17395 & ~n17397;
  assign n17399 = ~n14949 & ~n17398;
  assign n17400 = ~n14199 & ~n14443;
  assign n17401 = n14949 & n17400;
  assign n17402 = ~n17399 & ~n17401;
  assign n17403 = ~n14238 & n15389;
  assign n17404 = ~n15299 & ~n17403;
  assign n17405 = n15047 & ~n17404;
  assign n17406 = n15196 & n17394;
  assign n17407 = n17402 & n17406;
  assign n17408 = ~n17405 & n17407;
  assign n17409 = n15432 & ~n17408;
  assign n17410 = ~n17387 & ~n17409;
  assign n17411 = P2_STATE2_REG_2_ & ~n17410;
  assign n17412 = n15047 & n17411;
  assign n17413 = n14239 & n17412;
  assign n17414 = ~n17385 & n17413;
  assign n17415 = P2_INSTQUEUE_REG_0__7_ & n14560;
  assign n17416 = P2_INSTQUEUE_REG_1__7_ & n14563;
  assign n17417 = P2_INSTQUEUE_REG_2__7_ & n14566;
  assign n17418 = P2_INSTQUEUE_REG_3__7_ & n14568;
  assign n17419 = ~n17415 & ~n17416;
  assign n17420 = ~n17417 & n17419;
  assign n17421 = ~n17418 & n17420;
  assign n17422 = P2_INSTQUEUE_REG_4__7_ & n14574;
  assign n17423 = P2_INSTQUEUE_REG_5__7_ & n14577;
  assign n17424 = P2_INSTQUEUE_REG_6__7_ & n14579;
  assign n17425 = P2_INSTQUEUE_REG_7__7_ & n14581;
  assign n17426 = ~n17422 & ~n17423;
  assign n17427 = ~n17424 & n17426;
  assign n17428 = ~n17425 & n17427;
  assign n17429 = P2_INSTQUEUE_REG_15__7_ & n14587;
  assign n17430 = P2_INSTQUEUE_REG_14__7_ & n14589;
  assign n17431 = P2_INSTQUEUE_REG_13__7_ & n14592;
  assign n17432 = P2_INSTQUEUE_REG_12__7_ & n14594;
  assign n17433 = ~n17429 & ~n17430;
  assign n17434 = ~n17431 & n17433;
  assign n17435 = ~n17432 & n17434;
  assign n17436 = P2_INSTQUEUE_REG_11__7_ & n14599;
  assign n17437 = P2_INSTQUEUE_REG_10__7_ & n14601;
  assign n17438 = P2_INSTQUEUE_REG_9__7_ & n14603;
  assign n17439 = P2_INSTQUEUE_REG_8__7_ & n14605;
  assign n17440 = ~n17436 & ~n17437;
  assign n17441 = ~n17438 & n17440;
  assign n17442 = ~n17439 & n17441;
  assign n17443 = n17421 & n17428;
  assign n17444 = n17435 & n17443;
  assign n17445 = n17442 & n17444;
  assign n17446 = P2_EBX_REG_0_ & n14365;
  assign n17447 = ~n14365 & ~n14920;
  assign n17448 = ~n17446 & ~n17447;
  assign n17449 = n14365 & ~n17448;
  assign n17450 = ~n14365 & n17448;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = ~n17445 & ~n17451;
  assign n17453 = ~n17382 & n17445;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = ~P2_INSTADDRPOINTER_REG_0_ & ~n17454;
  assign n17456 = P2_INSTADDRPOINTER_REG_0_ & n17454;
  assign n17457 = ~n17455 & ~n17456;
  assign n17458 = n14244 & n17412;
  assign n17459 = ~n17457 & n17458;
  assign n17460 = P2_INSTADDRPOINTER_REG_0_ & n17410;
  assign n17461 = ~P2_STATE2_REG_2_ & ~n17410;
  assign n17462 = P2_REIP_REG_0_ & n17461;
  assign n17463 = ~n17460 & ~n17462;
  assign n17464 = n14979 & n17411;
  assign n17465 = ~P2_INSTADDRPOINTER_REG_0_ & n17464;
  assign n17466 = n14240 & n15047;
  assign n17467 = ~n14962 & ~n17466;
  assign n17468 = n15167 & n17467;
  assign n17469 = n17411 & ~n17468;
  assign n17470 = ~P2_INSTADDRPOINTER_REG_0_ & n17469;
  assign n17471 = ~n17465 & ~n17470;
  assign n17472 = n14239 & n14486;
  assign n17473 = ~n14990 & ~n17472;
  assign n17474 = ~n14967 & n17473;
  assign n17475 = ~n15172 & n17474;
  assign n17476 = n17411 & ~n17475;
  assign n17477 = ~n15277 & n17476;
  assign n17478 = ~n14978 & ~n15173;
  assign n17479 = ~n15178 & n17478;
  assign n17480 = n17411 & ~n17479;
  assign n17481 = ~n17339 & n17480;
  assign n17482 = ~n17477 & ~n17481;
  assign n17483 = ~n17414 & ~n17459;
  assign n17484 = n17463 & n17483;
  assign n17485 = n17471 & n17484;
  assign n3874 = ~n17482 | ~n17485;
  assign n17487 = P2_INSTADDRPOINTER_REG_0_ & ~n17382;
  assign n17488 = ~P2_INSTADDRPOINTER_REG_1_ & n17487;
  assign n17489 = P2_INSTADDRPOINTER_REG_1_ & ~n17487;
  assign n17490 = ~n17488 & ~n17489;
  assign n17491 = P2_INSTQUEUE_REG_15__1_ & n15580;
  assign n17492 = P2_INSTQUEUE_REG_14__1_ & n15778;
  assign n17493 = P2_INSTQUEUE_REG_13__1_ & n15875;
  assign n17494 = P2_INSTQUEUE_REG_12__1_ & n15969;
  assign n17495 = ~n17491 & ~n17492;
  assign n17496 = ~n17493 & n17495;
  assign n17497 = ~n17494 & n17496;
  assign n17498 = P2_INSTQUEUE_REG_11__1_ & n16067;
  assign n17499 = P2_INSTQUEUE_REG_10__1_ & n16158;
  assign n17500 = P2_INSTQUEUE_REG_9__1_ & n16252;
  assign n17501 = P2_INSTQUEUE_REG_8__1_ & n16343;
  assign n17502 = ~n17498 & ~n17499;
  assign n17503 = ~n17500 & n17502;
  assign n17504 = ~n17501 & n17503;
  assign n17505 = P2_INSTQUEUE_REG_7__1_ & n16438;
  assign n17506 = P2_INSTQUEUE_REG_6__1_ & n16529;
  assign n17507 = P2_INSTQUEUE_REG_5__1_ & n16623;
  assign n17508 = P2_INSTQUEUE_REG_4__1_ & n16714;
  assign n17509 = ~n17505 & ~n17506;
  assign n17510 = ~n17507 & n17509;
  assign n17511 = ~n17508 & n17510;
  assign n17512 = P2_INSTQUEUE_REG_3__1_ & n16813;
  assign n17513 = P2_INSTQUEUE_REG_2__1_ & n16904;
  assign n17514 = P2_INSTQUEUE_REG_1__1_ & n16998;
  assign n17515 = P2_INSTQUEUE_REG_0__1_ & n17089;
  assign n17516 = ~n17512 & ~n17513;
  assign n17517 = ~n17514 & n17516;
  assign n17518 = ~n17515 & n17517;
  assign n17519 = n17497 & n17504;
  assign n17520 = n17511 & n17519;
  assign n17521 = n17518 & n17520;
  assign n17522 = ~n14238 & ~n17521;
  assign n17523 = n14238 & ~n14802;
  assign n17524 = ~n17522 & ~n17523;
  assign n17525 = n14238 & ~n17379;
  assign n17526 = ~n17524 & n17525;
  assign n17527 = ~n14238 & n17526;
  assign n17528 = ~n17524 & ~n17525;
  assign n17529 = n14238 & n17528;
  assign n17530 = ~n17527 & ~n17529;
  assign n17531 = n14238 & n17525;
  assign n17532 = ~n14238 & ~n17525;
  assign n17533 = ~n17531 & ~n17532;
  assign n17534 = n17524 & ~n17533;
  assign n17535 = n17530 & ~n17534;
  assign n17536 = ~n17490 & n17535;
  assign n17537 = ~P2_INSTADDRPOINTER_REG_1_ & ~n17487;
  assign n17538 = ~n17535 & n17537;
  assign n17539 = n17487 & ~n17535;
  assign n17540 = P2_INSTADDRPOINTER_REG_1_ & n17539;
  assign n17541 = ~n17536 & ~n17538;
  assign n17542 = ~n17540 & n17541;
  assign n17543 = n17413 & ~n17542;
  assign n17544 = P2_INSTADDRPOINTER_REG_0_ & ~n17454;
  assign n17545 = ~P2_INSTADDRPOINTER_REG_1_ & n17544;
  assign n17546 = P2_INSTADDRPOINTER_REG_1_ & ~n17544;
  assign n17547 = ~n17545 & ~n17546;
  assign n17548 = P2_EBX_REG_1_ & n14365;
  assign n17549 = ~n14365 & ~n14910;
  assign n17550 = ~n17548 & ~n17549;
  assign n17551 = n17449 & n17550;
  assign n17552 = ~n17449 & ~n17550;
  assign n17553 = ~n17551 & ~n17552;
  assign n17554 = ~n17445 & ~n17553;
  assign n17555 = n17445 & ~n17535;
  assign n17556 = ~n17554 & ~n17555;
  assign n17557 = ~n17547 & n17556;
  assign n17558 = ~P2_INSTADDRPOINTER_REG_1_ & ~n17544;
  assign n17559 = ~n17556 & n17558;
  assign n17560 = n17544 & ~n17556;
  assign n17561 = P2_INSTADDRPOINTER_REG_1_ & n17560;
  assign n17562 = ~n17557 & ~n17559;
  assign n17563 = ~n17561 & n17562;
  assign n17564 = n17458 & ~n17563;
  assign n17565 = P2_INSTADDRPOINTER_REG_1_ & n17410;
  assign n17566 = P2_REIP_REG_1_ & n17461;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = P2_INSTADDRPOINTER_REG_0_ & ~P2_INSTADDRPOINTER_REG_1_;
  assign n17569 = ~P2_INSTADDRPOINTER_REG_0_ & P2_INSTADDRPOINTER_REG_1_;
  assign n17570 = ~n17568 & ~n17569;
  assign n17571 = n17464 & ~n17570;
  assign n17572 = n17469 & ~n17570;
  assign n17573 = ~n17571 & ~n17572;
  assign n17574 = ~n15263 & n17476;
  assign n17575 = ~n17326 & n17480;
  assign n17576 = ~n17574 & ~n17575;
  assign n17577 = ~n17543 & ~n17564;
  assign n17578 = n17567 & n17577;
  assign n17579 = n17573 & n17578;
  assign n3879 = ~n17576 | ~n17579;
  assign n17581 = ~n17487 & n17535;
  assign n17582 = P2_INSTADDRPOINTER_REG_1_ & ~n17581;
  assign n17583 = ~n17539 & ~n17582;
  assign n17584 = n17524 & ~n17525;
  assign n17585 = ~n14238 & ~n17584;
  assign n17586 = ~n17526 & ~n17585;
  assign n17587 = P2_INSTQUEUE_REG_15__2_ & n15580;
  assign n17588 = P2_INSTQUEUE_REG_14__2_ & n15778;
  assign n17589 = P2_INSTQUEUE_REG_13__2_ & n15875;
  assign n17590 = P2_INSTQUEUE_REG_12__2_ & n15969;
  assign n17591 = ~n17587 & ~n17588;
  assign n17592 = ~n17589 & n17591;
  assign n17593 = ~n17590 & n17592;
  assign n17594 = P2_INSTQUEUE_REG_11__2_ & n16067;
  assign n17595 = P2_INSTQUEUE_REG_10__2_ & n16158;
  assign n17596 = P2_INSTQUEUE_REG_9__2_ & n16252;
  assign n17597 = P2_INSTQUEUE_REG_8__2_ & n16343;
  assign n17598 = ~n17594 & ~n17595;
  assign n17599 = ~n17596 & n17598;
  assign n17600 = ~n17597 & n17599;
  assign n17601 = P2_INSTQUEUE_REG_7__2_ & n16438;
  assign n17602 = P2_INSTQUEUE_REG_6__2_ & n16529;
  assign n17603 = P2_INSTQUEUE_REG_5__2_ & n16623;
  assign n17604 = P2_INSTQUEUE_REG_4__2_ & n16714;
  assign n17605 = ~n17601 & ~n17602;
  assign n17606 = ~n17603 & n17605;
  assign n17607 = ~n17604 & n17606;
  assign n17608 = P2_INSTQUEUE_REG_3__2_ & n16813;
  assign n17609 = P2_INSTQUEUE_REG_2__2_ & n16904;
  assign n17610 = P2_INSTQUEUE_REG_1__2_ & n16998;
  assign n17611 = P2_INSTQUEUE_REG_0__2_ & n17089;
  assign n17612 = ~n17608 & ~n17609;
  assign n17613 = ~n17610 & n17612;
  assign n17614 = ~n17611 & n17613;
  assign n17615 = n17593 & n17600;
  assign n17616 = n17607 & n17615;
  assign n17617 = n17614 & n17616;
  assign n17618 = ~n14238 & ~n17617;
  assign n17619 = n14238 & ~n14722;
  assign n17620 = ~n17618 & ~n17619;
  assign n17621 = ~n14238 & ~n17620;
  assign n17622 = n14238 & n17620;
  assign n17623 = ~n17621 & ~n17622;
  assign n17624 = n17586 & ~n17623;
  assign n17625 = ~n17586 & n17623;
  assign n17626 = ~n17624 & ~n17625;
  assign n17627 = ~P2_INSTADDRPOINTER_REG_2_ & ~n17626;
  assign n17628 = P2_INSTADDRPOINTER_REG_2_ & n17626;
  assign n17629 = ~n17627 & ~n17628;
  assign n17630 = n17583 & ~n17629;
  assign n17631 = ~n17583 & n17629;
  assign n17632 = ~n17630 & ~n17631;
  assign n17633 = n17413 & ~n17632;
  assign n17634 = P2_INSTADDRPOINTER_REG_1_ & n17544;
  assign n17635 = P2_INSTADDRPOINTER_REG_1_ & ~n17556;
  assign n17636 = ~n17560 & ~n17634;
  assign n17637 = ~n17635 & n17636;
  assign n17638 = ~n17449 & n17550;
  assign n17639 = P2_EBX_REG_2_ & n14365;
  assign n17640 = ~n14365 & ~n14902;
  assign n17641 = ~n17639 & ~n17640;
  assign n17642 = n17638 & n17641;
  assign n17643 = ~n17638 & ~n17641;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = ~n17445 & n17644;
  assign n17646 = n17445 & ~n17626;
  assign n17647 = ~n17645 & ~n17646;
  assign n17648 = ~P2_INSTADDRPOINTER_REG_2_ & ~n17647;
  assign n17649 = P2_INSTADDRPOINTER_REG_2_ & n17647;
  assign n17650 = ~n17648 & ~n17649;
  assign n17651 = n17637 & ~n17650;
  assign n17652 = ~n17637 & n17650;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = n17458 & ~n17653;
  assign n17655 = P2_INSTADDRPOINTER_REG_2_ & n17410;
  assign n17656 = P2_REIP_REG_2_ & n17461;
  assign n17657 = ~n17655 & ~n17656;
  assign n17658 = P2_INSTADDRPOINTER_REG_0_ & P2_INSTADDRPOINTER_REG_1_;
  assign n17659 = ~P2_INSTADDRPOINTER_REG_2_ & ~n17658;
  assign n17660 = P2_INSTADDRPOINTER_REG_2_ & n17658;
  assign n17661 = ~n17659 & ~n17660;
  assign n17662 = n17464 & ~n17661;
  assign n17663 = ~P2_INSTADDRPOINTER_REG_2_ & n17658;
  assign n17664 = P2_INSTADDRPOINTER_REG_2_ & ~n17658;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = n17469 & ~n17665;
  assign n17667 = ~n17662 & ~n17666;
  assign n17668 = ~n15216 & n17476;
  assign n17669 = ~n17306 & n17480;
  assign n17670 = ~n17668 & ~n17669;
  assign n17671 = ~n17633 & ~n17654;
  assign n17672 = n17657 & n17671;
  assign n17673 = n17667 & n17672;
  assign n3884 = ~n17670 | ~n17673;
  assign n17675 = P2_INSTADDRPOINTER_REG_2_ & ~n17626;
  assign n17676 = ~P2_INSTADDRPOINTER_REG_2_ & n17626;
  assign n17677 = ~n17583 & ~n17676;
  assign n17678 = ~n17675 & ~n17677;
  assign n17679 = n14238 & ~n17620;
  assign n17680 = ~n14238 & n17620;
  assign n17681 = ~n17586 & ~n17680;
  assign n17682 = ~n17679 & ~n17681;
  assign n17683 = P2_INSTQUEUE_REG_15__3_ & n15580;
  assign n17684 = P2_INSTQUEUE_REG_14__3_ & n15778;
  assign n17685 = P2_INSTQUEUE_REG_13__3_ & n15875;
  assign n17686 = P2_INSTQUEUE_REG_12__3_ & n15969;
  assign n17687 = ~n17683 & ~n17684;
  assign n17688 = ~n17685 & n17687;
  assign n17689 = ~n17686 & n17688;
  assign n17690 = P2_INSTQUEUE_REG_11__3_ & n16067;
  assign n17691 = P2_INSTQUEUE_REG_10__3_ & n16158;
  assign n17692 = P2_INSTQUEUE_REG_9__3_ & n16252;
  assign n17693 = P2_INSTQUEUE_REG_8__3_ & n16343;
  assign n17694 = ~n17690 & ~n17691;
  assign n17695 = ~n17692 & n17694;
  assign n17696 = ~n17693 & n17695;
  assign n17697 = P2_INSTQUEUE_REG_7__3_ & n16438;
  assign n17698 = P2_INSTQUEUE_REG_6__3_ & n16529;
  assign n17699 = P2_INSTQUEUE_REG_5__3_ & n16623;
  assign n17700 = P2_INSTQUEUE_REG_4__3_ & n16714;
  assign n17701 = ~n17697 & ~n17698;
  assign n17702 = ~n17699 & n17701;
  assign n17703 = ~n17700 & n17702;
  assign n17704 = P2_INSTQUEUE_REG_3__3_ & n16813;
  assign n17705 = P2_INSTQUEUE_REG_2__3_ & n16904;
  assign n17706 = P2_INSTQUEUE_REG_1__3_ & n16998;
  assign n17707 = P2_INSTQUEUE_REG_0__3_ & n17089;
  assign n17708 = ~n17704 & ~n17705;
  assign n17709 = ~n17706 & n17708;
  assign n17710 = ~n17707 & n17709;
  assign n17711 = n17689 & n17696;
  assign n17712 = n17703 & n17711;
  assign n17713 = n17710 & n17712;
  assign n17714 = ~n14238 & ~n17713;
  assign n17715 = n14238 & ~n14685;
  assign n17716 = ~n17714 & ~n17715;
  assign n17717 = n17682 & n17716;
  assign n17718 = ~n17682 & ~n17716;
  assign n17719 = ~n17717 & ~n17718;
  assign n17720 = ~P2_INSTADDRPOINTER_REG_3_ & n17719;
  assign n17721 = P2_INSTADDRPOINTER_REG_3_ & ~n17719;
  assign n17722 = ~n17720 & ~n17721;
  assign n17723 = n17678 & ~n17722;
  assign n17724 = ~n17678 & n17722;
  assign n17725 = ~n17723 & ~n17724;
  assign n17726 = n17413 & ~n17725;
  assign n17727 = P2_INSTADDRPOINTER_REG_2_ & ~n17647;
  assign n17728 = ~P2_INSTADDRPOINTER_REG_2_ & n17647;
  assign n17729 = ~n17637 & ~n17728;
  assign n17730 = ~n17727 & ~n17729;
  assign n17731 = P2_EBX_REG_3_ & n14365;
  assign n17732 = ~n14365 & ~n14888;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = ~n17642 & ~n17733;
  assign n17735 = n17642 & n17733;
  assign n17736 = ~n17734 & ~n17735;
  assign n17737 = ~n17445 & n17736;
  assign n17738 = n17445 & n17719;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = ~P2_INSTADDRPOINTER_REG_3_ & ~n17739;
  assign n17741 = P2_INSTADDRPOINTER_REG_3_ & n17739;
  assign n17742 = ~n17740 & ~n17741;
  assign n17743 = n17730 & ~n17742;
  assign n17744 = ~n17730 & n17742;
  assign n17745 = ~n17743 & ~n17744;
  assign n17746 = n17458 & ~n17745;
  assign n17747 = P2_INSTADDRPOINTER_REG_3_ & n17410;
  assign n17748 = P2_REIP_REG_3_ & n17461;
  assign n17749 = ~n17747 & ~n17748;
  assign n17750 = ~P2_INSTADDRPOINTER_REG_3_ & n17659;
  assign n17751 = P2_INSTADDRPOINTER_REG_3_ & ~n17659;
  assign n17752 = ~n17750 & ~n17751;
  assign n17753 = n17464 & n17752;
  assign n17754 = ~P2_INSTADDRPOINTER_REG_3_ & n17660;
  assign n17755 = P2_INSTADDRPOINTER_REG_3_ & ~n17660;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = n17469 & ~n17756;
  assign n17758 = ~n17753 & ~n17757;
  assign n17759 = ~n15147 & n17476;
  assign n17760 = ~n17289 & n17480;
  assign n17761 = ~n17759 & ~n17760;
  assign n17762 = ~n17726 & ~n17746;
  assign n17763 = n17749 & n17762;
  assign n17764 = n17758 & n17763;
  assign n3889 = ~n17761 | ~n17764;
  assign n17766 = P2_INSTADDRPOINTER_REG_3_ & n17719;
  assign n17767 = ~P2_INSTADDRPOINTER_REG_3_ & ~n17719;
  assign n17768 = ~n17678 & ~n17767;
  assign n17769 = ~n17766 & ~n17768;
  assign n17770 = P2_INSTQUEUE_REG_15__4_ & n15580;
  assign n17771 = P2_INSTQUEUE_REG_14__4_ & n15778;
  assign n17772 = P2_INSTQUEUE_REG_13__4_ & n15875;
  assign n17773 = P2_INSTQUEUE_REG_12__4_ & n15969;
  assign n17774 = ~n17770 & ~n17771;
  assign n17775 = ~n17772 & n17774;
  assign n17776 = ~n17773 & n17775;
  assign n17777 = P2_INSTQUEUE_REG_11__4_ & n16067;
  assign n17778 = P2_INSTQUEUE_REG_10__4_ & n16158;
  assign n17779 = P2_INSTQUEUE_REG_9__4_ & n16252;
  assign n17780 = P2_INSTQUEUE_REG_8__4_ & n16343;
  assign n17781 = ~n17777 & ~n17778;
  assign n17782 = ~n17779 & n17781;
  assign n17783 = ~n17780 & n17782;
  assign n17784 = P2_INSTQUEUE_REG_7__4_ & n16438;
  assign n17785 = P2_INSTQUEUE_REG_6__4_ & n16529;
  assign n17786 = P2_INSTQUEUE_REG_5__4_ & n16623;
  assign n17787 = P2_INSTQUEUE_REG_4__4_ & n16714;
  assign n17788 = ~n17784 & ~n17785;
  assign n17789 = ~n17786 & n17788;
  assign n17790 = ~n17787 & n17789;
  assign n17791 = P2_INSTQUEUE_REG_3__4_ & n16813;
  assign n17792 = P2_INSTQUEUE_REG_2__4_ & n16904;
  assign n17793 = P2_INSTQUEUE_REG_1__4_ & n16998;
  assign n17794 = P2_INSTQUEUE_REG_0__4_ & n17089;
  assign n17795 = ~n17791 & ~n17792;
  assign n17796 = ~n17793 & n17795;
  assign n17797 = ~n17794 & n17796;
  assign n17798 = n17776 & n17783;
  assign n17799 = n17790 & n17798;
  assign n17800 = n17797 & n17799;
  assign n17801 = ~n14238 & ~n17800;
  assign n17802 = n14238 & ~n14760;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = n17718 & n17803;
  assign n17805 = ~n17718 & ~n17803;
  assign n17806 = ~n17804 & ~n17805;
  assign n17807 = ~P2_INSTADDRPOINTER_REG_4_ & ~n17806;
  assign n17808 = P2_INSTADDRPOINTER_REG_4_ & n17806;
  assign n17809 = ~n17807 & ~n17808;
  assign n17810 = n17769 & ~n17809;
  assign n17811 = ~n17769 & n17809;
  assign n17812 = ~n17810 & ~n17811;
  assign n17813 = n17413 & ~n17812;
  assign n17814 = ~P2_INSTADDRPOINTER_REG_3_ & n17739;
  assign n17815 = n17727 & ~n17814;
  assign n17816 = P2_INSTADDRPOINTER_REG_3_ & ~n17739;
  assign n17817 = ~n17815 & ~n17816;
  assign n17818 = ~n17728 & ~n17814;
  assign n17819 = ~n17637 & n17818;
  assign n17820 = n17817 & ~n17819;
  assign n17821 = P2_EBX_REG_4_ & n14365;
  assign n17822 = ~n14365 & ~n14880;
  assign n17823 = ~n17821 & ~n17822;
  assign n17824 = n17735 & n17823;
  assign n17825 = ~n17735 & ~n17823;
  assign n17826 = ~n17824 & ~n17825;
  assign n17827 = ~n17445 & n17826;
  assign n17828 = n17445 & ~n17806;
  assign n17829 = ~n17827 & ~n17828;
  assign n17830 = ~P2_INSTADDRPOINTER_REG_4_ & ~n17829;
  assign n17831 = P2_INSTADDRPOINTER_REG_4_ & n17829;
  assign n17832 = ~n17830 & ~n17831;
  assign n17833 = n17820 & ~n17832;
  assign n17834 = ~n17820 & n17832;
  assign n17835 = ~n17833 & ~n17834;
  assign n17836 = n17458 & ~n17835;
  assign n17837 = P2_INSTADDRPOINTER_REG_4_ & n17410;
  assign n17838 = P2_REIP_REG_4_ & n17461;
  assign n17839 = ~n17837 & ~n17838;
  assign n17840 = ~P2_INSTADDRPOINTER_REG_4_ & n17751;
  assign n17841 = P2_INSTADDRPOINTER_REG_4_ & ~n17751;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = n17464 & ~n17842;
  assign n17844 = P2_INSTADDRPOINTER_REG_3_ & n17660;
  assign n17845 = ~P2_INSTADDRPOINTER_REG_4_ & n17844;
  assign n17846 = P2_INSTADDRPOINTER_REG_4_ & ~n17844;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = n17469 & ~n17847;
  assign n17849 = ~n17843 & ~n17848;
  assign n17850 = ~n15134 & ~n15141;
  assign n17851 = n15134 & n15141;
  assign n17852 = ~n15131 & ~n17851;
  assign n17853 = ~n17850 & ~n17852;
  assign n17854 = P2_EBX_REG_4_ & n14995;
  assign n17855 = P2_REIP_REG_4_ & n14997;
  assign n17856 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_4_;
  assign n17857 = P2_INSTADDRPOINTER_REG_4_ & ~n15016;
  assign n17858 = ~n17854 & ~n17855;
  assign n17859 = ~n17856 & n17858;
  assign n17860 = ~n17857 & n17859;
  assign n17861 = n17853 & n17860;
  assign n17862 = ~n17853 & ~n17860;
  assign n17863 = ~n17861 & ~n17862;
  assign n17864 = n17476 & n17863;
  assign n17865 = ~n17278 & ~n17283;
  assign n17866 = n17278 & n17283;
  assign n17867 = ~n17275 & ~n17866;
  assign n17868 = ~n17865 & ~n17867;
  assign n17869 = ~n14760 & n17242;
  assign n17870 = P2_REIP_REG_4_ & n17226;
  assign n17871 = P2_EAX_REG_4_ & n17228;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = P2_INSTADDRPOINTER_REG_4_ & ~n17236;
  assign n17874 = n17872 & ~n17873;
  assign n17875 = n17869 & n17874;
  assign n17876 = ~n17869 & ~n17874;
  assign n17877 = ~n17875 & ~n17876;
  assign n17878 = n17868 & ~n17877;
  assign n17879 = ~n17868 & n17877;
  assign n17880 = ~n17878 & ~n17879;
  assign n17881 = n17480 & ~n17880;
  assign n17882 = ~n17864 & ~n17881;
  assign n17883 = ~n17813 & ~n17836;
  assign n17884 = n17839 & n17883;
  assign n17885 = n17849 & n17884;
  assign n3894 = ~n17882 | ~n17885;
  assign n17887 = P2_INSTADDRPOINTER_REG_4_ & ~n17806;
  assign n17888 = ~P2_INSTADDRPOINTER_REG_4_ & n17806;
  assign n17889 = ~n17769 & ~n17888;
  assign n17890 = ~n17887 & ~n17889;
  assign n17891 = n17718 & ~n17803;
  assign n17892 = P2_INSTQUEUE_REG_15__5_ & n15580;
  assign n17893 = P2_INSTQUEUE_REG_14__5_ & n15778;
  assign n17894 = P2_INSTQUEUE_REG_13__5_ & n15875;
  assign n17895 = P2_INSTQUEUE_REG_12__5_ & n15969;
  assign n17896 = ~n17892 & ~n17893;
  assign n17897 = ~n17894 & n17896;
  assign n17898 = ~n17895 & n17897;
  assign n17899 = P2_INSTQUEUE_REG_11__5_ & n16067;
  assign n17900 = P2_INSTQUEUE_REG_10__5_ & n16158;
  assign n17901 = P2_INSTQUEUE_REG_9__5_ & n16252;
  assign n17902 = P2_INSTQUEUE_REG_8__5_ & n16343;
  assign n17903 = ~n17899 & ~n17900;
  assign n17904 = ~n17901 & n17903;
  assign n17905 = ~n17902 & n17904;
  assign n17906 = P2_INSTQUEUE_REG_7__5_ & n16438;
  assign n17907 = P2_INSTQUEUE_REG_6__5_ & n16529;
  assign n17908 = P2_INSTQUEUE_REG_5__5_ & n16623;
  assign n17909 = P2_INSTQUEUE_REG_4__5_ & n16714;
  assign n17910 = ~n17906 & ~n17907;
  assign n17911 = ~n17908 & n17910;
  assign n17912 = ~n17909 & n17911;
  assign n17913 = P2_INSTQUEUE_REG_3__5_ & n16813;
  assign n17914 = P2_INSTQUEUE_REG_2__5_ & n16904;
  assign n17915 = P2_INSTQUEUE_REG_1__5_ & n16998;
  assign n17916 = P2_INSTQUEUE_REG_0__5_ & n17089;
  assign n17917 = ~n17913 & ~n17914;
  assign n17918 = ~n17915 & n17917;
  assign n17919 = ~n17916 & n17918;
  assign n17920 = n17898 & n17905;
  assign n17921 = n17912 & n17920;
  assign n17922 = n17919 & n17921;
  assign n17923 = ~n14238 & ~n17922;
  assign n17924 = n14238 & ~n14647;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = n17891 & n17925;
  assign n17927 = ~n17891 & ~n17925;
  assign n17928 = ~n17926 & ~n17927;
  assign n17929 = ~P2_INSTADDRPOINTER_REG_5_ & ~n17928;
  assign n17930 = P2_INSTADDRPOINTER_REG_5_ & n17928;
  assign n17931 = ~n17929 & ~n17930;
  assign n17932 = n17890 & ~n17931;
  assign n17933 = ~n17890 & n17931;
  assign n17934 = ~n17932 & ~n17933;
  assign n17935 = n17413 & ~n17934;
  assign n17936 = P2_INSTADDRPOINTER_REG_4_ & ~n17829;
  assign n17937 = ~P2_INSTADDRPOINTER_REG_4_ & n17829;
  assign n17938 = ~n17820 & ~n17937;
  assign n17939 = ~n17936 & ~n17938;
  assign n17940 = P2_EBX_REG_5_ & n14365;
  assign n17941 = ~n14365 & ~n14869;
  assign n17942 = ~n17940 & ~n17941;
  assign n17943 = ~n17824 & ~n17942;
  assign n17944 = n17824 & n17942;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = ~n17445 & n17945;
  assign n17947 = n17445 & ~n17928;
  assign n17948 = ~n17946 & ~n17947;
  assign n17949 = ~P2_INSTADDRPOINTER_REG_5_ & ~n17948;
  assign n17950 = P2_INSTADDRPOINTER_REG_5_ & n17948;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 = n17939 & ~n17951;
  assign n17953 = ~n17939 & n17951;
  assign n17954 = ~n17952 & ~n17953;
  assign n17955 = n17458 & ~n17954;
  assign n17956 = P2_INSTADDRPOINTER_REG_5_ & n17410;
  assign n17957 = P2_REIP_REG_5_ & n17461;
  assign n17958 = ~n17956 & ~n17957;
  assign n17959 = P2_INSTADDRPOINTER_REG_4_ & n17751;
  assign n17960 = ~P2_INSTADDRPOINTER_REG_5_ & n17959;
  assign n17961 = P2_INSTADDRPOINTER_REG_5_ & ~n17959;
  assign n17962 = ~n17960 & ~n17961;
  assign n17963 = n17464 & ~n17962;
  assign n17964 = P2_INSTADDRPOINTER_REG_4_ & n17844;
  assign n17965 = ~P2_INSTADDRPOINTER_REG_5_ & n17964;
  assign n17966 = P2_INSTADDRPOINTER_REG_5_ & ~n17964;
  assign n17967 = ~n17965 & ~n17966;
  assign n17968 = n17469 & ~n17967;
  assign n17969 = ~n17963 & ~n17968;
  assign n17970 = P2_EBX_REG_5_ & n14995;
  assign n17971 = P2_REIP_REG_5_ & n14997;
  assign n17972 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_5_;
  assign n17973 = P2_INSTADDRPOINTER_REG_5_ & ~n15016;
  assign n17974 = ~n17970 & ~n17971;
  assign n17975 = ~n17972 & n17974;
  assign n17976 = ~n17973 & n17975;
  assign n17977 = n17862 & n17976;
  assign n17978 = ~n17862 & ~n17976;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 = n17476 & ~n17979;
  assign n17981 = n17869 & ~n17874;
  assign n17982 = ~n17869 & n17874;
  assign n17983 = ~n17868 & ~n17982;
  assign n17984 = ~n17981 & ~n17983;
  assign n17985 = ~n14647 & n17242;
  assign n17986 = P2_REIP_REG_5_ & n17226;
  assign n17987 = P2_EAX_REG_5_ & n17228;
  assign n17988 = ~n17986 & ~n17987;
  assign n17989 = P2_INSTADDRPOINTER_REG_5_ & ~n17236;
  assign n17990 = n17988 & ~n17989;
  assign n17991 = n17985 & n17990;
  assign n17992 = ~n17985 & ~n17990;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 = n17984 & ~n17993;
  assign n17995 = ~n17984 & n17993;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = n17480 & ~n17996;
  assign n17998 = ~n17980 & ~n17997;
  assign n17999 = ~n17935 & ~n17955;
  assign n18000 = n17958 & n17999;
  assign n18001 = n17969 & n18000;
  assign n3899 = ~n17998 | ~n18001;
  assign n18003 = P2_INSTADDRPOINTER_REG_5_ & ~n17928;
  assign n18004 = ~P2_INSTADDRPOINTER_REG_5_ & n17928;
  assign n18005 = ~n17890 & ~n18004;
  assign n18006 = ~n18003 & ~n18005;
  assign n18007 = n17891 & ~n17925;
  assign n18008 = P2_INSTQUEUE_REG_15__6_ & n15580;
  assign n18009 = P2_INSTQUEUE_REG_14__6_ & n15778;
  assign n18010 = P2_INSTQUEUE_REG_13__6_ & n15875;
  assign n18011 = P2_INSTQUEUE_REG_12__6_ & n15969;
  assign n18012 = ~n18008 & ~n18009;
  assign n18013 = ~n18010 & n18012;
  assign n18014 = ~n18011 & n18013;
  assign n18015 = P2_INSTQUEUE_REG_11__6_ & n16067;
  assign n18016 = P2_INSTQUEUE_REG_10__6_ & n16158;
  assign n18017 = P2_INSTQUEUE_REG_9__6_ & n16252;
  assign n18018 = P2_INSTQUEUE_REG_8__6_ & n16343;
  assign n18019 = ~n18015 & ~n18016;
  assign n18020 = ~n18017 & n18019;
  assign n18021 = ~n18018 & n18020;
  assign n18022 = P2_INSTQUEUE_REG_7__6_ & n16438;
  assign n18023 = P2_INSTQUEUE_REG_6__6_ & n16529;
  assign n18024 = P2_INSTQUEUE_REG_5__6_ & n16623;
  assign n18025 = P2_INSTQUEUE_REG_4__6_ & n16714;
  assign n18026 = ~n18022 & ~n18023;
  assign n18027 = ~n18024 & n18026;
  assign n18028 = ~n18025 & n18027;
  assign n18029 = P2_INSTQUEUE_REG_3__6_ & n16813;
  assign n18030 = P2_INSTQUEUE_REG_2__6_ & n16904;
  assign n18031 = P2_INSTQUEUE_REG_1__6_ & n16998;
  assign n18032 = P2_INSTQUEUE_REG_0__6_ & n17089;
  assign n18033 = ~n18029 & ~n18030;
  assign n18034 = ~n18031 & n18033;
  assign n18035 = ~n18032 & n18034;
  assign n18036 = n18014 & n18021;
  assign n18037 = n18028 & n18036;
  assign n18038 = n18035 & n18037;
  assign n18039 = ~n14238 & ~n18038;
  assign n18040 = n14238 & ~n14612;
  assign n18041 = ~n18039 & ~n18040;
  assign n18042 = n18007 & n18041;
  assign n18043 = ~n18007 & ~n18041;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = ~P2_INSTADDRPOINTER_REG_6_ & ~n18044;
  assign n18046 = P2_INSTADDRPOINTER_REG_6_ & n18044;
  assign n18047 = ~n18045 & ~n18046;
  assign n18048 = n18006 & ~n18047;
  assign n18049 = ~n18006 & n18047;
  assign n18050 = ~n18048 & ~n18049;
  assign n18051 = n17413 & ~n18050;
  assign n18052 = ~P2_INSTADDRPOINTER_REG_5_ & n17948;
  assign n18053 = n17936 & ~n18052;
  assign n18054 = P2_INSTADDRPOINTER_REG_5_ & ~n17948;
  assign n18055 = ~n18053 & ~n18054;
  assign n18056 = ~n17937 & ~n18052;
  assign n18057 = ~n17820 & n18056;
  assign n18058 = n18055 & ~n18057;
  assign n18059 = P2_EBX_REG_6_ & n14365;
  assign n18060 = ~n14365 & ~n14855;
  assign n18061 = ~n18059 & ~n18060;
  assign n18062 = n17944 & n18061;
  assign n18063 = ~n17944 & ~n18061;
  assign n18064 = ~n18062 & ~n18063;
  assign n18065 = ~n17445 & n18064;
  assign n18066 = n17445 & ~n18044;
  assign n18067 = ~n18065 & ~n18066;
  assign n18068 = ~P2_INSTADDRPOINTER_REG_6_ & ~n18067;
  assign n18069 = P2_INSTADDRPOINTER_REG_6_ & n18067;
  assign n18070 = ~n18068 & ~n18069;
  assign n18071 = n18058 & ~n18070;
  assign n18072 = ~n18058 & n18070;
  assign n18073 = ~n18071 & ~n18072;
  assign n18074 = n17458 & ~n18073;
  assign n18075 = P2_INSTADDRPOINTER_REG_6_ & n17410;
  assign n18076 = P2_REIP_REG_6_ & n17461;
  assign n18077 = ~n18075 & ~n18076;
  assign n18078 = P2_INSTADDRPOINTER_REG_5_ & n17959;
  assign n18079 = ~P2_INSTADDRPOINTER_REG_6_ & n18078;
  assign n18080 = P2_INSTADDRPOINTER_REG_6_ & ~n18078;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = n17464 & ~n18081;
  assign n18083 = P2_INSTADDRPOINTER_REG_5_ & n17964;
  assign n18084 = ~P2_INSTADDRPOINTER_REG_6_ & n18083;
  assign n18085 = P2_INSTADDRPOINTER_REG_6_ & ~n18083;
  assign n18086 = ~n18084 & ~n18085;
  assign n18087 = n17469 & ~n18086;
  assign n18088 = ~n18082 & ~n18087;
  assign n18089 = n17862 & ~n17976;
  assign n18090 = P2_EBX_REG_6_ & n14995;
  assign n18091 = P2_REIP_REG_6_ & n14997;
  assign n18092 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_6_;
  assign n18093 = P2_INSTADDRPOINTER_REG_6_ & ~n15016;
  assign n18094 = ~n18090 & ~n18091;
  assign n18095 = ~n18092 & n18094;
  assign n18096 = ~n18093 & n18095;
  assign n18097 = n18089 & n18096;
  assign n18098 = ~n18089 & ~n18096;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = n17476 & ~n18099;
  assign n18101 = n17985 & ~n17990;
  assign n18102 = ~n17985 & n17990;
  assign n18103 = ~n17984 & ~n18102;
  assign n18104 = ~n18101 & ~n18103;
  assign n18105 = ~n14612 & n17242;
  assign n18106 = P2_REIP_REG_6_ & n17226;
  assign n18107 = P2_EAX_REG_6_ & n17228;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = P2_INSTADDRPOINTER_REG_6_ & ~n17236;
  assign n18110 = n18108 & ~n18109;
  assign n18111 = n18105 & n18110;
  assign n18112 = ~n18105 & ~n18110;
  assign n18113 = ~n18111 & ~n18112;
  assign n18114 = n18104 & ~n18113;
  assign n18115 = ~n18104 & n18113;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = n17480 & ~n18116;
  assign n18118 = ~n18100 & ~n18117;
  assign n18119 = ~n18051 & ~n18074;
  assign n18120 = n18077 & n18119;
  assign n18121 = n18088 & n18120;
  assign n3904 = ~n18118 | ~n18121;
  assign n18123 = P2_INSTADDRPOINTER_REG_6_ & ~n18044;
  assign n18124 = ~P2_INSTADDRPOINTER_REG_6_ & n18044;
  assign n18125 = ~n18006 & ~n18124;
  assign n18126 = ~n18123 & ~n18125;
  assign n18127 = n18007 & ~n18041;
  assign n18128 = P2_INSTQUEUE_REG_15__7_ & n15580;
  assign n18129 = P2_INSTQUEUE_REG_14__7_ & n15778;
  assign n18130 = P2_INSTQUEUE_REG_13__7_ & n15875;
  assign n18131 = P2_INSTQUEUE_REG_12__7_ & n15969;
  assign n18132 = ~n18128 & ~n18129;
  assign n18133 = ~n18130 & n18132;
  assign n18134 = ~n18131 & n18133;
  assign n18135 = P2_INSTQUEUE_REG_11__7_ & n16067;
  assign n18136 = P2_INSTQUEUE_REG_10__7_ & n16158;
  assign n18137 = P2_INSTQUEUE_REG_9__7_ & n16252;
  assign n18138 = P2_INSTQUEUE_REG_8__7_ & n16343;
  assign n18139 = ~n18135 & ~n18136;
  assign n18140 = ~n18137 & n18139;
  assign n18141 = ~n18138 & n18140;
  assign n18142 = P2_INSTQUEUE_REG_7__7_ & n16438;
  assign n18143 = P2_INSTQUEUE_REG_6__7_ & n16529;
  assign n18144 = P2_INSTQUEUE_REG_5__7_ & n16623;
  assign n18145 = P2_INSTQUEUE_REG_4__7_ & n16714;
  assign n18146 = ~n18142 & ~n18143;
  assign n18147 = ~n18144 & n18146;
  assign n18148 = ~n18145 & n18147;
  assign n18149 = P2_INSTQUEUE_REG_3__7_ & n16813;
  assign n18150 = P2_INSTQUEUE_REG_2__7_ & n16904;
  assign n18151 = P2_INSTQUEUE_REG_1__7_ & n16998;
  assign n18152 = P2_INSTQUEUE_REG_0__7_ & n17089;
  assign n18153 = ~n18149 & ~n18150;
  assign n18154 = ~n18151 & n18153;
  assign n18155 = ~n18152 & n18154;
  assign n18156 = n18134 & n18141;
  assign n18157 = n18148 & n18156;
  assign n18158 = n18155 & n18157;
  assign n18159 = ~n14238 & ~n18158;
  assign n18160 = n14238 & ~n17445;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = n18127 & n18161;
  assign n18163 = ~n18127 & ~n18161;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = ~P2_INSTADDRPOINTER_REG_7_ & ~n18164;
  assign n18166 = P2_INSTADDRPOINTER_REG_7_ & n18164;
  assign n18167 = ~n18165 & ~n18166;
  assign n18168 = n18126 & ~n18167;
  assign n18169 = ~n18126 & n18167;
  assign n18170 = ~n18168 & ~n18169;
  assign n18171 = n17413 & ~n18170;
  assign n18172 = P2_INSTADDRPOINTER_REG_6_ & ~n18067;
  assign n18173 = ~P2_INSTADDRPOINTER_REG_6_ & n18067;
  assign n18174 = ~n18058 & ~n18173;
  assign n18175 = ~n18172 & ~n18174;
  assign n18176 = P2_EBX_REG_7_ & n14365;
  assign n18177 = n14244 & ~n17445;
  assign n18178 = n14244 & ~n18177;
  assign n18179 = ~n14244 & n18177;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~n14615 & ~n14852;
  assign n18182 = ~n14614 & ~n18181;
  assign n18183 = ~n18180 & ~n18182;
  assign n18184 = n18180 & n18182;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 = ~n14365 & ~n18185;
  assign n18187 = ~n18176 & ~n18186;
  assign n18188 = ~n18062 & ~n18187;
  assign n18189 = n18062 & n18187;
  assign n18190 = ~n18188 & ~n18189;
  assign n18191 = ~n17445 & n18190;
  assign n18192 = n17445 & ~n18164;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = ~P2_INSTADDRPOINTER_REG_7_ & ~n18193;
  assign n18195 = P2_INSTADDRPOINTER_REG_7_ & n18193;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = n18175 & ~n18196;
  assign n18198 = ~n18175 & n18196;
  assign n18199 = ~n18197 & ~n18198;
  assign n18200 = n17458 & ~n18199;
  assign n18201 = P2_INSTADDRPOINTER_REG_7_ & n17410;
  assign n18202 = P2_REIP_REG_7_ & n17461;
  assign n18203 = ~n18201 & ~n18202;
  assign n18204 = P2_INSTADDRPOINTER_REG_6_ & n18078;
  assign n18205 = ~P2_INSTADDRPOINTER_REG_7_ & n18204;
  assign n18206 = P2_INSTADDRPOINTER_REG_7_ & ~n18204;
  assign n18207 = ~n18205 & ~n18206;
  assign n18208 = n17464 & ~n18207;
  assign n18209 = P2_INSTADDRPOINTER_REG_6_ & n18083;
  assign n18210 = ~P2_INSTADDRPOINTER_REG_7_ & n18209;
  assign n18211 = P2_INSTADDRPOINTER_REG_7_ & ~n18209;
  assign n18212 = ~n18210 & ~n18211;
  assign n18213 = n17469 & ~n18212;
  assign n18214 = ~n18208 & ~n18213;
  assign n18215 = n18089 & ~n18096;
  assign n18216 = P2_EBX_REG_7_ & n14995;
  assign n18217 = P2_REIP_REG_7_ & n14997;
  assign n18218 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_7_;
  assign n18219 = P2_INSTADDRPOINTER_REG_7_ & ~n15016;
  assign n18220 = ~n18216 & ~n18217;
  assign n18221 = ~n18218 & n18220;
  assign n18222 = ~n18219 & n18221;
  assign n18223 = n18215 & n18222;
  assign n18224 = ~n18215 & ~n18222;
  assign n18225 = ~n18223 & ~n18224;
  assign n18226 = n17476 & ~n18225;
  assign n18227 = n18105 & ~n18110;
  assign n18228 = ~n18105 & n18110;
  assign n18229 = ~n18104 & ~n18228;
  assign n18230 = ~n18227 & ~n18229;
  assign n18231 = n17242 & ~n17445;
  assign n18232 = P2_REIP_REG_7_ & n17226;
  assign n18233 = P2_EAX_REG_7_ & n17228;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = P2_INSTADDRPOINTER_REG_7_ & ~n17236;
  assign n18236 = n18234 & ~n18235;
  assign n18237 = n18231 & n18236;
  assign n18238 = ~n18231 & ~n18236;
  assign n18239 = ~n18237 & ~n18238;
  assign n18240 = n18230 & ~n18239;
  assign n18241 = ~n18230 & n18239;
  assign n18242 = ~n18240 & ~n18241;
  assign n18243 = n17480 & ~n18242;
  assign n18244 = ~n18226 & ~n18243;
  assign n18245 = ~n18171 & ~n18200;
  assign n18246 = n18203 & n18245;
  assign n18247 = n18214 & n18246;
  assign n3909 = ~n18244 | ~n18247;
  assign n18249 = P2_INSTADDRPOINTER_REG_7_ & ~n18164;
  assign n18250 = ~P2_INSTADDRPOINTER_REG_7_ & n18164;
  assign n18251 = ~n18126 & ~n18250;
  assign n18252 = ~n18249 & ~n18251;
  assign n18253 = ~n18041 & ~n18161;
  assign n18254 = n18007 & n18253;
  assign n18255 = ~P2_INSTADDRPOINTER_REG_8_ & n18254;
  assign n18256 = P2_INSTADDRPOINTER_REG_8_ & ~n18254;
  assign n18257 = ~n18255 & ~n18256;
  assign n18258 = n18252 & ~n18257;
  assign n18259 = ~n18252 & n18257;
  assign n18260 = ~n18258 & ~n18259;
  assign n18261 = n17413 & ~n18260;
  assign n18262 = ~P2_INSTADDRPOINTER_REG_7_ & n18193;
  assign n18263 = n18172 & ~n18262;
  assign n18264 = P2_INSTADDRPOINTER_REG_7_ & ~n18193;
  assign n18265 = ~n18263 & ~n18264;
  assign n18266 = ~n18173 & ~n18262;
  assign n18267 = ~n18058 & n18266;
  assign n18268 = n18265 & ~n18267;
  assign n18269 = ~n18179 & ~n18182;
  assign n18270 = ~n18178 & ~n18269;
  assign n18271 = ~n14365 & n18270;
  assign n18272 = P2_EBX_REG_8_ & n14365;
  assign n18273 = ~n18271 & ~n18272;
  assign n18274 = n18189 & n18273;
  assign n18275 = ~n18189 & ~n18273;
  assign n18276 = ~n18274 & ~n18275;
  assign n18277 = ~n17445 & n18276;
  assign n18278 = n17445 & n18254;
  assign n18279 = ~n18277 & ~n18278;
  assign n18280 = ~P2_INSTADDRPOINTER_REG_8_ & ~n18279;
  assign n18281 = P2_INSTADDRPOINTER_REG_8_ & n18279;
  assign n18282 = ~n18280 & ~n18281;
  assign n18283 = n18268 & ~n18282;
  assign n18284 = ~n18268 & n18282;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = n17458 & ~n18285;
  assign n18287 = P2_INSTADDRPOINTER_REG_8_ & n17410;
  assign n18288 = P2_REIP_REG_8_ & n17461;
  assign n18289 = ~n18287 & ~n18288;
  assign n18290 = P2_INSTADDRPOINTER_REG_7_ & n18204;
  assign n18291 = ~P2_INSTADDRPOINTER_REG_8_ & n18290;
  assign n18292 = P2_INSTADDRPOINTER_REG_8_ & ~n18290;
  assign n18293 = ~n18291 & ~n18292;
  assign n18294 = n17464 & ~n18293;
  assign n18295 = P2_INSTADDRPOINTER_REG_7_ & n18209;
  assign n18296 = ~P2_INSTADDRPOINTER_REG_8_ & n18295;
  assign n18297 = P2_INSTADDRPOINTER_REG_8_ & ~n18295;
  assign n18298 = ~n18296 & ~n18297;
  assign n18299 = n17469 & ~n18298;
  assign n18300 = ~n18294 & ~n18299;
  assign n18301 = n18215 & ~n18222;
  assign n18302 = P2_EBX_REG_8_ & n14995;
  assign n18303 = P2_REIP_REG_8_ & n14997;
  assign n18304 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_8_;
  assign n18305 = P2_INSTADDRPOINTER_REG_8_ & ~n15016;
  assign n18306 = ~n18302 & ~n18303;
  assign n18307 = ~n18304 & n18306;
  assign n18308 = ~n18305 & n18307;
  assign n18309 = n18301 & n18308;
  assign n18310 = ~n18301 & ~n18308;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = n17476 & ~n18311;
  assign n18313 = n18231 & ~n18236;
  assign n18314 = ~n18231 & n18236;
  assign n18315 = ~n18230 & ~n18314;
  assign n18316 = ~n18313 & ~n18315;
  assign n18317 = P2_REIP_REG_8_ & n17226;
  assign n18318 = P2_INSTADDRPOINTER_REG_8_ & ~n17236;
  assign n18319 = P2_INSTQUEUERD_ADDR_REG_1_ & n14986;
  assign n18320 = ~P2_INSTQUEUERD_ADDR_REG_0_ & n15208;
  assign n18321 = n18319 & n18320;
  assign n18322 = P2_INSTQUEUE_REG_0__0_ & n18321;
  assign n18323 = P2_INSTQUEUERD_ADDR_REG_0_ & n15208;
  assign n18324 = n18319 & n18323;
  assign n18325 = P2_INSTQUEUE_REG_1__0_ & n18324;
  assign n18326 = ~P2_INSTQUEUERD_ADDR_REG_1_ & n14986;
  assign n18327 = n18320 & n18326;
  assign n18328 = P2_INSTQUEUE_REG_2__0_ & n18327;
  assign n18329 = n18323 & n18326;
  assign n18330 = P2_INSTQUEUE_REG_3__0_ & n18329;
  assign n18331 = ~n18322 & ~n18325;
  assign n18332 = ~n18328 & n18331;
  assign n18333 = ~n18330 & n18332;
  assign n18334 = ~P2_INSTQUEUERD_ADDR_REG_0_ & ~n15208;
  assign n18335 = n18319 & n18334;
  assign n18336 = P2_INSTQUEUE_REG_4__0_ & n18335;
  assign n18337 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n15208;
  assign n18338 = n18319 & n18337;
  assign n18339 = P2_INSTQUEUE_REG_5__0_ & n18338;
  assign n18340 = n18326 & n18334;
  assign n18341 = P2_INSTQUEUE_REG_6__0_ & n18340;
  assign n18342 = n18326 & n18337;
  assign n18343 = P2_INSTQUEUE_REG_7__0_ & n18342;
  assign n18344 = ~n18336 & ~n18339;
  assign n18345 = ~n18341 & n18344;
  assign n18346 = ~n18343 & n18345;
  assign n18347 = P2_INSTQUEUERD_ADDR_REG_1_ & ~n14986;
  assign n18348 = n18320 & n18347;
  assign n18349 = P2_INSTQUEUE_REG_8__0_ & n18348;
  assign n18350 = n18323 & n18347;
  assign n18351 = P2_INSTQUEUE_REG_9__0_ & n18350;
  assign n18352 = ~P2_INSTQUEUERD_ADDR_REG_1_ & ~n14986;
  assign n18353 = n18320 & n18352;
  assign n18354 = P2_INSTQUEUE_REG_10__0_ & n18353;
  assign n18355 = n18323 & n18352;
  assign n18356 = P2_INSTQUEUE_REG_11__0_ & n18355;
  assign n18357 = ~n18349 & ~n18351;
  assign n18358 = ~n18354 & n18357;
  assign n18359 = ~n18356 & n18358;
  assign n18360 = n18334 & n18347;
  assign n18361 = P2_INSTQUEUE_REG_12__0_ & n18360;
  assign n18362 = n18337 & n18347;
  assign n18363 = P2_INSTQUEUE_REG_13__0_ & n18362;
  assign n18364 = n18334 & n18352;
  assign n18365 = P2_INSTQUEUE_REG_14__0_ & n18364;
  assign n18366 = n18337 & n18352;
  assign n18367 = P2_INSTQUEUE_REG_15__0_ & n18366;
  assign n18368 = ~n18361 & ~n18363;
  assign n18369 = ~n18365 & n18368;
  assign n18370 = ~n18367 & n18369;
  assign n18371 = n18333 & n18346;
  assign n18372 = n18359 & n18371;
  assign n18373 = n18370 & n18372;
  assign n18374 = n17242 & ~n18373;
  assign n18375 = P2_EAX_REG_8_ & n17228;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = ~n18317 & ~n18318;
  assign n18378 = n18376 & n18377;
  assign n18379 = n18316 & ~n18378;
  assign n18380 = ~n18316 & n18378;
  assign n18381 = ~n18379 & ~n18380;
  assign n18382 = n17480 & ~n18381;
  assign n18383 = ~n18312 & ~n18382;
  assign n18384 = ~n18261 & ~n18286;
  assign n18385 = n18289 & n18384;
  assign n18386 = n18300 & n18385;
  assign n3914 = ~n18383 | ~n18386;
  assign n18388 = ~P2_INSTADDRPOINTER_REG_8_ & ~n18254;
  assign n18389 = P2_INSTADDRPOINTER_REG_7_ & ~n18388;
  assign n18390 = ~n18164 & n18389;
  assign n18391 = P2_INSTADDRPOINTER_REG_8_ & n18254;
  assign n18392 = ~n18390 & ~n18391;
  assign n18393 = ~n18126 & ~n18388;
  assign n18394 = ~n18250 & n18393;
  assign n18395 = n18392 & ~n18394;
  assign n18396 = ~P2_INSTADDRPOINTER_REG_9_ & n18395;
  assign n18397 = P2_INSTADDRPOINTER_REG_9_ & ~n18395;
  assign n18398 = ~n18396 & ~n18397;
  assign n18399 = n17413 & n18398;
  assign n18400 = P2_INSTADDRPOINTER_REG_8_ & ~n18279;
  assign n18401 = ~P2_INSTADDRPOINTER_REG_8_ & n18279;
  assign n18402 = ~n18268 & ~n18401;
  assign n18403 = ~n18400 & ~n18402;
  assign n18404 = P2_EBX_REG_9_ & n14365;
  assign n18405 = ~n18271 & ~n18404;
  assign n18406 = ~n18274 & ~n18405;
  assign n18407 = n18273 & n18405;
  assign n18408 = n18189 & n18407;
  assign n18409 = ~n18406 & ~n18408;
  assign n18410 = ~n17445 & n18409;
  assign n18411 = ~P2_INSTADDRPOINTER_REG_9_ & n18410;
  assign n18412 = P2_INSTADDRPOINTER_REG_9_ & ~n18410;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = n18403 & ~n18413;
  assign n18415 = ~n18403 & n18413;
  assign n18416 = ~n18414 & ~n18415;
  assign n18417 = n17458 & ~n18416;
  assign n18418 = P2_INSTADDRPOINTER_REG_9_ & n17410;
  assign n18419 = P2_REIP_REG_9_ & n17461;
  assign n18420 = ~n18418 & ~n18419;
  assign n18421 = P2_INSTADDRPOINTER_REG_8_ & n18290;
  assign n18422 = ~P2_INSTADDRPOINTER_REG_9_ & n18421;
  assign n18423 = P2_INSTADDRPOINTER_REG_9_ & ~n18421;
  assign n18424 = ~n18422 & ~n18423;
  assign n18425 = n17464 & ~n18424;
  assign n18426 = P2_INSTADDRPOINTER_REG_8_ & n18295;
  assign n18427 = ~P2_INSTADDRPOINTER_REG_9_ & n18426;
  assign n18428 = P2_INSTADDRPOINTER_REG_9_ & ~n18426;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = n17469 & ~n18429;
  assign n18431 = ~n18425 & ~n18430;
  assign n18432 = n18301 & ~n18308;
  assign n18433 = P2_EBX_REG_9_ & n14995;
  assign n18434 = P2_REIP_REG_9_ & n14997;
  assign n18435 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_9_;
  assign n18436 = P2_INSTADDRPOINTER_REG_9_ & ~n15016;
  assign n18437 = ~n18433 & ~n18434;
  assign n18438 = ~n18435 & n18437;
  assign n18439 = ~n18436 & n18438;
  assign n18440 = n18432 & n18439;
  assign n18441 = ~n18432 & ~n18439;
  assign n18442 = ~n18440 & ~n18441;
  assign n18443 = n17476 & ~n18442;
  assign n18444 = ~n18316 & ~n18378;
  assign n18445 = P2_REIP_REG_9_ & n17226;
  assign n18446 = P2_INSTADDRPOINTER_REG_9_ & ~n17236;
  assign n18447 = P2_INSTQUEUE_REG_0__1_ & n18321;
  assign n18448 = P2_INSTQUEUE_REG_1__1_ & n18324;
  assign n18449 = P2_INSTQUEUE_REG_2__1_ & n18327;
  assign n18450 = P2_INSTQUEUE_REG_3__1_ & n18329;
  assign n18451 = ~n18447 & ~n18448;
  assign n18452 = ~n18449 & n18451;
  assign n18453 = ~n18450 & n18452;
  assign n18454 = P2_INSTQUEUE_REG_4__1_ & n18335;
  assign n18455 = P2_INSTQUEUE_REG_5__1_ & n18338;
  assign n18456 = P2_INSTQUEUE_REG_6__1_ & n18340;
  assign n18457 = P2_INSTQUEUE_REG_7__1_ & n18342;
  assign n18458 = ~n18454 & ~n18455;
  assign n18459 = ~n18456 & n18458;
  assign n18460 = ~n18457 & n18459;
  assign n18461 = P2_INSTQUEUE_REG_8__1_ & n18348;
  assign n18462 = P2_INSTQUEUE_REG_9__1_ & n18350;
  assign n18463 = P2_INSTQUEUE_REG_10__1_ & n18353;
  assign n18464 = P2_INSTQUEUE_REG_11__1_ & n18355;
  assign n18465 = ~n18461 & ~n18462;
  assign n18466 = ~n18463 & n18465;
  assign n18467 = ~n18464 & n18466;
  assign n18468 = P2_INSTQUEUE_REG_12__1_ & n18360;
  assign n18469 = P2_INSTQUEUE_REG_13__1_ & n18362;
  assign n18470 = P2_INSTQUEUE_REG_14__1_ & n18364;
  assign n18471 = P2_INSTQUEUE_REG_15__1_ & n18366;
  assign n18472 = ~n18468 & ~n18469;
  assign n18473 = ~n18470 & n18472;
  assign n18474 = ~n18471 & n18473;
  assign n18475 = n18453 & n18460;
  assign n18476 = n18467 & n18475;
  assign n18477 = n18474 & n18476;
  assign n18478 = n17242 & ~n18477;
  assign n18479 = P2_EAX_REG_9_ & n17228;
  assign n18480 = ~n18478 & ~n18479;
  assign n18481 = ~n18445 & ~n18446;
  assign n18482 = n18480 & n18481;
  assign n18483 = ~n18444 & ~n18482;
  assign n18484 = n18444 & n18482;
  assign n18485 = ~n18483 & ~n18484;
  assign n18486 = n17480 & ~n18485;
  assign n18487 = ~n18443 & ~n18486;
  assign n18488 = ~n18399 & ~n18417;
  assign n18489 = n18420 & n18488;
  assign n18490 = n18431 & n18489;
  assign n3919 = ~n18487 | ~n18490;
  assign n18492 = ~P2_INSTADDRPOINTER_REG_10_ & ~n18397;
  assign n18493 = P2_INSTADDRPOINTER_REG_9_ & P2_INSTADDRPOINTER_REG_10_;
  assign n18494 = ~n18395 & n18493;
  assign n18495 = ~n18492 & ~n18494;
  assign n18496 = n17413 & n18495;
  assign n18497 = ~P2_INSTADDRPOINTER_REG_9_ & ~n18410;
  assign n18498 = n18400 & ~n18497;
  assign n18499 = P2_INSTADDRPOINTER_REG_9_ & n18410;
  assign n18500 = ~n18498 & ~n18499;
  assign n18501 = ~n18401 & ~n18497;
  assign n18502 = ~n18268 & n18501;
  assign n18503 = n18500 & ~n18502;
  assign n18504 = P2_EBX_REG_10_ & n14365;
  assign n18505 = ~n18271 & ~n18504;
  assign n18506 = n18408 & n18505;
  assign n18507 = ~n18408 & ~n18505;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = ~n17445 & n18508;
  assign n18510 = ~P2_INSTADDRPOINTER_REG_10_ & n18509;
  assign n18511 = P2_INSTADDRPOINTER_REG_10_ & ~n18509;
  assign n18512 = ~n18510 & ~n18511;
  assign n18513 = n18503 & ~n18512;
  assign n18514 = ~n18503 & n18512;
  assign n18515 = ~n18513 & ~n18514;
  assign n18516 = n17458 & ~n18515;
  assign n18517 = P2_INSTADDRPOINTER_REG_10_ & n17410;
  assign n18518 = P2_REIP_REG_10_ & n17461;
  assign n18519 = ~n18517 & ~n18518;
  assign n18520 = P2_INSTADDRPOINTER_REG_9_ & n18421;
  assign n18521 = ~P2_INSTADDRPOINTER_REG_10_ & n18520;
  assign n18522 = P2_INSTADDRPOINTER_REG_10_ & ~n18520;
  assign n18523 = ~n18521 & ~n18522;
  assign n18524 = n17464 & ~n18523;
  assign n18525 = P2_INSTADDRPOINTER_REG_9_ & n18426;
  assign n18526 = ~P2_INSTADDRPOINTER_REG_10_ & n18525;
  assign n18527 = P2_INSTADDRPOINTER_REG_10_ & ~n18525;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = n17469 & ~n18528;
  assign n18530 = ~n18524 & ~n18529;
  assign n18531 = n18432 & ~n18439;
  assign n18532 = P2_EBX_REG_10_ & n14995;
  assign n18533 = P2_REIP_REG_10_ & n14997;
  assign n18534 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_10_;
  assign n18535 = P2_INSTADDRPOINTER_REG_10_ & ~n15016;
  assign n18536 = ~n18532 & ~n18533;
  assign n18537 = ~n18534 & n18536;
  assign n18538 = ~n18535 & n18537;
  assign n18539 = n18531 & n18538;
  assign n18540 = ~n18531 & ~n18538;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = n17476 & ~n18541;
  assign n18543 = n18444 & ~n18482;
  assign n18544 = P2_REIP_REG_10_ & n17226;
  assign n18545 = P2_INSTADDRPOINTER_REG_10_ & ~n17236;
  assign n18546 = P2_INSTQUEUE_REG_0__2_ & n18321;
  assign n18547 = P2_INSTQUEUE_REG_1__2_ & n18324;
  assign n18548 = P2_INSTQUEUE_REG_2__2_ & n18327;
  assign n18549 = P2_INSTQUEUE_REG_3__2_ & n18329;
  assign n18550 = ~n18546 & ~n18547;
  assign n18551 = ~n18548 & n18550;
  assign n18552 = ~n18549 & n18551;
  assign n18553 = P2_INSTQUEUE_REG_4__2_ & n18335;
  assign n18554 = P2_INSTQUEUE_REG_5__2_ & n18338;
  assign n18555 = P2_INSTQUEUE_REG_6__2_ & n18340;
  assign n18556 = P2_INSTQUEUE_REG_7__2_ & n18342;
  assign n18557 = ~n18553 & ~n18554;
  assign n18558 = ~n18555 & n18557;
  assign n18559 = ~n18556 & n18558;
  assign n18560 = P2_INSTQUEUE_REG_8__2_ & n18348;
  assign n18561 = P2_INSTQUEUE_REG_9__2_ & n18350;
  assign n18562 = P2_INSTQUEUE_REG_10__2_ & n18353;
  assign n18563 = P2_INSTQUEUE_REG_11__2_ & n18355;
  assign n18564 = ~n18560 & ~n18561;
  assign n18565 = ~n18562 & n18564;
  assign n18566 = ~n18563 & n18565;
  assign n18567 = P2_INSTQUEUE_REG_12__2_ & n18360;
  assign n18568 = P2_INSTQUEUE_REG_13__2_ & n18362;
  assign n18569 = P2_INSTQUEUE_REG_14__2_ & n18364;
  assign n18570 = P2_INSTQUEUE_REG_15__2_ & n18366;
  assign n18571 = ~n18567 & ~n18568;
  assign n18572 = ~n18569 & n18571;
  assign n18573 = ~n18570 & n18572;
  assign n18574 = n18552 & n18559;
  assign n18575 = n18566 & n18574;
  assign n18576 = n18573 & n18575;
  assign n18577 = n17242 & ~n18576;
  assign n18578 = P2_EAX_REG_10_ & n17228;
  assign n18579 = ~n18577 & ~n18578;
  assign n18580 = ~n18544 & ~n18545;
  assign n18581 = n18579 & n18580;
  assign n18582 = ~n18543 & ~n18581;
  assign n18583 = n18543 & n18581;
  assign n18584 = ~n18582 & ~n18583;
  assign n18585 = n17480 & ~n18584;
  assign n18586 = ~n18542 & ~n18585;
  assign n18587 = ~n18496 & ~n18516;
  assign n18588 = n18519 & n18587;
  assign n18589 = n18530 & n18588;
  assign n3924 = ~n18586 | ~n18589;
  assign n18591 = ~P2_INSTADDRPOINTER_REG_11_ & ~n18494;
  assign n18592 = P2_INSTADDRPOINTER_REG_11_ & n18493;
  assign n18593 = ~n18395 & n18592;
  assign n18594 = ~n18591 & ~n18593;
  assign n18595 = n17413 & n18594;
  assign n18596 = P2_INSTADDRPOINTER_REG_10_ & n18509;
  assign n18597 = ~P2_INSTADDRPOINTER_REG_10_ & ~n18509;
  assign n18598 = ~n18503 & ~n18597;
  assign n18599 = ~n18596 & ~n18598;
  assign n18600 = P2_EBX_REG_11_ & n14365;
  assign n18601 = ~n18271 & ~n18600;
  assign n18602 = ~n18506 & ~n18601;
  assign n18603 = n18505 & n18601;
  assign n18604 = n18408 & n18603;
  assign n18605 = ~n18602 & ~n18604;
  assign n18606 = ~n17445 & n18605;
  assign n18607 = ~P2_INSTADDRPOINTER_REG_11_ & n18606;
  assign n18608 = P2_INSTADDRPOINTER_REG_11_ & ~n18606;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = n18599 & ~n18609;
  assign n18611 = ~n18599 & n18609;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = n17458 & ~n18612;
  assign n18614 = P2_INSTADDRPOINTER_REG_11_ & n17410;
  assign n18615 = P2_REIP_REG_11_ & n17461;
  assign n18616 = ~n18614 & ~n18615;
  assign n18617 = P2_INSTADDRPOINTER_REG_10_ & n18520;
  assign n18618 = ~P2_INSTADDRPOINTER_REG_11_ & n18617;
  assign n18619 = P2_INSTADDRPOINTER_REG_11_ & ~n18617;
  assign n18620 = ~n18618 & ~n18619;
  assign n18621 = n17464 & ~n18620;
  assign n18622 = P2_INSTADDRPOINTER_REG_10_ & n18525;
  assign n18623 = ~P2_INSTADDRPOINTER_REG_11_ & n18622;
  assign n18624 = P2_INSTADDRPOINTER_REG_11_ & ~n18622;
  assign n18625 = ~n18623 & ~n18624;
  assign n18626 = n17469 & ~n18625;
  assign n18627 = ~n18621 & ~n18626;
  assign n18628 = n18531 & ~n18538;
  assign n18629 = P2_EBX_REG_11_ & n14995;
  assign n18630 = P2_REIP_REG_11_ & n14997;
  assign n18631 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_11_;
  assign n18632 = P2_INSTADDRPOINTER_REG_11_ & ~n15016;
  assign n18633 = ~n18629 & ~n18630;
  assign n18634 = ~n18631 & n18633;
  assign n18635 = ~n18632 & n18634;
  assign n18636 = n18628 & n18635;
  assign n18637 = ~n18628 & ~n18635;
  assign n18638 = ~n18636 & ~n18637;
  assign n18639 = n17476 & ~n18638;
  assign n18640 = n18543 & ~n18581;
  assign n18641 = P2_REIP_REG_11_ & n17226;
  assign n18642 = P2_INSTADDRPOINTER_REG_11_ & ~n17236;
  assign n18643 = P2_INSTQUEUE_REG_0__3_ & n18321;
  assign n18644 = P2_INSTQUEUE_REG_1__3_ & n18324;
  assign n18645 = P2_INSTQUEUE_REG_2__3_ & n18327;
  assign n18646 = P2_INSTQUEUE_REG_3__3_ & n18329;
  assign n18647 = ~n18643 & ~n18644;
  assign n18648 = ~n18645 & n18647;
  assign n18649 = ~n18646 & n18648;
  assign n18650 = P2_INSTQUEUE_REG_4__3_ & n18335;
  assign n18651 = P2_INSTQUEUE_REG_5__3_ & n18338;
  assign n18652 = P2_INSTQUEUE_REG_6__3_ & n18340;
  assign n18653 = P2_INSTQUEUE_REG_7__3_ & n18342;
  assign n18654 = ~n18650 & ~n18651;
  assign n18655 = ~n18652 & n18654;
  assign n18656 = ~n18653 & n18655;
  assign n18657 = P2_INSTQUEUE_REG_8__3_ & n18348;
  assign n18658 = P2_INSTQUEUE_REG_9__3_ & n18350;
  assign n18659 = P2_INSTQUEUE_REG_10__3_ & n18353;
  assign n18660 = P2_INSTQUEUE_REG_11__3_ & n18355;
  assign n18661 = ~n18657 & ~n18658;
  assign n18662 = ~n18659 & n18661;
  assign n18663 = ~n18660 & n18662;
  assign n18664 = P2_INSTQUEUE_REG_12__3_ & n18360;
  assign n18665 = P2_INSTQUEUE_REG_13__3_ & n18362;
  assign n18666 = P2_INSTQUEUE_REG_14__3_ & n18364;
  assign n18667 = P2_INSTQUEUE_REG_15__3_ & n18366;
  assign n18668 = ~n18664 & ~n18665;
  assign n18669 = ~n18666 & n18668;
  assign n18670 = ~n18667 & n18669;
  assign n18671 = n18649 & n18656;
  assign n18672 = n18663 & n18671;
  assign n18673 = n18670 & n18672;
  assign n18674 = n17242 & ~n18673;
  assign n18675 = P2_EAX_REG_11_ & n17228;
  assign n18676 = ~n18674 & ~n18675;
  assign n18677 = ~n18641 & ~n18642;
  assign n18678 = n18676 & n18677;
  assign n18679 = ~n18640 & ~n18678;
  assign n18680 = n18640 & n18678;
  assign n18681 = ~n18679 & ~n18680;
  assign n18682 = n17480 & ~n18681;
  assign n18683 = ~n18639 & ~n18682;
  assign n18684 = ~n18595 & ~n18613;
  assign n18685 = n18616 & n18684;
  assign n18686 = n18627 & n18685;
  assign n3929 = ~n18683 | ~n18686;
  assign n18688 = ~P2_INSTADDRPOINTER_REG_12_ & n18593;
  assign n18689 = P2_INSTADDRPOINTER_REG_12_ & ~n18593;
  assign n18690 = ~n18688 & ~n18689;
  assign n18691 = n17413 & ~n18690;
  assign n18692 = ~P2_INSTADDRPOINTER_REG_11_ & ~n18606;
  assign n18693 = n18596 & ~n18692;
  assign n18694 = P2_INSTADDRPOINTER_REG_11_ & n18606;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = ~n18597 & ~n18692;
  assign n18697 = ~n18503 & n18696;
  assign n18698 = n18695 & ~n18697;
  assign n18699 = P2_EBX_REG_12_ & n14365;
  assign n18700 = ~n18271 & ~n18699;
  assign n18701 = n18604 & n18700;
  assign n18702 = ~n18604 & ~n18700;
  assign n18703 = ~n18701 & ~n18702;
  assign n18704 = ~n17445 & n18703;
  assign n18705 = ~P2_INSTADDRPOINTER_REG_12_ & n18704;
  assign n18706 = P2_INSTADDRPOINTER_REG_12_ & ~n18704;
  assign n18707 = ~n18705 & ~n18706;
  assign n18708 = n18698 & ~n18707;
  assign n18709 = ~n18698 & n18707;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = n17458 & ~n18710;
  assign n18712 = P2_INSTADDRPOINTER_REG_12_ & n17410;
  assign n18713 = P2_REIP_REG_12_ & n17461;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = P2_INSTADDRPOINTER_REG_11_ & n18617;
  assign n18716 = ~P2_INSTADDRPOINTER_REG_12_ & n18715;
  assign n18717 = P2_INSTADDRPOINTER_REG_12_ & ~n18715;
  assign n18718 = ~n18716 & ~n18717;
  assign n18719 = n17464 & ~n18718;
  assign n18720 = P2_INSTADDRPOINTER_REG_11_ & n18622;
  assign n18721 = ~P2_INSTADDRPOINTER_REG_12_ & n18720;
  assign n18722 = P2_INSTADDRPOINTER_REG_12_ & ~n18720;
  assign n18723 = ~n18721 & ~n18722;
  assign n18724 = n17469 & ~n18723;
  assign n18725 = ~n18719 & ~n18724;
  assign n18726 = n18628 & ~n18635;
  assign n18727 = P2_EBX_REG_12_ & n14995;
  assign n18728 = P2_REIP_REG_12_ & n14997;
  assign n18729 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_12_;
  assign n18730 = P2_INSTADDRPOINTER_REG_12_ & ~n15016;
  assign n18731 = ~n18727 & ~n18728;
  assign n18732 = ~n18729 & n18731;
  assign n18733 = ~n18730 & n18732;
  assign n18734 = n18726 & n18733;
  assign n18735 = ~n18726 & ~n18733;
  assign n18736 = ~n18734 & ~n18735;
  assign n18737 = n17476 & ~n18736;
  assign n18738 = n18640 & ~n18678;
  assign n18739 = P2_REIP_REG_12_ & n17226;
  assign n18740 = P2_INSTADDRPOINTER_REG_12_ & ~n17236;
  assign n18741 = P2_INSTQUEUE_REG_0__4_ & n18321;
  assign n18742 = P2_INSTQUEUE_REG_1__4_ & n18324;
  assign n18743 = P2_INSTQUEUE_REG_2__4_ & n18327;
  assign n18744 = P2_INSTQUEUE_REG_3__4_ & n18329;
  assign n18745 = ~n18741 & ~n18742;
  assign n18746 = ~n18743 & n18745;
  assign n18747 = ~n18744 & n18746;
  assign n18748 = P2_INSTQUEUE_REG_4__4_ & n18335;
  assign n18749 = P2_INSTQUEUE_REG_5__4_ & n18338;
  assign n18750 = P2_INSTQUEUE_REG_6__4_ & n18340;
  assign n18751 = P2_INSTQUEUE_REG_7__4_ & n18342;
  assign n18752 = ~n18748 & ~n18749;
  assign n18753 = ~n18750 & n18752;
  assign n18754 = ~n18751 & n18753;
  assign n18755 = P2_INSTQUEUE_REG_8__4_ & n18348;
  assign n18756 = P2_INSTQUEUE_REG_9__4_ & n18350;
  assign n18757 = P2_INSTQUEUE_REG_10__4_ & n18353;
  assign n18758 = P2_INSTQUEUE_REG_11__4_ & n18355;
  assign n18759 = ~n18755 & ~n18756;
  assign n18760 = ~n18757 & n18759;
  assign n18761 = ~n18758 & n18760;
  assign n18762 = P2_INSTQUEUE_REG_12__4_ & n18360;
  assign n18763 = P2_INSTQUEUE_REG_13__4_ & n18362;
  assign n18764 = P2_INSTQUEUE_REG_14__4_ & n18364;
  assign n18765 = P2_INSTQUEUE_REG_15__4_ & n18366;
  assign n18766 = ~n18762 & ~n18763;
  assign n18767 = ~n18764 & n18766;
  assign n18768 = ~n18765 & n18767;
  assign n18769 = n18747 & n18754;
  assign n18770 = n18761 & n18769;
  assign n18771 = n18768 & n18770;
  assign n18772 = n17242 & ~n18771;
  assign n18773 = P2_EAX_REG_12_ & n17228;
  assign n18774 = ~n18772 & ~n18773;
  assign n18775 = ~n18739 & ~n18740;
  assign n18776 = n18774 & n18775;
  assign n18777 = ~n18738 & ~n18776;
  assign n18778 = n18738 & n18776;
  assign n18779 = ~n18777 & ~n18778;
  assign n18780 = n17480 & ~n18779;
  assign n18781 = ~n18737 & ~n18780;
  assign n18782 = ~n18691 & ~n18711;
  assign n18783 = n18714 & n18782;
  assign n18784 = n18725 & n18783;
  assign n3934 = ~n18781 | ~n18784;
  assign n18786 = P2_INSTADDRPOINTER_REG_11_ & P2_INSTADDRPOINTER_REG_12_;
  assign n18787 = P2_INSTADDRPOINTER_REG_10_ & n18786;
  assign n18788 = P2_INSTADDRPOINTER_REG_9_ & n18787;
  assign n18789 = ~n18395 & n18788;
  assign n18790 = ~P2_INSTADDRPOINTER_REG_13_ & ~n18789;
  assign n18791 = P2_INSTADDRPOINTER_REG_13_ & n18788;
  assign n18792 = ~n18395 & n18791;
  assign n18793 = ~n18790 & ~n18792;
  assign n18794 = n17413 & n18793;
  assign n18795 = P2_INSTADDRPOINTER_REG_12_ & n18704;
  assign n18796 = ~P2_INSTADDRPOINTER_REG_12_ & ~n18704;
  assign n18797 = ~n18698 & ~n18796;
  assign n18798 = ~n18795 & ~n18797;
  assign n18799 = P2_EBX_REG_13_ & n14365;
  assign n18800 = ~n18271 & ~n18799;
  assign n18801 = ~n18701 & ~n18800;
  assign n18802 = n18700 & n18800;
  assign n18803 = n18604 & n18802;
  assign n18804 = ~n18801 & ~n18803;
  assign n18805 = ~n17445 & n18804;
  assign n18806 = ~P2_INSTADDRPOINTER_REG_13_ & n18805;
  assign n18807 = P2_INSTADDRPOINTER_REG_13_ & ~n18805;
  assign n18808 = ~n18806 & ~n18807;
  assign n18809 = n18798 & ~n18808;
  assign n18810 = ~n18798 & n18808;
  assign n18811 = ~n18809 & ~n18810;
  assign n18812 = n17458 & ~n18811;
  assign n18813 = P2_INSTADDRPOINTER_REG_13_ & n17410;
  assign n18814 = P2_REIP_REG_13_ & n17461;
  assign n18815 = ~n18813 & ~n18814;
  assign n18816 = P2_INSTADDRPOINTER_REG_12_ & n18715;
  assign n18817 = ~P2_INSTADDRPOINTER_REG_13_ & n18816;
  assign n18818 = P2_INSTADDRPOINTER_REG_13_ & ~n18816;
  assign n18819 = ~n18817 & ~n18818;
  assign n18820 = n17464 & ~n18819;
  assign n18821 = P2_INSTADDRPOINTER_REG_12_ & n18720;
  assign n18822 = ~P2_INSTADDRPOINTER_REG_13_ & n18821;
  assign n18823 = P2_INSTADDRPOINTER_REG_13_ & ~n18821;
  assign n18824 = ~n18822 & ~n18823;
  assign n18825 = n17469 & ~n18824;
  assign n18826 = ~n18820 & ~n18825;
  assign n18827 = n18726 & ~n18733;
  assign n18828 = P2_EBX_REG_13_ & n14995;
  assign n18829 = P2_REIP_REG_13_ & n14997;
  assign n18830 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_13_;
  assign n18831 = P2_INSTADDRPOINTER_REG_13_ & ~n15016;
  assign n18832 = ~n18828 & ~n18829;
  assign n18833 = ~n18830 & n18832;
  assign n18834 = ~n18831 & n18833;
  assign n18835 = n18827 & n18834;
  assign n18836 = ~n18827 & ~n18834;
  assign n18837 = ~n18835 & ~n18836;
  assign n18838 = n17476 & ~n18837;
  assign n18839 = n18738 & ~n18776;
  assign n18840 = P2_REIP_REG_13_ & n17226;
  assign n18841 = P2_INSTADDRPOINTER_REG_13_ & ~n17236;
  assign n18842 = P2_INSTQUEUE_REG_0__5_ & n18321;
  assign n18843 = P2_INSTQUEUE_REG_1__5_ & n18324;
  assign n18844 = P2_INSTQUEUE_REG_2__5_ & n18327;
  assign n18845 = P2_INSTQUEUE_REG_3__5_ & n18329;
  assign n18846 = ~n18842 & ~n18843;
  assign n18847 = ~n18844 & n18846;
  assign n18848 = ~n18845 & n18847;
  assign n18849 = P2_INSTQUEUE_REG_4__5_ & n18335;
  assign n18850 = P2_INSTQUEUE_REG_5__5_ & n18338;
  assign n18851 = P2_INSTQUEUE_REG_6__5_ & n18340;
  assign n18852 = P2_INSTQUEUE_REG_7__5_ & n18342;
  assign n18853 = ~n18849 & ~n18850;
  assign n18854 = ~n18851 & n18853;
  assign n18855 = ~n18852 & n18854;
  assign n18856 = P2_INSTQUEUE_REG_8__5_ & n18348;
  assign n18857 = P2_INSTQUEUE_REG_9__5_ & n18350;
  assign n18858 = P2_INSTQUEUE_REG_10__5_ & n18353;
  assign n18859 = P2_INSTQUEUE_REG_11__5_ & n18355;
  assign n18860 = ~n18856 & ~n18857;
  assign n18861 = ~n18858 & n18860;
  assign n18862 = ~n18859 & n18861;
  assign n18863 = P2_INSTQUEUE_REG_12__5_ & n18360;
  assign n18864 = P2_INSTQUEUE_REG_13__5_ & n18362;
  assign n18865 = P2_INSTQUEUE_REG_14__5_ & n18364;
  assign n18866 = P2_INSTQUEUE_REG_15__5_ & n18366;
  assign n18867 = ~n18863 & ~n18864;
  assign n18868 = ~n18865 & n18867;
  assign n18869 = ~n18866 & n18868;
  assign n18870 = n18848 & n18855;
  assign n18871 = n18862 & n18870;
  assign n18872 = n18869 & n18871;
  assign n18873 = n17242 & ~n18872;
  assign n18874 = P2_EAX_REG_13_ & n17228;
  assign n18875 = ~n18873 & ~n18874;
  assign n18876 = ~n18840 & ~n18841;
  assign n18877 = n18875 & n18876;
  assign n18878 = ~n18839 & ~n18877;
  assign n18879 = n18839 & n18877;
  assign n18880 = ~n18878 & ~n18879;
  assign n18881 = n17480 & ~n18880;
  assign n18882 = ~n18838 & ~n18881;
  assign n18883 = ~n18794 & ~n18812;
  assign n18884 = n18815 & n18883;
  assign n18885 = n18826 & n18884;
  assign n3939 = ~n18882 | ~n18885;
  assign n18887 = ~P2_INSTADDRPOINTER_REG_14_ & ~n18792;
  assign n18888 = P2_INSTADDRPOINTER_REG_14_ & n18791;
  assign n18889 = ~n18395 & n18888;
  assign n18890 = ~n18887 & ~n18889;
  assign n18891 = n17413 & n18890;
  assign n18892 = ~P2_INSTADDRPOINTER_REG_13_ & ~n18805;
  assign n18893 = n18795 & ~n18892;
  assign n18894 = P2_INSTADDRPOINTER_REG_13_ & n18805;
  assign n18895 = ~n18893 & ~n18894;
  assign n18896 = ~n18796 & ~n18892;
  assign n18897 = ~n18698 & n18896;
  assign n18898 = n18895 & ~n18897;
  assign n18899 = P2_EBX_REG_14_ & n14365;
  assign n18900 = ~n18271 & ~n18899;
  assign n18901 = n18803 & n18900;
  assign n18902 = ~n18803 & ~n18900;
  assign n18903 = ~n18901 & ~n18902;
  assign n18904 = ~n17445 & n18903;
  assign n18905 = ~P2_INSTADDRPOINTER_REG_14_ & n18904;
  assign n18906 = P2_INSTADDRPOINTER_REG_14_ & ~n18904;
  assign n18907 = ~n18905 & ~n18906;
  assign n18908 = n18898 & ~n18907;
  assign n18909 = ~n18898 & n18907;
  assign n18910 = ~n18908 & ~n18909;
  assign n18911 = n17458 & ~n18910;
  assign n18912 = P2_INSTADDRPOINTER_REG_14_ & n17410;
  assign n18913 = P2_REIP_REG_14_ & n17461;
  assign n18914 = ~n18912 & ~n18913;
  assign n18915 = P2_INSTADDRPOINTER_REG_13_ & n18816;
  assign n18916 = ~P2_INSTADDRPOINTER_REG_14_ & n18915;
  assign n18917 = P2_INSTADDRPOINTER_REG_14_ & ~n18915;
  assign n18918 = ~n18916 & ~n18917;
  assign n18919 = n17464 & ~n18918;
  assign n18920 = P2_INSTADDRPOINTER_REG_13_ & n18821;
  assign n18921 = ~P2_INSTADDRPOINTER_REG_14_ & n18920;
  assign n18922 = P2_INSTADDRPOINTER_REG_14_ & ~n18920;
  assign n18923 = ~n18921 & ~n18922;
  assign n18924 = n17469 & ~n18923;
  assign n18925 = ~n18919 & ~n18924;
  assign n18926 = n18827 & ~n18834;
  assign n18927 = P2_EBX_REG_14_ & n14995;
  assign n18928 = P2_REIP_REG_14_ & n14997;
  assign n18929 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_14_;
  assign n18930 = P2_INSTADDRPOINTER_REG_14_ & ~n15016;
  assign n18931 = ~n18927 & ~n18928;
  assign n18932 = ~n18929 & n18931;
  assign n18933 = ~n18930 & n18932;
  assign n18934 = n18926 & n18933;
  assign n18935 = ~n18926 & ~n18933;
  assign n18936 = ~n18934 & ~n18935;
  assign n18937 = n17476 & ~n18936;
  assign n18938 = n18839 & ~n18877;
  assign n18939 = P2_REIP_REG_14_ & n17226;
  assign n18940 = P2_INSTADDRPOINTER_REG_14_ & ~n17236;
  assign n18941 = P2_INSTQUEUE_REG_0__6_ & n18321;
  assign n18942 = P2_INSTQUEUE_REG_1__6_ & n18324;
  assign n18943 = P2_INSTQUEUE_REG_2__6_ & n18327;
  assign n18944 = P2_INSTQUEUE_REG_3__6_ & n18329;
  assign n18945 = ~n18941 & ~n18942;
  assign n18946 = ~n18943 & n18945;
  assign n18947 = ~n18944 & n18946;
  assign n18948 = P2_INSTQUEUE_REG_4__6_ & n18335;
  assign n18949 = P2_INSTQUEUE_REG_5__6_ & n18338;
  assign n18950 = P2_INSTQUEUE_REG_6__6_ & n18340;
  assign n18951 = P2_INSTQUEUE_REG_7__6_ & n18342;
  assign n18952 = ~n18948 & ~n18949;
  assign n18953 = ~n18950 & n18952;
  assign n18954 = ~n18951 & n18953;
  assign n18955 = P2_INSTQUEUE_REG_8__6_ & n18348;
  assign n18956 = P2_INSTQUEUE_REG_9__6_ & n18350;
  assign n18957 = P2_INSTQUEUE_REG_10__6_ & n18353;
  assign n18958 = P2_INSTQUEUE_REG_11__6_ & n18355;
  assign n18959 = ~n18955 & ~n18956;
  assign n18960 = ~n18957 & n18959;
  assign n18961 = ~n18958 & n18960;
  assign n18962 = P2_INSTQUEUE_REG_12__6_ & n18360;
  assign n18963 = P2_INSTQUEUE_REG_13__6_ & n18362;
  assign n18964 = P2_INSTQUEUE_REG_14__6_ & n18364;
  assign n18965 = P2_INSTQUEUE_REG_15__6_ & n18366;
  assign n18966 = ~n18962 & ~n18963;
  assign n18967 = ~n18964 & n18966;
  assign n18968 = ~n18965 & n18967;
  assign n18969 = n18947 & n18954;
  assign n18970 = n18961 & n18969;
  assign n18971 = n18968 & n18970;
  assign n18972 = n17242 & ~n18971;
  assign n18973 = P2_EAX_REG_14_ & n17228;
  assign n18974 = ~n18972 & ~n18973;
  assign n18975 = ~n18939 & ~n18940;
  assign n18976 = n18974 & n18975;
  assign n18977 = ~n18938 & ~n18976;
  assign n18978 = n18938 & n18976;
  assign n18979 = ~n18977 & ~n18978;
  assign n18980 = n17480 & ~n18979;
  assign n18981 = ~n18937 & ~n18980;
  assign n18982 = ~n18891 & ~n18911;
  assign n18983 = n18914 & n18982;
  assign n18984 = n18925 & n18983;
  assign n3944 = ~n18981 | ~n18984;
  assign n18986 = ~P2_INSTADDRPOINTER_REG_15_ & n18889;
  assign n18987 = P2_INSTADDRPOINTER_REG_15_ & ~n18889;
  assign n18988 = ~n18986 & ~n18987;
  assign n18989 = n17413 & ~n18988;
  assign n18990 = P2_INSTADDRPOINTER_REG_14_ & n18904;
  assign n18991 = ~P2_INSTADDRPOINTER_REG_14_ & ~n18904;
  assign n18992 = ~n18898 & ~n18991;
  assign n18993 = ~n18990 & ~n18992;
  assign n18994 = P2_EBX_REG_15_ & n14365;
  assign n18995 = ~n18271 & ~n18994;
  assign n18996 = ~n18901 & ~n18995;
  assign n18997 = n18900 & n18995;
  assign n18998 = n18803 & n18997;
  assign n18999 = ~n18996 & ~n18998;
  assign n19000 = ~n17445 & n18999;
  assign n19001 = ~P2_INSTADDRPOINTER_REG_15_ & n19000;
  assign n19002 = P2_INSTADDRPOINTER_REG_15_ & ~n19000;
  assign n19003 = ~n19001 & ~n19002;
  assign n19004 = n18993 & ~n19003;
  assign n19005 = ~n18993 & n19003;
  assign n19006 = ~n19004 & ~n19005;
  assign n19007 = n17458 & ~n19006;
  assign n19008 = P2_INSTADDRPOINTER_REG_15_ & n17410;
  assign n19009 = P2_REIP_REG_15_ & n17461;
  assign n19010 = ~n19008 & ~n19009;
  assign n19011 = P2_INSTADDRPOINTER_REG_14_ & n18915;
  assign n19012 = ~P2_INSTADDRPOINTER_REG_15_ & n19011;
  assign n19013 = P2_INSTADDRPOINTER_REG_15_ & ~n19011;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = n17464 & ~n19014;
  assign n19016 = P2_INSTADDRPOINTER_REG_14_ & n18920;
  assign n19017 = ~P2_INSTADDRPOINTER_REG_15_ & n19016;
  assign n19018 = P2_INSTADDRPOINTER_REG_15_ & ~n19016;
  assign n19019 = ~n19017 & ~n19018;
  assign n19020 = n17469 & ~n19019;
  assign n19021 = ~n19015 & ~n19020;
  assign n19022 = n18926 & ~n18933;
  assign n19023 = P2_EBX_REG_15_ & n14995;
  assign n19024 = P2_REIP_REG_15_ & n14997;
  assign n19025 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_15_;
  assign n19026 = P2_INSTADDRPOINTER_REG_15_ & ~n15016;
  assign n19027 = ~n19023 & ~n19024;
  assign n19028 = ~n19025 & n19027;
  assign n19029 = ~n19026 & n19028;
  assign n19030 = n19022 & n19029;
  assign n19031 = ~n19022 & ~n19029;
  assign n19032 = ~n19030 & ~n19031;
  assign n19033 = n17476 & ~n19032;
  assign n19034 = n18938 & ~n18976;
  assign n19035 = P2_REIP_REG_15_ & n17226;
  assign n19036 = P2_INSTADDRPOINTER_REG_15_ & ~n17236;
  assign n19037 = P2_INSTQUEUE_REG_0__7_ & n18321;
  assign n19038 = P2_INSTQUEUE_REG_1__7_ & n18324;
  assign n19039 = P2_INSTQUEUE_REG_2__7_ & n18327;
  assign n19040 = P2_INSTQUEUE_REG_3__7_ & n18329;
  assign n19041 = ~n19037 & ~n19038;
  assign n19042 = ~n19039 & n19041;
  assign n19043 = ~n19040 & n19042;
  assign n19044 = P2_INSTQUEUE_REG_4__7_ & n18335;
  assign n19045 = P2_INSTQUEUE_REG_5__7_ & n18338;
  assign n19046 = P2_INSTQUEUE_REG_6__7_ & n18340;
  assign n19047 = P2_INSTQUEUE_REG_7__7_ & n18342;
  assign n19048 = ~n19044 & ~n19045;
  assign n19049 = ~n19046 & n19048;
  assign n19050 = ~n19047 & n19049;
  assign n19051 = P2_INSTQUEUE_REG_8__7_ & n18348;
  assign n19052 = P2_INSTQUEUE_REG_9__7_ & n18350;
  assign n19053 = P2_INSTQUEUE_REG_10__7_ & n18353;
  assign n19054 = P2_INSTQUEUE_REG_11__7_ & n18355;
  assign n19055 = ~n19051 & ~n19052;
  assign n19056 = ~n19053 & n19055;
  assign n19057 = ~n19054 & n19056;
  assign n19058 = P2_INSTQUEUE_REG_12__7_ & n18360;
  assign n19059 = P2_INSTQUEUE_REG_13__7_ & n18362;
  assign n19060 = P2_INSTQUEUE_REG_14__7_ & n18364;
  assign n19061 = P2_INSTQUEUE_REG_15__7_ & n18366;
  assign n19062 = ~n19058 & ~n19059;
  assign n19063 = ~n19060 & n19062;
  assign n19064 = ~n19061 & n19063;
  assign n19065 = n19043 & n19050;
  assign n19066 = n19057 & n19065;
  assign n19067 = n19064 & n19066;
  assign n19068 = n17242 & ~n19067;
  assign n19069 = P2_EAX_REG_15_ & n17228;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = ~n19035 & ~n19036;
  assign n19072 = n19070 & n19071;
  assign n19073 = ~n19034 & ~n19072;
  assign n19074 = n19034 & n19072;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = n17480 & ~n19075;
  assign n19077 = ~n19033 & ~n19076;
  assign n19078 = ~n18989 & ~n19007;
  assign n19079 = n19010 & n19078;
  assign n19080 = n19021 & n19079;
  assign n3949 = ~n19077 | ~n19080;
  assign n19082 = P2_INSTADDRPOINTER_REG_14_ & P2_INSTADDRPOINTER_REG_15_;
  assign n19083 = P2_INSTADDRPOINTER_REG_13_ & n19082;
  assign n19084 = n18788 & n19083;
  assign n19085 = ~n18395 & n19084;
  assign n19086 = ~P2_INSTADDRPOINTER_REG_16_ & ~n19085;
  assign n19087 = P2_INSTADDRPOINTER_REG_16_ & n19084;
  assign n19088 = ~n18395 & n19087;
  assign n19089 = ~n19086 & ~n19088;
  assign n19090 = n17413 & n19089;
  assign n19091 = ~P2_INSTADDRPOINTER_REG_15_ & ~n19000;
  assign n19092 = n18990 & ~n19091;
  assign n19093 = P2_INSTADDRPOINTER_REG_15_ & n19000;
  assign n19094 = ~n19092 & ~n19093;
  assign n19095 = ~n18991 & ~n19091;
  assign n19096 = ~n18898 & n19095;
  assign n19097 = n19094 & ~n19096;
  assign n19098 = P2_EBX_REG_16_ & n14365;
  assign n19099 = ~n18271 & ~n19098;
  assign n19100 = n18998 & n19099;
  assign n19101 = ~n18998 & ~n19099;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = ~n17445 & n19102;
  assign n19104 = ~P2_INSTADDRPOINTER_REG_16_ & n19103;
  assign n19105 = P2_INSTADDRPOINTER_REG_16_ & ~n19103;
  assign n19106 = ~n19104 & ~n19105;
  assign n19107 = n19097 & ~n19106;
  assign n19108 = ~n19097 & n19106;
  assign n19109 = ~n19107 & ~n19108;
  assign n19110 = n17458 & ~n19109;
  assign n19111 = P2_INSTADDRPOINTER_REG_16_ & n17410;
  assign n19112 = P2_REIP_REG_16_ & n17461;
  assign n19113 = ~n19111 & ~n19112;
  assign n19114 = P2_INSTADDRPOINTER_REG_15_ & n19011;
  assign n19115 = ~P2_INSTADDRPOINTER_REG_16_ & n19114;
  assign n19116 = P2_INSTADDRPOINTER_REG_16_ & ~n19114;
  assign n19117 = ~n19115 & ~n19116;
  assign n19118 = n17464 & ~n19117;
  assign n19119 = P2_INSTADDRPOINTER_REG_15_ & n19016;
  assign n19120 = ~P2_INSTADDRPOINTER_REG_16_ & n19119;
  assign n19121 = P2_INSTADDRPOINTER_REG_16_ & ~n19119;
  assign n19122 = ~n19120 & ~n19121;
  assign n19123 = n17469 & ~n19122;
  assign n19124 = ~n19118 & ~n19123;
  assign n19125 = n19022 & ~n19029;
  assign n19126 = P2_EBX_REG_16_ & n14995;
  assign n19127 = P2_REIP_REG_16_ & n14997;
  assign n19128 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_16_;
  assign n19129 = P2_INSTADDRPOINTER_REG_16_ & ~n15016;
  assign n19130 = ~n19126 & ~n19127;
  assign n19131 = ~n19128 & n19130;
  assign n19132 = ~n19129 & n19131;
  assign n19133 = n19125 & n19132;
  assign n19134 = ~n19125 & ~n19132;
  assign n19135 = ~n19133 & ~n19134;
  assign n19136 = n17476 & ~n19135;
  assign n19137 = n19034 & ~n19072;
  assign n19138 = P2_REIP_REG_16_ & n17226;
  assign n19139 = P2_EAX_REG_16_ & n17228;
  assign n19140 = ~n19138 & ~n19139;
  assign n19141 = P2_INSTADDRPOINTER_REG_16_ & ~n17236;
  assign n19142 = n19140 & ~n19141;
  assign n19143 = ~n19137 & ~n19142;
  assign n19144 = n19137 & n19142;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = n17480 & ~n19145;
  assign n19147 = ~n19136 & ~n19146;
  assign n19148 = ~n19090 & ~n19110;
  assign n19149 = n19113 & n19148;
  assign n19150 = n19124 & n19149;
  assign n3954 = ~n19147 | ~n19150;
  assign n19152 = ~P2_INSTADDRPOINTER_REG_17_ & n19088;
  assign n19153 = P2_INSTADDRPOINTER_REG_17_ & ~n19088;
  assign n19154 = ~n19152 & ~n19153;
  assign n19155 = n17413 & ~n19154;
  assign n19156 = P2_INSTADDRPOINTER_REG_16_ & n19103;
  assign n19157 = ~P2_INSTADDRPOINTER_REG_16_ & ~n19103;
  assign n19158 = ~n19097 & ~n19157;
  assign n19159 = ~n19156 & ~n19158;
  assign n19160 = P2_EBX_REG_17_ & n14365;
  assign n19161 = ~n18271 & ~n19160;
  assign n19162 = ~n19100 & ~n19161;
  assign n19163 = n19099 & n19161;
  assign n19164 = n18998 & n19163;
  assign n19165 = ~n19162 & ~n19164;
  assign n19166 = ~n17445 & n19165;
  assign n19167 = ~P2_INSTADDRPOINTER_REG_17_ & n19166;
  assign n19168 = P2_INSTADDRPOINTER_REG_17_ & ~n19166;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = n19159 & ~n19169;
  assign n19171 = ~n19159 & n19169;
  assign n19172 = ~n19170 & ~n19171;
  assign n19173 = n17458 & ~n19172;
  assign n19174 = P2_INSTADDRPOINTER_REG_17_ & n17410;
  assign n19175 = P2_REIP_REG_17_ & n17461;
  assign n19176 = ~n19174 & ~n19175;
  assign n19177 = P2_INSTADDRPOINTER_REG_16_ & n19114;
  assign n19178 = ~P2_INSTADDRPOINTER_REG_17_ & n19177;
  assign n19179 = P2_INSTADDRPOINTER_REG_17_ & ~n19177;
  assign n19180 = ~n19178 & ~n19179;
  assign n19181 = n17464 & ~n19180;
  assign n19182 = P2_INSTADDRPOINTER_REG_16_ & n19119;
  assign n19183 = ~P2_INSTADDRPOINTER_REG_17_ & n19182;
  assign n19184 = P2_INSTADDRPOINTER_REG_17_ & ~n19182;
  assign n19185 = ~n19183 & ~n19184;
  assign n19186 = n17469 & ~n19185;
  assign n19187 = ~n19181 & ~n19186;
  assign n19188 = n19125 & ~n19132;
  assign n19189 = P2_EBX_REG_17_ & n14995;
  assign n19190 = P2_REIP_REG_17_ & n14997;
  assign n19191 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_17_;
  assign n19192 = P2_INSTADDRPOINTER_REG_17_ & ~n15016;
  assign n19193 = ~n19189 & ~n19190;
  assign n19194 = ~n19191 & n19193;
  assign n19195 = ~n19192 & n19194;
  assign n19196 = n19188 & n19195;
  assign n19197 = ~n19188 & ~n19195;
  assign n19198 = ~n19196 & ~n19197;
  assign n19199 = n17476 & ~n19198;
  assign n19200 = n19137 & ~n19142;
  assign n19201 = P2_REIP_REG_17_ & n17226;
  assign n19202 = P2_EAX_REG_17_ & n17228;
  assign n19203 = ~n19201 & ~n19202;
  assign n19204 = P2_INSTADDRPOINTER_REG_17_ & ~n17236;
  assign n19205 = n19203 & ~n19204;
  assign n19206 = ~n19200 & ~n19205;
  assign n19207 = n19200 & n19205;
  assign n19208 = ~n19206 & ~n19207;
  assign n19209 = n17480 & ~n19208;
  assign n19210 = ~n19199 & ~n19209;
  assign n19211 = ~n19155 & ~n19173;
  assign n19212 = n19176 & n19211;
  assign n19213 = n19187 & n19212;
  assign n3959 = ~n19210 | ~n19213;
  assign n19215 = P2_INSTADDRPOINTER_REG_16_ & P2_INSTADDRPOINTER_REG_17_;
  assign n19216 = n19084 & n19215;
  assign n19217 = ~n18395 & n19216;
  assign n19218 = ~P2_INSTADDRPOINTER_REG_18_ & n19217;
  assign n19219 = P2_INSTADDRPOINTER_REG_18_ & ~n19217;
  assign n19220 = ~n19218 & ~n19219;
  assign n19221 = n17413 & ~n19220;
  assign n19222 = ~P2_INSTADDRPOINTER_REG_17_ & ~n19166;
  assign n19223 = n19156 & ~n19222;
  assign n19224 = P2_INSTADDRPOINTER_REG_17_ & n19166;
  assign n19225 = ~n19223 & ~n19224;
  assign n19226 = ~n19157 & ~n19222;
  assign n19227 = ~n19097 & n19226;
  assign n19228 = n19225 & ~n19227;
  assign n19229 = P2_EBX_REG_18_ & n14365;
  assign n19230 = ~n18271 & ~n19229;
  assign n19231 = n19164 & n19230;
  assign n19232 = ~n19164 & ~n19230;
  assign n19233 = ~n19231 & ~n19232;
  assign n19234 = ~n17445 & n19233;
  assign n19235 = ~P2_INSTADDRPOINTER_REG_18_ & n19234;
  assign n19236 = P2_INSTADDRPOINTER_REG_18_ & ~n19234;
  assign n19237 = ~n19235 & ~n19236;
  assign n19238 = n19228 & ~n19237;
  assign n19239 = ~n19228 & n19237;
  assign n19240 = ~n19238 & ~n19239;
  assign n19241 = n17458 & ~n19240;
  assign n19242 = P2_INSTADDRPOINTER_REG_18_ & n17410;
  assign n19243 = P2_REIP_REG_18_ & n17461;
  assign n19244 = ~n19242 & ~n19243;
  assign n19245 = P2_INSTADDRPOINTER_REG_17_ & n19177;
  assign n19246 = ~P2_INSTADDRPOINTER_REG_18_ & n19245;
  assign n19247 = P2_INSTADDRPOINTER_REG_18_ & ~n19245;
  assign n19248 = ~n19246 & ~n19247;
  assign n19249 = n17464 & ~n19248;
  assign n19250 = P2_INSTADDRPOINTER_REG_17_ & n19182;
  assign n19251 = ~P2_INSTADDRPOINTER_REG_18_ & n19250;
  assign n19252 = P2_INSTADDRPOINTER_REG_18_ & ~n19250;
  assign n19253 = ~n19251 & ~n19252;
  assign n19254 = n17469 & ~n19253;
  assign n19255 = ~n19249 & ~n19254;
  assign n19256 = n19188 & ~n19195;
  assign n19257 = P2_EBX_REG_18_ & n14995;
  assign n19258 = P2_REIP_REG_18_ & n14997;
  assign n19259 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_18_;
  assign n19260 = P2_INSTADDRPOINTER_REG_18_ & ~n15016;
  assign n19261 = ~n19257 & ~n19258;
  assign n19262 = ~n19259 & n19261;
  assign n19263 = ~n19260 & n19262;
  assign n19264 = n19256 & n19263;
  assign n19265 = ~n19256 & ~n19263;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = n17476 & ~n19266;
  assign n19268 = n19200 & ~n19205;
  assign n19269 = P2_REIP_REG_18_ & n17226;
  assign n19270 = P2_EAX_REG_18_ & n17228;
  assign n19271 = ~n19269 & ~n19270;
  assign n19272 = P2_INSTADDRPOINTER_REG_18_ & ~n17236;
  assign n19273 = n19271 & ~n19272;
  assign n19274 = ~n19268 & ~n19273;
  assign n19275 = n19268 & n19273;
  assign n19276 = ~n19274 & ~n19275;
  assign n19277 = n17480 & ~n19276;
  assign n19278 = ~n19267 & ~n19277;
  assign n19279 = ~n19221 & ~n19241;
  assign n19280 = n19244 & n19279;
  assign n19281 = n19255 & n19280;
  assign n3964 = ~n19278 | ~n19281;
  assign n19283 = P2_INSTADDRPOINTER_REG_17_ & P2_INSTADDRPOINTER_REG_18_;
  assign n19284 = P2_INSTADDRPOINTER_REG_16_ & n19283;
  assign n19285 = n19084 & n19284;
  assign n19286 = ~n18395 & n19285;
  assign n19287 = ~P2_INSTADDRPOINTER_REG_19_ & ~n19286;
  assign n19288 = P2_INSTADDRPOINTER_REG_19_ & n19285;
  assign n19289 = ~n18395 & n19288;
  assign n19290 = ~n19287 & ~n19289;
  assign n19291 = n17413 & n19290;
  assign n19292 = P2_INSTADDRPOINTER_REG_18_ & n19234;
  assign n19293 = ~P2_INSTADDRPOINTER_REG_18_ & ~n19234;
  assign n19294 = ~n19228 & ~n19293;
  assign n19295 = ~n19292 & ~n19294;
  assign n19296 = P2_EBX_REG_19_ & n14365;
  assign n19297 = ~n18271 & ~n19296;
  assign n19298 = ~n19231 & ~n19297;
  assign n19299 = n19230 & n19297;
  assign n19300 = n19164 & n19299;
  assign n19301 = ~n19298 & ~n19300;
  assign n19302 = ~n17445 & n19301;
  assign n19303 = ~P2_INSTADDRPOINTER_REG_19_ & n19302;
  assign n19304 = P2_INSTADDRPOINTER_REG_19_ & ~n19302;
  assign n19305 = ~n19303 & ~n19304;
  assign n19306 = n19295 & ~n19305;
  assign n19307 = ~n19295 & n19305;
  assign n19308 = ~n19306 & ~n19307;
  assign n19309 = n17458 & ~n19308;
  assign n19310 = P2_INSTADDRPOINTER_REG_19_ & n17410;
  assign n19311 = P2_REIP_REG_19_ & n17461;
  assign n19312 = ~n19310 & ~n19311;
  assign n19313 = P2_INSTADDRPOINTER_REG_18_ & n19245;
  assign n19314 = ~P2_INSTADDRPOINTER_REG_19_ & n19313;
  assign n19315 = P2_INSTADDRPOINTER_REG_19_ & ~n19313;
  assign n19316 = ~n19314 & ~n19315;
  assign n19317 = n17464 & ~n19316;
  assign n19318 = P2_INSTADDRPOINTER_REG_18_ & n19250;
  assign n19319 = ~P2_INSTADDRPOINTER_REG_19_ & n19318;
  assign n19320 = P2_INSTADDRPOINTER_REG_19_ & ~n19318;
  assign n19321 = ~n19319 & ~n19320;
  assign n19322 = n17469 & ~n19321;
  assign n19323 = ~n19317 & ~n19322;
  assign n19324 = n19256 & ~n19263;
  assign n19325 = P2_EBX_REG_19_ & n14995;
  assign n19326 = P2_REIP_REG_19_ & n14997;
  assign n19327 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_19_;
  assign n19328 = P2_INSTADDRPOINTER_REG_19_ & ~n15016;
  assign n19329 = ~n19325 & ~n19326;
  assign n19330 = ~n19327 & n19329;
  assign n19331 = ~n19328 & n19330;
  assign n19332 = n19324 & n19331;
  assign n19333 = ~n19324 & ~n19331;
  assign n19334 = ~n19332 & ~n19333;
  assign n19335 = n17476 & ~n19334;
  assign n19336 = n19268 & ~n19273;
  assign n19337 = P2_REIP_REG_19_ & n17226;
  assign n19338 = P2_EAX_REG_19_ & n17228;
  assign n19339 = ~n19337 & ~n19338;
  assign n19340 = P2_INSTADDRPOINTER_REG_19_ & ~n17236;
  assign n19341 = n19339 & ~n19340;
  assign n19342 = ~n19336 & ~n19341;
  assign n19343 = n19336 & n19341;
  assign n19344 = ~n19342 & ~n19343;
  assign n19345 = n17480 & ~n19344;
  assign n19346 = ~n19335 & ~n19345;
  assign n19347 = ~n19291 & ~n19309;
  assign n19348 = n19312 & n19347;
  assign n19349 = n19323 & n19348;
  assign n3969 = ~n19346 | ~n19349;
  assign n19351 = ~P2_INSTADDRPOINTER_REG_20_ & ~n19289;
  assign n19352 = P2_INSTADDRPOINTER_REG_19_ & P2_INSTADDRPOINTER_REG_20_;
  assign n19353 = n19285 & n19352;
  assign n19354 = ~n18395 & n19353;
  assign n19355 = ~n19351 & ~n19354;
  assign n19356 = n17413 & n19355;
  assign n19357 = ~P2_INSTADDRPOINTER_REG_19_ & ~n19302;
  assign n19358 = P2_INSTADDRPOINTER_REG_19_ & n19302;
  assign n19359 = ~n19292 & ~n19358;
  assign n19360 = ~n19357 & ~n19359;
  assign n19361 = ~n19293 & ~n19357;
  assign n19362 = ~n19228 & n19361;
  assign n19363 = ~n19360 & ~n19362;
  assign n19364 = P2_EBX_REG_20_ & n14365;
  assign n19365 = ~n18271 & ~n19364;
  assign n19366 = n19300 & n19365;
  assign n19367 = ~n19300 & ~n19365;
  assign n19368 = ~n19366 & ~n19367;
  assign n19369 = ~n17445 & n19368;
  assign n19370 = ~P2_INSTADDRPOINTER_REG_20_ & n19369;
  assign n19371 = P2_INSTADDRPOINTER_REG_20_ & ~n19369;
  assign n19372 = ~n19370 & ~n19371;
  assign n19373 = n19363 & ~n19372;
  assign n19374 = ~n19363 & n19372;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = n17458 & ~n19375;
  assign n19377 = P2_INSTADDRPOINTER_REG_20_ & n17410;
  assign n19378 = P2_REIP_REG_20_ & n17461;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = P2_INSTADDRPOINTER_REG_19_ & n19313;
  assign n19381 = ~P2_INSTADDRPOINTER_REG_20_ & n19380;
  assign n19382 = P2_INSTADDRPOINTER_REG_20_ & ~n19380;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = n17464 & ~n19383;
  assign n19385 = P2_INSTADDRPOINTER_REG_19_ & n19318;
  assign n19386 = ~P2_INSTADDRPOINTER_REG_20_ & n19385;
  assign n19387 = P2_INSTADDRPOINTER_REG_20_ & ~n19385;
  assign n19388 = ~n19386 & ~n19387;
  assign n19389 = n17469 & ~n19388;
  assign n19390 = ~n19384 & ~n19389;
  assign n19391 = n19324 & ~n19331;
  assign n19392 = P2_EBX_REG_20_ & n14995;
  assign n19393 = P2_REIP_REG_20_ & n14997;
  assign n19394 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_20_;
  assign n19395 = P2_INSTADDRPOINTER_REG_20_ & ~n15016;
  assign n19396 = ~n19392 & ~n19393;
  assign n19397 = ~n19394 & n19396;
  assign n19398 = ~n19395 & n19397;
  assign n19399 = n19391 & n19398;
  assign n19400 = ~n19391 & ~n19398;
  assign n19401 = ~n19399 & ~n19400;
  assign n19402 = n17476 & ~n19401;
  assign n19403 = n19336 & ~n19341;
  assign n19404 = P2_REIP_REG_20_ & n17226;
  assign n19405 = P2_EAX_REG_20_ & n17228;
  assign n19406 = ~n19404 & ~n19405;
  assign n19407 = P2_INSTADDRPOINTER_REG_20_ & ~n17236;
  assign n19408 = n19406 & ~n19407;
  assign n19409 = ~n19403 & ~n19408;
  assign n19410 = n19403 & n19408;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = n17480 & ~n19411;
  assign n19413 = ~n19402 & ~n19412;
  assign n19414 = ~n19356 & ~n19376;
  assign n19415 = n19379 & n19414;
  assign n19416 = n19390 & n19415;
  assign n3974 = ~n19413 | ~n19416;
  assign n19418 = ~P2_INSTADDRPOINTER_REG_21_ & n19354;
  assign n19419 = P2_INSTADDRPOINTER_REG_21_ & ~n19354;
  assign n19420 = ~n19418 & ~n19419;
  assign n19421 = n17413 & ~n19420;
  assign n19422 = ~P2_INSTADDRPOINTER_REG_20_ & ~n19369;
  assign n19423 = ~n19357 & ~n19422;
  assign n19424 = ~n19359 & n19423;
  assign n19425 = P2_INSTADDRPOINTER_REG_20_ & n19369;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = n19294 & n19423;
  assign n19428 = n19426 & ~n19427;
  assign n19429 = P2_EBX_REG_21_ & n14365;
  assign n19430 = ~n18271 & ~n19429;
  assign n19431 = ~n19366 & ~n19430;
  assign n19432 = n19365 & n19430;
  assign n19433 = n19300 & n19432;
  assign n19434 = ~n19431 & ~n19433;
  assign n19435 = ~n17445 & n19434;
  assign n19436 = ~P2_INSTADDRPOINTER_REG_21_ & n19435;
  assign n19437 = P2_INSTADDRPOINTER_REG_21_ & ~n19435;
  assign n19438 = ~n19436 & ~n19437;
  assign n19439 = n19428 & ~n19438;
  assign n19440 = ~n19428 & n19438;
  assign n19441 = ~n19439 & ~n19440;
  assign n19442 = n17458 & ~n19441;
  assign n19443 = P2_INSTADDRPOINTER_REG_21_ & n17410;
  assign n19444 = P2_REIP_REG_21_ & n17461;
  assign n19445 = ~n19443 & ~n19444;
  assign n19446 = P2_INSTADDRPOINTER_REG_20_ & n19380;
  assign n19447 = ~P2_INSTADDRPOINTER_REG_21_ & n19446;
  assign n19448 = P2_INSTADDRPOINTER_REG_21_ & ~n19446;
  assign n19449 = ~n19447 & ~n19448;
  assign n19450 = n17464 & ~n19449;
  assign n19451 = P2_INSTADDRPOINTER_REG_20_ & n19385;
  assign n19452 = ~P2_INSTADDRPOINTER_REG_21_ & n19451;
  assign n19453 = P2_INSTADDRPOINTER_REG_21_ & ~n19451;
  assign n19454 = ~n19452 & ~n19453;
  assign n19455 = n17469 & ~n19454;
  assign n19456 = ~n19450 & ~n19455;
  assign n19457 = n19391 & ~n19398;
  assign n19458 = P2_EBX_REG_21_ & n14995;
  assign n19459 = P2_REIP_REG_21_ & n14997;
  assign n19460 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_21_;
  assign n19461 = P2_INSTADDRPOINTER_REG_21_ & ~n15016;
  assign n19462 = ~n19458 & ~n19459;
  assign n19463 = ~n19460 & n19462;
  assign n19464 = ~n19461 & n19463;
  assign n19465 = n19457 & n19464;
  assign n19466 = ~n19457 & ~n19464;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = n17476 & ~n19467;
  assign n19469 = n19403 & ~n19408;
  assign n19470 = P2_REIP_REG_21_ & n17226;
  assign n19471 = P2_EAX_REG_21_ & n17228;
  assign n19472 = ~n19470 & ~n19471;
  assign n19473 = P2_INSTADDRPOINTER_REG_21_ & ~n17236;
  assign n19474 = n19472 & ~n19473;
  assign n19475 = ~n19469 & ~n19474;
  assign n19476 = n19469 & n19474;
  assign n19477 = ~n19475 & ~n19476;
  assign n19478 = n17480 & ~n19477;
  assign n19479 = ~n19468 & ~n19478;
  assign n19480 = ~n19421 & ~n19442;
  assign n19481 = n19445 & n19480;
  assign n19482 = n19456 & n19481;
  assign n3979 = ~n19479 | ~n19482;
  assign n19484 = P2_INSTADDRPOINTER_REG_21_ & n19353;
  assign n19485 = ~n18395 & n19484;
  assign n19486 = ~P2_INSTADDRPOINTER_REG_22_ & ~n19485;
  assign n19487 = P2_INSTADDRPOINTER_REG_21_ & P2_INSTADDRPOINTER_REG_22_;
  assign n19488 = n19353 & n19487;
  assign n19489 = ~n18395 & n19488;
  assign n19490 = ~n19486 & ~n19489;
  assign n19491 = n17413 & n19490;
  assign n19492 = P2_INSTADDRPOINTER_REG_21_ & n19435;
  assign n19493 = ~P2_INSTADDRPOINTER_REG_21_ & ~n19435;
  assign n19494 = ~n19428 & ~n19493;
  assign n19495 = ~n19492 & ~n19494;
  assign n19496 = P2_EBX_REG_22_ & n14365;
  assign n19497 = ~n18271 & ~n19496;
  assign n19498 = n19433 & n19497;
  assign n19499 = ~n19433 & ~n19497;
  assign n19500 = ~n19498 & ~n19499;
  assign n19501 = ~n17445 & n19500;
  assign n19502 = ~P2_INSTADDRPOINTER_REG_22_ & n19501;
  assign n19503 = P2_INSTADDRPOINTER_REG_22_ & ~n19501;
  assign n19504 = ~n19502 & ~n19503;
  assign n19505 = n19495 & ~n19504;
  assign n19506 = ~n19495 & n19504;
  assign n19507 = ~n19505 & ~n19506;
  assign n19508 = n17458 & ~n19507;
  assign n19509 = P2_INSTADDRPOINTER_REG_22_ & n17410;
  assign n19510 = P2_REIP_REG_22_ & n17461;
  assign n19511 = ~n19509 & ~n19510;
  assign n19512 = P2_INSTADDRPOINTER_REG_21_ & n19446;
  assign n19513 = ~P2_INSTADDRPOINTER_REG_22_ & n19512;
  assign n19514 = P2_INSTADDRPOINTER_REG_22_ & ~n19512;
  assign n19515 = ~n19513 & ~n19514;
  assign n19516 = n17464 & ~n19515;
  assign n19517 = P2_INSTADDRPOINTER_REG_21_ & n19451;
  assign n19518 = ~P2_INSTADDRPOINTER_REG_22_ & n19517;
  assign n19519 = P2_INSTADDRPOINTER_REG_22_ & ~n19517;
  assign n19520 = ~n19518 & ~n19519;
  assign n19521 = n17469 & ~n19520;
  assign n19522 = ~n19516 & ~n19521;
  assign n19523 = n19457 & ~n19464;
  assign n19524 = P2_EBX_REG_22_ & n14995;
  assign n19525 = P2_REIP_REG_22_ & n14997;
  assign n19526 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_22_;
  assign n19527 = P2_INSTADDRPOINTER_REG_22_ & ~n15016;
  assign n19528 = ~n19524 & ~n19525;
  assign n19529 = ~n19526 & n19528;
  assign n19530 = ~n19527 & n19529;
  assign n19531 = n19523 & n19530;
  assign n19532 = ~n19523 & ~n19530;
  assign n19533 = ~n19531 & ~n19532;
  assign n19534 = n17476 & ~n19533;
  assign n19535 = n19469 & ~n19474;
  assign n19536 = P2_REIP_REG_22_ & n17226;
  assign n19537 = P2_EAX_REG_22_ & n17228;
  assign n19538 = ~n19536 & ~n19537;
  assign n19539 = P2_INSTADDRPOINTER_REG_22_ & ~n17236;
  assign n19540 = n19538 & ~n19539;
  assign n19541 = ~n19535 & ~n19540;
  assign n19542 = n19535 & n19540;
  assign n19543 = ~n19541 & ~n19542;
  assign n19544 = n17480 & ~n19543;
  assign n19545 = ~n19534 & ~n19544;
  assign n19546 = ~n19491 & ~n19508;
  assign n19547 = n19511 & n19546;
  assign n19548 = n19522 & n19547;
  assign n3984 = ~n19545 | ~n19548;
  assign n19550 = ~P2_INSTADDRPOINTER_REG_23_ & ~n19489;
  assign n19551 = P2_INSTADDRPOINTER_REG_22_ & P2_INSTADDRPOINTER_REG_23_;
  assign n19552 = P2_INSTADDRPOINTER_REG_21_ & n19551;
  assign n19553 = n19353 & n19552;
  assign n19554 = ~n18395 & n19553;
  assign n19555 = ~n19550 & ~n19554;
  assign n19556 = n17413 & n19555;
  assign n19557 = ~P2_INSTADDRPOINTER_REG_22_ & ~n19501;
  assign n19558 = n19492 & ~n19557;
  assign n19559 = P2_INSTADDRPOINTER_REG_22_ & n19501;
  assign n19560 = ~n19558 & ~n19559;
  assign n19561 = ~n19493 & ~n19557;
  assign n19562 = ~n19428 & n19561;
  assign n19563 = n19560 & ~n19562;
  assign n19564 = P2_EBX_REG_23_ & n14365;
  assign n19565 = ~n18271 & ~n19564;
  assign n19566 = ~n19498 & ~n19565;
  assign n19567 = n19497 & n19565;
  assign n19568 = n19433 & n19567;
  assign n19569 = ~n19566 & ~n19568;
  assign n19570 = ~n17445 & n19569;
  assign n19571 = ~P2_INSTADDRPOINTER_REG_23_ & n19570;
  assign n19572 = P2_INSTADDRPOINTER_REG_23_ & ~n19570;
  assign n19573 = ~n19571 & ~n19572;
  assign n19574 = n19563 & ~n19573;
  assign n19575 = ~n19563 & n19573;
  assign n19576 = ~n19574 & ~n19575;
  assign n19577 = n17458 & ~n19576;
  assign n19578 = P2_INSTADDRPOINTER_REG_23_ & n17410;
  assign n19579 = P2_REIP_REG_23_ & n17461;
  assign n19580 = ~n19578 & ~n19579;
  assign n19581 = P2_INSTADDRPOINTER_REG_22_ & n19512;
  assign n19582 = ~P2_INSTADDRPOINTER_REG_23_ & n19581;
  assign n19583 = P2_INSTADDRPOINTER_REG_23_ & ~n19581;
  assign n19584 = ~n19582 & ~n19583;
  assign n19585 = n17464 & ~n19584;
  assign n19586 = P2_INSTADDRPOINTER_REG_22_ & n19517;
  assign n19587 = ~P2_INSTADDRPOINTER_REG_23_ & n19586;
  assign n19588 = P2_INSTADDRPOINTER_REG_23_ & ~n19586;
  assign n19589 = ~n19587 & ~n19588;
  assign n19590 = n17469 & ~n19589;
  assign n19591 = ~n19585 & ~n19590;
  assign n19592 = n19523 & ~n19530;
  assign n19593 = P2_EBX_REG_23_ & n14995;
  assign n19594 = P2_REIP_REG_23_ & n14997;
  assign n19595 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_23_;
  assign n19596 = P2_INSTADDRPOINTER_REG_23_ & ~n15016;
  assign n19597 = ~n19593 & ~n19594;
  assign n19598 = ~n19595 & n19597;
  assign n19599 = ~n19596 & n19598;
  assign n19600 = n19592 & n19599;
  assign n19601 = ~n19592 & ~n19599;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = n17476 & ~n19602;
  assign n19604 = n19535 & ~n19540;
  assign n19605 = P2_REIP_REG_23_ & n17226;
  assign n19606 = P2_EAX_REG_23_ & n17228;
  assign n19607 = ~n19605 & ~n19606;
  assign n19608 = P2_INSTADDRPOINTER_REG_23_ & ~n17236;
  assign n19609 = n19607 & ~n19608;
  assign n19610 = ~n19604 & ~n19609;
  assign n19611 = n19604 & n19609;
  assign n19612 = ~n19610 & ~n19611;
  assign n19613 = n17480 & ~n19612;
  assign n19614 = ~n19603 & ~n19613;
  assign n19615 = ~n19556 & ~n19577;
  assign n19616 = n19580 & n19615;
  assign n19617 = n19591 & n19616;
  assign n3989 = ~n19614 | ~n19617;
  assign n19619 = ~P2_INSTADDRPOINTER_REG_24_ & n19554;
  assign n19620 = P2_INSTADDRPOINTER_REG_24_ & ~n19554;
  assign n19621 = ~n19619 & ~n19620;
  assign n19622 = n17413 & ~n19621;
  assign n19623 = P2_INSTADDRPOINTER_REG_23_ & n19570;
  assign n19624 = ~P2_INSTADDRPOINTER_REG_23_ & ~n19570;
  assign n19625 = ~n19563 & ~n19624;
  assign n19626 = ~n19623 & ~n19625;
  assign n19627 = P2_EBX_REG_24_ & n14365;
  assign n19628 = ~n18271 & ~n19627;
  assign n19629 = n19568 & n19628;
  assign n19630 = ~n19568 & ~n19628;
  assign n19631 = ~n19629 & ~n19630;
  assign n19632 = ~n17445 & n19631;
  assign n19633 = ~P2_INSTADDRPOINTER_REG_24_ & n19632;
  assign n19634 = P2_INSTADDRPOINTER_REG_24_ & ~n19632;
  assign n19635 = ~n19633 & ~n19634;
  assign n19636 = n19626 & ~n19635;
  assign n19637 = ~n19626 & n19635;
  assign n19638 = ~n19636 & ~n19637;
  assign n19639 = n17458 & ~n19638;
  assign n19640 = P2_INSTADDRPOINTER_REG_24_ & n17410;
  assign n19641 = P2_REIP_REG_24_ & n17461;
  assign n19642 = ~n19640 & ~n19641;
  assign n19643 = P2_INSTADDRPOINTER_REG_23_ & n19581;
  assign n19644 = ~P2_INSTADDRPOINTER_REG_24_ & n19643;
  assign n19645 = P2_INSTADDRPOINTER_REG_24_ & ~n19643;
  assign n19646 = ~n19644 & ~n19645;
  assign n19647 = n17464 & ~n19646;
  assign n19648 = P2_INSTADDRPOINTER_REG_23_ & n19586;
  assign n19649 = ~P2_INSTADDRPOINTER_REG_24_ & n19648;
  assign n19650 = P2_INSTADDRPOINTER_REG_24_ & ~n19648;
  assign n19651 = ~n19649 & ~n19650;
  assign n19652 = n17469 & ~n19651;
  assign n19653 = ~n19647 & ~n19652;
  assign n19654 = n19592 & ~n19599;
  assign n19655 = P2_EBX_REG_24_ & n14995;
  assign n19656 = P2_REIP_REG_24_ & n14997;
  assign n19657 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_24_;
  assign n19658 = P2_INSTADDRPOINTER_REG_24_ & ~n15016;
  assign n19659 = ~n19655 & ~n19656;
  assign n19660 = ~n19657 & n19659;
  assign n19661 = ~n19658 & n19660;
  assign n19662 = n19654 & n19661;
  assign n19663 = ~n19654 & ~n19661;
  assign n19664 = ~n19662 & ~n19663;
  assign n19665 = n17476 & ~n19664;
  assign n19666 = n19604 & ~n19609;
  assign n19667 = P2_REIP_REG_24_ & n17226;
  assign n19668 = P2_EAX_REG_24_ & n17228;
  assign n19669 = ~n19667 & ~n19668;
  assign n19670 = P2_INSTADDRPOINTER_REG_24_ & ~n17236;
  assign n19671 = n19669 & ~n19670;
  assign n19672 = ~n19666 & ~n19671;
  assign n19673 = n19666 & n19671;
  assign n19674 = ~n19672 & ~n19673;
  assign n19675 = n17480 & ~n19674;
  assign n19676 = ~n19665 & ~n19675;
  assign n19677 = ~n19622 & ~n19639;
  assign n19678 = n19642 & n19677;
  assign n19679 = n19653 & n19678;
  assign n3994 = ~n19676 | ~n19679;
  assign n19681 = P2_INSTADDRPOINTER_REG_24_ & n19553;
  assign n19682 = ~n18395 & n19681;
  assign n19683 = ~P2_INSTADDRPOINTER_REG_25_ & n19682;
  assign n19684 = P2_INSTADDRPOINTER_REG_25_ & ~n19682;
  assign n19685 = ~n19683 & ~n19684;
  assign n19686 = n17413 & ~n19685;
  assign n19687 = ~P2_INSTADDRPOINTER_REG_24_ & ~n19632;
  assign n19688 = n19623 & ~n19687;
  assign n19689 = P2_INSTADDRPOINTER_REG_24_ & n19632;
  assign n19690 = ~n19688 & ~n19689;
  assign n19691 = ~n19624 & ~n19687;
  assign n19692 = ~n19563 & n19691;
  assign n19693 = n19690 & ~n19692;
  assign n19694 = ~P2_INSTADDRPOINTER_REG_25_ & n19693;
  assign n19695 = P2_INSTADDRPOINTER_REG_25_ & ~n19693;
  assign n19696 = ~n19694 & ~n19695;
  assign n19697 = P2_EBX_REG_25_ & n14365;
  assign n19698 = ~n18271 & ~n19697;
  assign n19699 = ~n19629 & ~n19698;
  assign n19700 = n19628 & n19698;
  assign n19701 = n19568 & n19700;
  assign n19702 = ~n19699 & ~n19701;
  assign n19703 = ~n17445 & n19702;
  assign n19704 = ~n19696 & n19703;
  assign n19705 = n19696 & ~n19703;
  assign n19706 = ~n19704 & ~n19705;
  assign n19707 = n17458 & ~n19706;
  assign n19708 = P2_INSTADDRPOINTER_REG_25_ & n17410;
  assign n19709 = P2_REIP_REG_25_ & n17461;
  assign n19710 = ~n19708 & ~n19709;
  assign n19711 = P2_INSTADDRPOINTER_REG_24_ & n19643;
  assign n19712 = ~P2_INSTADDRPOINTER_REG_25_ & n19711;
  assign n19713 = P2_INSTADDRPOINTER_REG_25_ & ~n19711;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = n17464 & ~n19714;
  assign n19716 = P2_INSTADDRPOINTER_REG_24_ & n19648;
  assign n19717 = ~P2_INSTADDRPOINTER_REG_25_ & n19716;
  assign n19718 = P2_INSTADDRPOINTER_REG_25_ & ~n19716;
  assign n19719 = ~n19717 & ~n19718;
  assign n19720 = n17469 & ~n19719;
  assign n19721 = ~n19715 & ~n19720;
  assign n19722 = n19654 & ~n19661;
  assign n19723 = P2_EBX_REG_25_ & n14995;
  assign n19724 = P2_REIP_REG_25_ & n14997;
  assign n19725 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_25_;
  assign n19726 = P2_INSTADDRPOINTER_REG_25_ & ~n15016;
  assign n19727 = ~n19723 & ~n19724;
  assign n19728 = ~n19725 & n19727;
  assign n19729 = ~n19726 & n19728;
  assign n19730 = n19722 & n19729;
  assign n19731 = ~n19722 & ~n19729;
  assign n19732 = ~n19730 & ~n19731;
  assign n19733 = n17476 & ~n19732;
  assign n19734 = n19666 & ~n19671;
  assign n19735 = P2_REIP_REG_25_ & n17226;
  assign n19736 = P2_EAX_REG_25_ & n17228;
  assign n19737 = ~n19735 & ~n19736;
  assign n19738 = P2_INSTADDRPOINTER_REG_25_ & ~n17236;
  assign n19739 = n19737 & ~n19738;
  assign n19740 = ~n19734 & ~n19739;
  assign n19741 = n19734 & n19739;
  assign n19742 = ~n19740 & ~n19741;
  assign n19743 = n17480 & ~n19742;
  assign n19744 = ~n19733 & ~n19743;
  assign n19745 = ~n19686 & ~n19707;
  assign n19746 = n19710 & n19745;
  assign n19747 = n19721 & n19746;
  assign n3999 = ~n19744 | ~n19747;
  assign n19749 = P2_INSTADDRPOINTER_REG_24_ & P2_INSTADDRPOINTER_REG_25_;
  assign n19750 = n19553 & n19749;
  assign n19751 = ~n18395 & n19750;
  assign n19752 = ~P2_INSTADDRPOINTER_REG_26_ & ~n19751;
  assign n19753 = P2_INSTADDRPOINTER_REG_25_ & P2_INSTADDRPOINTER_REG_26_;
  assign n19754 = P2_INSTADDRPOINTER_REG_24_ & n19753;
  assign n19755 = n19553 & n19754;
  assign n19756 = ~n18395 & n19755;
  assign n19757 = ~n19752 & ~n19756;
  assign n19758 = n17413 & n19757;
  assign n19759 = ~n19693 & n19703;
  assign n19760 = P2_INSTADDRPOINTER_REG_25_ & n19703;
  assign n19761 = ~n19695 & ~n19759;
  assign n19762 = ~n19760 & n19761;
  assign n19763 = P2_EBX_REG_26_ & n14365;
  assign n19764 = ~n18271 & ~n19763;
  assign n19765 = n19701 & n19764;
  assign n19766 = ~n19701 & ~n19764;
  assign n19767 = ~n19765 & ~n19766;
  assign n19768 = ~n17445 & n19767;
  assign n19769 = ~P2_INSTADDRPOINTER_REG_26_ & n19768;
  assign n19770 = P2_INSTADDRPOINTER_REG_26_ & ~n19768;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = n19762 & ~n19771;
  assign n19773 = ~n19762 & n19771;
  assign n19774 = ~n19772 & ~n19773;
  assign n19775 = n17458 & ~n19774;
  assign n19776 = P2_INSTADDRPOINTER_REG_26_ & n17410;
  assign n19777 = P2_REIP_REG_26_ & n17461;
  assign n19778 = ~n19776 & ~n19777;
  assign n19779 = P2_INSTADDRPOINTER_REG_25_ & n19711;
  assign n19780 = ~P2_INSTADDRPOINTER_REG_26_ & n19779;
  assign n19781 = P2_INSTADDRPOINTER_REG_26_ & ~n19779;
  assign n19782 = ~n19780 & ~n19781;
  assign n19783 = n17464 & ~n19782;
  assign n19784 = P2_INSTADDRPOINTER_REG_25_ & n19716;
  assign n19785 = ~P2_INSTADDRPOINTER_REG_26_ & n19784;
  assign n19786 = P2_INSTADDRPOINTER_REG_26_ & ~n19784;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = n17469 & ~n19787;
  assign n19789 = ~n19783 & ~n19788;
  assign n19790 = n19722 & ~n19729;
  assign n19791 = P2_EBX_REG_26_ & n14995;
  assign n19792 = P2_REIP_REG_26_ & n14997;
  assign n19793 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_26_;
  assign n19794 = P2_INSTADDRPOINTER_REG_26_ & ~n15016;
  assign n19795 = ~n19791 & ~n19792;
  assign n19796 = ~n19793 & n19795;
  assign n19797 = ~n19794 & n19796;
  assign n19798 = n19790 & n19797;
  assign n19799 = ~n19790 & ~n19797;
  assign n19800 = ~n19798 & ~n19799;
  assign n19801 = n17476 & ~n19800;
  assign n19802 = n19734 & ~n19739;
  assign n19803 = P2_REIP_REG_26_ & n17226;
  assign n19804 = P2_EAX_REG_26_ & n17228;
  assign n19805 = ~n19803 & ~n19804;
  assign n19806 = P2_INSTADDRPOINTER_REG_26_ & ~n17236;
  assign n19807 = n19805 & ~n19806;
  assign n19808 = ~n19802 & ~n19807;
  assign n19809 = n19802 & n19807;
  assign n19810 = ~n19808 & ~n19809;
  assign n19811 = n17480 & ~n19810;
  assign n19812 = ~n19801 & ~n19811;
  assign n19813 = ~n19758 & ~n19775;
  assign n19814 = n19778 & n19813;
  assign n19815 = n19789 & n19814;
  assign n4004 = ~n19812 | ~n19815;
  assign n19817 = ~P2_INSTADDRPOINTER_REG_27_ & n19756;
  assign n19818 = P2_INSTADDRPOINTER_REG_27_ & ~n19756;
  assign n19819 = ~n19817 & ~n19818;
  assign n19820 = n17413 & ~n19819;
  assign n19821 = P2_INSTADDRPOINTER_REG_26_ & n19768;
  assign n19822 = ~P2_INSTADDRPOINTER_REG_26_ & ~n19768;
  assign n19823 = ~n19762 & ~n19822;
  assign n19824 = ~n19821 & ~n19823;
  assign n19825 = P2_EBX_REG_27_ & n14365;
  assign n19826 = ~n18271 & ~n19825;
  assign n19827 = ~n19765 & ~n19826;
  assign n19828 = n19764 & n19826;
  assign n19829 = n19701 & n19828;
  assign n19830 = ~n19827 & ~n19829;
  assign n19831 = ~n17445 & n19830;
  assign n19832 = ~P2_INSTADDRPOINTER_REG_27_ & n19831;
  assign n19833 = P2_INSTADDRPOINTER_REG_27_ & ~n19831;
  assign n19834 = ~n19832 & ~n19833;
  assign n19835 = n19824 & ~n19834;
  assign n19836 = ~n19824 & n19834;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = n17458 & ~n19837;
  assign n19839 = P2_INSTADDRPOINTER_REG_27_ & n17410;
  assign n19840 = P2_REIP_REG_27_ & n17461;
  assign n19841 = ~n19839 & ~n19840;
  assign n19842 = P2_INSTADDRPOINTER_REG_26_ & n19779;
  assign n19843 = ~P2_INSTADDRPOINTER_REG_27_ & n19842;
  assign n19844 = P2_INSTADDRPOINTER_REG_27_ & ~n19842;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = n17464 & ~n19845;
  assign n19847 = P2_INSTADDRPOINTER_REG_26_ & n19784;
  assign n19848 = ~P2_INSTADDRPOINTER_REG_27_ & n19847;
  assign n19849 = P2_INSTADDRPOINTER_REG_27_ & ~n19847;
  assign n19850 = ~n19848 & ~n19849;
  assign n19851 = n17469 & ~n19850;
  assign n19852 = ~n19846 & ~n19851;
  assign n19853 = n19790 & ~n19797;
  assign n19854 = P2_EBX_REG_27_ & n14995;
  assign n19855 = P2_REIP_REG_27_ & n14997;
  assign n19856 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_27_;
  assign n19857 = P2_INSTADDRPOINTER_REG_27_ & ~n15016;
  assign n19858 = ~n19854 & ~n19855;
  assign n19859 = ~n19856 & n19858;
  assign n19860 = ~n19857 & n19859;
  assign n19861 = n19853 & n19860;
  assign n19862 = ~n19853 & ~n19860;
  assign n19863 = ~n19861 & ~n19862;
  assign n19864 = n17476 & ~n19863;
  assign n19865 = n19802 & ~n19807;
  assign n19866 = P2_REIP_REG_27_ & n17226;
  assign n19867 = P2_EAX_REG_27_ & n17228;
  assign n19868 = ~n19866 & ~n19867;
  assign n19869 = P2_INSTADDRPOINTER_REG_27_ & ~n17236;
  assign n19870 = n19868 & ~n19869;
  assign n19871 = ~n19865 & ~n19870;
  assign n19872 = n19865 & n19870;
  assign n19873 = ~n19871 & ~n19872;
  assign n19874 = n17480 & ~n19873;
  assign n19875 = ~n19864 & ~n19874;
  assign n19876 = ~n19820 & ~n19838;
  assign n19877 = n19841 & n19876;
  assign n19878 = n19852 & n19877;
  assign n4009 = ~n19875 | ~n19878;
  assign n19880 = P2_INSTADDRPOINTER_REG_27_ & n19755;
  assign n19881 = ~n18395 & n19880;
  assign n19882 = ~P2_INSTADDRPOINTER_REG_28_ & ~n19881;
  assign n19883 = P2_INSTADDRPOINTER_REG_27_ & P2_INSTADDRPOINTER_REG_28_;
  assign n19884 = n19755 & n19883;
  assign n19885 = ~n18395 & n19884;
  assign n19886 = ~n19882 & ~n19885;
  assign n19887 = n17413 & n19886;
  assign n19888 = ~P2_INSTADDRPOINTER_REG_27_ & ~n19831;
  assign n19889 = n19821 & ~n19888;
  assign n19890 = P2_INSTADDRPOINTER_REG_27_ & n19831;
  assign n19891 = ~n19889 & ~n19890;
  assign n19892 = ~n19822 & ~n19888;
  assign n19893 = ~n19762 & n19892;
  assign n19894 = n19891 & ~n19893;
  assign n19895 = P2_EBX_REG_28_ & n14365;
  assign n19896 = ~n18271 & ~n19895;
  assign n19897 = n19829 & n19896;
  assign n19898 = ~n19829 & ~n19896;
  assign n19899 = ~n19897 & ~n19898;
  assign n19900 = ~n17445 & n19899;
  assign n19901 = ~P2_INSTADDRPOINTER_REG_28_ & n19900;
  assign n19902 = P2_INSTADDRPOINTER_REG_28_ & ~n19900;
  assign n19903 = ~n19901 & ~n19902;
  assign n19904 = n19894 & ~n19903;
  assign n19905 = ~n19894 & n19903;
  assign n19906 = ~n19904 & ~n19905;
  assign n19907 = n17458 & ~n19906;
  assign n19908 = P2_INSTADDRPOINTER_REG_28_ & n17410;
  assign n19909 = P2_REIP_REG_28_ & n17461;
  assign n19910 = ~n19908 & ~n19909;
  assign n19911 = P2_INSTADDRPOINTER_REG_27_ & n19842;
  assign n19912 = ~P2_INSTADDRPOINTER_REG_28_ & n19911;
  assign n19913 = P2_INSTADDRPOINTER_REG_28_ & ~n19911;
  assign n19914 = ~n19912 & ~n19913;
  assign n19915 = n17464 & ~n19914;
  assign n19916 = P2_INSTADDRPOINTER_REG_27_ & n19847;
  assign n19917 = ~P2_INSTADDRPOINTER_REG_28_ & n19916;
  assign n19918 = P2_INSTADDRPOINTER_REG_28_ & ~n19916;
  assign n19919 = ~n19917 & ~n19918;
  assign n19920 = n17469 & ~n19919;
  assign n19921 = ~n19915 & ~n19920;
  assign n19922 = n19853 & ~n19860;
  assign n19923 = P2_EBX_REG_28_ & n14995;
  assign n19924 = P2_REIP_REG_28_ & n14997;
  assign n19925 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_28_;
  assign n19926 = P2_INSTADDRPOINTER_REG_28_ & ~n15016;
  assign n19927 = ~n19923 & ~n19924;
  assign n19928 = ~n19925 & n19927;
  assign n19929 = ~n19926 & n19928;
  assign n19930 = n19922 & n19929;
  assign n19931 = ~n19922 & ~n19929;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = n17476 & ~n19932;
  assign n19934 = n19865 & ~n19870;
  assign n19935 = P2_REIP_REG_28_ & n17226;
  assign n19936 = P2_EAX_REG_28_ & n17228;
  assign n19937 = ~n19935 & ~n19936;
  assign n19938 = P2_INSTADDRPOINTER_REG_28_ & ~n17236;
  assign n19939 = n19937 & ~n19938;
  assign n19940 = ~n19934 & ~n19939;
  assign n19941 = n19934 & n19939;
  assign n19942 = ~n19940 & ~n19941;
  assign n19943 = n17480 & ~n19942;
  assign n19944 = ~n19933 & ~n19943;
  assign n19945 = ~n19887 & ~n19907;
  assign n19946 = n19910 & n19945;
  assign n19947 = n19921 & n19946;
  assign n4014 = ~n19944 | ~n19947;
  assign n19949 = ~P2_INSTADDRPOINTER_REG_29_ & ~n19885;
  assign n19950 = P2_INSTADDRPOINTER_REG_28_ & P2_INSTADDRPOINTER_REG_29_;
  assign n19951 = P2_INSTADDRPOINTER_REG_27_ & n19950;
  assign n19952 = n19755 & n19951;
  assign n19953 = ~n18395 & n19952;
  assign n19954 = ~n19949 & ~n19953;
  assign n19955 = n17413 & n19954;
  assign n19956 = ~P2_INSTADDRPOINTER_REG_28_ & ~n19900;
  assign n19957 = ~n19891 & ~n19956;
  assign n19958 = P2_INSTADDRPOINTER_REG_28_ & n19900;
  assign n19959 = ~n19957 & ~n19958;
  assign n19960 = ~n19888 & ~n19956;
  assign n19961 = ~n19822 & n19960;
  assign n19962 = ~n19762 & n19961;
  assign n19963 = n19959 & ~n19962;
  assign n19964 = P2_EBX_REG_29_ & n14365;
  assign n19965 = ~n18271 & ~n19964;
  assign n19966 = ~n19897 & ~n19965;
  assign n19967 = n19896 & n19965;
  assign n19968 = n19829 & n19967;
  assign n19969 = ~n19966 & ~n19968;
  assign n19970 = ~n17445 & n19969;
  assign n19971 = ~P2_INSTADDRPOINTER_REG_29_ & n19970;
  assign n19972 = P2_INSTADDRPOINTER_REG_29_ & ~n19970;
  assign n19973 = ~n19971 & ~n19972;
  assign n19974 = n19963 & ~n19973;
  assign n19975 = ~n19963 & n19973;
  assign n19976 = ~n19974 & ~n19975;
  assign n19977 = n17458 & ~n19976;
  assign n19978 = P2_INSTADDRPOINTER_REG_29_ & n17410;
  assign n19979 = P2_REIP_REG_29_ & n17461;
  assign n19980 = ~n19978 & ~n19979;
  assign n19981 = P2_INSTADDRPOINTER_REG_28_ & n19911;
  assign n19982 = ~P2_INSTADDRPOINTER_REG_29_ & n19981;
  assign n19983 = P2_INSTADDRPOINTER_REG_29_ & ~n19981;
  assign n19984 = ~n19982 & ~n19983;
  assign n19985 = n17464 & ~n19984;
  assign n19986 = P2_INSTADDRPOINTER_REG_28_ & n19916;
  assign n19987 = ~P2_INSTADDRPOINTER_REG_29_ & n19986;
  assign n19988 = P2_INSTADDRPOINTER_REG_29_ & ~n19986;
  assign n19989 = ~n19987 & ~n19988;
  assign n19990 = n17469 & ~n19989;
  assign n19991 = n19922 & ~n19929;
  assign n19992 = P2_EBX_REG_29_ & n14995;
  assign n19993 = P2_REIP_REG_29_ & n14997;
  assign n19994 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_29_;
  assign n19995 = P2_INSTADDRPOINTER_REG_29_ & ~n15016;
  assign n19996 = ~n19992 & ~n19993;
  assign n19997 = ~n19994 & n19996;
  assign n19998 = ~n19995 & n19997;
  assign n19999 = n19991 & n19998;
  assign n20000 = ~n19991 & ~n19998;
  assign n20001 = ~n19999 & ~n20000;
  assign n20002 = n17476 & ~n20001;
  assign n20003 = n19934 & ~n19939;
  assign n20004 = P2_REIP_REG_29_ & n17226;
  assign n20005 = P2_EAX_REG_29_ & n17228;
  assign n20006 = ~n20004 & ~n20005;
  assign n20007 = P2_INSTADDRPOINTER_REG_29_ & ~n17236;
  assign n20008 = n20006 & ~n20007;
  assign n20009 = ~n20003 & ~n20008;
  assign n20010 = n20003 & n20008;
  assign n20011 = ~n20009 & ~n20010;
  assign n20012 = n17480 & ~n20011;
  assign n20013 = ~n19985 & ~n19990;
  assign n20014 = ~n20002 & n20013;
  assign n20015 = ~n20012 & n20014;
  assign n20016 = ~n19955 & ~n19977;
  assign n20017 = n19980 & n20016;
  assign n4019 = ~n20015 | ~n20017;
  assign n20019 = ~P2_INSTADDRPOINTER_REG_30_ & n19953;
  assign n20020 = P2_INSTADDRPOINTER_REG_30_ & ~n19953;
  assign n20021 = ~n20019 & ~n20020;
  assign n20022 = n17413 & ~n20021;
  assign n20023 = P2_INSTADDRPOINTER_REG_29_ & n19970;
  assign n20024 = ~P2_INSTADDRPOINTER_REG_29_ & ~n19970;
  assign n20025 = ~n19963 & ~n20024;
  assign n20026 = ~n20023 & ~n20025;
  assign n20027 = P2_EBX_REG_30_ & n14365;
  assign n20028 = ~n18271 & ~n20027;
  assign n20029 = ~n19968 & ~n20028;
  assign n20030 = n19968 & n20028;
  assign n20031 = ~n20029 & ~n20030;
  assign n20032 = ~n17445 & n20031;
  assign n20033 = ~P2_INSTADDRPOINTER_REG_30_ & n20032;
  assign n20034 = P2_INSTADDRPOINTER_REG_30_ & ~n20032;
  assign n20035 = ~n20033 & ~n20034;
  assign n20036 = n20026 & ~n20035;
  assign n20037 = ~n20026 & n20035;
  assign n20038 = ~n20036 & ~n20037;
  assign n20039 = n17458 & ~n20038;
  assign n20040 = P2_INSTADDRPOINTER_REG_30_ & n17410;
  assign n20041 = P2_REIP_REG_30_ & n17461;
  assign n20042 = ~n20040 & ~n20041;
  assign n20043 = P2_INSTADDRPOINTER_REG_29_ & n19981;
  assign n20044 = ~P2_INSTADDRPOINTER_REG_30_ & n20043;
  assign n20045 = P2_INSTADDRPOINTER_REG_30_ & ~n20043;
  assign n20046 = ~n20044 & ~n20045;
  assign n20047 = n17464 & ~n20046;
  assign n20048 = P2_INSTADDRPOINTER_REG_29_ & n19986;
  assign n20049 = ~P2_INSTADDRPOINTER_REG_30_ & n20048;
  assign n20050 = P2_INSTADDRPOINTER_REG_30_ & ~n20048;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = n17469 & ~n20051;
  assign n20053 = n19991 & ~n19998;
  assign n20054 = P2_EBX_REG_30_ & n14995;
  assign n20055 = P2_REIP_REG_30_ & n14997;
  assign n20056 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_30_;
  assign n20057 = P2_INSTADDRPOINTER_REG_30_ & ~n15016;
  assign n20058 = ~n20054 & ~n20055;
  assign n20059 = ~n20056 & n20058;
  assign n20060 = ~n20057 & n20059;
  assign n20061 = n20053 & n20060;
  assign n20062 = ~n20053 & ~n20060;
  assign n20063 = ~n20061 & ~n20062;
  assign n20064 = n17476 & ~n20063;
  assign n20065 = ~n20047 & ~n20052;
  assign n20066 = ~n20064 & n20065;
  assign n20067 = P2_REIP_REG_30_ & n17226;
  assign n20068 = P2_EAX_REG_30_ & n17228;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = P2_INSTADDRPOINTER_REG_30_ & ~n17236;
  assign n20071 = n20069 & ~n20070;
  assign n20072 = n20003 & ~n20008;
  assign n20073 = ~n20071 & ~n20072;
  assign n20074 = n20071 & n20072;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = n17480 & ~n20075;
  assign n20077 = ~n20022 & ~n20039;
  assign n20078 = n20042 & n20077;
  assign n20079 = n20066 & n20078;
  assign n4024 = n20076 | ~n20079;
  assign n20081 = P2_INSTADDRPOINTER_REG_30_ & n19952;
  assign n20082 = ~n18395 & n20081;
  assign n20083 = ~P2_INSTADDRPOINTER_REG_31_ & n20082;
  assign n20084 = P2_INSTADDRPOINTER_REG_31_ & ~n20082;
  assign n20085 = ~n20083 & ~n20084;
  assign n20086 = n17413 & ~n20085;
  assign n20087 = P2_EBX_REG_31_ & n14365;
  assign n20088 = ~n18271 & ~n20087;
  assign n20089 = n20030 & n20088;
  assign n20090 = ~n20030 & ~n20088;
  assign n20091 = ~n20089 & ~n20090;
  assign n20092 = ~n17445 & n20091;
  assign n20093 = ~P2_INSTADDRPOINTER_REG_31_ & n20092;
  assign n20094 = P2_INSTADDRPOINTER_REG_31_ & ~n20092;
  assign n20095 = ~n20093 & ~n20094;
  assign n20096 = n20032 & ~n20095;
  assign n20097 = P2_INSTADDRPOINTER_REG_30_ & n20096;
  assign n20098 = ~n20032 & n20095;
  assign n20099 = ~P2_INSTADDRPOINTER_REG_30_ & n20098;
  assign n20100 = ~n20097 & ~n20099;
  assign n20101 = P2_INSTADDRPOINTER_REG_30_ & n20032;
  assign n20102 = ~n20023 & ~n20101;
  assign n20103 = n20095 & n20102;
  assign n20104 = ~n20025 & n20103;
  assign n20105 = ~P2_INSTADDRPOINTER_REG_30_ & ~n20032;
  assign n20106 = ~n20024 & ~n20105;
  assign n20107 = ~n20095 & n20106;
  assign n20108 = ~n19958 & ~n20023;
  assign n20109 = ~n19957 & ~n19962;
  assign n20110 = n20108 & n20109;
  assign n20111 = n20107 & ~n20110;
  assign n20112 = n20100 & ~n20104;
  assign n20113 = ~n20111 & n20112;
  assign n20114 = n17458 & n20113;
  assign n20115 = P2_INSTADDRPOINTER_REG_31_ & n17410;
  assign n20116 = P2_REIP_REG_31_ & n17461;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = P2_INSTADDRPOINTER_REG_30_ & n20043;
  assign n20119 = ~P2_INSTADDRPOINTER_REG_31_ & n20118;
  assign n20120 = P2_INSTADDRPOINTER_REG_31_ & ~n20118;
  assign n20121 = ~n20119 & ~n20120;
  assign n20122 = n17464 & ~n20121;
  assign n20123 = P2_INSTADDRPOINTER_REG_30_ & n20048;
  assign n20124 = ~P2_INSTADDRPOINTER_REG_31_ & n20123;
  assign n20125 = P2_INSTADDRPOINTER_REG_31_ & ~n20123;
  assign n20126 = ~n20124 & ~n20125;
  assign n20127 = n17469 & ~n20126;
  assign n20128 = n20053 & ~n20060;
  assign n20129 = P2_EBX_REG_31_ & n14995;
  assign n20130 = P2_REIP_REG_31_ & n14997;
  assign n20131 = P2_STATE2_REG_1_ & P2_PHYADDRPOINTER_REG_31_;
  assign n20132 = P2_INSTADDRPOINTER_REG_31_ & ~n15016;
  assign n20133 = ~n20129 & ~n20130;
  assign n20134 = ~n20131 & n20133;
  assign n20135 = ~n20132 & n20134;
  assign n20136 = n20128 & n20135;
  assign n20137 = ~n20128 & ~n20135;
  assign n20138 = ~n20136 & ~n20137;
  assign n20139 = n17476 & ~n20138;
  assign n20140 = ~n20122 & ~n20127;
  assign n20141 = ~n20139 & n20140;
  assign n20142 = P2_REIP_REG_31_ & n17226;
  assign n20143 = P2_EAX_REG_31_ & n17228;
  assign n20144 = ~n20142 & ~n20143;
  assign n20145 = P2_INSTADDRPOINTER_REG_31_ & ~n17236;
  assign n20146 = n20144 & ~n20145;
  assign n20147 = ~n20071 & ~n20146;
  assign n20148 = n20072 & n20147;
  assign n20149 = ~n20071 & n20072;
  assign n20150 = n20146 & ~n20149;
  assign n20151 = ~n20148 & ~n20150;
  assign n20152 = n17480 & n20151;
  assign n20153 = ~n20086 & ~n20114;
  assign n20154 = n20117 & n20153;
  assign n20155 = n20141 & n20154;
  assign n4029 = n20152 | ~n20155;
  assign n20157 = ~P2_STATE2_REG_0_ & ~n17335;
  assign n20158 = n15047 & n15432;
  assign n20159 = ~n15391 & n20158;
  assign n20160 = ~n20157 & ~n20159;
  assign n20161 = n15482 & ~n20160;
  assign n20162 = ~n17457 & n20161;
  assign n20163 = n15446 & ~n20160;
  assign n20164 = P2_REIP_REG_0_ & n20163;
  assign n20165 = P2_PHYADDRPOINTER_REG_0_ & n20160;
  assign n20166 = ~n20162 & ~n20164;
  assign n20167 = ~n20165 & n20166;
  assign n20168 = n14857 & ~n20160;
  assign n20169 = ~n17385 & n20168;
  assign n20170 = ~n15440 & ~n15495;
  assign n20171 = ~n20160 & ~n20170;
  assign n20172 = P2_PHYADDRPOINTER_REG_0_ & n20171;
  assign n20173 = P2_STATE2_REG_1_ & P2_STATEBS16_REG;
  assign n20174 = ~n20160 & n20173;
  assign n20175 = ~n15277 & n20174;
  assign n20176 = ~n20169 & ~n20172;
  assign n20177 = ~n20175 & n20176;
  assign n4034 = ~n20167 | ~n20177;
  assign n20179 = ~n17563 & n20161;
  assign n20180 = P2_REIP_REG_1_ & n20163;
  assign n20181 = P2_PHYADDRPOINTER_REG_1_ & n20160;
  assign n20182 = ~n20179 & ~n20180;
  assign n20183 = ~n20181 & n20182;
  assign n20184 = ~n17542 & n20168;
  assign n20185 = ~P2_PHYADDRPOINTER_REG_1_ & n20171;
  assign n20186 = ~n15263 & n20174;
  assign n20187 = ~n20184 & ~n20185;
  assign n20188 = ~n20186 & n20187;
  assign n4039 = ~n20183 | ~n20188;
  assign n20190 = ~n17653 & n20161;
  assign n20191 = P2_REIP_REG_2_ & n20163;
  assign n20192 = P2_PHYADDRPOINTER_REG_2_ & n20160;
  assign n20193 = ~n20190 & ~n20191;
  assign n20194 = ~n20192 & n20193;
  assign n20195 = ~n17632 & n20168;
  assign n20196 = P2_PHYADDRPOINTER_REG_1_ & ~P2_PHYADDRPOINTER_REG_2_;
  assign n20197 = ~P2_PHYADDRPOINTER_REG_1_ & P2_PHYADDRPOINTER_REG_2_;
  assign n20198 = ~n20196 & ~n20197;
  assign n20199 = n20171 & ~n20198;
  assign n20200 = ~n15216 & n20174;
  assign n20201 = ~n20195 & ~n20199;
  assign n20202 = ~n20200 & n20201;
  assign n4044 = ~n20194 | ~n20202;
  assign n20204 = ~n17745 & n20161;
  assign n20205 = P2_REIP_REG_3_ & n20163;
  assign n20206 = P2_PHYADDRPOINTER_REG_3_ & n20160;
  assign n20207 = ~n20204 & ~n20205;
  assign n20208 = ~n20206 & n20207;
  assign n20209 = ~n17725 & n20168;
  assign n20210 = P2_PHYADDRPOINTER_REG_1_ & P2_PHYADDRPOINTER_REG_2_;
  assign n20211 = ~P2_PHYADDRPOINTER_REG_3_ & n20210;
  assign n20212 = P2_PHYADDRPOINTER_REG_3_ & ~n20210;
  assign n20213 = ~n20211 & ~n20212;
  assign n20214 = n20171 & ~n20213;
  assign n20215 = ~n15147 & n20174;
  assign n20216 = ~n20209 & ~n20214;
  assign n20217 = ~n20215 & n20216;
  assign n4049 = ~n20208 | ~n20217;
  assign n20219 = ~n17835 & n20161;
  assign n20220 = P2_REIP_REG_4_ & n20163;
  assign n20221 = P2_PHYADDRPOINTER_REG_4_ & n20160;
  assign n20222 = ~n20219 & ~n20220;
  assign n20223 = ~n20221 & n20222;
  assign n20224 = ~n17812 & n20168;
  assign n20225 = ~P2_PHYADDRPOINTER_REG_4_ & n15306;
  assign n20226 = P2_PHYADDRPOINTER_REG_4_ & ~n15306;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = n20171 & ~n20227;
  assign n20229 = n17863 & n20174;
  assign n20230 = ~n20224 & ~n20228;
  assign n20231 = ~n20229 & n20230;
  assign n4054 = ~n20223 | ~n20231;
  assign n20233 = ~n17954 & n20161;
  assign n20234 = P2_REIP_REG_5_ & n20163;
  assign n20235 = P2_PHYADDRPOINTER_REG_5_ & n20160;
  assign n20236 = ~n20233 & ~n20234;
  assign n20237 = ~n20235 & n20236;
  assign n20238 = ~n17934 & n20168;
  assign n20239 = ~P2_PHYADDRPOINTER_REG_5_ & n15307;
  assign n20240 = P2_PHYADDRPOINTER_REG_5_ & ~n15307;
  assign n20241 = ~n20239 & ~n20240;
  assign n20242 = n20171 & ~n20241;
  assign n20243 = ~n17979 & n20174;
  assign n20244 = ~n20238 & ~n20242;
  assign n20245 = ~n20243 & n20244;
  assign n4059 = ~n20237 | ~n20245;
  assign n20247 = ~n18073 & n20161;
  assign n20248 = P2_REIP_REG_6_ & n20163;
  assign n20249 = P2_PHYADDRPOINTER_REG_6_ & n20160;
  assign n20250 = ~n20247 & ~n20248;
  assign n20251 = ~n20249 & n20250;
  assign n20252 = ~n18050 & n20168;
  assign n20253 = ~P2_PHYADDRPOINTER_REG_6_ & n15308;
  assign n20254 = P2_PHYADDRPOINTER_REG_6_ & ~n15308;
  assign n20255 = ~n20253 & ~n20254;
  assign n20256 = n20171 & ~n20255;
  assign n20257 = ~n18099 & n20174;
  assign n20258 = ~n20252 & ~n20256;
  assign n20259 = ~n20257 & n20258;
  assign n4064 = ~n20251 | ~n20259;
  assign n20261 = ~n18199 & n20161;
  assign n20262 = P2_REIP_REG_7_ & n20163;
  assign n20263 = P2_PHYADDRPOINTER_REG_7_ & n20160;
  assign n20264 = ~n20261 & ~n20262;
  assign n20265 = ~n20263 & n20264;
  assign n20266 = ~n18170 & n20168;
  assign n20267 = ~P2_PHYADDRPOINTER_REG_7_ & n15309;
  assign n20268 = P2_PHYADDRPOINTER_REG_7_ & ~n15309;
  assign n20269 = ~n20267 & ~n20268;
  assign n20270 = n20171 & ~n20269;
  assign n20271 = ~n18225 & n20174;
  assign n20272 = ~n20266 & ~n20270;
  assign n20273 = ~n20271 & n20272;
  assign n4069 = ~n20265 | ~n20273;
  assign n20275 = ~n18285 & n20161;
  assign n20276 = P2_REIP_REG_8_ & n20163;
  assign n20277 = P2_PHYADDRPOINTER_REG_8_ & n20160;
  assign n20278 = ~n20275 & ~n20276;
  assign n20279 = ~n20277 & n20278;
  assign n20280 = ~n18260 & n20168;
  assign n20281 = ~P2_PHYADDRPOINTER_REG_8_ & n15310;
  assign n20282 = P2_PHYADDRPOINTER_REG_8_ & ~n15310;
  assign n20283 = ~n20281 & ~n20282;
  assign n20284 = n20171 & ~n20283;
  assign n20285 = ~n18311 & n20174;
  assign n20286 = ~n20280 & ~n20284;
  assign n20287 = ~n20285 & n20286;
  assign n4074 = ~n20279 | ~n20287;
  assign n20289 = ~n18416 & n20161;
  assign n20290 = P2_REIP_REG_9_ & n20163;
  assign n20291 = P2_PHYADDRPOINTER_REG_9_ & n20160;
  assign n20292 = ~n20289 & ~n20290;
  assign n20293 = ~n20291 & n20292;
  assign n20294 = n18398 & n20168;
  assign n20295 = ~P2_PHYADDRPOINTER_REG_9_ & n15311;
  assign n20296 = P2_PHYADDRPOINTER_REG_9_ & ~n15311;
  assign n20297 = ~n20295 & ~n20296;
  assign n20298 = n20171 & ~n20297;
  assign n20299 = ~n18442 & n20174;
  assign n20300 = ~n20294 & ~n20298;
  assign n20301 = ~n20299 & n20300;
  assign n4079 = ~n20293 | ~n20301;
  assign n20303 = ~n18515 & n20161;
  assign n20304 = P2_REIP_REG_10_ & n20163;
  assign n20305 = P2_PHYADDRPOINTER_REG_10_ & n20160;
  assign n20306 = ~n20303 & ~n20304;
  assign n20307 = ~n20305 & n20306;
  assign n20308 = n18495 & n20168;
  assign n20309 = ~P2_PHYADDRPOINTER_REG_10_ & n15312;
  assign n20310 = P2_PHYADDRPOINTER_REG_10_ & ~n15312;
  assign n20311 = ~n20309 & ~n20310;
  assign n20312 = n20171 & ~n20311;
  assign n20313 = ~n18541 & n20174;
  assign n20314 = ~n20308 & ~n20312;
  assign n20315 = ~n20313 & n20314;
  assign n4084 = ~n20307 | ~n20315;
  assign n20317 = ~n18612 & n20161;
  assign n20318 = P2_REIP_REG_11_ & n20163;
  assign n20319 = P2_PHYADDRPOINTER_REG_11_ & n20160;
  assign n20320 = ~n20317 & ~n20318;
  assign n20321 = ~n20319 & n20320;
  assign n20322 = n18594 & n20168;
  assign n20323 = ~P2_PHYADDRPOINTER_REG_11_ & n15313;
  assign n20324 = P2_PHYADDRPOINTER_REG_11_ & ~n15313;
  assign n20325 = ~n20323 & ~n20324;
  assign n20326 = n20171 & ~n20325;
  assign n20327 = ~n18638 & n20174;
  assign n20328 = ~n20322 & ~n20326;
  assign n20329 = ~n20327 & n20328;
  assign n4089 = ~n20321 | ~n20329;
  assign n20331 = ~n18710 & n20161;
  assign n20332 = P2_REIP_REG_12_ & n20163;
  assign n20333 = P2_PHYADDRPOINTER_REG_12_ & n20160;
  assign n20334 = ~n20331 & ~n20332;
  assign n20335 = ~n20333 & n20334;
  assign n20336 = ~n18690 & n20168;
  assign n20337 = ~P2_PHYADDRPOINTER_REG_12_ & n15314;
  assign n20338 = P2_PHYADDRPOINTER_REG_12_ & ~n15314;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = n20171 & ~n20339;
  assign n20341 = ~n18736 & n20174;
  assign n20342 = ~n20336 & ~n20340;
  assign n20343 = ~n20341 & n20342;
  assign n4094 = ~n20335 | ~n20343;
  assign n20345 = ~n18811 & n20161;
  assign n20346 = P2_REIP_REG_13_ & n20163;
  assign n20347 = P2_PHYADDRPOINTER_REG_13_ & n20160;
  assign n20348 = ~n20345 & ~n20346;
  assign n20349 = ~n20347 & n20348;
  assign n20350 = n18793 & n20168;
  assign n20351 = ~P2_PHYADDRPOINTER_REG_13_ & n15315;
  assign n20352 = P2_PHYADDRPOINTER_REG_13_ & ~n15315;
  assign n20353 = ~n20351 & ~n20352;
  assign n20354 = n20171 & ~n20353;
  assign n20355 = ~n18837 & n20174;
  assign n20356 = ~n20350 & ~n20354;
  assign n20357 = ~n20355 & n20356;
  assign n4099 = ~n20349 | ~n20357;
  assign n20359 = ~n18910 & n20161;
  assign n20360 = P2_REIP_REG_14_ & n20163;
  assign n20361 = P2_PHYADDRPOINTER_REG_14_ & n20160;
  assign n20362 = ~n20359 & ~n20360;
  assign n20363 = ~n20361 & n20362;
  assign n20364 = n18890 & n20168;
  assign n20365 = ~P2_PHYADDRPOINTER_REG_14_ & n15316;
  assign n20366 = P2_PHYADDRPOINTER_REG_14_ & ~n15316;
  assign n20367 = ~n20365 & ~n20366;
  assign n20368 = n20171 & ~n20367;
  assign n20369 = ~n18936 & n20174;
  assign n20370 = ~n20364 & ~n20368;
  assign n20371 = ~n20369 & n20370;
  assign n4104 = ~n20363 | ~n20371;
  assign n20373 = ~n19006 & n20161;
  assign n20374 = P2_REIP_REG_15_ & n20163;
  assign n20375 = P2_PHYADDRPOINTER_REG_15_ & n20160;
  assign n20376 = ~n20373 & ~n20374;
  assign n20377 = ~n20375 & n20376;
  assign n20378 = ~n18988 & n20168;
  assign n20379 = ~P2_PHYADDRPOINTER_REG_15_ & n15317;
  assign n20380 = P2_PHYADDRPOINTER_REG_15_ & ~n15317;
  assign n20381 = ~n20379 & ~n20380;
  assign n20382 = n20171 & ~n20381;
  assign n20383 = ~n19032 & n20174;
  assign n20384 = ~n20378 & ~n20382;
  assign n20385 = ~n20383 & n20384;
  assign n4109 = ~n20377 | ~n20385;
  assign n20387 = ~n19109 & n20161;
  assign n20388 = P2_REIP_REG_16_ & n20163;
  assign n20389 = P2_PHYADDRPOINTER_REG_16_ & n20160;
  assign n20390 = ~n20387 & ~n20388;
  assign n20391 = ~n20389 & n20390;
  assign n20392 = n19089 & n20168;
  assign n20393 = ~P2_PHYADDRPOINTER_REG_16_ & n15318;
  assign n20394 = P2_PHYADDRPOINTER_REG_16_ & ~n15318;
  assign n20395 = ~n20393 & ~n20394;
  assign n20396 = n20171 & ~n20395;
  assign n20397 = ~n19135 & n20174;
  assign n20398 = ~n20392 & ~n20396;
  assign n20399 = ~n20397 & n20398;
  assign n4114 = ~n20391 | ~n20399;
  assign n20401 = ~n19172 & n20161;
  assign n20402 = P2_REIP_REG_17_ & n20163;
  assign n20403 = P2_PHYADDRPOINTER_REG_17_ & n20160;
  assign n20404 = ~n20401 & ~n20402;
  assign n20405 = ~n20403 & n20404;
  assign n20406 = ~n19154 & n20168;
  assign n20407 = ~P2_PHYADDRPOINTER_REG_17_ & n15319;
  assign n20408 = P2_PHYADDRPOINTER_REG_17_ & ~n15319;
  assign n20409 = ~n20407 & ~n20408;
  assign n20410 = n20171 & ~n20409;
  assign n20411 = ~n19198 & n20174;
  assign n20412 = ~n20406 & ~n20410;
  assign n20413 = ~n20411 & n20412;
  assign n4119 = ~n20405 | ~n20413;
  assign n20415 = ~n19240 & n20161;
  assign n20416 = P2_REIP_REG_18_ & n20163;
  assign n20417 = P2_PHYADDRPOINTER_REG_18_ & n20160;
  assign n20418 = ~n20415 & ~n20416;
  assign n20419 = ~n20417 & n20418;
  assign n20420 = ~n19220 & n20168;
  assign n20421 = ~P2_PHYADDRPOINTER_REG_18_ & n15320;
  assign n20422 = P2_PHYADDRPOINTER_REG_18_ & ~n15320;
  assign n20423 = ~n20421 & ~n20422;
  assign n20424 = n20171 & ~n20423;
  assign n20425 = ~n19266 & n20174;
  assign n20426 = ~n20420 & ~n20424;
  assign n20427 = ~n20425 & n20426;
  assign n4124 = ~n20419 | ~n20427;
  assign n20429 = ~n19308 & n20161;
  assign n20430 = P2_REIP_REG_19_ & n20163;
  assign n20431 = P2_PHYADDRPOINTER_REG_19_ & n20160;
  assign n20432 = ~n20429 & ~n20430;
  assign n20433 = ~n20431 & n20432;
  assign n20434 = n19290 & n20168;
  assign n20435 = ~P2_PHYADDRPOINTER_REG_19_ & n15321;
  assign n20436 = P2_PHYADDRPOINTER_REG_19_ & ~n15321;
  assign n20437 = ~n20435 & ~n20436;
  assign n20438 = n20171 & ~n20437;
  assign n20439 = ~n19334 & n20174;
  assign n20440 = ~n20434 & ~n20438;
  assign n20441 = ~n20439 & n20440;
  assign n4129 = ~n20433 | ~n20441;
  assign n20443 = ~n19375 & n20161;
  assign n20444 = P2_REIP_REG_20_ & n20163;
  assign n20445 = P2_PHYADDRPOINTER_REG_20_ & n20160;
  assign n20446 = ~n20443 & ~n20444;
  assign n20447 = ~n20445 & n20446;
  assign n20448 = n19355 & n20168;
  assign n20449 = ~P2_PHYADDRPOINTER_REG_20_ & n15322;
  assign n20450 = P2_PHYADDRPOINTER_REG_20_ & ~n15322;
  assign n20451 = ~n20449 & ~n20450;
  assign n20452 = n20171 & ~n20451;
  assign n20453 = ~n19401 & n20174;
  assign n20454 = ~n20448 & ~n20452;
  assign n20455 = ~n20453 & n20454;
  assign n4134 = ~n20447 | ~n20455;
  assign n20457 = ~n19441 & n20161;
  assign n20458 = P2_REIP_REG_21_ & n20163;
  assign n20459 = P2_PHYADDRPOINTER_REG_21_ & n20160;
  assign n20460 = ~n20457 & ~n20458;
  assign n20461 = ~n20459 & n20460;
  assign n20462 = ~n19420 & n20168;
  assign n20463 = ~P2_PHYADDRPOINTER_REG_21_ & n15323;
  assign n20464 = P2_PHYADDRPOINTER_REG_21_ & ~n15323;
  assign n20465 = ~n20463 & ~n20464;
  assign n20466 = n20171 & ~n20465;
  assign n20467 = ~n19467 & n20174;
  assign n20468 = ~n20462 & ~n20466;
  assign n20469 = ~n20467 & n20468;
  assign n4139 = ~n20461 | ~n20469;
  assign n20471 = ~n19507 & n20161;
  assign n20472 = P2_REIP_REG_22_ & n20163;
  assign n20473 = P2_PHYADDRPOINTER_REG_22_ & n20160;
  assign n20474 = ~n20471 & ~n20472;
  assign n20475 = ~n20473 & n20474;
  assign n20476 = n19490 & n20168;
  assign n20477 = ~P2_PHYADDRPOINTER_REG_22_ & n15324;
  assign n20478 = P2_PHYADDRPOINTER_REG_22_ & ~n15324;
  assign n20479 = ~n20477 & ~n20478;
  assign n20480 = n20171 & ~n20479;
  assign n20481 = ~n19533 & n20174;
  assign n20482 = ~n20476 & ~n20480;
  assign n20483 = ~n20481 & n20482;
  assign n4144 = ~n20475 | ~n20483;
  assign n20485 = ~n19576 & n20161;
  assign n20486 = P2_REIP_REG_23_ & n20163;
  assign n20487 = P2_PHYADDRPOINTER_REG_23_ & n20160;
  assign n20488 = ~n20485 & ~n20486;
  assign n20489 = ~n20487 & n20488;
  assign n20490 = n19555 & n20168;
  assign n20491 = ~P2_PHYADDRPOINTER_REG_23_ & n15325;
  assign n20492 = P2_PHYADDRPOINTER_REG_23_ & ~n15325;
  assign n20493 = ~n20491 & ~n20492;
  assign n20494 = n20171 & ~n20493;
  assign n20495 = ~n19602 & n20174;
  assign n20496 = ~n20490 & ~n20494;
  assign n20497 = ~n20495 & n20496;
  assign n4149 = ~n20489 | ~n20497;
  assign n20499 = ~n19638 & n20161;
  assign n20500 = P2_REIP_REG_24_ & n20163;
  assign n20501 = P2_PHYADDRPOINTER_REG_24_ & n20160;
  assign n20502 = ~n20499 & ~n20500;
  assign n20503 = ~n20501 & n20502;
  assign n20504 = ~n19621 & n20168;
  assign n20505 = ~P2_PHYADDRPOINTER_REG_24_ & n15326;
  assign n20506 = P2_PHYADDRPOINTER_REG_24_ & ~n15326;
  assign n20507 = ~n20505 & ~n20506;
  assign n20508 = n20171 & ~n20507;
  assign n20509 = ~n19664 & n20174;
  assign n20510 = ~n20504 & ~n20508;
  assign n20511 = ~n20509 & n20510;
  assign n4154 = ~n20503 | ~n20511;
  assign n20513 = ~n19706 & n20161;
  assign n20514 = P2_REIP_REG_25_ & n20163;
  assign n20515 = P2_PHYADDRPOINTER_REG_25_ & n20160;
  assign n20516 = ~n20513 & ~n20514;
  assign n20517 = ~n20515 & n20516;
  assign n20518 = ~n19685 & n20168;
  assign n20519 = ~P2_PHYADDRPOINTER_REG_25_ & n15327;
  assign n20520 = P2_PHYADDRPOINTER_REG_25_ & ~n15327;
  assign n20521 = ~n20519 & ~n20520;
  assign n20522 = n20171 & ~n20521;
  assign n20523 = ~n19732 & n20174;
  assign n20524 = ~n20518 & ~n20522;
  assign n20525 = ~n20523 & n20524;
  assign n4159 = ~n20517 | ~n20525;
  assign n20527 = ~n19774 & n20161;
  assign n20528 = P2_REIP_REG_26_ & n20163;
  assign n20529 = P2_PHYADDRPOINTER_REG_26_ & n20160;
  assign n20530 = ~n20527 & ~n20528;
  assign n20531 = ~n20529 & n20530;
  assign n20532 = n19757 & n20168;
  assign n20533 = ~P2_PHYADDRPOINTER_REG_26_ & n15328;
  assign n20534 = P2_PHYADDRPOINTER_REG_26_ & ~n15328;
  assign n20535 = ~n20533 & ~n20534;
  assign n20536 = n20171 & ~n20535;
  assign n20537 = ~n19800 & n20174;
  assign n20538 = ~n20532 & ~n20536;
  assign n20539 = ~n20537 & n20538;
  assign n4164 = ~n20531 | ~n20539;
  assign n20541 = ~n19837 & n20161;
  assign n20542 = P2_REIP_REG_27_ & n20163;
  assign n20543 = P2_PHYADDRPOINTER_REG_27_ & n20160;
  assign n20544 = ~n20541 & ~n20542;
  assign n20545 = ~n20543 & n20544;
  assign n20546 = ~n19819 & n20168;
  assign n20547 = ~P2_PHYADDRPOINTER_REG_27_ & n15329;
  assign n20548 = P2_PHYADDRPOINTER_REG_27_ & ~n15329;
  assign n20549 = ~n20547 & ~n20548;
  assign n20550 = n20171 & ~n20549;
  assign n20551 = ~n19863 & n20174;
  assign n20552 = ~n20546 & ~n20550;
  assign n20553 = ~n20551 & n20552;
  assign n4169 = ~n20545 | ~n20553;
  assign n20555 = ~n19906 & n20161;
  assign n20556 = P2_REIP_REG_28_ & n20163;
  assign n20557 = P2_PHYADDRPOINTER_REG_28_ & n20160;
  assign n20558 = ~n20555 & ~n20556;
  assign n20559 = ~n20557 & n20558;
  assign n20560 = n19886 & n20168;
  assign n20561 = ~P2_PHYADDRPOINTER_REG_28_ & n15330;
  assign n20562 = P2_PHYADDRPOINTER_REG_28_ & ~n15330;
  assign n20563 = ~n20561 & ~n20562;
  assign n20564 = n20171 & ~n20563;
  assign n20565 = ~n19932 & n20174;
  assign n20566 = ~n20560 & ~n20564;
  assign n20567 = ~n20565 & n20566;
  assign n4174 = ~n20559 | ~n20567;
  assign n20569 = ~n19976 & n20161;
  assign n20570 = P2_REIP_REG_29_ & n20163;
  assign n20571 = P2_PHYADDRPOINTER_REG_29_ & n20160;
  assign n20572 = ~n20569 & ~n20570;
  assign n20573 = ~n20571 & n20572;
  assign n20574 = n19954 & n20168;
  assign n20575 = ~P2_PHYADDRPOINTER_REG_29_ & n15331;
  assign n20576 = P2_PHYADDRPOINTER_REG_29_ & ~n15331;
  assign n20577 = ~n20575 & ~n20576;
  assign n20578 = n20171 & ~n20577;
  assign n20579 = ~n20001 & n20174;
  assign n20580 = ~n20574 & ~n20578;
  assign n20581 = ~n20579 & n20580;
  assign n4179 = ~n20573 | ~n20581;
  assign n20583 = P2_PHYADDRPOINTER_REG_30_ & n20160;
  assign n20584 = P2_REIP_REG_30_ & n20163;
  assign n20585 = ~n20038 & n20161;
  assign n20586 = ~n20583 & ~n20584;
  assign n20587 = ~n20585 & n20586;
  assign n20588 = ~n20021 & n20168;
  assign n20589 = ~P2_PHYADDRPOINTER_REG_30_ & n15332;
  assign n20590 = P2_PHYADDRPOINTER_REG_30_ & ~n15332;
  assign n20591 = ~n20589 & ~n20590;
  assign n20592 = n20171 & ~n20591;
  assign n20593 = ~n20063 & n20174;
  assign n20594 = ~n20588 & ~n20592;
  assign n20595 = ~n20593 & n20594;
  assign n4184 = ~n20587 | ~n20595;
  assign n20597 = n20113 & n20161;
  assign n20598 = P2_REIP_REG_31_ & n20163;
  assign n20599 = P2_PHYADDRPOINTER_REG_31_ & n20160;
  assign n20600 = ~n20597 & ~n20598;
  assign n20601 = ~n20599 & n20600;
  assign n20602 = ~n20085 & n20168;
  assign n20603 = ~n15336 & n20171;
  assign n20604 = ~n20138 & n20174;
  assign n20605 = ~n20602 & ~n20603;
  assign n20606 = ~n20604 & n20605;
  assign n4189 = ~n20601 | ~n20606;
  assign n20608 = BUF1_REG_15_ & n4541;
  assign n20609 = BUF2_REG_15_ & ~n4541;
  assign n20610 = ~n20608 & ~n20609;
  assign n20611 = n14051 & ~n14238;
  assign n20612 = n15428 & ~n20611;
  assign n20613 = n14550 & n20612;
  assign n20614 = n15183 & n20613;
  assign n20615 = ~n14238 & n20614;
  assign n20616 = ~n20610 & n20615;
  assign n20617 = n14238 & n20614;
  assign n20618 = P2_EAX_REG_15_ & n20617;
  assign n20619 = P2_LWORD_REG_15_ & ~n20614;
  assign n20620 = ~n20616 & ~n20618;
  assign n4194 = n20619 | ~n20620;
  assign n20622 = BUF1_REG_14_ & n4541;
  assign n20623 = BUF2_REG_14_ & ~n4541;
  assign n20624 = ~n20622 & ~n20623;
  assign n20625 = n20615 & ~n20624;
  assign n20626 = P2_EAX_REG_14_ & n20617;
  assign n20627 = P2_LWORD_REG_14_ & ~n20614;
  assign n20628 = ~n20625 & ~n20626;
  assign n4199 = n20627 | ~n20628;
  assign n20630 = BUF1_REG_13_ & n4541;
  assign n20631 = BUF2_REG_13_ & ~n4541;
  assign n20632 = ~n20630 & ~n20631;
  assign n20633 = n20615 & ~n20632;
  assign n20634 = P2_EAX_REG_13_ & n20617;
  assign n20635 = P2_LWORD_REG_13_ & ~n20614;
  assign n20636 = ~n20633 & ~n20634;
  assign n4204 = n20635 | ~n20636;
  assign n20638 = BUF1_REG_12_ & n4541;
  assign n20639 = BUF2_REG_12_ & ~n4541;
  assign n20640 = ~n20638 & ~n20639;
  assign n20641 = n20615 & ~n20640;
  assign n20642 = P2_EAX_REG_12_ & n20617;
  assign n20643 = P2_LWORD_REG_12_ & ~n20614;
  assign n20644 = ~n20641 & ~n20642;
  assign n4209 = n20643 | ~n20644;
  assign n20646 = BUF1_REG_11_ & n4541;
  assign n20647 = BUF2_REG_11_ & ~n4541;
  assign n20648 = ~n20646 & ~n20647;
  assign n20649 = n20615 & ~n20648;
  assign n20650 = P2_EAX_REG_11_ & n20617;
  assign n20651 = P2_LWORD_REG_11_ & ~n20614;
  assign n20652 = ~n20649 & ~n20650;
  assign n4214 = n20651 | ~n20652;
  assign n20654 = BUF1_REG_10_ & n4541;
  assign n20655 = BUF2_REG_10_ & ~n4541;
  assign n20656 = ~n20654 & ~n20655;
  assign n20657 = n20615 & ~n20656;
  assign n20658 = P2_EAX_REG_10_ & n20617;
  assign n20659 = P2_LWORD_REG_10_ & ~n20614;
  assign n20660 = ~n20657 & ~n20658;
  assign n4219 = n20659 | ~n20660;
  assign n20662 = BUF1_REG_9_ & n4541;
  assign n20663 = BUF2_REG_9_ & ~n4541;
  assign n20664 = ~n20662 & ~n20663;
  assign n20665 = n20615 & ~n20664;
  assign n20666 = P2_EAX_REG_9_ & n20617;
  assign n20667 = P2_LWORD_REG_9_ & ~n20614;
  assign n20668 = ~n20665 & ~n20666;
  assign n4224 = n20667 | ~n20668;
  assign n20670 = BUF1_REG_8_ & n4541;
  assign n20671 = BUF2_REG_8_ & ~n4541;
  assign n20672 = ~n20670 & ~n20671;
  assign n20673 = n20615 & ~n20672;
  assign n20674 = P2_EAX_REG_8_ & n20617;
  assign n20675 = P2_LWORD_REG_8_ & ~n20614;
  assign n20676 = ~n20673 & ~n20674;
  assign n4229 = n20675 | ~n20676;
  assign n20678 = ~n15590 & n20615;
  assign n20679 = P2_EAX_REG_7_ & n20617;
  assign n20680 = P2_LWORD_REG_7_ & ~n20614;
  assign n20681 = ~n20678 & ~n20679;
  assign n4234 = n20680 | ~n20681;
  assign n20683 = ~n15618 & n20615;
  assign n20684 = P2_EAX_REG_6_ & n20617;
  assign n20685 = P2_LWORD_REG_6_ & ~n20614;
  assign n20686 = ~n20683 & ~n20684;
  assign n4239 = n20685 | ~n20686;
  assign n20688 = ~n15640 & n20615;
  assign n20689 = P2_EAX_REG_5_ & n20617;
  assign n20690 = P2_LWORD_REG_5_ & ~n20614;
  assign n20691 = ~n20688 & ~n20689;
  assign n4244 = n20690 | ~n20691;
  assign n20693 = ~n15662 & n20615;
  assign n20694 = P2_EAX_REG_4_ & n20617;
  assign n20695 = P2_LWORD_REG_4_ & ~n20614;
  assign n20696 = ~n20693 & ~n20694;
  assign n4249 = n20695 | ~n20696;
  assign n20698 = ~n15684 & n20615;
  assign n20699 = P2_EAX_REG_3_ & n20617;
  assign n20700 = P2_LWORD_REG_3_ & ~n20614;
  assign n20701 = ~n20698 & ~n20699;
  assign n4254 = n20700 | ~n20701;
  assign n20703 = ~n15706 & n20615;
  assign n20704 = P2_EAX_REG_2_ & n20617;
  assign n20705 = P2_LWORD_REG_2_ & ~n20614;
  assign n20706 = ~n20703 & ~n20704;
  assign n4259 = n20705 | ~n20706;
  assign n20708 = ~n15728 & n20615;
  assign n20709 = P2_EAX_REG_1_ & n20617;
  assign n20710 = P2_LWORD_REG_1_ & ~n20614;
  assign n20711 = ~n20708 & ~n20709;
  assign n4264 = n20710 | ~n20711;
  assign n20713 = ~n15750 & n20615;
  assign n20714 = P2_EAX_REG_0_ & n20617;
  assign n20715 = P2_LWORD_REG_0_ & ~n20614;
  assign n20716 = ~n20713 & ~n20714;
  assign n4269 = n20715 | ~n20716;
  assign n20718 = P2_EAX_REG_30_ & n20617;
  assign n20719 = P2_UWORD_REG_14_ & ~n20614;
  assign n20720 = ~n20625 & ~n20718;
  assign n4274 = n20719 | ~n20720;
  assign n20722 = P2_EAX_REG_29_ & n20617;
  assign n20723 = P2_UWORD_REG_13_ & ~n20614;
  assign n20724 = ~n20633 & ~n20722;
  assign n4279 = n20723 | ~n20724;
  assign n20726 = P2_EAX_REG_28_ & n20617;
  assign n20727 = P2_UWORD_REG_12_ & ~n20614;
  assign n20728 = ~n20641 & ~n20726;
  assign n4284 = n20727 | ~n20728;
  assign n20730 = P2_EAX_REG_27_ & n20617;
  assign n20731 = P2_UWORD_REG_11_ & ~n20614;
  assign n20732 = ~n20649 & ~n20730;
  assign n4289 = n20731 | ~n20732;
  assign n20734 = P2_EAX_REG_26_ & n20617;
  assign n20735 = P2_UWORD_REG_10_ & ~n20614;
  assign n20736 = ~n20657 & ~n20734;
  assign n4294 = n20735 | ~n20736;
  assign n20738 = P2_EAX_REG_25_ & n20617;
  assign n20739 = P2_UWORD_REG_9_ & ~n20614;
  assign n20740 = ~n20665 & ~n20738;
  assign n4299 = n20739 | ~n20740;
  assign n20742 = P2_EAX_REG_24_ & n20617;
  assign n20743 = P2_UWORD_REG_8_ & ~n20614;
  assign n20744 = ~n20673 & ~n20742;
  assign n4304 = n20743 | ~n20744;
  assign n20746 = P2_EAX_REG_23_ & n20617;
  assign n20747 = P2_UWORD_REG_7_ & ~n20614;
  assign n20748 = ~n20678 & ~n20746;
  assign n4309 = n20747 | ~n20748;
  assign n20750 = P2_EAX_REG_22_ & n20617;
  assign n20751 = P2_UWORD_REG_6_ & ~n20614;
  assign n20752 = ~n20683 & ~n20750;
  assign n4314 = n20751 | ~n20752;
  assign n20754 = P2_EAX_REG_21_ & n20617;
  assign n20755 = P2_UWORD_REG_5_ & ~n20614;
  assign n20756 = ~n20688 & ~n20754;
  assign n4319 = n20755 | ~n20756;
  assign n20758 = P2_EAX_REG_20_ & n20617;
  assign n20759 = P2_UWORD_REG_4_ & ~n20614;
  assign n20760 = ~n20693 & ~n20758;
  assign n4324 = n20759 | ~n20760;
  assign n20762 = P2_EAX_REG_19_ & n20617;
  assign n20763 = P2_UWORD_REG_3_ & ~n20614;
  assign n20764 = ~n20698 & ~n20762;
  assign n4329 = n20763 | ~n20764;
  assign n20766 = P2_EAX_REG_18_ & n20617;
  assign n20767 = P2_UWORD_REG_2_ & ~n20614;
  assign n20768 = ~n20703 & ~n20766;
  assign n4334 = n20767 | ~n20768;
  assign n20770 = P2_EAX_REG_17_ & n20617;
  assign n20771 = P2_UWORD_REG_1_ & ~n20614;
  assign n20772 = ~n20708 & ~n20770;
  assign n4339 = n20771 | ~n20772;
  assign n20774 = P2_EAX_REG_16_ & n20617;
  assign n20775 = P2_UWORD_REG_0_ & ~n20614;
  assign n20776 = ~n20713 & ~n20774;
  assign n4344 = n20775 | ~n20776;
  assign n20778 = P2_STATE2_REG_1_ & n15495;
  assign n20779 = n14239 & n15432;
  assign n20780 = n15183 & n20779;
  assign n20781 = ~n14238 & n15428;
  assign n20782 = n15013 & n20781;
  assign n20783 = ~n14949 & n20782;
  assign n20784 = ~n20780 & ~n20783;
  assign n20785 = n14144 & ~n20784;
  assign n20786 = ~n20778 & ~n20785;
  assign n20787 = ~P2_STATE2_REG_0_ & ~n20786;
  assign n20788 = P2_LWORD_REG_0_ & n20787;
  assign n20789 = P2_STATE2_REG_0_ & ~n20786;
  assign n20790 = P2_EAX_REG_0_ & n20789;
  assign n20791 = P2_DATAO_REG_0_ & n20786;
  assign n20792 = ~n20788 & ~n20790;
  assign n4349 = n20791 | ~n20792;
  assign n20794 = P2_LWORD_REG_1_ & n20787;
  assign n20795 = P2_EAX_REG_1_ & n20789;
  assign n20796 = P2_DATAO_REG_1_ & n20786;
  assign n20797 = ~n20794 & ~n20795;
  assign n4354 = n20796 | ~n20797;
  assign n20799 = P2_LWORD_REG_2_ & n20787;
  assign n20800 = P2_EAX_REG_2_ & n20789;
  assign n20801 = P2_DATAO_REG_2_ & n20786;
  assign n20802 = ~n20799 & ~n20800;
  assign n4359 = n20801 | ~n20802;
  assign n20804 = P2_LWORD_REG_3_ & n20787;
  assign n20805 = P2_EAX_REG_3_ & n20789;
  assign n20806 = P2_DATAO_REG_3_ & n20786;
  assign n20807 = ~n20804 & ~n20805;
  assign n4364 = n20806 | ~n20807;
  assign n20809 = P2_LWORD_REG_4_ & n20787;
  assign n20810 = P2_EAX_REG_4_ & n20789;
  assign n20811 = P2_DATAO_REG_4_ & n20786;
  assign n20812 = ~n20809 & ~n20810;
  assign n4369 = n20811 | ~n20812;
  assign n20814 = P2_LWORD_REG_5_ & n20787;
  assign n20815 = P2_EAX_REG_5_ & n20789;
  assign n20816 = P2_DATAO_REG_5_ & n20786;
  assign n20817 = ~n20814 & ~n20815;
  assign n4374 = n20816 | ~n20817;
  assign n20819 = P2_LWORD_REG_6_ & n20787;
  assign n20820 = P2_EAX_REG_6_ & n20789;
  assign n20821 = P2_DATAO_REG_6_ & n20786;
  assign n20822 = ~n20819 & ~n20820;
  assign n4379 = n20821 | ~n20822;
  assign n20824 = P2_LWORD_REG_7_ & n20787;
  assign n20825 = P2_EAX_REG_7_ & n20789;
  assign n20826 = P2_DATAO_REG_7_ & n20786;
  assign n20827 = ~n20824 & ~n20825;
  assign n4384 = n20826 | ~n20827;
  assign n20829 = P2_LWORD_REG_8_ & n20787;
  assign n20830 = P2_EAX_REG_8_ & n20789;
  assign n20831 = P2_DATAO_REG_8_ & n20786;
  assign n20832 = ~n20829 & ~n20830;
  assign n4389 = n20831 | ~n20832;
  assign n20834 = P2_LWORD_REG_9_ & n20787;
  assign n20835 = P2_EAX_REG_9_ & n20789;
  assign n20836 = P2_DATAO_REG_9_ & n20786;
  assign n20837 = ~n20834 & ~n20835;
  assign n4394 = n20836 | ~n20837;
  assign n20839 = P2_LWORD_REG_10_ & n20787;
  assign n20840 = P2_EAX_REG_10_ & n20789;
  assign n20841 = P2_DATAO_REG_10_ & n20786;
  assign n20842 = ~n20839 & ~n20840;
  assign n4399 = n20841 | ~n20842;
  assign n20844 = P2_LWORD_REG_11_ & n20787;
  assign n20845 = P2_EAX_REG_11_ & n20789;
  assign n20846 = P2_DATAO_REG_11_ & n20786;
  assign n20847 = ~n20844 & ~n20845;
  assign n4404 = n20846 | ~n20847;
  assign n20849 = P2_LWORD_REG_12_ & n20787;
  assign n20850 = P2_EAX_REG_12_ & n20789;
  assign n20851 = P2_DATAO_REG_12_ & n20786;
  assign n20852 = ~n20849 & ~n20850;
  assign n4409 = n20851 | ~n20852;
  assign n20854 = P2_LWORD_REG_13_ & n20787;
  assign n20855 = P2_EAX_REG_13_ & n20789;
  assign n20856 = P2_DATAO_REG_13_ & n20786;
  assign n20857 = ~n20854 & ~n20855;
  assign n4414 = n20856 | ~n20857;
  assign n20859 = P2_LWORD_REG_14_ & n20787;
  assign n20860 = P2_EAX_REG_14_ & n20789;
  assign n20861 = P2_DATAO_REG_14_ & n20786;
  assign n20862 = ~n20859 & ~n20860;
  assign n4419 = n20861 | ~n20862;
  assign n20864 = P2_LWORD_REG_15_ & n20787;
  assign n20865 = P2_EAX_REG_15_ & n20789;
  assign n20866 = P2_DATAO_REG_15_ & n20786;
  assign n20867 = ~n20864 & ~n20865;
  assign n4424 = n20866 | ~n20867;
  assign n20869 = P2_UWORD_REG_0_ & n20787;
  assign n20870 = n14550 & ~n20786;
  assign n20871 = P2_EAX_REG_16_ & n20870;
  assign n20872 = P2_DATAO_REG_16_ & n20786;
  assign n20873 = ~n20869 & ~n20871;
  assign n4429 = n20872 | ~n20873;
  assign n20875 = P2_UWORD_REG_1_ & n20787;
  assign n20876 = P2_EAX_REG_17_ & n20870;
  assign n20877 = P2_DATAO_REG_17_ & n20786;
  assign n20878 = ~n20875 & ~n20876;
  assign n4434 = n20877 | ~n20878;
  assign n20880 = P2_UWORD_REG_2_ & n20787;
  assign n20881 = P2_EAX_REG_18_ & n20870;
  assign n20882 = P2_DATAO_REG_18_ & n20786;
  assign n20883 = ~n20880 & ~n20881;
  assign n4439 = n20882 | ~n20883;
  assign n20885 = P2_UWORD_REG_3_ & n20787;
  assign n20886 = P2_EAX_REG_19_ & n20870;
  assign n20887 = P2_DATAO_REG_19_ & n20786;
  assign n20888 = ~n20885 & ~n20886;
  assign n4444 = n20887 | ~n20888;
  assign n20890 = P2_UWORD_REG_4_ & n20787;
  assign n20891 = P2_EAX_REG_20_ & n20870;
  assign n20892 = P2_DATAO_REG_20_ & n20786;
  assign n20893 = ~n20890 & ~n20891;
  assign n4449 = n20892 | ~n20893;
  assign n20895 = P2_UWORD_REG_5_ & n20787;
  assign n20896 = P2_EAX_REG_21_ & n20870;
  assign n20897 = P2_DATAO_REG_21_ & n20786;
  assign n20898 = ~n20895 & ~n20896;
  assign n4454 = n20897 | ~n20898;
  assign n20900 = P2_UWORD_REG_6_ & n20787;
  assign n20901 = P2_EAX_REG_22_ & n20870;
  assign n20902 = P2_DATAO_REG_22_ & n20786;
  assign n20903 = ~n20900 & ~n20901;
  assign n4459 = n20902 | ~n20903;
  assign n20905 = P2_UWORD_REG_7_ & n20787;
  assign n20906 = P2_EAX_REG_23_ & n20870;
  assign n20907 = P2_DATAO_REG_23_ & n20786;
  assign n20908 = ~n20905 & ~n20906;
  assign n4464 = n20907 | ~n20908;
  assign n20910 = P2_UWORD_REG_8_ & n20787;
  assign n20911 = P2_EAX_REG_24_ & n20870;
  assign n20912 = P2_DATAO_REG_24_ & n20786;
  assign n20913 = ~n20910 & ~n20911;
  assign n4469 = n20912 | ~n20913;
  assign n20915 = P2_UWORD_REG_9_ & n20787;
  assign n20916 = P2_EAX_REG_25_ & n20870;
  assign n20917 = P2_DATAO_REG_25_ & n20786;
  assign n20918 = ~n20915 & ~n20916;
  assign n4474 = n20917 | ~n20918;
  assign n20920 = P2_UWORD_REG_10_ & n20787;
  assign n20921 = P2_EAX_REG_26_ & n20870;
  assign n20922 = P2_DATAO_REG_26_ & n20786;
  assign n20923 = ~n20920 & ~n20921;
  assign n4479 = n20922 | ~n20923;
  assign n20925 = P2_UWORD_REG_11_ & n20787;
  assign n20926 = P2_EAX_REG_27_ & n20870;
  assign n20927 = P2_DATAO_REG_27_ & n20786;
  assign n20928 = ~n20925 & ~n20926;
  assign n4484 = n20927 | ~n20928;
  assign n20930 = P2_UWORD_REG_12_ & n20787;
  assign n20931 = P2_EAX_REG_28_ & n20870;
  assign n20932 = P2_DATAO_REG_28_ & n20786;
  assign n20933 = ~n20930 & ~n20931;
  assign n4489 = n20932 | ~n20933;
  assign n20935 = P2_UWORD_REG_13_ & n20787;
  assign n20936 = P2_EAX_REG_29_ & n20870;
  assign n20937 = P2_DATAO_REG_29_ & n20786;
  assign n20938 = ~n20935 & ~n20936;
  assign n4494 = n20937 | ~n20938;
  assign n20940 = P2_UWORD_REG_14_ & n20787;
  assign n20941 = P2_EAX_REG_30_ & n20870;
  assign n20942 = P2_DATAO_REG_30_ & n20786;
  assign n20943 = ~n20940 & ~n20941;
  assign n4499 = n20942 | ~n20943;
  assign n4504 = P2_DATAO_REG_31_ & n20786;
  assign n20946 = n15513 & ~n17339;
  assign n20947 = ~n15513 & n17339;
  assign n20948 = ~n20946 & ~n20947;
  assign n20949 = ~n15061 & n15177;
  assign n20950 = n15432 & ~n20949;
  assign n20951 = n14974 & n20950;
  assign n20952 = ~n20948 & n20951;
  assign n20953 = ~n14286 & n20950;
  assign n20954 = ~n14974 & n20953;
  assign n20955 = ~n15750 & n20954;
  assign n20956 = P2_EAX_REG_0_ & ~n20950;
  assign n20957 = n14286 & n20950;
  assign n20958 = ~n17339 & n20957;
  assign n20959 = ~n20956 & ~n20958;
  assign n20960 = ~n20952 & ~n20955;
  assign n4509 = ~n20959 | ~n20960;
  assign n20962 = ~n15513 & ~n17339;
  assign n20963 = ~n17326 & n20962;
  assign n20964 = ~n15510 & n20963;
  assign n20965 = ~n17326 & ~n20962;
  assign n20966 = n15510 & n20965;
  assign n20967 = ~n20964 & ~n20966;
  assign n20968 = n15510 & n20962;
  assign n20969 = ~n15510 & ~n20962;
  assign n20970 = ~n20968 & ~n20969;
  assign n20971 = n17326 & ~n20970;
  assign n20972 = n20967 & ~n20971;
  assign n20973 = n20951 & ~n20972;
  assign n20974 = ~n15728 & n20954;
  assign n20975 = P2_EAX_REG_1_ & ~n20950;
  assign n20976 = ~n17326 & n20957;
  assign n20977 = ~n20975 & ~n20976;
  assign n20978 = ~n20973 & ~n20974;
  assign n4514 = ~n20977 | ~n20978;
  assign n20980 = n17326 & ~n20962;
  assign n20981 = ~n15510 & ~n20980;
  assign n20982 = ~n20963 & ~n20981;
  assign n20983 = n15539 & n17306;
  assign n20984 = ~n15539 & ~n17306;
  assign n20985 = ~n20983 & ~n20984;
  assign n20986 = n20982 & ~n20985;
  assign n20987 = ~n20982 & n20985;
  assign n20988 = ~n20986 & ~n20987;
  assign n20989 = n20951 & ~n20988;
  assign n20990 = ~n15706 & n20954;
  assign n20991 = P2_EAX_REG_2_ & ~n20950;
  assign n20992 = ~n17306 & n20957;
  assign n20993 = ~n20991 & ~n20992;
  assign n20994 = ~n20989 & ~n20990;
  assign n4519 = ~n20993 | ~n20994;
  assign n20996 = n15539 & ~n17306;
  assign n20997 = ~n15539 & n17306;
  assign n20998 = ~n20982 & ~n20997;
  assign n20999 = ~n20996 & ~n20998;
  assign n21000 = ~n15557 & n17289;
  assign n21001 = n15557 & ~n17289;
  assign n21002 = ~n21000 & ~n21001;
  assign n21003 = n20999 & ~n21002;
  assign n21004 = ~n20999 & n21002;
  assign n21005 = ~n21003 & ~n21004;
  assign n21006 = n20951 & ~n21005;
  assign n21007 = ~n15684 & n20954;
  assign n21008 = P2_EAX_REG_3_ & ~n20950;
  assign n21009 = ~n17289 & n20957;
  assign n21010 = ~n21008 & ~n21009;
  assign n21011 = ~n21006 & ~n21007;
  assign n4524 = ~n21010 | ~n21011;
  assign n21013 = ~n15557 & ~n17289;
  assign n21014 = n15557 & n17289;
  assign n21015 = ~n20999 & ~n21014;
  assign n21016 = ~n21013 & ~n21015;
  assign n21017 = ~n15550 & n15551;
  assign n21018 = n15550 & ~n15551;
  assign n21019 = ~n15545 & ~n21018;
  assign n21020 = ~n21017 & ~n21019;
  assign n21021 = P2_INSTQUEUERD_ADDR_REG_4_ & ~n15491;
  assign n21022 = P2_INSTQUEUE_REG_0__4_ & n15483;
  assign n21023 = n21021 & ~n21022;
  assign n21024 = ~n21021 & n21022;
  assign n21025 = ~n21023 & ~n21024;
  assign n21026 = n21020 & ~n21025;
  assign n21027 = ~n21020 & n21025;
  assign n21028 = ~n21026 & ~n21027;
  assign n21029 = n17880 & ~n21028;
  assign n21030 = ~n17880 & n21028;
  assign n21031 = ~n21029 & ~n21030;
  assign n21032 = n21016 & ~n21031;
  assign n21033 = ~n21016 & n21031;
  assign n21034 = ~n21032 & ~n21033;
  assign n21035 = n20951 & ~n21034;
  assign n21036 = ~n15662 & n20954;
  assign n21037 = P2_EAX_REG_4_ & ~n20950;
  assign n21038 = ~n17880 & n20957;
  assign n21039 = ~n21037 & ~n21038;
  assign n21040 = ~n21035 & ~n21036;
  assign n4529 = ~n21039 | ~n21040;
  assign n21042 = ~n17880 & ~n21028;
  assign n21043 = n17880 & n21028;
  assign n21044 = ~n21016 & ~n21043;
  assign n21045 = ~n21042 & ~n21044;
  assign n21046 = n21021 & n21022;
  assign n21047 = ~n21021 & ~n21022;
  assign n21048 = ~n21020 & ~n21047;
  assign n21049 = ~n21046 & ~n21048;
  assign n21050 = P2_INSTQUEUE_REG_0__5_ & n15483;
  assign n21051 = n21049 & n21050;
  assign n21052 = ~n21049 & ~n21050;
  assign n21053 = ~n21051 & ~n21052;
  assign n21054 = n17996 & n21053;
  assign n21055 = ~n21045 & ~n21054;
  assign n21056 = ~n17996 & ~n21053;
  assign n21057 = n21055 & ~n21056;
  assign n21058 = n17996 & ~n21053;
  assign n21059 = ~n17996 & n21053;
  assign n21060 = ~n21058 & ~n21059;
  assign n21061 = n21045 & n21060;
  assign n21062 = ~n21057 & ~n21061;
  assign n21063 = n20951 & n21062;
  assign n21064 = ~n15640 & n20954;
  assign n21065 = P2_EAX_REG_5_ & ~n20950;
  assign n21066 = ~n17996 & n20957;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = ~n21063 & ~n21064;
  assign n4534 = ~n21067 | ~n21068;
  assign n21070 = ~n21049 & n21050;
  assign n21071 = P2_INSTQUEUE_REG_0__6_ & n15483;
  assign n21072 = ~n21070 & n21071;
  assign n21073 = n21070 & ~n21071;
  assign n21074 = ~n21072 & ~n21073;
  assign n21075 = n18116 & ~n21074;
  assign n21076 = ~n18116 & n21074;
  assign n21077 = ~n21075 & ~n21076;
  assign n21078 = ~n21055 & ~n21056;
  assign n21079 = ~n21077 & n21078;
  assign n21080 = n18116 & n21074;
  assign n21081 = ~n18116 & ~n21074;
  assign n21082 = ~n21080 & ~n21081;
  assign n21083 = ~n21078 & ~n21082;
  assign n21084 = ~n21079 & ~n21083;
  assign n21085 = n20951 & ~n21084;
  assign n21086 = ~n15618 & n20954;
  assign n21087 = P2_EAX_REG_6_ & ~n20950;
  assign n21088 = ~n18116 & n20957;
  assign n21089 = ~n21087 & ~n21088;
  assign n21090 = ~n21085 & ~n21086;
  assign n4539 = ~n21089 | ~n21090;
  assign n21092 = P2_EAX_REG_7_ & ~n20950;
  assign n21093 = ~n18242 & n20957;
  assign n21094 = ~n21092 & ~n21093;
  assign n21095 = ~n15590 & n20954;
  assign n21096 = n21078 & ~n21081;
  assign n21097 = n21070 & n21071;
  assign n21098 = P2_INSTQUEUE_REG_0__7_ & n15483;
  assign n21099 = ~n21097 & n21098;
  assign n21100 = n21097 & ~n21098;
  assign n21101 = ~n21099 & ~n21100;
  assign n21102 = n18242 & n21101;
  assign n21103 = ~n21080 & ~n21096;
  assign n21104 = ~n21102 & n21103;
  assign n21105 = ~n18242 & ~n21101;
  assign n21106 = n21104 & ~n21105;
  assign n21107 = ~n21078 & ~n21080;
  assign n21108 = n18242 & ~n21101;
  assign n21109 = ~n18242 & n21101;
  assign n21110 = ~n21108 & ~n21109;
  assign n21111 = ~n21081 & ~n21107;
  assign n21112 = n21110 & n21111;
  assign n21113 = ~n21106 & ~n21112;
  assign n21114 = n20951 & n21113;
  assign n21115 = n21094 & ~n21095;
  assign n4544 = n21114 | ~n21115;
  assign n21117 = P2_EAX_REG_8_ & ~n20950;
  assign n21118 = ~n18381 & n20957;
  assign n21119 = ~n21117 & ~n21118;
  assign n21120 = ~n20672 & n20954;
  assign n21121 = ~n21104 & ~n21105;
  assign n21122 = n21097 & n21098;
  assign n21123 = n15483 & ~n18373;
  assign n21124 = ~n21122 & n21123;
  assign n21125 = n21122 & ~n21123;
  assign n21126 = ~n21124 & ~n21125;
  assign n21127 = n18381 & ~n21126;
  assign n21128 = ~n18381 & n21126;
  assign n21129 = ~n21127 & ~n21128;
  assign n21130 = n21121 & ~n21129;
  assign n21131 = ~n21121 & n21129;
  assign n21132 = ~n21130 & ~n21131;
  assign n21133 = n20951 & ~n21132;
  assign n21134 = n21119 & ~n21120;
  assign n4549 = n21133 | ~n21134;
  assign n21136 = P2_EAX_REG_9_ & ~n20950;
  assign n21137 = ~n18485 & n20957;
  assign n21138 = ~n21136 & ~n21137;
  assign n21139 = ~n20664 & n20954;
  assign n21140 = ~n18381 & ~n21126;
  assign n21141 = n18381 & n21126;
  assign n21142 = ~n21121 & ~n21141;
  assign n21143 = ~n21140 & ~n21142;
  assign n21144 = n21122 & n21123;
  assign n21145 = n15483 & ~n18477;
  assign n21146 = ~n21144 & n21145;
  assign n21147 = n21144 & ~n21145;
  assign n21148 = ~n21146 & ~n21147;
  assign n21149 = n18485 & n21148;
  assign n21150 = ~n21143 & ~n21149;
  assign n21151 = ~n18485 & ~n21148;
  assign n21152 = n21150 & ~n21151;
  assign n21153 = n18485 & ~n21148;
  assign n21154 = ~n18485 & n21148;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = n21143 & n21155;
  assign n21157 = ~n21152 & ~n21156;
  assign n21158 = n20951 & n21157;
  assign n21159 = n21138 & ~n21139;
  assign n4554 = n21158 | ~n21159;
  assign n21161 = P2_EAX_REG_10_ & ~n20950;
  assign n21162 = ~n20656 & n20954;
  assign n21163 = ~n18584 & n20957;
  assign n21164 = n21144 & n21145;
  assign n21165 = n15483 & ~n18576;
  assign n21166 = ~n21164 & n21165;
  assign n21167 = n21164 & ~n21165;
  assign n21168 = ~n21166 & ~n21167;
  assign n21169 = n18584 & ~n21168;
  assign n21170 = ~n18584 & n21168;
  assign n21171 = ~n21169 & ~n21170;
  assign n21172 = ~n21150 & ~n21151;
  assign n21173 = ~n21171 & n21172;
  assign n21174 = n18584 & n21168;
  assign n21175 = ~n18584 & ~n21168;
  assign n21176 = ~n21174 & ~n21175;
  assign n21177 = ~n21172 & ~n21176;
  assign n21178 = ~n21173 & ~n21177;
  assign n21179 = n20951 & ~n21178;
  assign n21180 = ~n21161 & ~n21162;
  assign n21181 = ~n21163 & n21180;
  assign n4559 = n21179 | ~n21181;
  assign n21183 = P2_EAX_REG_11_ & ~n20950;
  assign n21184 = ~n20648 & n20954;
  assign n21185 = ~n18681 & n20957;
  assign n21186 = n21172 & ~n21175;
  assign n21187 = n21164 & n21165;
  assign n21188 = n15483 & ~n18673;
  assign n21189 = ~n21187 & n21188;
  assign n21190 = n21187 & ~n21188;
  assign n21191 = ~n21189 & ~n21190;
  assign n21192 = n18681 & n21191;
  assign n21193 = ~n21174 & ~n21186;
  assign n21194 = ~n21192 & n21193;
  assign n21195 = ~n18681 & ~n21191;
  assign n21196 = n21194 & ~n21195;
  assign n21197 = ~n21172 & ~n21174;
  assign n21198 = n18681 & ~n21191;
  assign n21199 = ~n18681 & n21191;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = ~n21175 & ~n21197;
  assign n21202 = n21200 & n21201;
  assign n21203 = ~n21196 & ~n21202;
  assign n21204 = n20951 & n21203;
  assign n21205 = ~n21183 & ~n21184;
  assign n21206 = ~n21185 & n21205;
  assign n4564 = n21204 | ~n21206;
  assign n21208 = P2_EAX_REG_12_ & ~n20950;
  assign n21209 = ~n20640 & n20954;
  assign n21210 = ~n18779 & n20957;
  assign n21211 = ~n21194 & ~n21195;
  assign n21212 = n21187 & n21188;
  assign n21213 = n15483 & ~n18771;
  assign n21214 = ~n21212 & n21213;
  assign n21215 = n21212 & ~n21213;
  assign n21216 = ~n21214 & ~n21215;
  assign n21217 = n18779 & ~n21216;
  assign n21218 = ~n18779 & n21216;
  assign n21219 = ~n21217 & ~n21218;
  assign n21220 = n21211 & ~n21219;
  assign n21221 = ~n21211 & n21219;
  assign n21222 = ~n21220 & ~n21221;
  assign n21223 = n20951 & ~n21222;
  assign n21224 = ~n21208 & ~n21209;
  assign n21225 = ~n21210 & n21224;
  assign n4569 = n21223 | ~n21225;
  assign n21227 = P2_EAX_REG_13_ & ~n20950;
  assign n21228 = ~n20632 & n20954;
  assign n21229 = ~n18880 & n20957;
  assign n21230 = ~n18779 & ~n21216;
  assign n21231 = n18779 & n21216;
  assign n21232 = ~n21211 & ~n21231;
  assign n21233 = ~n21230 & ~n21232;
  assign n21234 = n21212 & n21213;
  assign n21235 = n15483 & ~n18872;
  assign n21236 = ~n21234 & n21235;
  assign n21237 = n21234 & ~n21235;
  assign n21238 = ~n21236 & ~n21237;
  assign n21239 = n18880 & n21238;
  assign n21240 = ~n21233 & ~n21239;
  assign n21241 = ~n18880 & ~n21238;
  assign n21242 = n21240 & ~n21241;
  assign n21243 = n18880 & ~n21238;
  assign n21244 = ~n18880 & n21238;
  assign n21245 = ~n21243 & ~n21244;
  assign n21246 = n21233 & n21245;
  assign n21247 = ~n21242 & ~n21246;
  assign n21248 = n20951 & n21247;
  assign n21249 = ~n21227 & ~n21228;
  assign n21250 = ~n21229 & n21249;
  assign n4574 = n21248 | ~n21250;
  assign n21252 = P2_EAX_REG_14_ & ~n20950;
  assign n21253 = ~n20624 & n20954;
  assign n21254 = ~n18979 & n20957;
  assign n21255 = n21234 & n21235;
  assign n21256 = n15483 & ~n18971;
  assign n21257 = ~n21255 & n21256;
  assign n21258 = n21255 & ~n21256;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = n18979 & ~n21259;
  assign n21261 = ~n18979 & n21259;
  assign n21262 = ~n21260 & ~n21261;
  assign n21263 = ~n21240 & ~n21241;
  assign n21264 = ~n21262 & n21263;
  assign n21265 = n18979 & n21259;
  assign n21266 = ~n18979 & ~n21259;
  assign n21267 = ~n21265 & ~n21266;
  assign n21268 = ~n21263 & ~n21267;
  assign n21269 = ~n21264 & ~n21268;
  assign n21270 = n20951 & ~n21269;
  assign n21271 = ~n21252 & ~n21253;
  assign n21272 = ~n21254 & n21271;
  assign n4579 = n21270 | ~n21272;
  assign n21274 = P2_EAX_REG_15_ & ~n20950;
  assign n21275 = ~n20610 & n20954;
  assign n21276 = ~n19075 & n20957;
  assign n21277 = n21263 & ~n21266;
  assign n21278 = n21255 & n21256;
  assign n21279 = n15483 & ~n19067;
  assign n21280 = ~n21278 & n21279;
  assign n21281 = n21278 & ~n21279;
  assign n21282 = ~n21280 & ~n21281;
  assign n21283 = n19075 & n21282;
  assign n21284 = ~n21265 & ~n21277;
  assign n21285 = ~n21283 & n21284;
  assign n21286 = ~n19075 & ~n21282;
  assign n21287 = n21285 & ~n21286;
  assign n21288 = ~n21263 & ~n21265;
  assign n21289 = n19075 & ~n21282;
  assign n21290 = ~n19075 & n21282;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = ~n21266 & ~n21288;
  assign n21293 = n21291 & n21292;
  assign n21294 = ~n21287 & ~n21293;
  assign n21295 = n20951 & n21294;
  assign n21296 = ~n21274 & ~n21275;
  assign n21297 = ~n21276 & n21296;
  assign n4584 = n21295 | ~n21297;
  assign n21299 = ~n14404 & n20953;
  assign n21300 = ~n15755 & n21299;
  assign n21301 = n14365 & n20953;
  assign n21302 = ~n15750 & n21301;
  assign n21303 = P2_EAX_REG_16_ & ~n20950;
  assign n21304 = ~n19145 & n20957;
  assign n21305 = ~n21285 & ~n21286;
  assign n21306 = n21278 & n21279;
  assign n21307 = P2_INSTQUEUERD_ADDR_REG_2_ & ~n14175;
  assign n21308 = ~n14187 & ~n21307;
  assign n21309 = ~P2_INSTQUEUERD_ADDR_REG_3_ & n21307;
  assign n21310 = P2_INSTQUEUERD_ADDR_REG_3_ & ~n21307;
  assign n21311 = ~n21309 & ~n21310;
  assign n21312 = n21308 & ~n21311;
  assign n21313 = ~P2_INSTQUEUERD_ADDR_REG_0_ & n14555;
  assign n21314 = n21312 & n21313;
  assign n21315 = P2_INSTQUEUE_REG_15__0_ & n21314;
  assign n21316 = P2_INSTQUEUERD_ADDR_REG_0_ & n14555;
  assign n21317 = n21312 & n21316;
  assign n21318 = P2_INSTQUEUE_REG_14__0_ & n21317;
  assign n21319 = ~P2_INSTQUEUERD_ADDR_REG_0_ & ~n14555;
  assign n21320 = n21312 & n21319;
  assign n21321 = P2_INSTQUEUE_REG_13__0_ & n21320;
  assign n21322 = P2_INSTQUEUERD_ADDR_REG_0_ & ~n14555;
  assign n21323 = n21312 & n21322;
  assign n21324 = P2_INSTQUEUE_REG_12__0_ & n21323;
  assign n21325 = ~n21315 & ~n21318;
  assign n21326 = ~n21321 & n21325;
  assign n21327 = ~n21324 & n21326;
  assign n21328 = ~n21308 & ~n21311;
  assign n21329 = n21313 & n21328;
  assign n21330 = P2_INSTQUEUE_REG_11__0_ & n21329;
  assign n21331 = n21316 & n21328;
  assign n21332 = P2_INSTQUEUE_REG_10__0_ & n21331;
  assign n21333 = n21319 & n21328;
  assign n21334 = P2_INSTQUEUE_REG_9__0_ & n21333;
  assign n21335 = n21322 & n21328;
  assign n21336 = P2_INSTQUEUE_REG_8__0_ & n21335;
  assign n21337 = ~n21330 & ~n21332;
  assign n21338 = ~n21334 & n21337;
  assign n21339 = ~n21336 & n21338;
  assign n21340 = n21308 & n21311;
  assign n21341 = n21313 & n21340;
  assign n21342 = P2_INSTQUEUE_REG_7__0_ & n21341;
  assign n21343 = n21316 & n21340;
  assign n21344 = P2_INSTQUEUE_REG_6__0_ & n21343;
  assign n21345 = n21319 & n21340;
  assign n21346 = P2_INSTQUEUE_REG_5__0_ & n21345;
  assign n21347 = n21322 & n21340;
  assign n21348 = P2_INSTQUEUE_REG_4__0_ & n21347;
  assign n21349 = ~n21342 & ~n21344;
  assign n21350 = ~n21346 & n21349;
  assign n21351 = ~n21348 & n21350;
  assign n21352 = ~n21308 & n21311;
  assign n21353 = n21313 & n21352;
  assign n21354 = P2_INSTQUEUE_REG_3__0_ & n21353;
  assign n21355 = n21316 & n21352;
  assign n21356 = P2_INSTQUEUE_REG_2__0_ & n21355;
  assign n21357 = n21319 & n21352;
  assign n21358 = P2_INSTQUEUE_REG_1__0_ & n21357;
  assign n21359 = n21322 & n21352;
  assign n21360 = P2_INSTQUEUE_REG_0__0_ & n21359;
  assign n21361 = ~n21354 & ~n21356;
  assign n21362 = ~n21358 & n21361;
  assign n21363 = ~n21360 & n21362;
  assign n21364 = n21327 & n21339;
  assign n21365 = n21351 & n21364;
  assign n21366 = n21363 & n21365;
  assign n21367 = n15007 & ~n21366;
  assign n21368 = n15483 & ~n21366;
  assign n21369 = ~n21367 & ~n21368;
  assign n21370 = ~n21306 & ~n21369;
  assign n21371 = n21306 & n21369;
  assign n21372 = ~n21370 & ~n21371;
  assign n21373 = n19145 & ~n21372;
  assign n21374 = ~n19145 & n21372;
  assign n21375 = ~n21373 & ~n21374;
  assign n21376 = n21305 & ~n21375;
  assign n21377 = ~n21305 & n21375;
  assign n21378 = ~n21376 & ~n21377;
  assign n21379 = n20951 & ~n21378;
  assign n21380 = ~n21300 & ~n21302;
  assign n21381 = ~n21303 & n21380;
  assign n21382 = ~n21304 & n21381;
  assign n4589 = n21379 | ~n21382;
  assign n21384 = ~n15733 & n21299;
  assign n21385 = ~n15728 & n21301;
  assign n21386 = P2_EAX_REG_17_ & ~n20950;
  assign n21387 = ~n19208 & n20957;
  assign n21388 = ~n19145 & ~n21372;
  assign n21389 = n19145 & n21372;
  assign n21390 = ~n21305 & ~n21389;
  assign n21391 = ~n21388 & ~n21390;
  assign n21392 = n21306 & ~n21369;
  assign n21393 = P2_INSTQUEUE_REG_15__1_ & n21314;
  assign n21394 = P2_INSTQUEUE_REG_14__1_ & n21317;
  assign n21395 = P2_INSTQUEUE_REG_13__1_ & n21320;
  assign n21396 = P2_INSTQUEUE_REG_12__1_ & n21323;
  assign n21397 = ~n21393 & ~n21394;
  assign n21398 = ~n21395 & n21397;
  assign n21399 = ~n21396 & n21398;
  assign n21400 = P2_INSTQUEUE_REG_11__1_ & n21329;
  assign n21401 = P2_INSTQUEUE_REG_10__1_ & n21331;
  assign n21402 = P2_INSTQUEUE_REG_9__1_ & n21333;
  assign n21403 = P2_INSTQUEUE_REG_8__1_ & n21335;
  assign n21404 = ~n21400 & ~n21401;
  assign n21405 = ~n21402 & n21404;
  assign n21406 = ~n21403 & n21405;
  assign n21407 = P2_INSTQUEUE_REG_7__1_ & n21341;
  assign n21408 = P2_INSTQUEUE_REG_6__1_ & n21343;
  assign n21409 = P2_INSTQUEUE_REG_5__1_ & n21345;
  assign n21410 = P2_INSTQUEUE_REG_4__1_ & n21347;
  assign n21411 = ~n21407 & ~n21408;
  assign n21412 = ~n21409 & n21411;
  assign n21413 = ~n21410 & n21412;
  assign n21414 = P2_INSTQUEUE_REG_3__1_ & n21353;
  assign n21415 = P2_INSTQUEUE_REG_2__1_ & n21355;
  assign n21416 = P2_INSTQUEUE_REG_1__1_ & n21357;
  assign n21417 = P2_INSTQUEUE_REG_0__1_ & n21359;
  assign n21418 = ~n21414 & ~n21415;
  assign n21419 = ~n21416 & n21418;
  assign n21420 = ~n21417 & n21419;
  assign n21421 = n21399 & n21406;
  assign n21422 = n21413 & n21421;
  assign n21423 = n21420 & n21422;
  assign n21424 = n15007 & ~n21423;
  assign n21425 = n15483 & ~n21423;
  assign n21426 = ~n21424 & ~n21425;
  assign n21427 = ~n21392 & ~n21426;
  assign n21428 = n21392 & n21426;
  assign n21429 = ~n21427 & ~n21428;
  assign n21430 = n19208 & ~n21429;
  assign n21431 = ~n19208 & n21429;
  assign n21432 = ~n21430 & ~n21431;
  assign n21433 = n21391 & ~n21432;
  assign n21434 = ~n21391 & n21432;
  assign n21435 = ~n21433 & ~n21434;
  assign n21436 = n20951 & ~n21435;
  assign n21437 = ~n21384 & ~n21385;
  assign n21438 = ~n21386 & n21437;
  assign n21439 = ~n21387 & n21438;
  assign n4594 = n21436 | ~n21439;
  assign n21441 = ~n15711 & n21299;
  assign n21442 = ~n15706 & n21301;
  assign n21443 = P2_EAX_REG_18_ & ~n20950;
  assign n21444 = ~n19276 & n20957;
  assign n21445 = ~n19208 & ~n21429;
  assign n21446 = n19208 & n21429;
  assign n21447 = ~n21391 & ~n21446;
  assign n21448 = ~n21445 & ~n21447;
  assign n21449 = n21392 & ~n21426;
  assign n21450 = P2_INSTQUEUE_REG_15__2_ & n21314;
  assign n21451 = P2_INSTQUEUE_REG_14__2_ & n21317;
  assign n21452 = P2_INSTQUEUE_REG_13__2_ & n21320;
  assign n21453 = P2_INSTQUEUE_REG_12__2_ & n21323;
  assign n21454 = ~n21450 & ~n21451;
  assign n21455 = ~n21452 & n21454;
  assign n21456 = ~n21453 & n21455;
  assign n21457 = P2_INSTQUEUE_REG_11__2_ & n21329;
  assign n21458 = P2_INSTQUEUE_REG_10__2_ & n21331;
  assign n21459 = P2_INSTQUEUE_REG_9__2_ & n21333;
  assign n21460 = P2_INSTQUEUE_REG_8__2_ & n21335;
  assign n21461 = ~n21457 & ~n21458;
  assign n21462 = ~n21459 & n21461;
  assign n21463 = ~n21460 & n21462;
  assign n21464 = P2_INSTQUEUE_REG_7__2_ & n21341;
  assign n21465 = P2_INSTQUEUE_REG_6__2_ & n21343;
  assign n21466 = P2_INSTQUEUE_REG_5__2_ & n21345;
  assign n21467 = P2_INSTQUEUE_REG_4__2_ & n21347;
  assign n21468 = ~n21464 & ~n21465;
  assign n21469 = ~n21466 & n21468;
  assign n21470 = ~n21467 & n21469;
  assign n21471 = P2_INSTQUEUE_REG_3__2_ & n21353;
  assign n21472 = P2_INSTQUEUE_REG_2__2_ & n21355;
  assign n21473 = P2_INSTQUEUE_REG_1__2_ & n21357;
  assign n21474 = P2_INSTQUEUE_REG_0__2_ & n21359;
  assign n21475 = ~n21471 & ~n21472;
  assign n21476 = ~n21473 & n21475;
  assign n21477 = ~n21474 & n21476;
  assign n21478 = n21456 & n21463;
  assign n21479 = n21470 & n21478;
  assign n21480 = n21477 & n21479;
  assign n21481 = n15007 & ~n21480;
  assign n21482 = n15483 & ~n21480;
  assign n21483 = ~n21481 & ~n21482;
  assign n21484 = ~n21449 & ~n21483;
  assign n21485 = n21449 & n21483;
  assign n21486 = ~n21484 & ~n21485;
  assign n21487 = n19276 & ~n21486;
  assign n21488 = ~n19276 & n21486;
  assign n21489 = ~n21487 & ~n21488;
  assign n21490 = n21448 & ~n21489;
  assign n21491 = ~n21448 & n21489;
  assign n21492 = ~n21490 & ~n21491;
  assign n21493 = n20951 & ~n21492;
  assign n21494 = ~n21441 & ~n21442;
  assign n21495 = ~n21443 & n21494;
  assign n21496 = ~n21444 & n21495;
  assign n4599 = n21493 | ~n21496;
  assign n21498 = ~n15689 & n21299;
  assign n21499 = ~n15684 & n21301;
  assign n21500 = P2_EAX_REG_19_ & ~n20950;
  assign n21501 = ~n19344 & n20957;
  assign n21502 = ~n19276 & ~n21486;
  assign n21503 = n19276 & n21486;
  assign n21504 = ~n21448 & ~n21503;
  assign n21505 = ~n21502 & ~n21504;
  assign n21506 = n21449 & ~n21483;
  assign n21507 = P2_INSTQUEUE_REG_15__3_ & n21314;
  assign n21508 = P2_INSTQUEUE_REG_14__3_ & n21317;
  assign n21509 = P2_INSTQUEUE_REG_13__3_ & n21320;
  assign n21510 = P2_INSTQUEUE_REG_12__3_ & n21323;
  assign n21511 = ~n21507 & ~n21508;
  assign n21512 = ~n21509 & n21511;
  assign n21513 = ~n21510 & n21512;
  assign n21514 = P2_INSTQUEUE_REG_11__3_ & n21329;
  assign n21515 = P2_INSTQUEUE_REG_10__3_ & n21331;
  assign n21516 = P2_INSTQUEUE_REG_9__3_ & n21333;
  assign n21517 = P2_INSTQUEUE_REG_8__3_ & n21335;
  assign n21518 = ~n21514 & ~n21515;
  assign n21519 = ~n21516 & n21518;
  assign n21520 = ~n21517 & n21519;
  assign n21521 = P2_INSTQUEUE_REG_7__3_ & n21341;
  assign n21522 = P2_INSTQUEUE_REG_6__3_ & n21343;
  assign n21523 = P2_INSTQUEUE_REG_5__3_ & n21345;
  assign n21524 = P2_INSTQUEUE_REG_4__3_ & n21347;
  assign n21525 = ~n21521 & ~n21522;
  assign n21526 = ~n21523 & n21525;
  assign n21527 = ~n21524 & n21526;
  assign n21528 = P2_INSTQUEUE_REG_3__3_ & n21353;
  assign n21529 = P2_INSTQUEUE_REG_2__3_ & n21355;
  assign n21530 = P2_INSTQUEUE_REG_1__3_ & n21357;
  assign n21531 = P2_INSTQUEUE_REG_0__3_ & n21359;
  assign n21532 = ~n21528 & ~n21529;
  assign n21533 = ~n21530 & n21532;
  assign n21534 = ~n21531 & n21533;
  assign n21535 = n21513 & n21520;
  assign n21536 = n21527 & n21535;
  assign n21537 = n21534 & n21536;
  assign n21538 = n15007 & ~n21537;
  assign n21539 = n15483 & ~n21537;
  assign n21540 = ~n21538 & ~n21539;
  assign n21541 = ~n21506 & ~n21540;
  assign n21542 = n21506 & n21540;
  assign n21543 = ~n21541 & ~n21542;
  assign n21544 = n19344 & ~n21543;
  assign n21545 = ~n19344 & n21543;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = n21505 & ~n21546;
  assign n21548 = ~n21505 & n21546;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = n20951 & ~n21549;
  assign n21551 = ~n21498 & ~n21499;
  assign n21552 = ~n21500 & n21551;
  assign n21553 = ~n21501 & n21552;
  assign n4604 = n21550 | ~n21553;
  assign n21555 = ~n15667 & n21299;
  assign n21556 = ~n15662 & n21301;
  assign n21557 = P2_EAX_REG_20_ & ~n20950;
  assign n21558 = ~n19411 & n20957;
  assign n21559 = ~n19344 & ~n21543;
  assign n21560 = n19344 & n21543;
  assign n21561 = ~n21505 & ~n21560;
  assign n21562 = ~n21559 & ~n21561;
  assign n21563 = n21506 & ~n21540;
  assign n21564 = P2_INSTQUEUE_REG_15__4_ & n21314;
  assign n21565 = P2_INSTQUEUE_REG_14__4_ & n21317;
  assign n21566 = P2_INSTQUEUE_REG_13__4_ & n21320;
  assign n21567 = P2_INSTQUEUE_REG_12__4_ & n21323;
  assign n21568 = ~n21564 & ~n21565;
  assign n21569 = ~n21566 & n21568;
  assign n21570 = ~n21567 & n21569;
  assign n21571 = P2_INSTQUEUE_REG_11__4_ & n21329;
  assign n21572 = P2_INSTQUEUE_REG_10__4_ & n21331;
  assign n21573 = P2_INSTQUEUE_REG_9__4_ & n21333;
  assign n21574 = P2_INSTQUEUE_REG_8__4_ & n21335;
  assign n21575 = ~n21571 & ~n21572;
  assign n21576 = ~n21573 & n21575;
  assign n21577 = ~n21574 & n21576;
  assign n21578 = P2_INSTQUEUE_REG_7__4_ & n21341;
  assign n21579 = P2_INSTQUEUE_REG_6__4_ & n21343;
  assign n21580 = P2_INSTQUEUE_REG_5__4_ & n21345;
  assign n21581 = P2_INSTQUEUE_REG_4__4_ & n21347;
  assign n21582 = ~n21578 & ~n21579;
  assign n21583 = ~n21580 & n21582;
  assign n21584 = ~n21581 & n21583;
  assign n21585 = P2_INSTQUEUE_REG_3__4_ & n21353;
  assign n21586 = P2_INSTQUEUE_REG_2__4_ & n21355;
  assign n21587 = P2_INSTQUEUE_REG_1__4_ & n21357;
  assign n21588 = P2_INSTQUEUE_REG_0__4_ & n21359;
  assign n21589 = ~n21585 & ~n21586;
  assign n21590 = ~n21587 & n21589;
  assign n21591 = ~n21588 & n21590;
  assign n21592 = n21570 & n21577;
  assign n21593 = n21584 & n21592;
  assign n21594 = n21591 & n21593;
  assign n21595 = n15007 & ~n21594;
  assign n21596 = n15483 & ~n21594;
  assign n21597 = ~n21595 & ~n21596;
  assign n21598 = ~n21563 & ~n21597;
  assign n21599 = n21563 & n21597;
  assign n21600 = ~n21598 & ~n21599;
  assign n21601 = n19411 & ~n21600;
  assign n21602 = ~n19411 & n21600;
  assign n21603 = ~n21601 & ~n21602;
  assign n21604 = n21562 & ~n21603;
  assign n21605 = ~n21562 & n21603;
  assign n21606 = ~n21604 & ~n21605;
  assign n21607 = n20951 & ~n21606;
  assign n21608 = ~n21555 & ~n21556;
  assign n21609 = ~n21557 & n21608;
  assign n21610 = ~n21558 & n21609;
  assign n4609 = n21607 | ~n21610;
  assign n21612 = ~n15645 & n21299;
  assign n21613 = ~n15640 & n21301;
  assign n21614 = P2_EAX_REG_21_ & ~n20950;
  assign n21615 = ~n19477 & n20957;
  assign n21616 = ~n19411 & ~n21600;
  assign n21617 = n19411 & n21600;
  assign n21618 = ~n21562 & ~n21617;
  assign n21619 = ~n21616 & ~n21618;
  assign n21620 = n21563 & ~n21597;
  assign n21621 = P2_INSTQUEUE_REG_15__5_ & n21314;
  assign n21622 = P2_INSTQUEUE_REG_14__5_ & n21317;
  assign n21623 = P2_INSTQUEUE_REG_13__5_ & n21320;
  assign n21624 = P2_INSTQUEUE_REG_12__5_ & n21323;
  assign n21625 = ~n21621 & ~n21622;
  assign n21626 = ~n21623 & n21625;
  assign n21627 = ~n21624 & n21626;
  assign n21628 = P2_INSTQUEUE_REG_11__5_ & n21329;
  assign n21629 = P2_INSTQUEUE_REG_10__5_ & n21331;
  assign n21630 = P2_INSTQUEUE_REG_9__5_ & n21333;
  assign n21631 = P2_INSTQUEUE_REG_8__5_ & n21335;
  assign n21632 = ~n21628 & ~n21629;
  assign n21633 = ~n21630 & n21632;
  assign n21634 = ~n21631 & n21633;
  assign n21635 = P2_INSTQUEUE_REG_7__5_ & n21341;
  assign n21636 = P2_INSTQUEUE_REG_6__5_ & n21343;
  assign n21637 = P2_INSTQUEUE_REG_5__5_ & n21345;
  assign n21638 = P2_INSTQUEUE_REG_4__5_ & n21347;
  assign n21639 = ~n21635 & ~n21636;
  assign n21640 = ~n21637 & n21639;
  assign n21641 = ~n21638 & n21640;
  assign n21642 = P2_INSTQUEUE_REG_3__5_ & n21353;
  assign n21643 = P2_INSTQUEUE_REG_2__5_ & n21355;
  assign n21644 = P2_INSTQUEUE_REG_1__5_ & n21357;
  assign n21645 = P2_INSTQUEUE_REG_0__5_ & n21359;
  assign n21646 = ~n21642 & ~n21643;
  assign n21647 = ~n21644 & n21646;
  assign n21648 = ~n21645 & n21647;
  assign n21649 = n21627 & n21634;
  assign n21650 = n21641 & n21649;
  assign n21651 = n21648 & n21650;
  assign n21652 = n15007 & ~n21651;
  assign n21653 = n15483 & ~n21651;
  assign n21654 = ~n21652 & ~n21653;
  assign n21655 = ~n21620 & ~n21654;
  assign n21656 = n21620 & n21654;
  assign n21657 = ~n21655 & ~n21656;
  assign n21658 = n19477 & ~n21657;
  assign n21659 = ~n19477 & n21657;
  assign n21660 = ~n21658 & ~n21659;
  assign n21661 = n21619 & ~n21660;
  assign n21662 = ~n21619 & n21660;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = n20951 & ~n21663;
  assign n21665 = ~n21612 & ~n21613;
  assign n21666 = ~n21614 & n21665;
  assign n21667 = ~n21615 & n21666;
  assign n4614 = n21664 | ~n21667;
  assign n21669 = ~n15623 & n21299;
  assign n21670 = ~n15618 & n21301;
  assign n21671 = P2_EAX_REG_22_ & ~n20950;
  assign n21672 = ~n19543 & n20957;
  assign n21673 = ~n19477 & ~n21657;
  assign n21674 = n19477 & n21657;
  assign n21675 = ~n21619 & ~n21674;
  assign n21676 = ~n21673 & ~n21675;
  assign n21677 = n21620 & ~n21654;
  assign n21678 = P2_INSTQUEUE_REG_15__6_ & n21314;
  assign n21679 = P2_INSTQUEUE_REG_14__6_ & n21317;
  assign n21680 = P2_INSTQUEUE_REG_13__6_ & n21320;
  assign n21681 = P2_INSTQUEUE_REG_12__6_ & n21323;
  assign n21682 = ~n21678 & ~n21679;
  assign n21683 = ~n21680 & n21682;
  assign n21684 = ~n21681 & n21683;
  assign n21685 = P2_INSTQUEUE_REG_11__6_ & n21329;
  assign n21686 = P2_INSTQUEUE_REG_10__6_ & n21331;
  assign n21687 = P2_INSTQUEUE_REG_9__6_ & n21333;
  assign n21688 = P2_INSTQUEUE_REG_8__6_ & n21335;
  assign n21689 = ~n21685 & ~n21686;
  assign n21690 = ~n21687 & n21689;
  assign n21691 = ~n21688 & n21690;
  assign n21692 = P2_INSTQUEUE_REG_7__6_ & n21341;
  assign n21693 = P2_INSTQUEUE_REG_6__6_ & n21343;
  assign n21694 = P2_INSTQUEUE_REG_5__6_ & n21345;
  assign n21695 = P2_INSTQUEUE_REG_4__6_ & n21347;
  assign n21696 = ~n21692 & ~n21693;
  assign n21697 = ~n21694 & n21696;
  assign n21698 = ~n21695 & n21697;
  assign n21699 = P2_INSTQUEUE_REG_3__6_ & n21353;
  assign n21700 = P2_INSTQUEUE_REG_2__6_ & n21355;
  assign n21701 = P2_INSTQUEUE_REG_1__6_ & n21357;
  assign n21702 = P2_INSTQUEUE_REG_0__6_ & n21359;
  assign n21703 = ~n21699 & ~n21700;
  assign n21704 = ~n21701 & n21703;
  assign n21705 = ~n21702 & n21704;
  assign n21706 = n21684 & n21691;
  assign n21707 = n21698 & n21706;
  assign n21708 = n21705 & n21707;
  assign n21709 = n15007 & ~n21708;
  assign n21710 = n15483 & ~n21708;
  assign n21711 = ~n21709 & ~n21710;
  assign n21712 = ~n21677 & ~n21711;
  assign n21713 = n21677 & n21711;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = n19543 & ~n21714;
  assign n21716 = ~n19543 & n21714;
  assign n21717 = ~n21715 & ~n21716;
  assign n21718 = n21676 & ~n21717;
  assign n21719 = ~n21676 & n21717;
  assign n21720 = ~n21718 & ~n21719;
  assign n21721 = n20951 & ~n21720;
  assign n21722 = ~n21669 & ~n21670;
  assign n21723 = ~n21671 & n21722;
  assign n21724 = ~n21672 & n21723;
  assign n4619 = n21721 | ~n21724;
  assign n21726 = ~n15600 & n21299;
  assign n21727 = ~n15590 & n21301;
  assign n21728 = P2_EAX_REG_23_ & ~n20950;
  assign n21729 = ~n19612 & n20957;
  assign n21730 = ~n19543 & ~n21714;
  assign n21731 = n19543 & n21714;
  assign n21732 = ~n21676 & ~n21731;
  assign n21733 = ~n21730 & ~n21732;
  assign n21734 = n21677 & ~n21711;
  assign n21735 = P2_INSTQUEUE_REG_15__7_ & n21314;
  assign n21736 = P2_INSTQUEUE_REG_14__7_ & n21317;
  assign n21737 = P2_INSTQUEUE_REG_13__7_ & n21320;
  assign n21738 = P2_INSTQUEUE_REG_12__7_ & n21323;
  assign n21739 = ~n21735 & ~n21736;
  assign n21740 = ~n21737 & n21739;
  assign n21741 = ~n21738 & n21740;
  assign n21742 = P2_INSTQUEUE_REG_11__7_ & n21329;
  assign n21743 = P2_INSTQUEUE_REG_10__7_ & n21331;
  assign n21744 = P2_INSTQUEUE_REG_9__7_ & n21333;
  assign n21745 = P2_INSTQUEUE_REG_8__7_ & n21335;
  assign n21746 = ~n21742 & ~n21743;
  assign n21747 = ~n21744 & n21746;
  assign n21748 = ~n21745 & n21747;
  assign n21749 = P2_INSTQUEUE_REG_7__7_ & n21341;
  assign n21750 = P2_INSTQUEUE_REG_6__7_ & n21343;
  assign n21751 = P2_INSTQUEUE_REG_5__7_ & n21345;
  assign n21752 = P2_INSTQUEUE_REG_4__7_ & n21347;
  assign n21753 = ~n21749 & ~n21750;
  assign n21754 = ~n21751 & n21753;
  assign n21755 = ~n21752 & n21754;
  assign n21756 = P2_INSTQUEUE_REG_3__7_ & n21353;
  assign n21757 = P2_INSTQUEUE_REG_2__7_ & n21355;
  assign n21758 = P2_INSTQUEUE_REG_1__7_ & n21357;
  assign n21759 = P2_INSTQUEUE_REG_0__7_ & n21359;
  assign n21760 = ~n21756 & ~n21757;
  assign n21761 = ~n21758 & n21760;
  assign n21762 = ~n21759 & n21761;
  assign n21763 = n21741 & n21748;
  assign n21764 = n21755 & n21763;
  assign n21765 = n21762 & n21764;
  assign n21766 = n15007 & ~n21765;
  assign n21767 = P2_INSTQUEUERD_ADDR_REG_3_ & ~P2_INSTQUEUERD_ADDR_REG_2_;
  assign n21768 = ~P2_INSTQUEUERD_ADDR_REG_3_ & P2_INSTQUEUERD_ADDR_REG_2_;
  assign n21769 = ~n21767 & ~n21768;
  assign n21770 = ~P2_INSTQUEUE_REG_6__0_ & n21769;
  assign n21771 = ~P2_INSTQUEUE_REG_14__0_ & ~n21769;
  assign n21772 = ~n21770 & ~n21771;
  assign n21773 = n14149 & n21772;
  assign n21774 = ~P2_INSTQUEUE_REG_2__0_ & n21769;
  assign n21775 = ~P2_INSTQUEUE_REG_10__0_ & ~n21769;
  assign n21776 = ~n21774 & ~n21775;
  assign n21777 = n14155 & n21776;
  assign n21778 = ~P2_INSTQUEUE_REG_1__0_ & n21769;
  assign n21779 = ~P2_INSTQUEUE_REG_9__0_ & ~n21769;
  assign n21780 = ~n21778 & ~n21779;
  assign n21781 = n14161 & n21780;
  assign n21782 = ~P2_INSTQUEUE_REG_3__0_ & n21769;
  assign n21783 = ~P2_INSTQUEUE_REG_11__0_ & ~n21769;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = n14167 & n21784;
  assign n21786 = ~n21773 & ~n21777;
  assign n21787 = ~n21781 & n21786;
  assign n21788 = ~n21785 & n21787;
  assign n21789 = ~P2_INSTQUEUE_REG_0__0_ & n21769;
  assign n21790 = ~P2_INSTQUEUE_REG_8__0_ & ~n21769;
  assign n21791 = ~n21789 & ~n21790;
  assign n21792 = n14176 & n21791;
  assign n21793 = ~P2_INSTQUEUE_REG_5__0_ & n21769;
  assign n21794 = ~P2_INSTQUEUE_REG_13__0_ & ~n21769;
  assign n21795 = ~n21793 & ~n21794;
  assign n21796 = n14182 & n21795;
  assign n21797 = ~P2_INSTQUEUE_REG_4__0_ & n21769;
  assign n21798 = ~P2_INSTQUEUE_REG_12__0_ & ~n21769;
  assign n21799 = ~n21797 & ~n21798;
  assign n21800 = n14187 & n21799;
  assign n21801 = ~P2_INSTQUEUE_REG_7__0_ & n21769;
  assign n21802 = ~P2_INSTQUEUE_REG_15__0_ & ~n21769;
  assign n21803 = ~n21801 & ~n21802;
  assign n21804 = n14193 & n21803;
  assign n21805 = ~n21792 & ~n21796;
  assign n21806 = ~n21800 & n21805;
  assign n21807 = ~n21804 & n21806;
  assign n21808 = n21788 & n21807;
  assign n21809 = ~n21765 & n21808;
  assign n21810 = n21765 & ~n21808;
  assign n21811 = ~n21809 & ~n21810;
  assign n21812 = n15483 & ~n21811;
  assign n21813 = ~n21766 & ~n21812;
  assign n21814 = n15007 & ~n21808;
  assign n21815 = ~n21813 & ~n21814;
  assign n21816 = n21813 & n21814;
  assign n21817 = ~n21815 & ~n21816;
  assign n21818 = ~n21734 & ~n21817;
  assign n21819 = n21734 & n21817;
  assign n21820 = ~n21818 & ~n21819;
  assign n21821 = n19612 & ~n21820;
  assign n21822 = ~n19612 & n21820;
  assign n21823 = ~n21821 & ~n21822;
  assign n21824 = n21733 & ~n21823;
  assign n21825 = ~n21733 & n21823;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = n20951 & ~n21826;
  assign n21828 = ~n21726 & ~n21727;
  assign n21829 = ~n21728 & n21828;
  assign n21830 = ~n21729 & n21829;
  assign n4624 = n21827 | ~n21830;
  assign n21832 = ~n15762 & n21299;
  assign n21833 = ~n20672 & n21301;
  assign n21834 = P2_EAX_REG_24_ & ~n20950;
  assign n21835 = ~n19674 & n20957;
  assign n21836 = ~n19612 & ~n21820;
  assign n21837 = n19612 & n21820;
  assign n21838 = ~n21733 & ~n21837;
  assign n21839 = ~n21836 & ~n21838;
  assign n21840 = ~n21813 & n21814;
  assign n21841 = n21813 & ~n21814;
  assign n21842 = n21734 & ~n21841;
  assign n21843 = ~n21840 & ~n21842;
  assign n21844 = ~n21765 & ~n21808;
  assign n21845 = ~P2_INSTQUEUE_REG_6__1_ & n21769;
  assign n21846 = ~P2_INSTQUEUE_REG_14__1_ & ~n21769;
  assign n21847 = ~n21845 & ~n21846;
  assign n21848 = n14149 & n21847;
  assign n21849 = ~P2_INSTQUEUE_REG_2__1_ & n21769;
  assign n21850 = ~P2_INSTQUEUE_REG_10__1_ & ~n21769;
  assign n21851 = ~n21849 & ~n21850;
  assign n21852 = n14155 & n21851;
  assign n21853 = ~P2_INSTQUEUE_REG_1__1_ & n21769;
  assign n21854 = ~P2_INSTQUEUE_REG_9__1_ & ~n21769;
  assign n21855 = ~n21853 & ~n21854;
  assign n21856 = n14161 & n21855;
  assign n21857 = ~P2_INSTQUEUE_REG_3__1_ & n21769;
  assign n21858 = ~P2_INSTQUEUE_REG_11__1_ & ~n21769;
  assign n21859 = ~n21857 & ~n21858;
  assign n21860 = n14167 & n21859;
  assign n21861 = ~n21848 & ~n21852;
  assign n21862 = ~n21856 & n21861;
  assign n21863 = ~n21860 & n21862;
  assign n21864 = ~P2_INSTQUEUE_REG_0__1_ & n21769;
  assign n21865 = ~P2_INSTQUEUE_REG_8__1_ & ~n21769;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = n14176 & n21866;
  assign n21868 = ~P2_INSTQUEUE_REG_5__1_ & n21769;
  assign n21869 = ~P2_INSTQUEUE_REG_13__1_ & ~n21769;
  assign n21870 = ~n21868 & ~n21869;
  assign n21871 = n14182 & n21870;
  assign n21872 = ~P2_INSTQUEUE_REG_4__1_ & n21769;
  assign n21873 = ~P2_INSTQUEUE_REG_12__1_ & ~n21769;
  assign n21874 = ~n21872 & ~n21873;
  assign n21875 = n14187 & n21874;
  assign n21876 = ~P2_INSTQUEUE_REG_7__1_ & n21769;
  assign n21877 = ~P2_INSTQUEUE_REG_15__1_ & ~n21769;
  assign n21878 = ~n21876 & ~n21877;
  assign n21879 = n14193 & n21878;
  assign n21880 = ~n21867 & ~n21871;
  assign n21881 = ~n21875 & n21880;
  assign n21882 = ~n21879 & n21881;
  assign n21883 = n21863 & n21882;
  assign n21884 = n21844 & n21883;
  assign n21885 = ~n21844 & ~n21883;
  assign n21886 = ~n21884 & ~n21885;
  assign n21887 = n15483 & ~n21886;
  assign n21888 = n15007 & ~n21883;
  assign n21889 = n21887 & ~n21888;
  assign n21890 = ~n21887 & n21888;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 = n21843 & ~n21891;
  assign n21893 = ~n21843 & n21891;
  assign n21894 = ~n21892 & ~n21893;
  assign n21895 = n19674 & ~n21894;
  assign n21896 = ~n19674 & n21894;
  assign n21897 = ~n21895 & ~n21896;
  assign n21898 = n21839 & ~n21897;
  assign n21899 = ~n21839 & n21897;
  assign n21900 = ~n21898 & ~n21899;
  assign n21901 = n20951 & ~n21900;
  assign n21902 = ~n21832 & ~n21833;
  assign n21903 = ~n21834 & n21902;
  assign n21904 = ~n21835 & n21903;
  assign n4629 = n21901 | ~n21904;
  assign n21906 = ~n15740 & n21299;
  assign n21907 = ~n20664 & n21301;
  assign n21908 = P2_EAX_REG_25_ & ~n20950;
  assign n21909 = ~n19742 & n20957;
  assign n21910 = ~n19674 & ~n21894;
  assign n21911 = n19674 & n21894;
  assign n21912 = ~n21839 & ~n21911;
  assign n21913 = ~n21910 & ~n21912;
  assign n21914 = n21887 & n21888;
  assign n21915 = ~n21887 & ~n21888;
  assign n21916 = ~n21843 & ~n21915;
  assign n21917 = ~n21914 & ~n21916;
  assign n21918 = n21844 & ~n21883;
  assign n21919 = ~P2_INSTQUEUE_REG_6__2_ & n21769;
  assign n21920 = ~P2_INSTQUEUE_REG_14__2_ & ~n21769;
  assign n21921 = ~n21919 & ~n21920;
  assign n21922 = n14149 & n21921;
  assign n21923 = ~P2_INSTQUEUE_REG_2__2_ & n21769;
  assign n21924 = ~P2_INSTQUEUE_REG_10__2_ & ~n21769;
  assign n21925 = ~n21923 & ~n21924;
  assign n21926 = n14155 & n21925;
  assign n21927 = ~P2_INSTQUEUE_REG_1__2_ & n21769;
  assign n21928 = ~P2_INSTQUEUE_REG_9__2_ & ~n21769;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = n14161 & n21929;
  assign n21931 = ~P2_INSTQUEUE_REG_3__2_ & n21769;
  assign n21932 = ~P2_INSTQUEUE_REG_11__2_ & ~n21769;
  assign n21933 = ~n21931 & ~n21932;
  assign n21934 = n14167 & n21933;
  assign n21935 = ~n21922 & ~n21926;
  assign n21936 = ~n21930 & n21935;
  assign n21937 = ~n21934 & n21936;
  assign n21938 = ~P2_INSTQUEUE_REG_0__2_ & n21769;
  assign n21939 = ~P2_INSTQUEUE_REG_8__2_ & ~n21769;
  assign n21940 = ~n21938 & ~n21939;
  assign n21941 = n14176 & n21940;
  assign n21942 = ~P2_INSTQUEUE_REG_5__2_ & n21769;
  assign n21943 = ~P2_INSTQUEUE_REG_13__2_ & ~n21769;
  assign n21944 = ~n21942 & ~n21943;
  assign n21945 = n14182 & n21944;
  assign n21946 = ~P2_INSTQUEUE_REG_4__2_ & n21769;
  assign n21947 = ~P2_INSTQUEUE_REG_12__2_ & ~n21769;
  assign n21948 = ~n21946 & ~n21947;
  assign n21949 = n14187 & n21948;
  assign n21950 = ~P2_INSTQUEUE_REG_7__2_ & n21769;
  assign n21951 = ~P2_INSTQUEUE_REG_15__2_ & ~n21769;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = n14193 & n21952;
  assign n21954 = ~n21941 & ~n21945;
  assign n21955 = ~n21949 & n21954;
  assign n21956 = ~n21953 & n21955;
  assign n21957 = n21937 & n21956;
  assign n21958 = n21918 & n21957;
  assign n21959 = ~n21918 & ~n21957;
  assign n21960 = ~n21958 & ~n21959;
  assign n21961 = n15483 & ~n21960;
  assign n21962 = n15007 & ~n21957;
  assign n21963 = n21961 & ~n21962;
  assign n21964 = ~n21961 & n21962;
  assign n21965 = ~n21963 & ~n21964;
  assign n21966 = n21917 & ~n21965;
  assign n21967 = ~n21917 & n21965;
  assign n21968 = ~n21966 & ~n21967;
  assign n21969 = n19742 & ~n21968;
  assign n21970 = ~n19742 & n21968;
  assign n21971 = ~n21969 & ~n21970;
  assign n21972 = n21913 & ~n21971;
  assign n21973 = ~n21913 & n21971;
  assign n21974 = ~n21972 & ~n21973;
  assign n21975 = n20951 & ~n21974;
  assign n21976 = ~n21906 & ~n21907;
  assign n21977 = ~n21908 & n21976;
  assign n21978 = ~n21909 & n21977;
  assign n4634 = n21975 | ~n21978;
  assign n21980 = ~n15718 & n21299;
  assign n21981 = ~n20656 & n21301;
  assign n21982 = P2_EAX_REG_26_ & ~n20950;
  assign n21983 = ~n19810 & n20957;
  assign n21984 = ~n19742 & ~n21968;
  assign n21985 = n19742 & n21968;
  assign n21986 = ~n21913 & ~n21985;
  assign n21987 = ~n21984 & ~n21986;
  assign n21988 = n21961 & n21962;
  assign n21989 = ~n21961 & ~n21962;
  assign n21990 = ~n21917 & ~n21989;
  assign n21991 = ~n21988 & ~n21990;
  assign n21992 = n21918 & ~n21957;
  assign n21993 = ~P2_INSTQUEUE_REG_6__3_ & n21769;
  assign n21994 = ~P2_INSTQUEUE_REG_14__3_ & ~n21769;
  assign n21995 = ~n21993 & ~n21994;
  assign n21996 = n14149 & n21995;
  assign n21997 = ~P2_INSTQUEUE_REG_2__3_ & n21769;
  assign n21998 = ~P2_INSTQUEUE_REG_10__3_ & ~n21769;
  assign n21999 = ~n21997 & ~n21998;
  assign n22000 = n14155 & n21999;
  assign n22001 = ~P2_INSTQUEUE_REG_1__3_ & n21769;
  assign n22002 = ~P2_INSTQUEUE_REG_9__3_ & ~n21769;
  assign n22003 = ~n22001 & ~n22002;
  assign n22004 = n14161 & n22003;
  assign n22005 = ~P2_INSTQUEUE_REG_3__3_ & n21769;
  assign n22006 = ~P2_INSTQUEUE_REG_11__3_ & ~n21769;
  assign n22007 = ~n22005 & ~n22006;
  assign n22008 = n14167 & n22007;
  assign n22009 = ~n21996 & ~n22000;
  assign n22010 = ~n22004 & n22009;
  assign n22011 = ~n22008 & n22010;
  assign n22012 = ~P2_INSTQUEUE_REG_0__3_ & n21769;
  assign n22013 = ~P2_INSTQUEUE_REG_8__3_ & ~n21769;
  assign n22014 = ~n22012 & ~n22013;
  assign n22015 = n14176 & n22014;
  assign n22016 = ~P2_INSTQUEUE_REG_5__3_ & n21769;
  assign n22017 = ~P2_INSTQUEUE_REG_13__3_ & ~n21769;
  assign n22018 = ~n22016 & ~n22017;
  assign n22019 = n14182 & n22018;
  assign n22020 = ~P2_INSTQUEUE_REG_4__3_ & n21769;
  assign n22021 = ~P2_INSTQUEUE_REG_12__3_ & ~n21769;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = n14187 & n22022;
  assign n22024 = ~P2_INSTQUEUE_REG_7__3_ & n21769;
  assign n22025 = ~P2_INSTQUEUE_REG_15__3_ & ~n21769;
  assign n22026 = ~n22024 & ~n22025;
  assign n22027 = n14193 & n22026;
  assign n22028 = ~n22015 & ~n22019;
  assign n22029 = ~n22023 & n22028;
  assign n22030 = ~n22027 & n22029;
  assign n22031 = n22011 & n22030;
  assign n22032 = n21992 & n22031;
  assign n22033 = ~n21992 & ~n22031;
  assign n22034 = ~n22032 & ~n22033;
  assign n22035 = n15483 & ~n22034;
  assign n22036 = n15007 & ~n22031;
  assign n22037 = n22035 & ~n22036;
  assign n22038 = ~n22035 & n22036;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = n21991 & ~n22039;
  assign n22041 = ~n21991 & n22039;
  assign n22042 = ~n22040 & ~n22041;
  assign n22043 = n19810 & ~n22042;
  assign n22044 = ~n19810 & n22042;
  assign n22045 = ~n22043 & ~n22044;
  assign n22046 = n21987 & ~n22045;
  assign n22047 = ~n21987 & n22045;
  assign n22048 = ~n22046 & ~n22047;
  assign n22049 = n20951 & ~n22048;
  assign n22050 = ~n21980 & ~n21981;
  assign n22051 = ~n21982 & n22050;
  assign n22052 = ~n21983 & n22051;
  assign n4639 = n22049 | ~n22052;
  assign n22054 = ~n15696 & n21299;
  assign n22055 = ~n20648 & n21301;
  assign n22056 = P2_EAX_REG_27_ & ~n20950;
  assign n22057 = ~n19873 & n20957;
  assign n22058 = ~n19810 & ~n22042;
  assign n22059 = n19810 & n22042;
  assign n22060 = ~n21987 & ~n22059;
  assign n22061 = ~n22058 & ~n22060;
  assign n22062 = n22035 & n22036;
  assign n22063 = ~n22035 & ~n22036;
  assign n22064 = ~n21991 & ~n22063;
  assign n22065 = ~n22062 & ~n22064;
  assign n22066 = n21992 & ~n22031;
  assign n22067 = ~P2_INSTQUEUE_REG_6__4_ & n21769;
  assign n22068 = ~P2_INSTQUEUE_REG_14__4_ & ~n21769;
  assign n22069 = ~n22067 & ~n22068;
  assign n22070 = n14149 & n22069;
  assign n22071 = ~P2_INSTQUEUE_REG_2__4_ & n21769;
  assign n22072 = ~P2_INSTQUEUE_REG_10__4_ & ~n21769;
  assign n22073 = ~n22071 & ~n22072;
  assign n22074 = n14155 & n22073;
  assign n22075 = ~P2_INSTQUEUE_REG_1__4_ & n21769;
  assign n22076 = ~P2_INSTQUEUE_REG_9__4_ & ~n21769;
  assign n22077 = ~n22075 & ~n22076;
  assign n22078 = n14161 & n22077;
  assign n22079 = ~P2_INSTQUEUE_REG_3__4_ & n21769;
  assign n22080 = ~P2_INSTQUEUE_REG_11__4_ & ~n21769;
  assign n22081 = ~n22079 & ~n22080;
  assign n22082 = n14167 & n22081;
  assign n22083 = ~n22070 & ~n22074;
  assign n22084 = ~n22078 & n22083;
  assign n22085 = ~n22082 & n22084;
  assign n22086 = ~P2_INSTQUEUE_REG_0__4_ & n21769;
  assign n22087 = ~P2_INSTQUEUE_REG_8__4_ & ~n21769;
  assign n22088 = ~n22086 & ~n22087;
  assign n22089 = n14176 & n22088;
  assign n22090 = ~P2_INSTQUEUE_REG_5__4_ & n21769;
  assign n22091 = ~P2_INSTQUEUE_REG_13__4_ & ~n21769;
  assign n22092 = ~n22090 & ~n22091;
  assign n22093 = n14182 & n22092;
  assign n22094 = ~P2_INSTQUEUE_REG_4__4_ & n21769;
  assign n22095 = ~P2_INSTQUEUE_REG_12__4_ & ~n21769;
  assign n22096 = ~n22094 & ~n22095;
  assign n22097 = n14187 & n22096;
  assign n22098 = ~P2_INSTQUEUE_REG_7__4_ & n21769;
  assign n22099 = ~P2_INSTQUEUE_REG_15__4_ & ~n21769;
  assign n22100 = ~n22098 & ~n22099;
  assign n22101 = n14193 & n22100;
  assign n22102 = ~n22089 & ~n22093;
  assign n22103 = ~n22097 & n22102;
  assign n22104 = ~n22101 & n22103;
  assign n22105 = n22085 & n22104;
  assign n22106 = n22066 & n22105;
  assign n22107 = ~n22066 & ~n22105;
  assign n22108 = ~n22106 & ~n22107;
  assign n22109 = n15483 & ~n22108;
  assign n22110 = n15007 & ~n22105;
  assign n22111 = n22109 & ~n22110;
  assign n22112 = ~n22109 & n22110;
  assign n22113 = ~n22111 & ~n22112;
  assign n22114 = n22065 & ~n22113;
  assign n22115 = ~n22065 & n22113;
  assign n22116 = ~n22114 & ~n22115;
  assign n22117 = n19873 & ~n22116;
  assign n22118 = ~n19873 & n22116;
  assign n22119 = ~n22117 & ~n22118;
  assign n22120 = n22061 & ~n22119;
  assign n22121 = ~n22061 & n22119;
  assign n22122 = ~n22120 & ~n22121;
  assign n22123 = n20951 & ~n22122;
  assign n22124 = ~n22054 & ~n22055;
  assign n22125 = ~n22056 & n22124;
  assign n22126 = ~n22057 & n22125;
  assign n4644 = n22123 | ~n22126;
  assign n22128 = ~n15674 & n21299;
  assign n22129 = ~n20640 & n21301;
  assign n22130 = P2_EAX_REG_28_ & ~n20950;
  assign n22131 = ~n19942 & n20957;
  assign n22132 = ~n19873 & ~n22116;
  assign n22133 = n19873 & n22116;
  assign n22134 = ~n22061 & ~n22133;
  assign n22135 = ~n22132 & ~n22134;
  assign n22136 = n22109 & n22110;
  assign n22137 = ~n22109 & ~n22110;
  assign n22138 = ~n22065 & ~n22137;
  assign n22139 = ~n22136 & ~n22138;
  assign n22140 = n22066 & ~n22105;
  assign n22141 = ~P2_INSTQUEUE_REG_6__5_ & n21769;
  assign n22142 = ~P2_INSTQUEUE_REG_14__5_ & ~n21769;
  assign n22143 = ~n22141 & ~n22142;
  assign n22144 = n14149 & n22143;
  assign n22145 = ~P2_INSTQUEUE_REG_2__5_ & n21769;
  assign n22146 = ~P2_INSTQUEUE_REG_10__5_ & ~n21769;
  assign n22147 = ~n22145 & ~n22146;
  assign n22148 = n14155 & n22147;
  assign n22149 = ~P2_INSTQUEUE_REG_1__5_ & n21769;
  assign n22150 = ~P2_INSTQUEUE_REG_9__5_ & ~n21769;
  assign n22151 = ~n22149 & ~n22150;
  assign n22152 = n14161 & n22151;
  assign n22153 = ~P2_INSTQUEUE_REG_3__5_ & n21769;
  assign n22154 = ~P2_INSTQUEUE_REG_11__5_ & ~n21769;
  assign n22155 = ~n22153 & ~n22154;
  assign n22156 = n14167 & n22155;
  assign n22157 = ~n22144 & ~n22148;
  assign n22158 = ~n22152 & n22157;
  assign n22159 = ~n22156 & n22158;
  assign n22160 = ~P2_INSTQUEUE_REG_0__5_ & n21769;
  assign n22161 = ~P2_INSTQUEUE_REG_8__5_ & ~n21769;
  assign n22162 = ~n22160 & ~n22161;
  assign n22163 = n14176 & n22162;
  assign n22164 = ~P2_INSTQUEUE_REG_5__5_ & n21769;
  assign n22165 = ~P2_INSTQUEUE_REG_13__5_ & ~n21769;
  assign n22166 = ~n22164 & ~n22165;
  assign n22167 = n14182 & n22166;
  assign n22168 = ~P2_INSTQUEUE_REG_4__5_ & n21769;
  assign n22169 = ~P2_INSTQUEUE_REG_12__5_ & ~n21769;
  assign n22170 = ~n22168 & ~n22169;
  assign n22171 = n14187 & n22170;
  assign n22172 = ~P2_INSTQUEUE_REG_7__5_ & n21769;
  assign n22173 = ~P2_INSTQUEUE_REG_15__5_ & ~n21769;
  assign n22174 = ~n22172 & ~n22173;
  assign n22175 = n14193 & n22174;
  assign n22176 = ~n22163 & ~n22167;
  assign n22177 = ~n22171 & n22176;
  assign n22178 = ~n22175 & n22177;
  assign n22179 = n22159 & n22178;
  assign n22180 = n22140 & n22179;
  assign n22181 = ~n22140 & ~n22179;
  assign n22182 = ~n22180 & ~n22181;
  assign n22183 = n15483 & ~n22182;
  assign n22184 = n15007 & ~n22179;
  assign n22185 = n22183 & ~n22184;
  assign n22186 = ~n22183 & n22184;
  assign n22187 = ~n22185 & ~n22186;
  assign n22188 = n22139 & ~n22187;
  assign n22189 = ~n22139 & n22187;
  assign n22190 = ~n22188 & ~n22189;
  assign n22191 = ~n19942 & n22190;
  assign n22192 = n19942 & ~n22190;
  assign n22193 = ~n22191 & ~n22192;
  assign n22194 = n22135 & ~n22193;
  assign n22195 = ~n22135 & n22193;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = n20951 & ~n22196;
  assign n22198 = ~n22128 & ~n22129;
  assign n22199 = ~n22130 & n22198;
  assign n22200 = ~n22131 & n22199;
  assign n4649 = n22197 | ~n22200;
  assign n22202 = ~n15652 & n21299;
  assign n22203 = ~n20632 & n21301;
  assign n22204 = P2_EAX_REG_29_ & ~n20950;
  assign n22205 = ~n20011 & n20957;
  assign n22206 = n22140 & ~n22179;
  assign n22207 = ~P2_INSTQUEUE_REG_6__6_ & n21769;
  assign n22208 = ~P2_INSTQUEUE_REG_14__6_ & ~n21769;
  assign n22209 = ~n22207 & ~n22208;
  assign n22210 = n14149 & n22209;
  assign n22211 = ~P2_INSTQUEUE_REG_2__6_ & n21769;
  assign n22212 = ~P2_INSTQUEUE_REG_10__6_ & ~n21769;
  assign n22213 = ~n22211 & ~n22212;
  assign n22214 = n14155 & n22213;
  assign n22215 = ~P2_INSTQUEUE_REG_1__6_ & n21769;
  assign n22216 = ~P2_INSTQUEUE_REG_9__6_ & ~n21769;
  assign n22217 = ~n22215 & ~n22216;
  assign n22218 = n14161 & n22217;
  assign n22219 = ~P2_INSTQUEUE_REG_3__6_ & n21769;
  assign n22220 = ~P2_INSTQUEUE_REG_11__6_ & ~n21769;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = n14167 & n22221;
  assign n22223 = ~n22210 & ~n22214;
  assign n22224 = ~n22218 & n22223;
  assign n22225 = ~n22222 & n22224;
  assign n22226 = ~P2_INSTQUEUE_REG_0__6_ & n21769;
  assign n22227 = ~P2_INSTQUEUE_REG_8__6_ & ~n21769;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = n14176 & n22228;
  assign n22230 = ~P2_INSTQUEUE_REG_5__6_ & n21769;
  assign n22231 = ~P2_INSTQUEUE_REG_13__6_ & ~n21769;
  assign n22232 = ~n22230 & ~n22231;
  assign n22233 = n14182 & n22232;
  assign n22234 = ~P2_INSTQUEUE_REG_4__6_ & n21769;
  assign n22235 = ~P2_INSTQUEUE_REG_12__6_ & ~n21769;
  assign n22236 = ~n22234 & ~n22235;
  assign n22237 = n14187 & n22236;
  assign n22238 = ~P2_INSTQUEUE_REG_7__6_ & n21769;
  assign n22239 = ~P2_INSTQUEUE_REG_15__6_ & ~n21769;
  assign n22240 = ~n22238 & ~n22239;
  assign n22241 = n14193 & n22240;
  assign n22242 = ~n22229 & ~n22233;
  assign n22243 = ~n22237 & n22242;
  assign n22244 = ~n22241 & n22243;
  assign n22245 = n22225 & n22244;
  assign n22246 = n22206 & n22245;
  assign n22247 = ~n22206 & ~n22245;
  assign n22248 = ~n22246 & ~n22247;
  assign n22249 = n15483 & ~n22248;
  assign n22250 = n15007 & ~n22245;
  assign n22251 = n22249 & ~n22250;
  assign n22252 = ~n22249 & n22250;
  assign n22253 = ~n22251 & ~n22252;
  assign n22254 = n22183 & n22184;
  assign n22255 = ~n22183 & ~n22184;
  assign n22256 = ~n22139 & ~n22255;
  assign n22257 = ~n22254 & ~n22256;
  assign n22258 = ~n22253 & n22257;
  assign n22259 = n22253 & ~n22257;
  assign n22260 = ~n22258 & ~n22259;
  assign n22261 = ~n20011 & n22260;
  assign n22262 = n20011 & ~n22260;
  assign n22263 = ~n22261 & ~n22262;
  assign n22264 = ~n19942 & ~n22190;
  assign n22265 = n19942 & n22190;
  assign n22266 = ~n22135 & ~n22265;
  assign n22267 = ~n22264 & ~n22266;
  assign n22268 = ~n22263 & n22267;
  assign n22269 = n22263 & ~n22267;
  assign n22270 = ~n22268 & ~n22269;
  assign n22271 = n20951 & ~n22270;
  assign n22272 = ~n22202 & ~n22203;
  assign n22273 = ~n22204 & n22272;
  assign n22274 = ~n22205 & n22273;
  assign n4654 = n22271 | ~n22274;
  assign n22276 = ~n15630 & n21299;
  assign n22277 = ~n20624 & n21301;
  assign n22278 = P2_EAX_REG_30_ & ~n20950;
  assign n22279 = ~n20075 & n20957;
  assign n22280 = n20011 & n22260;
  assign n22281 = ~n20011 & ~n22260;
  assign n22282 = n22267 & ~n22281;
  assign n22283 = ~n22249 & ~n22250;
  assign n22284 = n22206 & ~n22245;
  assign n22285 = ~P2_INSTQUEUE_REG_6__7_ & n21769;
  assign n22286 = ~P2_INSTQUEUE_REG_14__7_ & ~n21769;
  assign n22287 = ~n22285 & ~n22286;
  assign n22288 = n14149 & n22287;
  assign n22289 = ~P2_INSTQUEUE_REG_2__7_ & n21769;
  assign n22290 = ~P2_INSTQUEUE_REG_10__7_ & ~n21769;
  assign n22291 = ~n22289 & ~n22290;
  assign n22292 = n14155 & n22291;
  assign n22293 = ~P2_INSTQUEUE_REG_1__7_ & n21769;
  assign n22294 = ~P2_INSTQUEUE_REG_9__7_ & ~n21769;
  assign n22295 = ~n22293 & ~n22294;
  assign n22296 = n14161 & n22295;
  assign n22297 = ~P2_INSTQUEUE_REG_3__7_ & n21769;
  assign n22298 = ~P2_INSTQUEUE_REG_11__7_ & ~n21769;
  assign n22299 = ~n22297 & ~n22298;
  assign n22300 = n14167 & n22299;
  assign n22301 = ~n22288 & ~n22292;
  assign n22302 = ~n22296 & n22301;
  assign n22303 = ~n22300 & n22302;
  assign n22304 = ~P2_INSTQUEUE_REG_0__7_ & n21769;
  assign n22305 = ~P2_INSTQUEUE_REG_8__7_ & ~n21769;
  assign n22306 = ~n22304 & ~n22305;
  assign n22307 = n14176 & n22306;
  assign n22308 = ~P2_INSTQUEUE_REG_5__7_ & n21769;
  assign n22309 = ~P2_INSTQUEUE_REG_13__7_ & ~n21769;
  assign n22310 = ~n22308 & ~n22309;
  assign n22311 = n14182 & n22310;
  assign n22312 = ~P2_INSTQUEUE_REG_4__7_ & n21769;
  assign n22313 = ~P2_INSTQUEUE_REG_12__7_ & ~n21769;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = n14187 & n22314;
  assign n22316 = ~P2_INSTQUEUE_REG_7__7_ & n21769;
  assign n22317 = ~P2_INSTQUEUE_REG_15__7_ & ~n21769;
  assign n22318 = ~n22316 & ~n22317;
  assign n22319 = n14193 & n22318;
  assign n22320 = ~n22307 & ~n22311;
  assign n22321 = ~n22315 & n22320;
  assign n22322 = ~n22319 & n22321;
  assign n22323 = n22303 & n22322;
  assign n22324 = n22284 & n22323;
  assign n22325 = ~n22284 & ~n22323;
  assign n22326 = ~n22324 & ~n22325;
  assign n22327 = n15483 & ~n22326;
  assign n22328 = n15007 & ~n22323;
  assign n22329 = n22327 & ~n22328;
  assign n22330 = ~n22327 & n22328;
  assign n22331 = ~n22329 & ~n22330;
  assign n22332 = ~n22283 & ~n22331;
  assign n22333 = n22249 & n22250;
  assign n22334 = n22257 & ~n22333;
  assign n22335 = n22332 & ~n22334;
  assign n22336 = n22331 & ~n22333;
  assign n22337 = ~n22257 & ~n22283;
  assign n22338 = n22336 & ~n22337;
  assign n22339 = ~n22335 & ~n22338;
  assign n22340 = ~n20075 & ~n22339;
  assign n22341 = n20075 & n22339;
  assign n22342 = ~n22340 & ~n22341;
  assign n22343 = ~n22280 & ~n22282;
  assign n22344 = ~n22342 & n22343;
  assign n22345 = ~n22267 & ~n22280;
  assign n22346 = ~n22281 & ~n22345;
  assign n22347 = n22342 & n22346;
  assign n22348 = ~n22344 & ~n22347;
  assign n22349 = n20951 & n22348;
  assign n22350 = ~n22276 & ~n22277;
  assign n22351 = ~n22278 & n22350;
  assign n22352 = ~n22279 & n22351;
  assign n4659 = n22349 | ~n22352;
  assign n22354 = P2_EAX_REG_31_ & ~n20950;
  assign n22355 = ~n15608 & n21299;
  assign n22356 = n20151 & n20957;
  assign n22357 = ~n22354 & ~n22355;
  assign n4664 = n22356 | ~n22357;
  assign n22359 = ~n14962 & ~n15181;
  assign n22360 = n15432 & ~n22359;
  assign n22361 = n14286 & n22360;
  assign n22362 = ~n15277 & n22361;
  assign n22363 = ~n14286 & n22360;
  assign n22364 = ~n15513 & n22363;
  assign n22365 = P2_EBX_REG_0_ & ~n22360;
  assign n22366 = ~n22362 & ~n22364;
  assign n4669 = n22365 | ~n22366;
  assign n22368 = ~n15263 & n22361;
  assign n22369 = ~n15510 & n22363;
  assign n22370 = P2_EBX_REG_1_ & ~n22360;
  assign n22371 = ~n22368 & ~n22369;
  assign n4674 = n22370 | ~n22371;
  assign n22373 = ~n15216 & n22361;
  assign n22374 = n15539 & n22363;
  assign n22375 = P2_EBX_REG_2_ & ~n22360;
  assign n22376 = ~n22373 & ~n22374;
  assign n4679 = n22375 | ~n22376;
  assign n22378 = ~n15147 & n22361;
  assign n22379 = ~n15557 & n22363;
  assign n22380 = P2_EBX_REG_3_ & ~n22360;
  assign n22381 = ~n22378 & ~n22379;
  assign n4684 = n22380 | ~n22381;
  assign n22383 = n17863 & n22361;
  assign n22384 = ~n21028 & n22363;
  assign n22385 = P2_EBX_REG_4_ & ~n22360;
  assign n22386 = ~n22383 & ~n22384;
  assign n4689 = n22385 | ~n22386;
  assign n22388 = ~n17979 & n22361;
  assign n22389 = ~n21053 & n22363;
  assign n22390 = P2_EBX_REG_5_ & ~n22360;
  assign n22391 = ~n22388 & ~n22389;
  assign n4694 = n22390 | ~n22391;
  assign n22393 = ~n18099 & n22361;
  assign n22394 = ~n21074 & n22363;
  assign n22395 = P2_EBX_REG_6_ & ~n22360;
  assign n22396 = ~n22393 & ~n22394;
  assign n4699 = n22395 | ~n22396;
  assign n22398 = ~n18225 & n22361;
  assign n22399 = ~n21101 & n22363;
  assign n22400 = P2_EBX_REG_7_ & ~n22360;
  assign n22401 = ~n22398 & ~n22399;
  assign n4704 = n22400 | ~n22401;
  assign n22403 = ~n18311 & n22361;
  assign n22404 = P2_EBX_REG_8_ & ~n22360;
  assign n22405 = ~n21126 & n22363;
  assign n22406 = ~n22403 & ~n22404;
  assign n4709 = n22405 | ~n22406;
  assign n22408 = ~n18442 & n22361;
  assign n22409 = P2_EBX_REG_9_ & ~n22360;
  assign n22410 = ~n21148 & n22363;
  assign n22411 = ~n22408 & ~n22409;
  assign n4714 = n22410 | ~n22411;
  assign n22413 = ~n18541 & n22361;
  assign n22414 = P2_EBX_REG_10_ & ~n22360;
  assign n22415 = ~n21168 & n22363;
  assign n22416 = ~n22413 & ~n22414;
  assign n4719 = n22415 | ~n22416;
  assign n22418 = ~n18638 & n22361;
  assign n22419 = P2_EBX_REG_11_ & ~n22360;
  assign n22420 = ~n21191 & n22363;
  assign n22421 = ~n22418 & ~n22419;
  assign n4724 = n22420 | ~n22421;
  assign n22423 = ~n18736 & n22361;
  assign n22424 = P2_EBX_REG_12_ & ~n22360;
  assign n22425 = ~n21216 & n22363;
  assign n22426 = ~n22423 & ~n22424;
  assign n4729 = n22425 | ~n22426;
  assign n22428 = ~n18837 & n22361;
  assign n22429 = P2_EBX_REG_13_ & ~n22360;
  assign n22430 = ~n21238 & n22363;
  assign n22431 = ~n22428 & ~n22429;
  assign n4734 = n22430 | ~n22431;
  assign n22433 = ~n18936 & n22361;
  assign n22434 = P2_EBX_REG_14_ & ~n22360;
  assign n22435 = ~n21259 & n22363;
  assign n22436 = ~n22433 & ~n22434;
  assign n4739 = n22435 | ~n22436;
  assign n22438 = ~n19032 & n22361;
  assign n22439 = P2_EBX_REG_15_ & ~n22360;
  assign n22440 = ~n21282 & n22363;
  assign n22441 = ~n22438 & ~n22439;
  assign n4744 = n22440 | ~n22441;
  assign n22443 = ~n19135 & n22361;
  assign n22444 = P2_EBX_REG_16_ & ~n22360;
  assign n22445 = ~n21372 & n22363;
  assign n22446 = ~n22443 & ~n22444;
  assign n4749 = n22445 | ~n22446;
  assign n22448 = ~n19198 & n22361;
  assign n22449 = P2_EBX_REG_17_ & ~n22360;
  assign n22450 = ~n21429 & n22363;
  assign n22451 = ~n22448 & ~n22449;
  assign n4754 = n22450 | ~n22451;
  assign n22453 = ~n19266 & n22361;
  assign n22454 = P2_EBX_REG_18_ & ~n22360;
  assign n22455 = ~n21486 & n22363;
  assign n22456 = ~n22453 & ~n22454;
  assign n4759 = n22455 | ~n22456;
  assign n22458 = ~n19334 & n22361;
  assign n22459 = P2_EBX_REG_19_ & ~n22360;
  assign n22460 = ~n21543 & n22363;
  assign n22461 = ~n22458 & ~n22459;
  assign n4764 = n22460 | ~n22461;
  assign n22463 = ~n19401 & n22361;
  assign n22464 = P2_EBX_REG_20_ & ~n22360;
  assign n22465 = ~n21600 & n22363;
  assign n22466 = ~n22463 & ~n22464;
  assign n4769 = n22465 | ~n22466;
  assign n22468 = ~n19467 & n22361;
  assign n22469 = P2_EBX_REG_21_ & ~n22360;
  assign n22470 = ~n21657 & n22363;
  assign n22471 = ~n22468 & ~n22469;
  assign n4774 = n22470 | ~n22471;
  assign n22473 = ~n19533 & n22361;
  assign n22474 = P2_EBX_REG_22_ & ~n22360;
  assign n22475 = ~n21714 & n22363;
  assign n22476 = ~n22473 & ~n22474;
  assign n4779 = n22475 | ~n22476;
  assign n22478 = ~n19602 & n22361;
  assign n22479 = P2_EBX_REG_23_ & ~n22360;
  assign n22480 = ~n21820 & n22363;
  assign n22481 = ~n22478 & ~n22479;
  assign n4784 = n22480 | ~n22481;
  assign n22483 = ~n19664 & n22361;
  assign n22484 = P2_EBX_REG_24_ & ~n22360;
  assign n22485 = ~n21894 & n22363;
  assign n22486 = ~n22483 & ~n22484;
  assign n4789 = n22485 | ~n22486;
  assign n22488 = ~n19732 & n22361;
  assign n22489 = P2_EBX_REG_25_ & ~n22360;
  assign n22490 = ~n21968 & n22363;
  assign n22491 = ~n22488 & ~n22489;
  assign n4794 = n22490 | ~n22491;
  assign n22493 = ~n19800 & n22361;
  assign n22494 = P2_EBX_REG_26_ & ~n22360;
  assign n22495 = ~n22042 & n22363;
  assign n22496 = ~n22493 & ~n22494;
  assign n4799 = n22495 | ~n22496;
  assign n22498 = ~n19863 & n22361;
  assign n22499 = P2_EBX_REG_27_ & ~n22360;
  assign n22500 = ~n22116 & n22363;
  assign n22501 = ~n22498 & ~n22499;
  assign n4804 = n22500 | ~n22501;
  assign n22503 = ~n19932 & n22361;
  assign n22504 = P2_EBX_REG_28_ & ~n22360;
  assign n22505 = ~n22190 & n22363;
  assign n22506 = ~n22503 & ~n22504;
  assign n4809 = n22505 | ~n22506;
  assign n22508 = ~n20001 & n22361;
  assign n22509 = P2_EBX_REG_29_ & ~n22360;
  assign n22510 = ~n22260 & n22363;
  assign n22511 = ~n22508 & ~n22509;
  assign n4814 = n22510 | ~n22511;
  assign n22513 = ~n20063 & n22361;
  assign n22514 = P2_EBX_REG_30_ & ~n22360;
  assign n22515 = n22339 & n22363;
  assign n22516 = ~n22513 & ~n22514;
  assign n4819 = n22515 | ~n22516;
  assign n22518 = P2_EBX_REG_31_ & ~n22360;
  assign n22519 = ~n20138 & n22361;
  assign n4824 = n22518 | n22519;
  assign n22521 = ~n15442 & ~n15455;
  assign n22522 = ~n17387 & n22521;
  assign n22523 = ~n14949 & n15178;
  assign n22524 = n14548 & ~n15396;
  assign n22525 = ~n22523 & ~n22524;
  assign n22526 = n15432 & ~n22525;
  assign n22527 = n22522 & ~n22526;
  assign n22528 = P2_STATE2_REG_2_ & ~n22527;
  assign n22529 = n14244 & n22528;
  assign n22530 = ~n15413 & n22529;
  assign n22531 = ~P2_EBX_REG_31_ & n22530;
  assign n22532 = n14239 & n22528;
  assign n22533 = ~n14144 & n22532;
  assign n22534 = n14144 & n22532;
  assign n22535 = ~n15413 & n22534;
  assign n22536 = ~n22531 & ~n22533;
  assign n22537 = ~n22535 & n22536;
  assign n22538 = P2_EBX_REG_0_ & ~n22537;
  assign n22539 = n15413 & n22534;
  assign n22540 = ~n17339 & n22539;
  assign n22541 = P2_EBX_REG_31_ & n22530;
  assign n22542 = ~n17451 & n22541;
  assign n22543 = n15413 & n22529;
  assign n22544 = ~n15277 & n22543;
  assign n22545 = n14199 & n22528;
  assign n22546 = ~n15513 & n22545;
  assign n22547 = ~n22544 & ~n22546;
  assign n22548 = ~n22540 & ~n22542;
  assign n22549 = n22547 & n22548;
  assign n22550 = P2_STATE2_REG_1_ & ~n22527;
  assign n22551 = ~n15338 & n22550;
  assign n22552 = ~n15341 & n22551;
  assign n22553 = P2_REIP_REG_0_ & n22527;
  assign n22554 = P2_STATE2_REG_3_ & ~n22527;
  assign n22555 = P2_PHYADDRPOINTER_REG_0_ & n22554;
  assign n22556 = ~n22553 & ~n22555;
  assign n22557 = n15338 & n22550;
  assign n22558 = P2_PHYADDRPOINTER_REG_0_ & n22557;
  assign n22559 = n22556 & ~n22558;
  assign n22560 = ~n22538 & n22549;
  assign n22561 = ~n22552 & n22560;
  assign n4829 = ~n22559 | ~n22561;
  assign n22563 = P2_EBX_REG_1_ & ~n22537;
  assign n22564 = ~n17326 & n22539;
  assign n22565 = ~n17553 & n22541;
  assign n22566 = ~n15263 & n22543;
  assign n22567 = ~n15510 & n22545;
  assign n22568 = ~n22566 & ~n22567;
  assign n22569 = ~n22564 & ~n22565;
  assign n22570 = n22568 & n22569;
  assign n22571 = ~n15356 & n22551;
  assign n22572 = P2_REIP_REG_1_ & n22527;
  assign n22573 = P2_PHYADDRPOINTER_REG_1_ & n22554;
  assign n22574 = ~n22572 & ~n22573;
  assign n22575 = ~P2_PHYADDRPOINTER_REG_1_ & n22557;
  assign n22576 = n22574 & ~n22575;
  assign n22577 = ~n22563 & n22570;
  assign n22578 = ~n22571 & n22577;
  assign n4834 = ~n22576 | ~n22578;
  assign n22580 = P2_EBX_REG_2_ & ~n22537;
  assign n22581 = ~n17306 & n22539;
  assign n22582 = n17644 & n22541;
  assign n22583 = ~n15216 & n22543;
  assign n22584 = n15539 & n22545;
  assign n22585 = ~n22583 & ~n22584;
  assign n22586 = ~n22581 & ~n22582;
  assign n22587 = n22585 & n22586;
  assign n22588 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_2_;
  assign n22589 = ~P2_STATE2_REG_0_ & ~n20198;
  assign n22590 = ~n22588 & ~n22589;
  assign n22591 = n15341 & n15353;
  assign n22592 = ~n22590 & ~n22591;
  assign n22593 = n22590 & n22591;
  assign n22594 = ~n22592 & ~n22593;
  assign n22595 = n22551 & n22594;
  assign n22596 = P2_REIP_REG_2_ & n22527;
  assign n22597 = P2_PHYADDRPOINTER_REG_2_ & n22554;
  assign n22598 = ~n22596 & ~n22597;
  assign n22599 = ~n20198 & n22557;
  assign n22600 = n22598 & ~n22599;
  assign n22601 = ~n22580 & n22587;
  assign n22602 = ~n22595 & n22601;
  assign n4839 = ~n22600 | ~n22602;
  assign n22604 = P2_EBX_REG_3_ & ~n22537;
  assign n22605 = ~n17289 & n22539;
  assign n22606 = n17736 & n22541;
  assign n22607 = ~n15147 & n22543;
  assign n22608 = ~n15557 & n22545;
  assign n22609 = ~n22607 & ~n22608;
  assign n22610 = ~n22605 & ~n22606;
  assign n22611 = n22609 & n22610;
  assign n22612 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_3_;
  assign n22613 = ~P2_STATE2_REG_0_ & ~n20213;
  assign n22614 = ~n22612 & ~n22613;
  assign n22615 = n22593 & n22614;
  assign n22616 = ~n22593 & ~n22614;
  assign n22617 = ~n22615 & ~n22616;
  assign n22618 = n22551 & n22617;
  assign n22619 = P2_REIP_REG_3_ & n22527;
  assign n22620 = P2_PHYADDRPOINTER_REG_3_ & n22554;
  assign n22621 = ~n22619 & ~n22620;
  assign n22622 = ~n20213 & n22557;
  assign n22623 = n22621 & ~n22622;
  assign n22624 = ~n22604 & n22611;
  assign n22625 = ~n22618 & n22624;
  assign n4844 = ~n22623 | ~n22625;
  assign n22627 = ~n21028 & n22545;
  assign n22628 = P2_EBX_REG_4_ & ~n22537;
  assign n22629 = n17826 & n22541;
  assign n22630 = n17386 & ~n22527;
  assign n22631 = ~n17880 & n22539;
  assign n22632 = ~n22629 & ~n22630;
  assign n22633 = ~n22631 & n22632;
  assign n22634 = n17863 & n22543;
  assign n22635 = ~n20227 & n22557;
  assign n22636 = ~n22627 & ~n22628;
  assign n22637 = n22633 & n22636;
  assign n22638 = ~n22634 & n22637;
  assign n22639 = ~n22635 & n22638;
  assign n22640 = P2_REIP_REG_4_ & n22527;
  assign n22641 = P2_PHYADDRPOINTER_REG_4_ & n22554;
  assign n22642 = ~n22640 & ~n22641;
  assign n22643 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_4_;
  assign n22644 = ~P2_STATE2_REG_0_ & ~n20227;
  assign n22645 = ~n22643 & ~n22644;
  assign n22646 = ~n22615 & ~n22645;
  assign n22647 = n22614 & n22645;
  assign n22648 = n22593 & n22647;
  assign n22649 = ~n22646 & ~n22648;
  assign n22650 = n22551 & n22649;
  assign n22651 = n22642 & ~n22650;
  assign n4849 = ~n22639 | ~n22651;
  assign n22653 = ~n21053 & n22545;
  assign n22654 = P2_EBX_REG_5_ & ~n22537;
  assign n22655 = n17945 & n22541;
  assign n22656 = ~n17996 & n22539;
  assign n22657 = ~n22630 & ~n22655;
  assign n22658 = ~n22656 & n22657;
  assign n22659 = ~n17979 & n22543;
  assign n22660 = ~n20241 & n22557;
  assign n22661 = ~n22653 & ~n22654;
  assign n22662 = n22658 & n22661;
  assign n22663 = ~n22659 & n22662;
  assign n22664 = ~n22660 & n22663;
  assign n22665 = P2_REIP_REG_5_ & n22527;
  assign n22666 = P2_PHYADDRPOINTER_REG_5_ & n22554;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_5_;
  assign n22669 = ~P2_STATE2_REG_0_ & ~n20241;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = n22648 & n22670;
  assign n22672 = ~n22648 & ~n22670;
  assign n22673 = ~n22671 & ~n22672;
  assign n22674 = n22551 & n22673;
  assign n22675 = n22667 & ~n22674;
  assign n4854 = ~n22664 | ~n22675;
  assign n22677 = ~n18099 & n22543;
  assign n22678 = P2_EBX_REG_6_ & ~n22537;
  assign n22679 = n18064 & n22541;
  assign n22680 = ~n18116 & n22539;
  assign n22681 = ~n22630 & ~n22679;
  assign n22682 = ~n22680 & n22681;
  assign n22683 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_6_;
  assign n22684 = ~P2_STATE2_REG_0_ & ~n20255;
  assign n22685 = ~n22683 & ~n22684;
  assign n22686 = ~n22671 & ~n22685;
  assign n22687 = n22671 & n22685;
  assign n22688 = ~n22686 & ~n22687;
  assign n22689 = n22551 & n22688;
  assign n22690 = P2_REIP_REG_6_ & n22527;
  assign n22691 = P2_PHYADDRPOINTER_REG_6_ & n22554;
  assign n22692 = ~n22690 & ~n22691;
  assign n22693 = ~n20255 & n22557;
  assign n22694 = n22692 & ~n22693;
  assign n22695 = ~n22677 & ~n22678;
  assign n22696 = n22682 & n22695;
  assign n22697 = ~n22689 & n22696;
  assign n4859 = ~n22694 | ~n22697;
  assign n22699 = ~n18225 & n22543;
  assign n22700 = P2_EBX_REG_7_ & ~n22537;
  assign n22701 = n18190 & n22541;
  assign n22702 = ~n18242 & n22539;
  assign n22703 = ~n22630 & ~n22701;
  assign n22704 = ~n22702 & n22703;
  assign n22705 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_7_;
  assign n22706 = ~P2_STATE2_REG_0_ & ~n20269;
  assign n22707 = ~n22705 & ~n22706;
  assign n22708 = n22687 & n22707;
  assign n22709 = ~n22687 & ~n22707;
  assign n22710 = ~n22708 & ~n22709;
  assign n22711 = n22551 & n22710;
  assign n22712 = P2_REIP_REG_7_ & n22527;
  assign n22713 = P2_PHYADDRPOINTER_REG_7_ & n22554;
  assign n22714 = ~n22712 & ~n22713;
  assign n22715 = ~n20269 & n22557;
  assign n22716 = n22714 & ~n22715;
  assign n22717 = ~n22699 & ~n22700;
  assign n22718 = n22704 & n22717;
  assign n22719 = ~n22711 & n22718;
  assign n4864 = ~n22716 | ~n22719;
  assign n22721 = ~n18311 & n22543;
  assign n22722 = P2_EBX_REG_8_ & ~n22537;
  assign n22723 = n18276 & n22541;
  assign n22724 = ~n18381 & n22539;
  assign n22725 = ~n22630 & ~n22723;
  assign n22726 = ~n22724 & n22725;
  assign n22727 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_8_;
  assign n22728 = ~P2_STATE2_REG_0_ & ~n20283;
  assign n22729 = ~n22727 & ~n22728;
  assign n22730 = ~n22708 & ~n22729;
  assign n22731 = n22708 & n22729;
  assign n22732 = ~n22730 & ~n22731;
  assign n22733 = n22551 & n22732;
  assign n22734 = P2_REIP_REG_8_ & n22527;
  assign n22735 = P2_PHYADDRPOINTER_REG_8_ & n22554;
  assign n22736 = ~n22734 & ~n22735;
  assign n22737 = ~n20283 & n22557;
  assign n22738 = n22736 & ~n22737;
  assign n22739 = ~n22721 & ~n22722;
  assign n22740 = n22726 & n22739;
  assign n22741 = ~n22733 & n22740;
  assign n4869 = ~n22738 | ~n22741;
  assign n22743 = ~n18442 & n22543;
  assign n22744 = P2_EBX_REG_9_ & ~n22537;
  assign n22745 = n18409 & n22541;
  assign n22746 = ~n18485 & n22539;
  assign n22747 = ~n22630 & ~n22745;
  assign n22748 = ~n22746 & n22747;
  assign n22749 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_9_;
  assign n22750 = ~P2_STATE2_REG_0_ & ~n20297;
  assign n22751 = ~n22749 & ~n22750;
  assign n22752 = n22731 & n22751;
  assign n22753 = ~n22731 & ~n22751;
  assign n22754 = ~n22752 & ~n22753;
  assign n22755 = n22551 & n22754;
  assign n22756 = P2_REIP_REG_9_ & n22527;
  assign n22757 = P2_PHYADDRPOINTER_REG_9_ & n22554;
  assign n22758 = ~n22756 & ~n22757;
  assign n22759 = ~n20297 & n22557;
  assign n22760 = n22758 & ~n22759;
  assign n22761 = ~n22743 & ~n22744;
  assign n22762 = n22748 & n22761;
  assign n22763 = ~n22755 & n22762;
  assign n4874 = ~n22760 | ~n22763;
  assign n22765 = ~n18541 & n22543;
  assign n22766 = P2_EBX_REG_10_ & ~n22537;
  assign n22767 = n18508 & n22541;
  assign n22768 = ~n18584 & n22539;
  assign n22769 = ~n22630 & ~n22767;
  assign n22770 = ~n22768 & n22769;
  assign n22771 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_10_;
  assign n22772 = ~P2_STATE2_REG_0_ & ~n20311;
  assign n22773 = ~n22771 & ~n22772;
  assign n22774 = ~n22752 & ~n22773;
  assign n22775 = n22752 & n22773;
  assign n22776 = ~n22774 & ~n22775;
  assign n22777 = n22551 & n22776;
  assign n22778 = P2_REIP_REG_10_ & n22527;
  assign n22779 = P2_PHYADDRPOINTER_REG_10_ & n22554;
  assign n22780 = ~n22778 & ~n22779;
  assign n22781 = ~n20311 & n22557;
  assign n22782 = n22780 & ~n22781;
  assign n22783 = ~n22765 & ~n22766;
  assign n22784 = n22770 & n22783;
  assign n22785 = ~n22777 & n22784;
  assign n4879 = ~n22782 | ~n22785;
  assign n22787 = ~n18638 & n22543;
  assign n22788 = P2_EBX_REG_11_ & ~n22537;
  assign n22789 = n18605 & n22541;
  assign n22790 = ~n18681 & n22539;
  assign n22791 = ~n22630 & ~n22789;
  assign n22792 = ~n22790 & n22791;
  assign n22793 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_11_;
  assign n22794 = ~P2_STATE2_REG_0_ & ~n20325;
  assign n22795 = ~n22793 & ~n22794;
  assign n22796 = n22775 & n22795;
  assign n22797 = ~n22775 & ~n22795;
  assign n22798 = ~n22796 & ~n22797;
  assign n22799 = n22551 & n22798;
  assign n22800 = P2_REIP_REG_11_ & n22527;
  assign n22801 = P2_PHYADDRPOINTER_REG_11_ & n22554;
  assign n22802 = ~n22800 & ~n22801;
  assign n22803 = ~n20325 & n22557;
  assign n22804 = n22802 & ~n22803;
  assign n22805 = ~n22787 & ~n22788;
  assign n22806 = n22792 & n22805;
  assign n22807 = ~n22799 & n22806;
  assign n4884 = ~n22804 | ~n22807;
  assign n22809 = P2_EBX_REG_12_ & ~n22537;
  assign n22810 = n18703 & n22541;
  assign n22811 = ~n18736 & n22543;
  assign n22812 = ~n22630 & ~n22810;
  assign n22813 = ~n22811 & n22812;
  assign n22814 = ~n18779 & n22539;
  assign n22815 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_12_;
  assign n22816 = ~P2_STATE2_REG_0_ & ~n20339;
  assign n22817 = ~n22815 & ~n22816;
  assign n22818 = ~n22796 & ~n22817;
  assign n22819 = n22796 & n22817;
  assign n22820 = ~n22818 & ~n22819;
  assign n22821 = n22551 & n22820;
  assign n22822 = P2_REIP_REG_12_ & n22527;
  assign n22823 = P2_PHYADDRPOINTER_REG_12_ & n22554;
  assign n22824 = ~n22822 & ~n22823;
  assign n22825 = ~n20339 & n22557;
  assign n22826 = n22824 & ~n22825;
  assign n22827 = ~n22809 & n22813;
  assign n22828 = ~n22814 & n22827;
  assign n22829 = ~n22821 & n22828;
  assign n4889 = ~n22826 | ~n22829;
  assign n22831 = P2_EBX_REG_13_ & ~n22537;
  assign n22832 = n18804 & n22541;
  assign n22833 = ~n18837 & n22543;
  assign n22834 = ~n22630 & ~n22832;
  assign n22835 = ~n22833 & n22834;
  assign n22836 = ~n18880 & n22539;
  assign n22837 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_13_;
  assign n22838 = ~P2_STATE2_REG_0_ & ~n20353;
  assign n22839 = ~n22837 & ~n22838;
  assign n22840 = n22819 & n22839;
  assign n22841 = ~n22819 & ~n22839;
  assign n22842 = ~n22840 & ~n22841;
  assign n22843 = n22551 & n22842;
  assign n22844 = P2_REIP_REG_13_ & n22527;
  assign n22845 = P2_PHYADDRPOINTER_REG_13_ & n22554;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = ~n20353 & n22557;
  assign n22848 = n22846 & ~n22847;
  assign n22849 = ~n22831 & n22835;
  assign n22850 = ~n22836 & n22849;
  assign n22851 = ~n22843 & n22850;
  assign n4894 = ~n22848 | ~n22851;
  assign n22853 = P2_EBX_REG_14_ & ~n22537;
  assign n22854 = n18903 & n22541;
  assign n22855 = ~n18936 & n22543;
  assign n22856 = ~n22630 & ~n22854;
  assign n22857 = ~n22855 & n22856;
  assign n22858 = ~n18979 & n22539;
  assign n22859 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_14_;
  assign n22860 = ~P2_STATE2_REG_0_ & ~n20367;
  assign n22861 = ~n22859 & ~n22860;
  assign n22862 = ~n22840 & ~n22861;
  assign n22863 = n22840 & n22861;
  assign n22864 = ~n22862 & ~n22863;
  assign n22865 = n22551 & n22864;
  assign n22866 = P2_REIP_REG_14_ & n22527;
  assign n22867 = P2_PHYADDRPOINTER_REG_14_ & n22554;
  assign n22868 = ~n22866 & ~n22867;
  assign n22869 = ~n20367 & n22557;
  assign n22870 = n22868 & ~n22869;
  assign n22871 = ~n22853 & n22857;
  assign n22872 = ~n22858 & n22871;
  assign n22873 = ~n22865 & n22872;
  assign n4899 = ~n22870 | ~n22873;
  assign n22875 = n18999 & n22541;
  assign n22876 = ~n22630 & ~n22875;
  assign n22877 = P2_EBX_REG_15_ & ~n22537;
  assign n22878 = ~n19032 & n22543;
  assign n22879 = ~n19075 & n22539;
  assign n22880 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_15_;
  assign n22881 = ~P2_STATE2_REG_0_ & ~n20381;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = n22863 & n22882;
  assign n22884 = ~n22863 & ~n22882;
  assign n22885 = ~n22883 & ~n22884;
  assign n22886 = n22551 & n22885;
  assign n22887 = n22876 & ~n22877;
  assign n22888 = ~n22878 & n22887;
  assign n22889 = ~n22879 & n22888;
  assign n22890 = ~n22886 & n22889;
  assign n22891 = P2_REIP_REG_15_ & n22527;
  assign n22892 = P2_PHYADDRPOINTER_REG_15_ & n22554;
  assign n22893 = ~n22891 & ~n22892;
  assign n22894 = ~n20381 & n22557;
  assign n22895 = n22893 & ~n22894;
  assign n4904 = ~n22890 | ~n22895;
  assign n22897 = n19102 & n22541;
  assign n22898 = ~n22630 & ~n22897;
  assign n22899 = P2_EBX_REG_16_ & ~n22537;
  assign n22900 = ~n19135 & n22543;
  assign n22901 = ~n19145 & n22539;
  assign n22902 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_16_;
  assign n22903 = ~P2_STATE2_REG_0_ & ~n20395;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~n22883 & ~n22904;
  assign n22906 = n22883 & n22904;
  assign n22907 = ~n22905 & ~n22906;
  assign n22908 = n22551 & n22907;
  assign n22909 = n22898 & ~n22899;
  assign n22910 = ~n22900 & n22909;
  assign n22911 = ~n22901 & n22910;
  assign n22912 = ~n22908 & n22911;
  assign n22913 = P2_REIP_REG_16_ & n22527;
  assign n22914 = P2_PHYADDRPOINTER_REG_16_ & n22554;
  assign n22915 = ~n22913 & ~n22914;
  assign n22916 = ~n20395 & n22557;
  assign n22917 = n22915 & ~n22916;
  assign n4909 = ~n22912 | ~n22917;
  assign n22919 = n19165 & n22541;
  assign n22920 = ~n22630 & ~n22919;
  assign n22921 = P2_EBX_REG_17_ & ~n22537;
  assign n22922 = ~n19198 & n22543;
  assign n22923 = ~n19208 & n22539;
  assign n22924 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_17_;
  assign n22925 = ~P2_STATE2_REG_0_ & ~n20409;
  assign n22926 = ~n22924 & ~n22925;
  assign n22927 = n22906 & n22926;
  assign n22928 = ~n22906 & ~n22926;
  assign n22929 = ~n22927 & ~n22928;
  assign n22930 = n22551 & n22929;
  assign n22931 = n22920 & ~n22921;
  assign n22932 = ~n22922 & n22931;
  assign n22933 = ~n22923 & n22932;
  assign n22934 = ~n22930 & n22933;
  assign n22935 = P2_REIP_REG_17_ & n22527;
  assign n22936 = P2_PHYADDRPOINTER_REG_17_ & n22554;
  assign n22937 = ~n22935 & ~n22936;
  assign n22938 = ~n20409 & n22557;
  assign n22939 = n22937 & ~n22938;
  assign n4914 = ~n22934 | ~n22939;
  assign n22941 = n19233 & n22541;
  assign n22942 = ~n22630 & ~n22941;
  assign n22943 = P2_EBX_REG_18_ & ~n22537;
  assign n22944 = ~n19266 & n22543;
  assign n22945 = ~n19276 & n22539;
  assign n22946 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_18_;
  assign n22947 = ~P2_STATE2_REG_0_ & ~n20423;
  assign n22948 = ~n22946 & ~n22947;
  assign n22949 = ~n22927 & ~n22948;
  assign n22950 = n22927 & n22948;
  assign n22951 = ~n22949 & ~n22950;
  assign n22952 = n22551 & n22951;
  assign n22953 = n22942 & ~n22943;
  assign n22954 = ~n22944 & n22953;
  assign n22955 = ~n22945 & n22954;
  assign n22956 = ~n22952 & n22955;
  assign n22957 = P2_REIP_REG_18_ & n22527;
  assign n22958 = P2_PHYADDRPOINTER_REG_18_ & n22554;
  assign n22959 = ~n22957 & ~n22958;
  assign n22960 = ~n20423 & n22557;
  assign n22961 = n22959 & ~n22960;
  assign n4919 = ~n22956 | ~n22961;
  assign n22963 = n19301 & n22541;
  assign n22964 = ~n22630 & ~n22963;
  assign n22965 = P2_EBX_REG_19_ & ~n22537;
  assign n22966 = ~n19334 & n22543;
  assign n22967 = ~n19344 & n22539;
  assign n22968 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_19_;
  assign n22969 = ~P2_STATE2_REG_0_ & ~n20437;
  assign n22970 = ~n22968 & ~n22969;
  assign n22971 = n22950 & n22970;
  assign n22972 = ~n22950 & ~n22970;
  assign n22973 = ~n22971 & ~n22972;
  assign n22974 = n22551 & n22973;
  assign n22975 = n22964 & ~n22965;
  assign n22976 = ~n22966 & n22975;
  assign n22977 = ~n22967 & n22976;
  assign n22978 = ~n22974 & n22977;
  assign n22979 = P2_REIP_REG_19_ & n22527;
  assign n22980 = P2_PHYADDRPOINTER_REG_19_ & n22554;
  assign n22981 = ~n22979 & ~n22980;
  assign n22982 = ~n20437 & n22557;
  assign n22983 = n22981 & ~n22982;
  assign n4924 = ~n22978 | ~n22983;
  assign n22985 = n19368 & n22541;
  assign n22986 = P2_EBX_REG_20_ & ~n22537;
  assign n22987 = ~n19401 & n22543;
  assign n22988 = ~n19411 & n22539;
  assign n22989 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_20_;
  assign n22990 = ~P2_STATE2_REG_0_ & ~n20451;
  assign n22991 = ~n22989 & ~n22990;
  assign n22992 = ~n22971 & ~n22991;
  assign n22993 = n22971 & n22991;
  assign n22994 = ~n22992 & ~n22993;
  assign n22995 = n22551 & n22994;
  assign n22996 = ~n22985 & ~n22986;
  assign n22997 = ~n22987 & n22996;
  assign n22998 = ~n22988 & n22997;
  assign n22999 = ~n22995 & n22998;
  assign n23000 = P2_REIP_REG_20_ & n22527;
  assign n23001 = P2_PHYADDRPOINTER_REG_20_ & n22554;
  assign n23002 = ~n23000 & ~n23001;
  assign n23003 = ~n20451 & n22557;
  assign n23004 = n23002 & ~n23003;
  assign n4929 = ~n22999 | ~n23004;
  assign n23006 = n19434 & n22541;
  assign n23007 = P2_EBX_REG_21_ & ~n22537;
  assign n23008 = ~n19467 & n22543;
  assign n23009 = ~n19477 & n22539;
  assign n23010 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_21_;
  assign n23011 = ~P2_STATE2_REG_0_ & ~n20465;
  assign n23012 = ~n23010 & ~n23011;
  assign n23013 = n22993 & n23012;
  assign n23014 = ~n22993 & ~n23012;
  assign n23015 = ~n23013 & ~n23014;
  assign n23016 = n22551 & n23015;
  assign n23017 = ~n23006 & ~n23007;
  assign n23018 = ~n23008 & n23017;
  assign n23019 = ~n23009 & n23018;
  assign n23020 = ~n23016 & n23019;
  assign n23021 = P2_REIP_REG_21_ & n22527;
  assign n23022 = P2_PHYADDRPOINTER_REG_21_ & n22554;
  assign n23023 = ~n23021 & ~n23022;
  assign n23024 = ~n20465 & n22557;
  assign n23025 = n23023 & ~n23024;
  assign n4934 = ~n23020 | ~n23025;
  assign n23027 = n19500 & n22541;
  assign n23028 = P2_EBX_REG_22_ & ~n22537;
  assign n23029 = ~n19533 & n22543;
  assign n23030 = ~n19543 & n22539;
  assign n23031 = P2_REIP_REG_22_ & n22527;
  assign n23032 = P2_PHYADDRPOINTER_REG_22_ & n22554;
  assign n23033 = ~n23031 & ~n23032;
  assign n23034 = ~n20479 & n22557;
  assign n23035 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_22_;
  assign n23036 = ~P2_STATE2_REG_0_ & ~n20479;
  assign n23037 = ~n23035 & ~n23036;
  assign n23038 = ~n23013 & ~n23037;
  assign n23039 = n23013 & n23037;
  assign n23040 = ~n23038 & ~n23039;
  assign n23041 = n22551 & n23040;
  assign n23042 = n23033 & ~n23034;
  assign n23043 = ~n23041 & n23042;
  assign n23044 = ~n23027 & ~n23028;
  assign n23045 = ~n23029 & n23044;
  assign n23046 = ~n23030 & n23045;
  assign n4939 = ~n23043 | ~n23046;
  assign n23048 = ~n19612 & n22539;
  assign n23049 = n19569 & n22541;
  assign n23050 = P2_EBX_REG_23_ & ~n22537;
  assign n23051 = ~n19602 & n22543;
  assign n23052 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_23_;
  assign n23053 = ~P2_STATE2_REG_0_ & ~n20493;
  assign n23054 = ~n23052 & ~n23053;
  assign n23055 = n23039 & n23054;
  assign n23056 = ~n23039 & ~n23054;
  assign n23057 = ~n23055 & ~n23056;
  assign n23058 = n22551 & n23057;
  assign n23059 = P2_REIP_REG_23_ & n22527;
  assign n23060 = P2_PHYADDRPOINTER_REG_23_ & n22554;
  assign n23061 = ~n23059 & ~n23060;
  assign n23062 = ~n20493 & n22557;
  assign n23063 = n23061 & ~n23062;
  assign n23064 = ~n23049 & ~n23050;
  assign n23065 = ~n23051 & n23064;
  assign n23066 = ~n23058 & n23065;
  assign n23067 = n23063 & n23066;
  assign n4944 = n23048 | ~n23067;
  assign n23069 = ~n19674 & n22539;
  assign n23070 = n19631 & n22541;
  assign n23071 = P2_EBX_REG_24_ & ~n22537;
  assign n23072 = ~n19664 & n22543;
  assign n23073 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_24_;
  assign n23074 = ~P2_STATE2_REG_0_ & ~n20507;
  assign n23075 = ~n23073 & ~n23074;
  assign n23076 = ~n23055 & ~n23075;
  assign n23077 = n23055 & n23075;
  assign n23078 = ~n23076 & ~n23077;
  assign n23079 = n22551 & n23078;
  assign n23080 = P2_REIP_REG_24_ & n22527;
  assign n23081 = P2_PHYADDRPOINTER_REG_24_ & n22554;
  assign n23082 = ~n23080 & ~n23081;
  assign n23083 = ~n20507 & n22557;
  assign n23084 = n23082 & ~n23083;
  assign n23085 = ~n23070 & ~n23071;
  assign n23086 = ~n23072 & n23085;
  assign n23087 = ~n23079 & n23086;
  assign n23088 = n23084 & n23087;
  assign n4949 = n23069 | ~n23088;
  assign n23090 = n19702 & n22541;
  assign n23091 = P2_EBX_REG_25_ & ~n22537;
  assign n23092 = ~n19732 & n22543;
  assign n23093 = P2_REIP_REG_25_ & n22527;
  assign n23094 = P2_PHYADDRPOINTER_REG_25_ & n22554;
  assign n23095 = ~n23093 & ~n23094;
  assign n23096 = ~n20521 & n22557;
  assign n23097 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_25_;
  assign n23098 = ~P2_STATE2_REG_0_ & ~n20521;
  assign n23099 = ~n23097 & ~n23098;
  assign n23100 = n23077 & n23099;
  assign n23101 = ~n23077 & ~n23099;
  assign n23102 = ~n23100 & ~n23101;
  assign n23103 = n22551 & n23102;
  assign n23104 = n23095 & ~n23096;
  assign n23105 = ~n23103 & n23104;
  assign n23106 = ~n19742 & n22539;
  assign n23107 = ~n23090 & ~n23091;
  assign n23108 = ~n23092 & n23107;
  assign n23109 = n23105 & n23108;
  assign n4954 = n23106 | ~n23109;
  assign n23111 = n19767 & n22541;
  assign n23112 = P2_EBX_REG_26_ & ~n22537;
  assign n23113 = P2_REIP_REG_26_ & n22527;
  assign n23114 = P2_PHYADDRPOINTER_REG_26_ & n22554;
  assign n23115 = ~n23113 & ~n23114;
  assign n23116 = ~n20535 & n22557;
  assign n23117 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_26_;
  assign n23118 = ~P2_STATE2_REG_0_ & ~n20535;
  assign n23119 = ~n23117 & ~n23118;
  assign n23120 = ~n23100 & ~n23119;
  assign n23121 = n23100 & n23119;
  assign n23122 = ~n23120 & ~n23121;
  assign n23123 = n22551 & n23122;
  assign n23124 = n23115 & ~n23116;
  assign n23125 = ~n23123 & n23124;
  assign n23126 = ~n19800 & n22543;
  assign n23127 = ~n19810 & n22539;
  assign n23128 = ~n23111 & ~n23112;
  assign n23129 = n23125 & n23128;
  assign n23130 = ~n23126 & n23129;
  assign n4959 = n23127 | ~n23130;
  assign n23132 = n19830 & n22541;
  assign n23133 = P2_EBX_REG_27_ & ~n22537;
  assign n23134 = P2_REIP_REG_27_ & n22527;
  assign n23135 = P2_PHYADDRPOINTER_REG_27_ & n22554;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n20549 & n22557;
  assign n23138 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_27_;
  assign n23139 = ~P2_STATE2_REG_0_ & ~n20549;
  assign n23140 = ~n23138 & ~n23139;
  assign n23141 = n23121 & n23140;
  assign n23142 = ~n23121 & ~n23140;
  assign n23143 = ~n23141 & ~n23142;
  assign n23144 = n22551 & n23143;
  assign n23145 = n23136 & ~n23137;
  assign n23146 = ~n23144 & n23145;
  assign n23147 = ~n19863 & n22543;
  assign n23148 = ~n19873 & n22539;
  assign n23149 = ~n23132 & ~n23133;
  assign n23150 = n23146 & n23149;
  assign n23151 = ~n23147 & n23150;
  assign n4964 = n23148 | ~n23151;
  assign n23153 = n19899 & n22541;
  assign n23154 = P2_EBX_REG_28_ & ~n22537;
  assign n23155 = P2_REIP_REG_28_ & n22527;
  assign n23156 = P2_PHYADDRPOINTER_REG_28_ & n22554;
  assign n23157 = ~n23155 & ~n23156;
  assign n23158 = ~n20563 & n22557;
  assign n23159 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_28_;
  assign n23160 = ~P2_STATE2_REG_0_ & ~n20563;
  assign n23161 = ~n23159 & ~n23160;
  assign n23162 = ~n23141 & ~n23161;
  assign n23163 = n23141 & n23161;
  assign n23164 = ~n23162 & ~n23163;
  assign n23165 = n22551 & n23164;
  assign n23166 = n23157 & ~n23158;
  assign n23167 = ~n23165 & n23166;
  assign n23168 = ~n19932 & n22543;
  assign n23169 = ~n19942 & n22539;
  assign n23170 = ~n23153 & ~n23154;
  assign n23171 = n23167 & n23170;
  assign n23172 = ~n23168 & n23171;
  assign n4969 = n23169 | ~n23172;
  assign n23174 = n19969 & n22541;
  assign n23175 = P2_EBX_REG_29_ & ~n22537;
  assign n23176 = P2_REIP_REG_29_ & n22527;
  assign n23177 = P2_PHYADDRPOINTER_REG_29_ & n22554;
  assign n23178 = ~n23176 & ~n23177;
  assign n23179 = ~n20577 & n22557;
  assign n23180 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_29_;
  assign n23181 = ~P2_STATE2_REG_0_ & ~n20577;
  assign n23182 = ~n23180 & ~n23181;
  assign n23183 = ~n23163 & ~n23182;
  assign n23184 = n23163 & n23182;
  assign n23185 = ~n23183 & ~n23184;
  assign n23186 = n22551 & n23185;
  assign n23187 = n23178 & ~n23179;
  assign n23188 = ~n23186 & n23187;
  assign n23189 = ~n20001 & n22543;
  assign n23190 = ~n20011 & n22539;
  assign n23191 = ~n23174 & ~n23175;
  assign n23192 = n23188 & n23191;
  assign n23193 = ~n23189 & n23192;
  assign n4974 = n23190 | ~n23193;
  assign n23195 = n20031 & n22541;
  assign n23196 = P2_EBX_REG_30_ & ~n22537;
  assign n23197 = P2_REIP_REG_30_ & n22527;
  assign n23198 = P2_PHYADDRPOINTER_REG_30_ & n22554;
  assign n23199 = ~n23197 & ~n23198;
  assign n23200 = ~n20591 & n22557;
  assign n23201 = P2_STATE2_REG_0_ & P2_INSTADDRPOINTER_REG_30_;
  assign n23202 = ~P2_STATE2_REG_0_ & ~n20591;
  assign n23203 = ~n23201 & ~n23202;
  assign n23204 = n23184 & n23203;
  assign n23205 = ~n23184 & ~n23203;
  assign n23206 = ~n23204 & ~n23205;
  assign n23207 = n22551 & n23206;
  assign n23208 = n23199 & ~n23200;
  assign n23209 = ~n23207 & n23208;
  assign n23210 = ~n20063 & n22543;
  assign n23211 = ~n20075 & n22539;
  assign n23212 = ~n23195 & ~n23196;
  assign n23213 = n23209 & n23212;
  assign n23214 = ~n23210 & n23213;
  assign n4979 = n23211 | ~n23214;
  assign n23216 = n20091 & n22541;
  assign n23217 = P2_EBX_REG_31_ & ~n22537;
  assign n23218 = P2_REIP_REG_31_ & n22527;
  assign n23219 = P2_PHYADDRPOINTER_REG_31_ & n22554;
  assign n23220 = ~n23218 & ~n23219;
  assign n23221 = ~n15336 & n22557;
  assign n23222 = ~n15338 & n23204;
  assign n23223 = n15338 & ~n23204;
  assign n23224 = ~n23222 & ~n23223;
  assign n23225 = n22551 & ~n23224;
  assign n23226 = n23220 & ~n23221;
  assign n23227 = ~n23225 & n23226;
  assign n23228 = ~n20138 & n22543;
  assign n23229 = n20151 & n22539;
  assign n23230 = ~n23216 & ~n23217;
  assign n23231 = n23227 & n23230;
  assign n23232 = ~n23228 & n23231;
  assign n4984 = n23229 | ~n23232;
  assign n23234 = ~P2_DATAWIDTH_REG_1_ & ~P2_REIP_REG_1_;
  assign n23235 = ~P2_DATAWIDTH_REG_30_ & ~P2_DATAWIDTH_REG_31_;
  assign n23236 = P2_DATAWIDTH_REG_0_ & P2_DATAWIDTH_REG_1_;
  assign n23237 = ~P2_DATAWIDTH_REG_28_ & ~P2_DATAWIDTH_REG_29_;
  assign n23238 = ~P2_DATAWIDTH_REG_26_ & ~P2_DATAWIDTH_REG_27_;
  assign n23239 = n23235 & ~n23236;
  assign n23240 = n23237 & n23239;
  assign n23241 = n23238 & n23240;
  assign n23242 = ~P2_DATAWIDTH_REG_22_ & ~P2_DATAWIDTH_REG_23_;
  assign n23243 = ~P2_DATAWIDTH_REG_24_ & n23242;
  assign n23244 = ~P2_DATAWIDTH_REG_25_ & n23243;
  assign n23245 = ~P2_DATAWIDTH_REG_18_ & ~P2_DATAWIDTH_REG_19_;
  assign n23246 = ~P2_DATAWIDTH_REG_20_ & n23245;
  assign n23247 = ~P2_DATAWIDTH_REG_21_ & n23246;
  assign n23248 = n23244 & n23247;
  assign n23249 = ~P2_DATAWIDTH_REG_14_ & ~P2_DATAWIDTH_REG_15_;
  assign n23250 = ~P2_DATAWIDTH_REG_16_ & n23249;
  assign n23251 = ~P2_DATAWIDTH_REG_17_ & n23250;
  assign n23252 = ~P2_DATAWIDTH_REG_10_ & ~P2_DATAWIDTH_REG_11_;
  assign n23253 = ~P2_DATAWIDTH_REG_12_ & n23252;
  assign n23254 = ~P2_DATAWIDTH_REG_13_ & n23253;
  assign n23255 = n23251 & n23254;
  assign n23256 = ~P2_DATAWIDTH_REG_6_ & ~P2_DATAWIDTH_REG_7_;
  assign n23257 = ~P2_DATAWIDTH_REG_8_ & n23256;
  assign n23258 = ~P2_DATAWIDTH_REG_9_ & n23257;
  assign n23259 = ~P2_DATAWIDTH_REG_2_ & ~P2_DATAWIDTH_REG_3_;
  assign n23260 = ~P2_DATAWIDTH_REG_4_ & n23259;
  assign n23261 = ~P2_DATAWIDTH_REG_5_ & n23260;
  assign n23262 = n23258 & n23261;
  assign n23263 = n23241 & n23248;
  assign n23264 = n23255 & n23263;
  assign n23265 = n23262 & n23264;
  assign n23266 = n23234 & n23265;
  assign n23267 = P2_BYTEENABLE_REG_3_ & ~n23265;
  assign n23268 = ~P2_DATAWIDTH_REG_1_ & ~P2_REIP_REG_0_;
  assign n23269 = ~P2_DATAWIDTH_REG_0_ & n23268;
  assign n23270 = n23265 & n23269;
  assign n23271 = ~n23266 & ~n23267;
  assign n4989 = n23270 | ~n23271;
  assign n23273 = P2_DATAWIDTH_REG_0_ & P2_REIP_REG_0_;
  assign n23274 = n23234 & ~n23273;
  assign n23275 = n23265 & n23274;
  assign n23276 = P2_BYTEENABLE_REG_2_ & ~n23265;
  assign n23277 = ~n23275 & ~n23276;
  assign n23278 = P2_REIP_REG_1_ & n23265;
  assign n23279 = P2_REIP_REG_0_ & n23278;
  assign n4994 = ~n23277 | n23279;
  assign n23281 = P2_BYTEENABLE_REG_1_ & ~n23265;
  assign n23282 = ~n23270 & ~n23278;
  assign n4999 = n23281 | ~n23282;
  assign n23284 = P2_REIP_REG_0_ & n23265;
  assign n23285 = P2_BYTEENABLE_REG_0_ & ~n23265;
  assign n23286 = ~n23284 & ~n23285;
  assign n5004 = n23278 | ~n23286;
  assign n23288 = P2_W_R_N_REG & ~n13883;
  assign n23289 = ~P2_READREQUEST_REG & n13883;
  assign n5009 = n23288 | n23289;
  assign n23291 = ~n14954 & n15432;
  assign n23292 = P2_FLUSH_REG & ~n23291;
  assign n23293 = ~n14238 & ~n15389;
  assign n23294 = n14238 & ~n15298;
  assign n23295 = ~n23293 & ~n23294;
  assign n23296 = n15048 & n15428;
  assign n23297 = n23295 & n23296;
  assign n5014 = n23292 | n23297;
  assign n23299 = P2_MORE_REG & ~n23291;
  assign n23300 = ~n15404 & n23291;
  assign n5019 = n23299 | n23300;
  assign n23302 = BS16 & ~n14104;
  assign n23303 = P2_STATEBS16_REG & n14104;
  assign n23304 = ~P2_STATE_REG_0_ & n14054;
  assign n23305 = ~n23302 & ~n23303;
  assign n5024 = n23304 | ~n23305;
  assign n23307 = ~n14857 & ~n14922;
  assign n23308 = n14051 & ~n23307;
  assign n23309 = P2_STATEBS16_REG & n14144;
  assign n23310 = n14238 & ~n23309;
  assign n23311 = n14550 & n23310;
  assign n23312 = ~n15424 & ~n23311;
  assign n23313 = ~n14145 & n14856;
  assign n23314 = n23312 & ~n23313;
  assign n23315 = ~n15446 & ~n23308;
  assign n23316 = n23314 & n23315;
  assign n23317 = ~P2_STATE2_REG_0_ & n15437;
  assign n23318 = P2_STATE2_REG_1_ & ~n14051;
  assign n23319 = n15495 & n23318;
  assign n23320 = ~n15480 & ~n23317;
  assign n23321 = ~n23319 & n23320;
  assign n23322 = ~n22526 & n23321;
  assign n23323 = ~n23316 & ~n23322;
  assign n23324 = P2_REQUESTPENDING_REG & n23322;
  assign n5029 = n23323 | n23324;
  assign n23326 = P2_D_C_N_REG & ~n13883;
  assign n23327 = ~P2_CODEFETCH_REG & n13883;
  assign n23328 = ~n23326 & ~n23327;
  assign n5034 = n23304 | ~n23328;
  assign n23330 = P2_MEMORYFETCH_REG & n13883;
  assign n23331 = P2_M_IO_N_REG & ~n13883;
  assign n5039 = n23330 | n23331;
  assign n23333 = P2_STATE2_REG_0_ & n17386;
  assign n23334 = n14953 & n15432;
  assign n23335 = P2_CODEFETCH_REG & ~n23334;
  assign n5044 = n23333 | n23335;
  assign n23337 = P2_STATE_REG_0_ & P2_ADS_N_REG;
  assign n5049 = ~n14104 | n23337;
  assign n23339 = P2_STATE2_REG_2_ & ~n14244;
  assign n23340 = ~n14243 & n23339;
  assign n23341 = ~n17386 & ~n22526;
  assign n23342 = ~n23340 & ~n23341;
  assign n23343 = P2_READREQUEST_REG & n23341;
  assign n5054 = n23342 | n23343;
  assign n23345 = ~n14199 & n15432;
  assign n23346 = n15183 & n23345;
  assign n23347 = ~n17386 & ~n23346;
  assign n23348 = ~n14238 & n14949;
  assign n23349 = n14238 & ~n14548;
  assign n23350 = ~n23348 & ~n23349;
  assign n23351 = n15013 & n15428;
  assign n23352 = n23350 & n23351;
  assign n23353 = P2_MEMORYFETCH_REG & ~n23352;
  assign n5059 = ~n23347 | n23353;
  assign n23355 = P1_STATE_REG_1_ & ~P1_STATE_REG_0_;
  assign n23356 = P1_BYTEENABLE_REG_3_ & n23355;
  assign n23357 = P1_BE_N_REG_3_ & ~n23355;
  assign n5064 = n23356 | n23357;
  assign n23359 = P1_BYTEENABLE_REG_2_ & n23355;
  assign n23360 = P1_BE_N_REG_2_ & ~n23355;
  assign n5069 = n23359 | n23360;
  assign n23362 = P1_BYTEENABLE_REG_1_ & n23355;
  assign n23363 = P1_BE_N_REG_1_ & ~n23355;
  assign n5074 = n23362 | n23363;
  assign n23365 = P1_BYTEENABLE_REG_0_ & n23355;
  assign n23366 = P1_BE_N_REG_0_ & ~n23355;
  assign n5079 = n23365 | n23366;
  assign n23368 = P1_STATE_REG_2_ & n23355;
  assign n23369 = P1_REIP_REG_30_ & n23368;
  assign n23370 = ~P1_STATE_REG_2_ & n23355;
  assign n23371 = P1_REIP_REG_31_ & n23370;
  assign n23372 = P1_ADDRESS_REG_29_ & ~n23355;
  assign n23373 = ~n23369 & ~n23371;
  assign n5084 = n23372 | ~n23373;
  assign n23375 = P1_REIP_REG_29_ & n23368;
  assign n23376 = P1_REIP_REG_30_ & n23370;
  assign n23377 = P1_ADDRESS_REG_28_ & ~n23355;
  assign n23378 = ~n23375 & ~n23376;
  assign n5088 = n23377 | ~n23378;
  assign n23380 = P1_REIP_REG_28_ & n23368;
  assign n23381 = P1_REIP_REG_29_ & n23370;
  assign n23382 = P1_ADDRESS_REG_27_ & ~n23355;
  assign n23383 = ~n23380 & ~n23381;
  assign n5092 = n23382 | ~n23383;
  assign n23385 = P1_REIP_REG_27_ & n23368;
  assign n23386 = P1_REIP_REG_28_ & n23370;
  assign n23387 = P1_ADDRESS_REG_26_ & ~n23355;
  assign n23388 = ~n23385 & ~n23386;
  assign n5096 = n23387 | ~n23388;
  assign n23390 = P1_REIP_REG_26_ & n23368;
  assign n23391 = P1_REIP_REG_27_ & n23370;
  assign n23392 = P1_ADDRESS_REG_25_ & ~n23355;
  assign n23393 = ~n23390 & ~n23391;
  assign n5100 = n23392 | ~n23393;
  assign n23395 = P1_REIP_REG_25_ & n23368;
  assign n23396 = P1_REIP_REG_26_ & n23370;
  assign n23397 = P1_ADDRESS_REG_24_ & ~n23355;
  assign n23398 = ~n23395 & ~n23396;
  assign n5104 = n23397 | ~n23398;
  assign n23400 = P1_REIP_REG_24_ & n23368;
  assign n23401 = P1_REIP_REG_25_ & n23370;
  assign n23402 = P1_ADDRESS_REG_23_ & ~n23355;
  assign n23403 = ~n23400 & ~n23401;
  assign n5108 = n23402 | ~n23403;
  assign n23405 = P1_REIP_REG_23_ & n23368;
  assign n23406 = P1_REIP_REG_24_ & n23370;
  assign n23407 = P1_ADDRESS_REG_22_ & ~n23355;
  assign n23408 = ~n23405 & ~n23406;
  assign n5112 = n23407 | ~n23408;
  assign n23410 = P1_REIP_REG_22_ & n23368;
  assign n23411 = P1_REIP_REG_23_ & n23370;
  assign n23412 = P1_ADDRESS_REG_21_ & ~n23355;
  assign n23413 = ~n23410 & ~n23411;
  assign n5116 = n23412 | ~n23413;
  assign n23415 = P1_REIP_REG_21_ & n23368;
  assign n23416 = P1_REIP_REG_22_ & n23370;
  assign n23417 = P1_ADDRESS_REG_20_ & ~n23355;
  assign n23418 = ~n23415 & ~n23416;
  assign n5120 = n23417 | ~n23418;
  assign n23420 = P1_REIP_REG_20_ & n23368;
  assign n23421 = P1_REIP_REG_21_ & n23370;
  assign n23422 = P1_ADDRESS_REG_19_ & ~n23355;
  assign n23423 = ~n23420 & ~n23421;
  assign n5124 = n23422 | ~n23423;
  assign n23425 = P1_REIP_REG_19_ & n23368;
  assign n23426 = P1_REIP_REG_20_ & n23370;
  assign n23427 = P1_ADDRESS_REG_18_ & ~n23355;
  assign n23428 = ~n23425 & ~n23426;
  assign n5128 = n23427 | ~n23428;
  assign n23430 = P1_REIP_REG_18_ & n23368;
  assign n23431 = P1_REIP_REG_19_ & n23370;
  assign n23432 = P1_ADDRESS_REG_17_ & ~n23355;
  assign n23433 = ~n23430 & ~n23431;
  assign n5132 = n23432 | ~n23433;
  assign n23435 = P1_REIP_REG_17_ & n23368;
  assign n23436 = P1_REIP_REG_18_ & n23370;
  assign n23437 = P1_ADDRESS_REG_16_ & ~n23355;
  assign n23438 = ~n23435 & ~n23436;
  assign n5136 = n23437 | ~n23438;
  assign n23440 = P1_REIP_REG_16_ & n23368;
  assign n23441 = P1_REIP_REG_17_ & n23370;
  assign n23442 = P1_ADDRESS_REG_15_ & ~n23355;
  assign n23443 = ~n23440 & ~n23441;
  assign n5140 = n23442 | ~n23443;
  assign n23445 = P1_REIP_REG_15_ & n23368;
  assign n23446 = P1_REIP_REG_16_ & n23370;
  assign n23447 = P1_ADDRESS_REG_14_ & ~n23355;
  assign n23448 = ~n23445 & ~n23446;
  assign n5144 = n23447 | ~n23448;
  assign n23450 = P1_REIP_REG_14_ & n23368;
  assign n23451 = P1_REIP_REG_15_ & n23370;
  assign n23452 = P1_ADDRESS_REG_13_ & ~n23355;
  assign n23453 = ~n23450 & ~n23451;
  assign n5148 = n23452 | ~n23453;
  assign n23455 = P1_REIP_REG_13_ & n23368;
  assign n23456 = P1_REIP_REG_14_ & n23370;
  assign n23457 = P1_ADDRESS_REG_12_ & ~n23355;
  assign n23458 = ~n23455 & ~n23456;
  assign n5152 = n23457 | ~n23458;
  assign n23460 = P1_REIP_REG_12_ & n23368;
  assign n23461 = P1_REIP_REG_13_ & n23370;
  assign n23462 = P1_ADDRESS_REG_11_ & ~n23355;
  assign n23463 = ~n23460 & ~n23461;
  assign n5156 = n23462 | ~n23463;
  assign n23465 = P1_REIP_REG_11_ & n23368;
  assign n23466 = P1_REIP_REG_12_ & n23370;
  assign n23467 = P1_ADDRESS_REG_10_ & ~n23355;
  assign n23468 = ~n23465 & ~n23466;
  assign n5160 = n23467 | ~n23468;
  assign n23470 = P1_REIP_REG_10_ & n23368;
  assign n23471 = P1_REIP_REG_11_ & n23370;
  assign n23472 = P1_ADDRESS_REG_9_ & ~n23355;
  assign n23473 = ~n23470 & ~n23471;
  assign n5164 = n23472 | ~n23473;
  assign n23475 = P1_REIP_REG_9_ & n23368;
  assign n23476 = P1_REIP_REG_10_ & n23370;
  assign n23477 = P1_ADDRESS_REG_8_ & ~n23355;
  assign n23478 = ~n23475 & ~n23476;
  assign n5168 = n23477 | ~n23478;
  assign n23480 = P1_REIP_REG_8_ & n23368;
  assign n23481 = P1_REIP_REG_9_ & n23370;
  assign n23482 = P1_ADDRESS_REG_7_ & ~n23355;
  assign n23483 = ~n23480 & ~n23481;
  assign n5172 = n23482 | ~n23483;
  assign n23485 = P1_REIP_REG_7_ & n23368;
  assign n23486 = P1_REIP_REG_8_ & n23370;
  assign n23487 = P1_ADDRESS_REG_6_ & ~n23355;
  assign n23488 = ~n23485 & ~n23486;
  assign n5176 = n23487 | ~n23488;
  assign n23490 = P1_REIP_REG_6_ & n23368;
  assign n23491 = P1_REIP_REG_7_ & n23370;
  assign n23492 = P1_ADDRESS_REG_5_ & ~n23355;
  assign n23493 = ~n23490 & ~n23491;
  assign n5180 = n23492 | ~n23493;
  assign n23495 = P1_REIP_REG_5_ & n23368;
  assign n23496 = P1_REIP_REG_6_ & n23370;
  assign n23497 = P1_ADDRESS_REG_4_ & ~n23355;
  assign n23498 = ~n23495 & ~n23496;
  assign n5184 = n23497 | ~n23498;
  assign n23500 = P1_REIP_REG_4_ & n23368;
  assign n23501 = P1_REIP_REG_5_ & n23370;
  assign n23502 = P1_ADDRESS_REG_3_ & ~n23355;
  assign n23503 = ~n23500 & ~n23501;
  assign n5188 = n23502 | ~n23503;
  assign n23505 = P1_REIP_REG_3_ & n23368;
  assign n23506 = P1_REIP_REG_4_ & n23370;
  assign n23507 = P1_ADDRESS_REG_2_ & ~n23355;
  assign n23508 = ~n23505 & ~n23506;
  assign n5192 = n23507 | ~n23508;
  assign n23510 = P1_REIP_REG_2_ & n23368;
  assign n23511 = P1_REIP_REG_3_ & n23370;
  assign n23512 = P1_ADDRESS_REG_1_ & ~n23355;
  assign n23513 = ~n23510 & ~n23511;
  assign n5196 = n23512 | ~n23513;
  assign n23515 = P1_REIP_REG_1_ & n23368;
  assign n23516 = P1_REIP_REG_2_ & n23370;
  assign n23517 = P1_ADDRESS_REG_0_ & ~n23355;
  assign n23518 = ~n23515 & ~n23516;
  assign n5200 = n23517 | ~n23518;
  assign n23520 = ~P1_STATE_REG_2_ & P1_STATE_REG_1_;
  assign n23521 = NA & n23520;
  assign n23522 = ~HOLD & ~P1_REQUESTPENDING_REG;
  assign n23523 = READY1 & READY11_REG;
  assign n23524 = P1_STATE_REG_1_ & ~n23522;
  assign n23525 = n23523 & n23524;
  assign n23526 = ~P1_STATE_REG_2_ & ~P1_STATE_REG_1_;
  assign n23527 = HOLD & ~P1_REQUESTPENDING_REG;
  assign n23528 = n23526 & n23527;
  assign n23529 = ~n23525 & ~n23528;
  assign n23530 = P1_STATE_REG_0_ & ~n23521;
  assign n23531 = ~n23529 & n23530;
  assign n23532 = ~n23368 & ~n23531;
  assign n23533 = ~HOLD & P1_REQUESTPENDING_REG;
  assign n23534 = P1_STATE_REG_0_ & ~n23533;
  assign n23535 = ~n23522 & n23534;
  assign n23536 = ~NA & ~P1_STATE_REG_0_;
  assign n23537 = n23522 & ~n23523;
  assign n23538 = ~n23523 & n23533;
  assign n23539 = P1_STATE_REG_1_ & ~n23537;
  assign n23540 = ~n23538 & n23539;
  assign n23541 = ~n23535 & ~n23536;
  assign n23542 = ~n23540 & n23541;
  assign n23543 = P1_STATE_REG_2_ & ~n23542;
  assign n5204 = ~n23532 | n23543;
  assign n23545 = P1_STATE_REG_2_ & ~n23534;
  assign n23546 = P1_STATE_REG_0_ & P1_REQUESTPENDING_REG;
  assign n23547 = ~P1_STATE_REG_2_ & n23546;
  assign n23548 = ~n23545 & ~n23547;
  assign n23549 = ~P1_STATE_REG_1_ & ~n23548;
  assign n23550 = HOLD & ~n23523;
  assign n23551 = P1_STATE_REG_0_ & ~n23550;
  assign n23552 = P1_STATE_REG_2_ & ~n23551;
  assign n23553 = ~n23537 & ~n23552;
  assign n23554 = P1_STATE_REG_1_ & n23553;
  assign n23555 = n23355 & n23523;
  assign n23556 = ~n23370 & ~n23555;
  assign n23557 = ~n23549 & ~n23554;
  assign n5209 = ~n23556 | ~n23557;
  assign n23559 = P1_STATE_REG_1_ & ~n23538;
  assign n23560 = n23546 & ~n23559;
  assign n23561 = ~P1_STATE_REG_2_ & ~n23560;
  assign n23562 = P1_STATE_REG_2_ & n23534;
  assign n23563 = NA & ~P1_STATE_REG_0_;
  assign n23564 = P1_STATE_REG_2_ & ~n23533;
  assign n23565 = ~n23563 & ~n23564;
  assign n23566 = ~P1_STATE_REG_1_ & ~n23565;
  assign n23567 = ~n23561 & ~n23562;
  assign n5214 = n23566 | ~n23567;
  assign n23569 = ~BS16 & ~n23526;
  assign n23570 = P1_STATE_REG_0_ & n23520;
  assign n23571 = ~P1_STATE_REG_1_ & ~P1_STATE_REG_0_;
  assign n23572 = ~n23570 & ~n23571;
  assign n23573 = n23569 & ~n23572;
  assign n23574 = P1_DATAWIDTH_REG_0_ & n23572;
  assign n5219 = n23573 | n23574;
  assign n23576 = P1_DATAWIDTH_REG_1_ & n23572;
  assign n23577 = ~n23569 & ~n23572;
  assign n5224 = n23576 | n23577;
  assign n5229 = P1_DATAWIDTH_REG_2_ & n23572;
  assign n5234 = P1_DATAWIDTH_REG_3_ & n23572;
  assign n5239 = P1_DATAWIDTH_REG_4_ & n23572;
  assign n5244 = P1_DATAWIDTH_REG_5_ & n23572;
  assign n5249 = P1_DATAWIDTH_REG_6_ & n23572;
  assign n5254 = P1_DATAWIDTH_REG_7_ & n23572;
  assign n5259 = P1_DATAWIDTH_REG_8_ & n23572;
  assign n5264 = P1_DATAWIDTH_REG_9_ & n23572;
  assign n5269 = P1_DATAWIDTH_REG_10_ & n23572;
  assign n5274 = P1_DATAWIDTH_REG_11_ & n23572;
  assign n5279 = P1_DATAWIDTH_REG_12_ & n23572;
  assign n5284 = P1_DATAWIDTH_REG_13_ & n23572;
  assign n5289 = P1_DATAWIDTH_REG_14_ & n23572;
  assign n5294 = P1_DATAWIDTH_REG_15_ & n23572;
  assign n5299 = P1_DATAWIDTH_REG_16_ & n23572;
  assign n5304 = P1_DATAWIDTH_REG_17_ & n23572;
  assign n5309 = P1_DATAWIDTH_REG_18_ & n23572;
  assign n5314 = P1_DATAWIDTH_REG_19_ & n23572;
  assign n5319 = P1_DATAWIDTH_REG_20_ & n23572;
  assign n5324 = P1_DATAWIDTH_REG_21_ & n23572;
  assign n5329 = P1_DATAWIDTH_REG_22_ & n23572;
  assign n5334 = P1_DATAWIDTH_REG_23_ & n23572;
  assign n5339 = P1_DATAWIDTH_REG_24_ & n23572;
  assign n5344 = P1_DATAWIDTH_REG_25_ & n23572;
  assign n5349 = P1_DATAWIDTH_REG_26_ & n23572;
  assign n5354 = P1_DATAWIDTH_REG_27_ & n23572;
  assign n5359 = P1_DATAWIDTH_REG_28_ & n23572;
  assign n5364 = P1_DATAWIDTH_REG_29_ & n23572;
  assign n5369 = P1_DATAWIDTH_REG_30_ & n23572;
  assign n5374 = P1_DATAWIDTH_REG_31_ & n23572;
  assign n23609 = P1_STATE2_REG_2_ & P1_STATE2_REG_1_;
  assign n23610 = P1_STATE2_REG_1_ & n23523;
  assign n23611 = ~P1_STATE2_REG_0_ & ~n23610;
  assign n23612 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23613 = P1_INSTQUEUERD_ADDR_REG_1_ & n23612;
  assign n23614 = P1_INSTQUEUERD_ADDR_REG_2_ & n23613;
  assign n23615 = P1_INSTQUEUE_REG_15__0_ & n23614;
  assign n23616 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23617 = P1_INSTQUEUERD_ADDR_REG_2_ & n23616;
  assign n23618 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23617;
  assign n23619 = P1_INSTQUEUE_REG_14__0_ & n23618;
  assign n23620 = P1_INSTQUEUERD_ADDR_REG_2_ & n23612;
  assign n23621 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23620;
  assign n23622 = P1_INSTQUEUE_REG_13__0_ & n23621;
  assign n23623 = P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23624 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23625 = n23623 & n23624;
  assign n23626 = P1_INSTQUEUE_REG_12__0_ & n23625;
  assign n23627 = ~n23615 & ~n23619;
  assign n23628 = ~n23622 & n23627;
  assign n23629 = ~n23626 & n23628;
  assign n23630 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23613;
  assign n23631 = P1_INSTQUEUE_REG_11__0_ & n23630;
  assign n23632 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23633 = n23616 & n23632;
  assign n23634 = P1_INSTQUEUE_REG_10__0_ & n23633;
  assign n23635 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23636 = n23612 & n23635;
  assign n23637 = P1_INSTQUEUE_REG_9__0_ & n23636;
  assign n23638 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23624;
  assign n23639 = P1_INSTQUEUERD_ADDR_REG_3_ & n23638;
  assign n23640 = P1_INSTQUEUE_REG_8__0_ & n23639;
  assign n23641 = ~n23631 & ~n23634;
  assign n23642 = ~n23637 & n23641;
  assign n23643 = ~n23640 & n23642;
  assign n23644 = P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23645 = ~P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23646 = n23644 & n23645;
  assign n23647 = P1_INSTQUEUE_REG_6__0_ & n23646;
  assign n23648 = P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23649 = ~P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23650 = n23648 & n23649;
  assign n23651 = P1_INSTQUEUE_REG_5__0_ & n23650;
  assign n23652 = ~P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23653 = n23624 & n23652;
  assign n23654 = P1_INSTQUEUE_REG_4__0_ & n23653;
  assign n23655 = P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23656 = ~P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23657 = n23655 & n23656;
  assign n23658 = P1_INSTQUEUE_REG_3__0_ & n23657;
  assign n23659 = ~n23647 & ~n23651;
  assign n23660 = ~n23654 & n23659;
  assign n23661 = ~n23658 & n23660;
  assign n23662 = P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23663 = n23656 & n23662;
  assign n23664 = P1_INSTQUEUE_REG_2__0_ & n23663;
  assign n23665 = ~P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23666 = n23656 & n23665;
  assign n23667 = P1_INSTQUEUE_REG_1__0_ & n23666;
  assign n23668 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23638;
  assign n23669 = P1_INSTQUEUE_REG_0__0_ & n23668;
  assign n23670 = P1_INSTQUEUERD_ADDR_REG_2_ & n23655;
  assign n23671 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23670;
  assign n23672 = P1_INSTQUEUE_REG_7__0_ & n23671;
  assign n23673 = ~n23664 & ~n23667;
  assign n23674 = ~n23669 & n23673;
  assign n23675 = ~n23672 & n23674;
  assign n23676 = n23629 & n23643;
  assign n23677 = n23661 & n23676;
  assign n23678 = n23675 & n23677;
  assign n23679 = P1_INSTQUEUE_REG_15__1_ & n23614;
  assign n23680 = P1_INSTQUEUE_REG_14__1_ & n23618;
  assign n23681 = P1_INSTQUEUE_REG_13__1_ & n23621;
  assign n23682 = P1_INSTQUEUE_REG_12__1_ & n23625;
  assign n23683 = ~n23679 & ~n23680;
  assign n23684 = ~n23681 & n23683;
  assign n23685 = ~n23682 & n23684;
  assign n23686 = P1_INSTQUEUE_REG_11__1_ & n23630;
  assign n23687 = P1_INSTQUEUE_REG_10__1_ & n23633;
  assign n23688 = P1_INSTQUEUE_REG_9__1_ & n23636;
  assign n23689 = P1_INSTQUEUE_REG_8__1_ & n23639;
  assign n23690 = ~n23686 & ~n23687;
  assign n23691 = ~n23688 & n23690;
  assign n23692 = ~n23689 & n23691;
  assign n23693 = P1_INSTQUEUE_REG_6__1_ & n23646;
  assign n23694 = P1_INSTQUEUE_REG_5__1_ & n23650;
  assign n23695 = P1_INSTQUEUE_REG_4__1_ & n23653;
  assign n23696 = P1_INSTQUEUE_REG_3__1_ & n23657;
  assign n23697 = ~n23693 & ~n23694;
  assign n23698 = ~n23695 & n23697;
  assign n23699 = ~n23696 & n23698;
  assign n23700 = P1_INSTQUEUE_REG_2__1_ & n23663;
  assign n23701 = P1_INSTQUEUE_REG_1__1_ & n23666;
  assign n23702 = P1_INSTQUEUE_REG_0__1_ & n23668;
  assign n23703 = P1_INSTQUEUE_REG_7__1_ & n23671;
  assign n23704 = ~n23700 & ~n23701;
  assign n23705 = ~n23702 & n23704;
  assign n23706 = ~n23703 & n23705;
  assign n23707 = n23685 & n23692;
  assign n23708 = n23699 & n23707;
  assign n23709 = n23706 & n23708;
  assign n23710 = n23678 & n23709;
  assign n23711 = P1_INSTQUEUE_REG_15__3_ & n23614;
  assign n23712 = P1_INSTQUEUE_REG_14__3_ & n23618;
  assign n23713 = P1_INSTQUEUE_REG_13__3_ & n23621;
  assign n23714 = P1_INSTQUEUE_REG_12__3_ & n23625;
  assign n23715 = ~n23711 & ~n23712;
  assign n23716 = ~n23713 & n23715;
  assign n23717 = ~n23714 & n23716;
  assign n23718 = P1_INSTQUEUE_REG_11__3_ & n23630;
  assign n23719 = P1_INSTQUEUE_REG_10__3_ & n23633;
  assign n23720 = P1_INSTQUEUE_REG_9__3_ & n23636;
  assign n23721 = P1_INSTQUEUE_REG_8__3_ & n23639;
  assign n23722 = ~n23718 & ~n23719;
  assign n23723 = ~n23720 & n23722;
  assign n23724 = ~n23721 & n23723;
  assign n23725 = P1_INSTQUEUE_REG_6__3_ & n23646;
  assign n23726 = P1_INSTQUEUE_REG_5__3_ & n23650;
  assign n23727 = P1_INSTQUEUE_REG_4__3_ & n23653;
  assign n23728 = P1_INSTQUEUE_REG_3__3_ & n23657;
  assign n23729 = ~n23725 & ~n23726;
  assign n23730 = ~n23727 & n23729;
  assign n23731 = ~n23728 & n23730;
  assign n23732 = P1_INSTQUEUE_REG_2__3_ & n23663;
  assign n23733 = P1_INSTQUEUE_REG_1__3_ & n23666;
  assign n23734 = P1_INSTQUEUE_REG_0__3_ & n23668;
  assign n23735 = P1_INSTQUEUE_REG_7__3_ & n23671;
  assign n23736 = ~n23732 & ~n23733;
  assign n23737 = ~n23734 & n23736;
  assign n23738 = ~n23735 & n23737;
  assign n23739 = n23717 & n23724;
  assign n23740 = n23731 & n23739;
  assign n23741 = n23738 & n23740;
  assign n23742 = n23710 & ~n23741;
  assign n23743 = P1_INSTQUEUE_REG_8__6_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23744 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23743;
  assign n23745 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23744;
  assign n23746 = P1_INSTQUEUERD_ADDR_REG_3_ & n23745;
  assign n23747 = P1_INSTQUEUE_REG_0__6_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23748 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23747;
  assign n23749 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23748;
  assign n23750 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23749;
  assign n23751 = P1_INSTQUEUE_REG_11__6_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23752 = P1_INSTQUEUERD_ADDR_REG_1_ & n23751;
  assign n23753 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23752;
  assign n23754 = P1_INSTQUEUERD_ADDR_REG_0_ & n23753;
  assign n23755 = P1_INSTQUEUE_REG_10__6_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23756 = P1_INSTQUEUERD_ADDR_REG_1_ & n23755;
  assign n23757 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23756;
  assign n23758 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23757;
  assign n23759 = ~n23746 & ~n23750;
  assign n23760 = ~n23754 & n23759;
  assign n23761 = ~n23758 & n23760;
  assign n23762 = P1_INSTQUEUE_REG_3__6_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23763 = n23656 & n23762;
  assign n23764 = P1_INSTQUEUERD_ADDR_REG_1_ & n23763;
  assign n23765 = P1_INSTQUEUE_REG_9__6_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23766 = P1_INSTQUEUERD_ADDR_REG_0_ & n23765;
  assign n23767 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23766;
  assign n23768 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23767;
  assign n23769 = ~n23764 & ~n23768;
  assign n23770 = n23623 & n23662;
  assign n23771 = P1_INSTQUEUE_REG_14__6_ & n23770;
  assign n23772 = n23623 & n23665;
  assign n23773 = P1_INSTQUEUE_REG_13__6_ & n23772;
  assign n23774 = n23623 & n23655;
  assign n23775 = P1_INSTQUEUE_REG_15__6_ & n23774;
  assign n23776 = ~n23771 & ~n23773;
  assign n23777 = ~n23775 & n23776;
  assign n23778 = n23652 & n23662;
  assign n23779 = P1_INSTQUEUE_REG_6__6_ & n23778;
  assign n23780 = n23652 & n23665;
  assign n23781 = P1_INSTQUEUE_REG_5__6_ & n23780;
  assign n23782 = P1_INSTQUEUE_REG_12__6_ & n23624;
  assign n23783 = n23623 & n23782;
  assign n23784 = ~n23779 & ~n23781;
  assign n23785 = ~n23783 & n23784;
  assign n23786 = P1_INSTQUEUE_REG_4__6_ & n23624;
  assign n23787 = n23652 & n23786;
  assign n23788 = P1_INSTQUEUE_REG_2__6_ & n23656;
  assign n23789 = n23662 & n23788;
  assign n23790 = P1_INSTQUEUE_REG_1__6_ & n23656;
  assign n23791 = n23665 & n23790;
  assign n23792 = n23652 & n23655;
  assign n23793 = P1_INSTQUEUE_REG_7__6_ & n23792;
  assign n23794 = ~n23787 & ~n23789;
  assign n23795 = ~n23791 & n23794;
  assign n23796 = ~n23793 & n23795;
  assign n23797 = n23761 & n23769;
  assign n23798 = n23777 & n23797;
  assign n23799 = n23785 & n23798;
  assign n23800 = n23796 & n23799;
  assign n23801 = P1_INSTQUEUE_REG_15__7_ & n23614;
  assign n23802 = P1_INSTQUEUE_REG_14__7_ & n23618;
  assign n23803 = P1_INSTQUEUE_REG_13__7_ & n23621;
  assign n23804 = P1_INSTQUEUE_REG_12__7_ & n23625;
  assign n23805 = ~n23801 & ~n23802;
  assign n23806 = ~n23803 & n23805;
  assign n23807 = ~n23804 & n23806;
  assign n23808 = P1_INSTQUEUE_REG_11__7_ & n23630;
  assign n23809 = P1_INSTQUEUE_REG_10__7_ & n23633;
  assign n23810 = P1_INSTQUEUE_REG_9__7_ & n23636;
  assign n23811 = P1_INSTQUEUE_REG_8__7_ & n23639;
  assign n23812 = ~n23808 & ~n23809;
  assign n23813 = ~n23810 & n23812;
  assign n23814 = ~n23811 & n23813;
  assign n23815 = P1_INSTQUEUE_REG_6__7_ & n23646;
  assign n23816 = P1_INSTQUEUE_REG_5__7_ & n23650;
  assign n23817 = P1_INSTQUEUE_REG_4__7_ & n23653;
  assign n23818 = P1_INSTQUEUE_REG_3__7_ & n23657;
  assign n23819 = ~n23815 & ~n23816;
  assign n23820 = ~n23817 & n23819;
  assign n23821 = ~n23818 & n23820;
  assign n23822 = P1_INSTQUEUE_REG_2__7_ & n23663;
  assign n23823 = P1_INSTQUEUE_REG_1__7_ & n23666;
  assign n23824 = P1_INSTQUEUE_REG_0__7_ & n23668;
  assign n23825 = P1_INSTQUEUE_REG_7__7_ & n23671;
  assign n23826 = ~n23822 & ~n23823;
  assign n23827 = ~n23824 & n23826;
  assign n23828 = ~n23825 & n23827;
  assign n23829 = n23807 & n23814;
  assign n23830 = n23821 & n23829;
  assign n23831 = n23828 & n23830;
  assign n23832 = P1_INSTQUEUERD_ADDR_REG_0_ & n23644;
  assign n23833 = P1_INSTQUEUE_REG_15__5_ & n23832;
  assign n23834 = P1_INSTQUEUERD_ADDR_REG_3_ & n23833;
  assign n23835 = P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23836 = P1_INSTQUEUERD_ADDR_REG_1_ & n23835;
  assign n23837 = P1_INSTQUEUE_REG_14__5_ & n23836;
  assign n23838 = P1_INSTQUEUERD_ADDR_REG_3_ & n23837;
  assign n23839 = ~n23834 & ~n23838;
  assign n23840 = P1_INSTQUEUE_REG_9__5_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23841 = n23635 & n23840;
  assign n23842 = P1_INSTQUEUERD_ADDR_REG_3_ & n23841;
  assign n23843 = P1_INSTQUEUE_REG_3__5_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23844 = P1_INSTQUEUERD_ADDR_REG_1_ & n23843;
  assign n23845 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23844;
  assign n23846 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23845;
  assign n23847 = ~n23842 & ~n23846;
  assign n23848 = P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23849 = P1_INSTQUEUERD_ADDR_REG_0_ & n23848;
  assign n23850 = P1_INSTQUEUE_REG_13__5_ & n23849;
  assign n23851 = P1_INSTQUEUERD_ADDR_REG_3_ & n23850;
  assign n23852 = P1_INSTQUEUE_REG_12__5_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23853 = P1_INSTQUEUERD_ADDR_REG_2_ & n23624;
  assign n23854 = n23852 & n23853;
  assign n23855 = ~P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23856 = P1_INSTQUEUERD_ADDR_REG_0_ & n23855;
  assign n23857 = P1_INSTQUEUE_REG_11__5_ & n23856;
  assign n23858 = P1_INSTQUEUERD_ADDR_REG_3_ & n23857;
  assign n23859 = P1_INSTQUEUE_REG_10__5_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23860 = P1_INSTQUEUERD_ADDR_REG_1_ & n23632;
  assign n23861 = n23859 & n23860;
  assign n23862 = ~n23851 & ~n23854;
  assign n23863 = ~n23858 & n23862;
  assign n23864 = ~n23861 & n23863;
  assign n23865 = P1_INSTQUEUE_REG_8__5_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23866 = n23638 & n23865;
  assign n23867 = P1_INSTQUEUE_REG_6__5_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign n23868 = P1_INSTQUEUERD_ADDR_REG_2_ & n23645;
  assign n23869 = n23867 & n23868;
  assign n23870 = P1_INSTQUEUE_REG_5__5_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23871 = P1_INSTQUEUERD_ADDR_REG_2_ & n23649;
  assign n23872 = n23870 & n23871;
  assign n23873 = P1_INSTQUEUE_REG_4__5_ & n23624;
  assign n23874 = P1_INSTQUEUERD_ADDR_REG_2_ & n23873;
  assign n23875 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23874;
  assign n23876 = ~n23866 & ~n23869;
  assign n23877 = ~n23872 & n23876;
  assign n23878 = ~n23875 & n23877;
  assign n23879 = P1_INSTQUEUE_REG_2__5_ & n23656;
  assign n23880 = P1_INSTQUEUERD_ADDR_REG_1_ & n23879;
  assign n23881 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23880;
  assign n23882 = P1_INSTQUEUE_REG_1__5_ & n23656;
  assign n23883 = P1_INSTQUEUERD_ADDR_REG_0_ & n23882;
  assign n23884 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23883;
  assign n23885 = P1_INSTQUEUE_REG_0__5_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23886 = n23638 & n23885;
  assign n23887 = P1_INSTQUEUERD_ADDR_REG_1_ & n23652;
  assign n23888 = P1_INSTQUEUE_REG_7__5_ & n23887;
  assign n23889 = P1_INSTQUEUERD_ADDR_REG_0_ & n23888;
  assign n23890 = ~n23881 & ~n23884;
  assign n23891 = ~n23886 & n23890;
  assign n23892 = ~n23889 & n23891;
  assign n23893 = n23839 & n23847;
  assign n23894 = n23864 & n23893;
  assign n23895 = n23878 & n23894;
  assign n23896 = n23892 & n23895;
  assign n23897 = P1_INSTQUEUE_REG_11__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23898 = P1_INSTQUEUERD_ADDR_REG_1_ & n23897;
  assign n23899 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23898;
  assign n23900 = P1_INSTQUEUERD_ADDR_REG_3_ & n23899;
  assign n23901 = P1_INSTQUEUE_REG_3__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23902 = P1_INSTQUEUERD_ADDR_REG_1_ & n23901;
  assign n23903 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23902;
  assign n23904 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23903;
  assign n23905 = P1_INSTQUEUE_REG_9__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23906 = n23635 & n23905;
  assign n23907 = P1_INSTQUEUERD_ADDR_REG_0_ & n23906;
  assign n23908 = P1_INSTQUEUE_REG_10__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23909 = P1_INSTQUEUERD_ADDR_REG_1_ & n23908;
  assign n23910 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23909;
  assign n23911 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23910;
  assign n23912 = ~n23900 & ~n23904;
  assign n23913 = ~n23907 & n23912;
  assign n23914 = ~n23911 & n23913;
  assign n23915 = P1_INSTQUEUE_REG_8__4_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23916 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23915;
  assign n23917 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23916;
  assign n23918 = P1_INSTQUEUERD_ADDR_REG_3_ & n23917;
  assign n23919 = P1_INSTQUEUE_REG_0__4_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23920 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23919;
  assign n23921 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23920;
  assign n23922 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23921;
  assign n23923 = P1_INSTQUEUE_REG_15__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23924 = P1_INSTQUEUERD_ADDR_REG_1_ & n23923;
  assign n23925 = P1_INSTQUEUERD_ADDR_REG_2_ & n23924;
  assign n23926 = P1_INSTQUEUERD_ADDR_REG_0_ & n23925;
  assign n23927 = P1_INSTQUEUE_REG_14__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23928 = n23644 & n23927;
  assign n23929 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23928;
  assign n23930 = ~n23918 & ~n23922;
  assign n23931 = ~n23926 & n23930;
  assign n23932 = ~n23929 & n23931;
  assign n23933 = P1_INSTQUEUE_REG_6__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23934 = n23645 & n23933;
  assign n23935 = P1_INSTQUEUERD_ADDR_REG_1_ & n23934;
  assign n23936 = P1_INSTQUEUE_REG_13__4_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23937 = n23648 & n23936;
  assign n23938 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23937;
  assign n23939 = P1_INSTQUEUE_REG_12__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23940 = n23624 & n23939;
  assign n23941 = P1_INSTQUEUERD_ADDR_REG_3_ & n23940;
  assign n23942 = P1_INSTQUEUE_REG_4__4_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n23943 = n23624 & n23942;
  assign n23944 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23943;
  assign n23945 = ~n23935 & ~n23938;
  assign n23946 = ~n23941 & n23945;
  assign n23947 = ~n23944 & n23946;
  assign n23948 = P1_INSTQUEUE_REG_2__4_ & ~P1_INSTQUEUERD_ADDR_REG_3_;
  assign n23949 = ~P1_INSTQUEUERD_ADDR_REG_2_ & n23948;
  assign n23950 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n23949;
  assign n23951 = P1_INSTQUEUERD_ADDR_REG_1_ & n23950;
  assign n23952 = P1_INSTQUEUE_REG_5__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23953 = P1_INSTQUEUERD_ADDR_REG_2_ & n23952;
  assign n23954 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23953;
  assign n23955 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23954;
  assign n23956 = P1_INSTQUEUE_REG_7__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23957 = P1_INSTQUEUERD_ADDR_REG_2_ & n23956;
  assign n23958 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n23957;
  assign n23959 = P1_INSTQUEUERD_ADDR_REG_1_ & n23958;
  assign n23960 = P1_INSTQUEUE_REG_1__4_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n23961 = n23656 & n23960;
  assign n23962 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n23961;
  assign n23963 = ~n23951 & ~n23955;
  assign n23964 = ~n23959 & n23963;
  assign n23965 = ~n23962 & n23964;
  assign n23966 = n23914 & n23932;
  assign n23967 = n23947 & n23966;
  assign n23968 = n23965 & n23967;
  assign n23969 = n23800 & ~n23831;
  assign n23970 = ~n23896 & n23969;
  assign n23971 = ~n23968 & n23970;
  assign n23972 = P1_INSTQUEUE_REG_15__2_ & n23614;
  assign n23973 = P1_INSTQUEUE_REG_14__2_ & n23618;
  assign n23974 = P1_INSTQUEUE_REG_13__2_ & n23621;
  assign n23975 = P1_INSTQUEUE_REG_12__2_ & n23625;
  assign n23976 = ~n23972 & ~n23973;
  assign n23977 = ~n23974 & n23976;
  assign n23978 = ~n23975 & n23977;
  assign n23979 = P1_INSTQUEUE_REG_11__2_ & n23630;
  assign n23980 = P1_INSTQUEUE_REG_10__2_ & n23633;
  assign n23981 = P1_INSTQUEUE_REG_9__2_ & n23636;
  assign n23982 = P1_INSTQUEUE_REG_8__2_ & n23639;
  assign n23983 = ~n23979 & ~n23980;
  assign n23984 = ~n23981 & n23983;
  assign n23985 = ~n23982 & n23984;
  assign n23986 = P1_INSTQUEUE_REG_6__2_ & n23646;
  assign n23987 = P1_INSTQUEUE_REG_5__2_ & n23650;
  assign n23988 = P1_INSTQUEUE_REG_4__2_ & n23653;
  assign n23989 = P1_INSTQUEUE_REG_3__2_ & n23657;
  assign n23990 = ~n23986 & ~n23987;
  assign n23991 = ~n23988 & n23990;
  assign n23992 = ~n23989 & n23991;
  assign n23993 = P1_INSTQUEUE_REG_2__2_ & n23663;
  assign n23994 = P1_INSTQUEUE_REG_1__2_ & n23666;
  assign n23995 = P1_INSTQUEUE_REG_0__2_ & n23668;
  assign n23996 = P1_INSTQUEUE_REG_7__2_ & n23671;
  assign n23997 = ~n23993 & ~n23994;
  assign n23998 = ~n23995 & n23997;
  assign n23999 = ~n23996 & n23998;
  assign n24000 = n23978 & n23985;
  assign n24001 = n23992 & n24000;
  assign n24002 = n23999 & n24001;
  assign n24003 = n23971 & n24002;
  assign n24004 = n23742 & n24003;
  assign n24005 = n23678 & ~n23709;
  assign n24006 = n23741 & ~n24002;
  assign n24007 = ~n23800 & n23968;
  assign n24008 = ~n23831 & n24007;
  assign n24009 = ~n23896 & n24008;
  assign n24010 = n24006 & n24009;
  assign n24011 = n24005 & n24010;
  assign n24012 = ~n24004 & ~n24011;
  assign n24013 = n23800 & n23896;
  assign n24014 = n24002 & n24009;
  assign n24015 = ~n23741 & n24014;
  assign n24016 = ~n24013 & ~n24015;
  assign n24017 = ~n23678 & ~n23741;
  assign n24018 = n23968 & n24017;
  assign n24019 = n24002 & n24018;
  assign n24020 = ~n24016 & n24019;
  assign n24021 = n24012 & ~n24020;
  assign n24022 = P1_INSTQUEUERD_ADDR_REG_4_ & ~P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n24023 = ~P1_INSTQUEUERD_ADDR_REG_3_ & P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n24024 = P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUEWR_ADDR_REG_3_;
  assign n24025 = ~P1_INSTQUEUERD_ADDR_REG_2_ & P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n24026 = P1_INSTQUEUERD_ADDR_REG_2_ & ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n24027 = P1_INSTQUEUERD_ADDR_REG_0_ & ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n24028 = P1_INSTQUEUEWR_ADDR_REG_1_ & ~n24027;
  assign n24029 = ~P1_INSTQUEUEWR_ADDR_REG_1_ & n24027;
  assign n24030 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~n24029;
  assign n24031 = ~n24028 & ~n24030;
  assign n24032 = ~n24026 & ~n24031;
  assign n24033 = ~n24025 & ~n24032;
  assign n24034 = ~n24024 & ~n24033;
  assign n24035 = ~n24023 & ~n24034;
  assign n24036 = ~P1_INSTQUEUERD_ADDR_REG_4_ & P1_INSTQUEUEWR_ADDR_REG_4_;
  assign n24037 = n24035 & ~n24036;
  assign n24038 = ~n24022 & ~n24037;
  assign n24039 = P1_STATE2_REG_0_ & ~n23968;
  assign n24040 = ~n23678 & n24039;
  assign n24041 = ~n24038 & n24040;
  assign n24042 = P1_STATE2_REG_0_ & n23896;
  assign n24043 = n23709 & n24042;
  assign n24044 = ~n24038 & n24043;
  assign n24045 = P1_STATE2_REG_0_ & n23678;
  assign n24046 = n23709 & n24045;
  assign n24047 = ~n23709 & n24045;
  assign n24048 = ~n23709 & n24042;
  assign n24049 = ~n23896 & n23968;
  assign n24050 = P1_STATE2_REG_0_ & n24049;
  assign n24051 = ~n23678 & ~n23709;
  assign n24052 = n24050 & n24051;
  assign n24053 = P1_STATE2_REG_0_ & ~n23896;
  assign n24054 = ~n23678 & n23709;
  assign n24055 = n24053 & n24054;
  assign n24056 = ~n24046 & ~n24047;
  assign n24057 = ~n24048 & n24056;
  assign n24058 = ~n24052 & n24057;
  assign n24059 = ~n24055 & n24058;
  assign n24060 = ~n24038 & ~n24059;
  assign n24061 = ~n24044 & ~n24060;
  assign n24062 = ~P1_STATE2_REG_0_ & P1_INSTQUEUERD_ADDR_REG_4_;
  assign n24063 = ~n24022 & ~n24036;
  assign n24064 = ~n24035 & ~n24063;
  assign n24065 = n24035 & n24063;
  assign n24066 = ~n24064 & ~n24065;
  assign n24067 = n24040 & ~n24066;
  assign n24068 = ~n24062 & ~n24067;
  assign n24069 = n24043 & ~n24066;
  assign n24070 = ~n24059 & ~n24066;
  assign n24071 = ~n24069 & ~n24070;
  assign n24072 = ~n24068 & n24071;
  assign n24073 = n24041 & n24061;
  assign n24074 = ~n24072 & ~n24073;
  assign n24075 = ~n24023 & ~n24024;
  assign n24076 = ~n24033 & ~n24075;
  assign n24077 = n24033 & n24075;
  assign n24078 = ~n24076 & ~n24077;
  assign n24079 = n24043 & ~n24078;
  assign n24080 = P1_STATE2_REG_0_ & ~n24079;
  assign n24081 = ~n24059 & ~n24078;
  assign n24082 = n24080 & ~n24081;
  assign n24083 = ~P1_STATE2_REG_0_ & P1_INSTQUEUERD_ADDR_REG_3_;
  assign n24084 = n24040 & ~n24078;
  assign n24085 = ~n24083 & ~n24084;
  assign n24086 = ~n24082 & n24085;
  assign n24087 = n24068 & ~n24071;
  assign n24088 = ~n24086 & ~n24087;
  assign n24089 = ~n24025 & ~n24026;
  assign n24090 = ~n24031 & ~n24089;
  assign n24091 = n24031 & n24089;
  assign n24092 = ~n24090 & ~n24091;
  assign n24093 = n24040 & ~n24092;
  assign n24094 = ~P1_STATE2_REG_0_ & P1_INSTQUEUERD_ADDR_REG_2_;
  assign n24095 = ~n24093 & ~n24094;
  assign n24096 = ~n24046 & ~n24053;
  assign n24097 = n23709 & ~n24096;
  assign n24098 = n24095 & ~n24097;
  assign n24099 = n24043 & ~n24092;
  assign n24100 = ~n23678 & ~n23968;
  assign n24101 = P1_STATE2_REG_0_ & ~n24100;
  assign n24102 = ~n24099 & n24101;
  assign n24103 = ~n24059 & ~n24092;
  assign n24104 = n24102 & ~n24103;
  assign n24105 = ~n24098 & n24104;
  assign n24106 = n24082 & ~n24085;
  assign n24107 = ~n24105 & ~n24106;
  assign n24108 = ~P1_INSTQUEUERD_ADDR_REG_1_ & P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n24109 = P1_INSTQUEUERD_ADDR_REG_1_ & ~P1_INSTQUEUEWR_ADDR_REG_1_;
  assign n24110 = ~n24108 & ~n24109;
  assign n24111 = ~n24027 & ~n24110;
  assign n24112 = n24027 & n24110;
  assign n24113 = ~n24111 & ~n24112;
  assign n24114 = n24043 & ~n24113;
  assign n24115 = P1_STATE2_REG_0_ & ~n24114;
  assign n24116 = ~n24059 & ~n24113;
  assign n24117 = n24115 & ~n24116;
  assign n24118 = ~P1_STATE2_REG_0_ & P1_INSTQUEUERD_ADDR_REG_1_;
  assign n24119 = n24040 & ~n24113;
  assign n24120 = P1_STATE2_REG_0_ & n23968;
  assign n24121 = ~n23709 & n24120;
  assign n24122 = ~n24042 & ~n24121;
  assign n24123 = ~n24118 & ~n24119;
  assign n24124 = n24122 & n24123;
  assign n24125 = ~n24047 & n24124;
  assign n24126 = ~n24117 & n24125;
  assign n24127 = n24098 & ~n24104;
  assign n24128 = ~n24126 & ~n24127;
  assign n24129 = n24117 & ~n24125;
  assign n24130 = ~P1_INSTQUEUERD_ADDR_REG_0_ & P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n24131 = ~n24027 & ~n24130;
  assign n24132 = n24043 & ~n24131;
  assign n24133 = n24101 & ~n24132;
  assign n24134 = ~n24059 & ~n24131;
  assign n24135 = n24133 & ~n24134;
  assign n24136 = ~n23709 & ~n23896;
  assign n24137 = n24040 & n24136;
  assign n24138 = n24135 & n24137;
  assign n24139 = ~P1_STATE2_REG_0_ & P1_INSTQUEUERD_ADDR_REG_0_;
  assign n24140 = n24040 & ~n24131;
  assign n24141 = ~n23678 & n24050;
  assign n24142 = ~n24139 & ~n24140;
  assign n24143 = ~n24141 & n24142;
  assign n24144 = ~n24097 & n24143;
  assign n24145 = n24135 & ~n24144;
  assign n24146 = n24137 & ~n24144;
  assign n24147 = ~n24129 & ~n24138;
  assign n24148 = ~n24145 & n24147;
  assign n24149 = ~n24146 & n24148;
  assign n24150 = n24128 & ~n24149;
  assign n24151 = n24107 & ~n24150;
  assign n24152 = n24088 & ~n24151;
  assign n24153 = n24074 & ~n24152;
  assign n24154 = ~n24041 & ~n24061;
  assign n24155 = ~n24153 & ~n24154;
  assign n24156 = ~n24061 & ~n24155;
  assign n24157 = P1_STATE2_REG_0_ & n24061;
  assign n24158 = ~n24156 & ~n24157;
  assign n24159 = n24041 & ~n24158;
  assign n24160 = n24061 & ~n24155;
  assign n24161 = ~P1_STATE2_REG_0_ & ~n24061;
  assign n24162 = ~n24160 & ~n24161;
  assign n24163 = ~n24041 & ~n24162;
  assign n24164 = ~n24159 & ~n24163;
  assign n24165 = ~n24021 & n24164;
  assign n24166 = ~n23709 & ~n23741;
  assign n24167 = ~n23678 & n24166;
  assign n24168 = n24003 & n24167;
  assign n24169 = ~n24164 & n24168;
  assign n24170 = n23710 & n24010;
  assign n24171 = n24066 & n24078;
  assign n24172 = n24113 & n24171;
  assign n24173 = n24092 & n24172;
  assign n24174 = n24038 & ~n24173;
  assign n24175 = n24170 & ~n24174;
  assign n24176 = ~n24165 & ~n24169;
  assign n24177 = ~n24175 & n24176;
  assign n24178 = ~n23831 & ~n24177;
  assign n24179 = ~n23678 & ~n24164;
  assign n24180 = n24015 & n24179;
  assign n24181 = n23968 & n24013;
  assign n24182 = ~n23741 & ~n23831;
  assign n24183 = n24002 & n24182;
  assign n24184 = n24181 & n24183;
  assign n24185 = ~n24164 & n24184;
  assign n24186 = ~n23678 & ~n24185;
  assign n24187 = n23709 & ~n24174;
  assign n24188 = n24010 & ~n24187;
  assign n24189 = n23678 & ~n24188;
  assign n24190 = ~n23709 & n24164;
  assign n24191 = ~n24186 & ~n24189;
  assign n24192 = ~n24190 & n24191;
  assign n24193 = P1_STATE_REG_2_ & ~P1_STATE_REG_1_;
  assign n24194 = ~n23520 & ~n24193;
  assign n24195 = ~P1_STATE_REG_0_ & ~n24194;
  assign n24196 = ~n24051 & ~n24195;
  assign n24197 = ~n23710 & n24196;
  assign n24198 = ~n23523 & ~n24197;
  assign n24199 = n24192 & ~n24198;
  assign n24200 = ~P1_FLUSH_REG & ~P1_MORE_REG;
  assign n24201 = n24199 & ~n24200;
  assign n24202 = P1_STATE2_REG_1_ & ~P1_FLUSH_REG;
  assign n24203 = P1_INSTQUEUERD_ADDR_REG_2_ & n24202;
  assign n24204 = P1_INSTADDRPOINTER_REG_0_ & P1_INSTADDRPOINTER_REG_31_;
  assign n24205 = P1_INSTADDRPOINTER_REG_0_ & ~P1_INSTADDRPOINTER_REG_31_;
  assign n24206 = ~n24204 & ~n24205;
  assign n24207 = P1_STATE2_REG_1_ & ~n24206;
  assign n24208 = P1_INSTADDRPOINTER_REG_0_ & ~P1_INSTADDRPOINTER_REG_1_;
  assign n24209 = ~P1_INSTADDRPOINTER_REG_0_ & P1_INSTADDRPOINTER_REG_1_;
  assign n24210 = ~n24208 & ~n24209;
  assign n24211 = P1_INSTADDRPOINTER_REG_31_ & ~n24210;
  assign n24212 = P1_INSTADDRPOINTER_REG_1_ & ~P1_INSTADDRPOINTER_REG_31_;
  assign n24213 = ~n24211 & ~n24212;
  assign n24214 = P1_FLUSH_REG & n24207;
  assign n24215 = ~n24213 & n24214;
  assign n24216 = ~n24203 & ~n24215;
  assign n24217 = n23741 & n24002;
  assign n24218 = n23678 & n24217;
  assign n24219 = n23709 & n23971;
  assign n24220 = n24218 & n24219;
  assign n24221 = P1_INSTQUEUERD_ADDR_REG_2_ & ~n23655;
  assign n24222 = ~n23856 & ~n24221;
  assign n24223 = n24220 & ~n24222;
  assign n24224 = ~n24004 & ~n24168;
  assign n24225 = n24222 & ~n24224;
  assign n24226 = ~n23848 & ~n23855;
  assign n24227 = n24011 & ~n24226;
  assign n24228 = ~n24223 & ~n24225;
  assign n24229 = ~n24227 & n24228;
  assign n24230 = P1_STATE2_REG_0_ & ~n23678;
  assign n24231 = n23709 & ~n24194;
  assign n24232 = n24230 & n24231;
  assign n24233 = P1_STATE2_REG_0_ & n24051;
  assign n24234 = ~n24232 & ~n24233;
  assign n24235 = n24184 & ~n24234;
  assign n24236 = P1_STATE2_REG_0_ & n23710;
  assign n24237 = n24006 & n24236;
  assign n24238 = n24009 & n24237;
  assign n24239 = ~n24235 & ~n24238;
  assign n24240 = ~n23800 & ~n23831;
  assign n24241 = n24043 & n24240;
  assign n24242 = n24218 & n24241;
  assign n24243 = n24239 & ~n24242;
  assign n24244 = ~n24002 & n24013;
  assign n24245 = n23831 & n24244;
  assign n24246 = n23968 & n24245;
  assign n24247 = P1_STATE2_REG_0_ & n24246;
  assign n24248 = n23896 & n23968;
  assign n24249 = n23831 & ~n24248;
  assign n24250 = ~n23800 & n23896;
  assign n24251 = n23800 & ~n23968;
  assign n24252 = ~n24250 & ~n24251;
  assign n24253 = n24002 & n24252;
  assign n24254 = ~n23741 & ~n23971;
  assign n24255 = ~n24249 & ~n24253;
  assign n24256 = ~n24254 & n24255;
  assign n24257 = n24046 & ~n24256;
  assign n24258 = ~n23968 & n23969;
  assign n24259 = n24217 & n24258;
  assign n24260 = n24046 & n24259;
  assign n24261 = ~n24235 & ~n24247;
  assign n24262 = ~n24257 & n24261;
  assign n24263 = ~n24260 & n24262;
  assign n24264 = n23968 & ~n24250;
  assign n24265 = ~n23969 & n24264;
  assign n24266 = ~n24002 & ~n24265;
  assign n24267 = n24046 & n24266;
  assign n24268 = n23678 & ~n24166;
  assign n24269 = ~n24002 & ~n24268;
  assign n24270 = ~n23869 & ~n23872;
  assign n24271 = ~n23866 & n24270;
  assign n24272 = ~n23875 & ~n23881;
  assign n24273 = ~n23884 & n24272;
  assign n24274 = ~n23889 & n24273;
  assign n24275 = n23894 & n24271;
  assign n24276 = n24274 & n24275;
  assign n24277 = n23800 & ~n24276;
  assign n24278 = ~n23831 & n23968;
  assign n24279 = ~n24250 & ~n24277;
  assign n24280 = n24278 & n24279;
  assign n24281 = n24054 & ~n24280;
  assign n24282 = ~n24269 & ~n24281;
  assign n24283 = P1_STATE2_REG_0_ & ~n24282;
  assign n24284 = n24009 & n24166;
  assign n24285 = P1_STATE2_REG_0_ & n24284;
  assign n24286 = n23709 & n24002;
  assign n24287 = n23896 & n24286;
  assign n24288 = n23678 & n24287;
  assign n24289 = n23741 & n24288;
  assign n24290 = ~n23968 & n24240;
  assign n24291 = n24289 & n24290;
  assign n24292 = P1_STATE2_REG_0_ & n24291;
  assign n24293 = ~n24267 & ~n24283;
  assign n24294 = ~n24285 & n24293;
  assign n24295 = ~n24292 & n24294;
  assign n24296 = P1_STATE2_REG_0_ & n24167;
  assign n24297 = n23800 & ~n23896;
  assign n24298 = ~n23968 & ~n24297;
  assign n24299 = n23800 & n24049;
  assign n24300 = ~n23831 & ~n24250;
  assign n24301 = ~n24299 & n24300;
  assign n24302 = ~n24298 & n24301;
  assign n24303 = n24296 & ~n24302;
  assign n24304 = ~n23678 & n23741;
  assign n24305 = P1_STATE2_REG_0_ & n24304;
  assign n24306 = ~n24238 & ~n24305;
  assign n24307 = ~P1_STATE2_REG_3_ & ~P1_STATE2_REG_1_;
  assign n24308 = ~P1_STATE2_REG_0_ & n24307;
  assign n24309 = ~P1_INSTQUEUEWR_ADDR_REG_1_ & P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n24310 = P1_INSTQUEUEWR_ADDR_REG_1_ & ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = n24308 & ~n24311;
  assign n24313 = P1_STATE2_REG_2_ & ~P1_STATE2_REG_1_;
  assign n24314 = P1_INSTQUEUEWR_ADDR_REG_1_ & ~n24313;
  assign n24315 = ~n24312 & ~n24314;
  assign n24316 = n23831 & n23968;
  assign n24317 = n24250 & n24316;
  assign n24318 = n24218 & n24317;
  assign n24319 = P1_STATE2_REG_0_ & n24318;
  assign n24320 = n23968 & n24240;
  assign n24321 = n24289 & n24320;
  assign n24322 = P1_STATE2_REG_0_ & n24321;
  assign n24323 = n24315 & ~n24319;
  assign n24324 = ~n24322 & n24323;
  assign n24325 = ~n24047 & ~n24303;
  assign n24326 = n24306 & n24325;
  assign n24327 = n24324 & n24326;
  assign n24328 = n24263 & n24295;
  assign n24329 = n24327 & n24328;
  assign n24330 = ~P1_INSTQUEUERD_ADDR_REG_1_ & ~n24314;
  assign n24331 = ~n24312 & n24330;
  assign n24332 = ~n24329 & ~n24331;
  assign n24333 = ~n24243 & n24332;
  assign n24334 = n24256 & ~n24266;
  assign n24335 = n23709 & ~n24334;
  assign n24336 = ~n23709 & ~n24049;
  assign n24337 = ~n24335 & ~n24336;
  assign n24338 = n23678 & ~n24337;
  assign n24339 = ~n23678 & ~n24002;
  assign n24340 = P1_STATE2_REG_0_ & n24307;
  assign n24341 = n23968 & ~n24297;
  assign n24342 = n24182 & n24341;
  assign n24343 = ~n24250 & n24342;
  assign n24344 = n24054 & ~n24343;
  assign n24345 = n24340 & ~n24344;
  assign n24346 = ~n24258 & ~n24317;
  assign n24347 = n24218 & ~n24346;
  assign n24348 = n23741 & n24246;
  assign n24349 = ~n24284 & ~n24347;
  assign n24350 = ~n24348 & n24349;
  assign n24351 = ~n23678 & ~n24217;
  assign n24352 = n24302 & n24351;
  assign n24353 = ~n23709 & ~n24352;
  assign n24354 = n24350 & ~n24353;
  assign n24355 = ~n24338 & ~n24339;
  assign n24356 = n24345 & n24355;
  assign n24357 = n24354 & n24356;
  assign n24358 = ~n24303 & ~n24305;
  assign n24359 = ~n24259 & ~n24266;
  assign n24360 = n24256 & n24359;
  assign n24361 = n24046 & ~n24360;
  assign n24362 = ~n24047 & ~n24319;
  assign n24363 = ~n24322 & n24362;
  assign n24364 = P1_INSTQUEUEWR_ADDR_REG_0_ & ~n24313;
  assign n24365 = ~P1_INSTQUEUEWR_ADDR_REG_0_ & n24308;
  assign n24366 = ~n24364 & ~n24365;
  assign n24367 = ~n24247 & ~n24285;
  assign n24368 = ~n24292 & n24367;
  assign n24369 = ~n24283 & n24366;
  assign n24370 = n24239 & n24369;
  assign n24371 = n24368 & n24370;
  assign n24372 = n24358 & ~n24361;
  assign n24373 = n24363 & n24372;
  assign n24374 = n24371 & n24373;
  assign n24375 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n24366;
  assign n24376 = ~n24374 & ~n24375;
  assign n24377 = ~n24357 & n24376;
  assign n24378 = n24243 & ~n24332;
  assign n24379 = n24377 & ~n24378;
  assign n24380 = ~n24333 & ~n24379;
  assign n24381 = P1_INSTQUEUEWR_ADDR_REG_1_ & P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n24382 = ~P1_INSTQUEUEWR_ADDR_REG_2_ & n24381;
  assign n24383 = P1_INSTQUEUEWR_ADDR_REG_2_ & ~n24381;
  assign n24384 = ~n24382 & ~n24383;
  assign n24385 = n24308 & ~n24384;
  assign n24386 = P1_INSTQUEUEWR_ADDR_REG_2_ & ~n24313;
  assign n24387 = ~n24385 & ~n24386;
  assign n24388 = n24239 & ~n24283;
  assign n24389 = n24368 & n24388;
  assign n24390 = n24373 & n24389;
  assign n24391 = n24387 & n24390;
  assign n24392 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~n24386;
  assign n24393 = ~n24385 & n24392;
  assign n24394 = ~n24391 & ~n24393;
  assign n24395 = n24380 & ~n24394;
  assign n24396 = ~n24380 & n24394;
  assign n24397 = ~n24395 & ~n24396;
  assign n24398 = ~n24289 & ~n24348;
  assign n24399 = ~n23709 & n23831;
  assign n24400 = ~n24318 & ~n24399;
  assign n24401 = ~n24170 & ~n24284;
  assign n24402 = n24398 & n24401;
  assign n24403 = n24400 & n24402;
  assign n24404 = ~n24184 & n24403;
  assign n24405 = n24166 & ~n24301;
  assign n24406 = ~n24297 & n24300;
  assign n24407 = n24054 & ~n24406;
  assign n24408 = ~n24304 & ~n24407;
  assign n24409 = n23800 & ~n24002;
  assign n24410 = ~n24218 & ~n24409;
  assign n24411 = ~n23709 & ~n24410;
  assign n24412 = n24100 & ~n24297;
  assign n24413 = ~n24411 & ~n24412;
  assign n24414 = ~n24269 & ~n24405;
  assign n24415 = n24408 & n24414;
  assign n24416 = n24413 & n24415;
  assign n24417 = ~n24338 & n24416;
  assign n24418 = n24404 & n24417;
  assign n24419 = n24397 & ~n24418;
  assign n24420 = n24229 & ~n24419;
  assign n24421 = ~n23523 & n24051;
  assign n24422 = n24184 & n24421;
  assign n24423 = ~n24004 & ~n24422;
  assign n24424 = ~n23523 & n24195;
  assign n24425 = ~n24011 & ~n24184;
  assign n24426 = n24424 & ~n24425;
  assign n24427 = n24423 & ~n24426;
  assign n24428 = ~n24164 & ~n24427;
  assign n24429 = n24164 & n24168;
  assign n24430 = n24002 & n24005;
  assign n24431 = ~n24412 & ~n24430;
  assign n24432 = ~n23523 & n24170;
  assign n24433 = n24174 & n24432;
  assign n24434 = n24431 & ~n24433;
  assign n24435 = n23678 & n23741;
  assign n24436 = n24009 & n24435;
  assign n24437 = ~n24002 & ~n24436;
  assign n24438 = n23678 & ~n23971;
  assign n24439 = ~n23741 & ~n24438;
  assign n24440 = n24301 & n24439;
  assign n24441 = n24002 & ~n24440;
  assign n24442 = ~n24437 & ~n24441;
  assign n24443 = ~n24407 & n24442;
  assign n24444 = n24434 & n24443;
  assign n24445 = ~n24428 & ~n24429;
  assign n24446 = n24444 & n24445;
  assign n24447 = ~n24420 & ~n24446;
  assign n24448 = P1_INSTQUEUERD_ADDR_REG_2_ & n24446;
  assign n24449 = ~n24447 & ~n24448;
  assign n24450 = ~P1_STATE2_REG_1_ & ~n24449;
  assign n24451 = n24216 & ~n24450;
  assign n24452 = P1_INSTQUEUERD_ADDR_REG_4_ & n24446;
  assign n24453 = P1_STATE2_REG_0_ & n24005;
  assign n24454 = n24010 & n24453;
  assign n24455 = ~n24238 & ~n24454;
  assign n24456 = P1_INSTQUEUERD_ADDR_REG_4_ & ~n24455;
  assign n24457 = P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n24458 = P1_INSTQUEUEWR_ADDR_REG_3_ & ~n24381;
  assign n24459 = ~P1_INSTQUEUEWR_ADDR_REG_3_ & P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n24460 = n24381 & n24459;
  assign n24461 = ~n24457 & ~n24458;
  assign n24462 = ~n24460 & n24461;
  assign n24463 = n24308 & ~n24462;
  assign n24464 = P1_INSTQUEUEWR_ADDR_REG_3_ & ~n24313;
  assign n24465 = ~n24463 & ~n24464;
  assign n24466 = P1_INSTQUEUERD_ADDR_REG_3_ & ~n24390;
  assign n24467 = n24465 & ~n24466;
  assign n24468 = n24394 & ~n24467;
  assign n24469 = ~n24380 & n24468;
  assign n24470 = n24456 & ~n24469;
  assign n24471 = ~n24456 & n24469;
  assign n24472 = ~n24470 & ~n24471;
  assign n24473 = n24170 & ~n24472;
  assign n24474 = ~n24446 & n24473;
  assign n24475 = ~n24452 & ~n24474;
  assign n24476 = ~P1_STATE2_REG_1_ & ~n24475;
  assign n24477 = P1_INSTQUEUERD_ADDR_REG_4_ & n24202;
  assign n24478 = ~n24476 & ~n24477;
  assign n24479 = n24451 & n24478;
  assign n24480 = n24396 & n24467;
  assign n24481 = ~n24396 & ~n24467;
  assign n24482 = ~n24480 & ~n24481;
  assign n24483 = ~n24418 & ~n24482;
  assign n24484 = P1_INSTQUEUERD_ADDR_REG_3_ & ~n23644;
  assign n24485 = ~n23887 & ~n24484;
  assign n24486 = n24011 & ~n24485;
  assign n24487 = P1_INSTQUEUERD_ADDR_REG_3_ & ~n23670;
  assign n24488 = ~n23671 & ~n24487;
  assign n24489 = n24220 & ~n24488;
  assign n24490 = ~n24486 & ~n24489;
  assign n24491 = ~n23655 & n23656;
  assign n24492 = ~P1_INSTQUEUERD_ADDR_REG_2_ & ~n23655;
  assign n24493 = P1_INSTQUEUERD_ADDR_REG_3_ & ~n24492;
  assign n24494 = ~n24491 & ~n24493;
  assign n24495 = ~n24224 & n24494;
  assign n24496 = n24490 & ~n24495;
  assign n24497 = ~n24483 & n24496;
  assign n24498 = ~n24446 & ~n24497;
  assign n24499 = P1_INSTQUEUERD_ADDR_REG_3_ & n24446;
  assign n24500 = ~n24498 & ~n24499;
  assign n24501 = ~P1_STATE2_REG_1_ & ~n24500;
  assign n24502 = P1_INSTQUEUERD_ADDR_REG_3_ & n24202;
  assign n24503 = ~n24501 & ~n24502;
  assign n24504 = n24478 & n24503;
  assign n24505 = ~n24479 & ~n24504;
  assign n24506 = ~P1_INSTQUEUEWR_ADDR_REG_4_ & ~n24475;
  assign n24507 = P1_INSTQUEUEWR_ADDR_REG_3_ & n24500;
  assign n24508 = P1_INSTQUEUEWR_ADDR_REG_4_ & n24475;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = ~P1_INSTQUEUEWR_ADDR_REG_2_ & ~n24449;
  assign n24511 = ~P1_INSTQUEUEWR_ADDR_REG_3_ & ~n24500;
  assign n24512 = ~n24510 & ~n24511;
  assign n24513 = n23710 & n24003;
  assign n24514 = ~n24168 & ~n24513;
  assign n24515 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~n24514;
  assign n24516 = P1_INSTQUEUERD_ADDR_REG_0_ & n24011;
  assign n24517 = ~n24515 & ~n24516;
  assign n24518 = n24357 & n24376;
  assign n24519 = ~n24357 & ~n24376;
  assign n24520 = ~n24518 & ~n24519;
  assign n24521 = ~n24418 & ~n24520;
  assign n24522 = n24517 & ~n24521;
  assign n24523 = ~n24446 & ~n24522;
  assign n24524 = P1_INSTQUEUERD_ADDR_REG_0_ & n24446;
  assign n24525 = ~n24523 & ~n24524;
  assign n24526 = n24381 & n24525;
  assign n24527 = P1_INSTQUEUEWR_ADDR_REG_2_ & n24449;
  assign n24528 = ~P1_INSTQUEUERD_ADDR_REG_1_ & n24011;
  assign n24529 = ~n23624 & ~n23655;
  assign n24530 = ~n24514 & n24529;
  assign n24531 = ~n24528 & ~n24530;
  assign n24532 = ~n24333 & ~n24378;
  assign n24533 = ~n24377 & n24532;
  assign n24534 = n24377 & ~n24532;
  assign n24535 = ~n24533 & ~n24534;
  assign n24536 = ~n24418 & ~n24535;
  assign n24537 = n24531 & ~n24536;
  assign n24538 = ~n24446 & ~n24537;
  assign n24539 = P1_INSTQUEUERD_ADDR_REG_1_ & n24446;
  assign n24540 = ~n24538 & ~n24539;
  assign n24541 = P1_INSTQUEUEWR_ADDR_REG_1_ & n24540;
  assign n24542 = n24525 & n24540;
  assign n24543 = P1_INSTQUEUEWR_ADDR_REG_0_ & n24542;
  assign n24544 = ~n24526 & ~n24527;
  assign n24545 = ~n24541 & n24544;
  assign n24546 = ~n24543 & n24545;
  assign n24547 = n24512 & ~n24546;
  assign n24548 = n24509 & ~n24547;
  assign n24549 = ~n24506 & ~n24548;
  assign n24550 = ~n24178 & ~n24180;
  assign n24551 = ~n24201 & n24550;
  assign n24552 = ~n24505 & n24551;
  assign n24553 = n24549 & n24552;
  assign n24554 = ~P1_STATE2_REG_1_ & n24553;
  assign n24555 = P1_STATE2_REG_0_ & ~n24554;
  assign n24556 = ~P1_STATEBS16_REG & ~n23523;
  assign n24557 = n24054 & n24556;
  assign n24558 = ~n24164 & n24195;
  assign n24559 = n24184 & n24557;
  assign n24560 = n24558 & n24559;
  assign n24561 = P1_STATE2_REG_2_ & ~n24560;
  assign n24562 = ~n23611 & ~n24555;
  assign n24563 = n24561 & n24562;
  assign n24564 = P1_STATE2_REG_0_ & ~n24563;
  assign n24565 = n23609 & n24564;
  assign n24566 = P1_STATE2_REG_3_ & ~n24564;
  assign n5379 = n24565 | n24566;
  assign n24568 = ~P1_STATE2_REG_2_ & ~n23523;
  assign n24569 = P1_STATE2_REG_0_ & ~n24568;
  assign n24570 = ~P1_STATE2_REG_0_ & ~P1_STATEBS16_REG;
  assign n24571 = ~n24569 & ~n24570;
  assign n24572 = P1_STATE2_REG_1_ & n24571;
  assign n24573 = ~n24313 & ~n24572;
  assign n24574 = P1_STATE2_REG_2_ & ~n24564;
  assign n5384 = ~n24573 | n24574;
  assign n24576 = P1_STATE2_REG_0_ & n24313;
  assign n24577 = ~n24563 & n24576;
  assign n24578 = ~P1_STATE2_REG_2_ & P1_STATE2_REG_0_;
  assign n24579 = n23523 & n24578;
  assign n24580 = ~n24563 & ~n24579;
  assign n24581 = P1_STATE2_REG_1_ & ~n24580;
  assign n24582 = ~n23523 & n24307;
  assign n24583 = n24564 & n24582;
  assign n24584 = ~P1_STATE2_REG_2_ & ~P1_STATEBS16_REG;
  assign n24585 = P1_STATE2_REG_1_ & ~P1_STATE2_REG_0_;
  assign n24586 = n24584 & n24585;
  assign n24587 = ~n24577 & ~n24581;
  assign n24588 = ~n24583 & n24587;
  assign n5389 = n24586 | ~n24588;
  assign n24590 = P1_STATE2_REG_3_ & ~n24164;
  assign n24591 = ~P1_STATE2_REG_2_ & ~P1_STATE2_REG_1_;
  assign n24592 = n24590 & n24591;
  assign n24593 = ~n24563 & ~n24592;
  assign n24594 = ~P1_STATE2_REG_0_ & n24593;
  assign n24595 = P1_FLUSH_REG & n24206;
  assign n24596 = P1_STATE2_REG_1_ & n24595;
  assign n24597 = ~P1_STATE2_REG_1_ & ~n24525;
  assign n24598 = P1_INSTQUEUERD_ADDR_REG_0_ & n24202;
  assign n24599 = ~n24596 & ~n24597;
  assign n24600 = ~n24598 & n24599;
  assign n24601 = P1_INSTQUEUERD_ADDR_REG_1_ & n24202;
  assign n24602 = n24213 & n24214;
  assign n24603 = ~n24601 & ~n24602;
  assign n24604 = ~P1_STATE2_REG_1_ & ~n24540;
  assign n24605 = n24603 & ~n24604;
  assign n24606 = n24600 & n24605;
  assign n24607 = ~n24451 & ~n24606;
  assign n24608 = ~n24503 & n24607;
  assign n24609 = n24478 & ~n24608;
  assign n24610 = n23609 & n24609;
  assign n24611 = ~n24563 & ~n24610;
  assign n24612 = P1_STATE2_REG_0_ & ~n24611;
  assign n24613 = P1_STATE2_REG_3_ & P1_STATE2_REG_0_;
  assign n24614 = n24591 & n24613;
  assign n24615 = ~n24579 & ~n24614;
  assign n24616 = ~n24553 & n24576;
  assign n24617 = n24615 & ~n24616;
  assign n24618 = ~n24594 & ~n24612;
  assign n5394 = ~n24617 | ~n24618;
  assign n24620 = P1_INSTQUEUEWR_ADDR_REG_3_ & P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n24621 = n24381 & n24620;
  assign n24622 = n24397 & ~n24482;
  assign n24623 = ~n24520 & ~n24535;
  assign n24624 = n24622 & n24623;
  assign n24625 = ~n24621 & ~n24624;
  assign n24626 = ~P1_STATE2_REG_3_ & ~P1_STATE2_REG_2_;
  assign n24627 = ~P1_STATEBS16_REG & n24626;
  assign n24628 = n24222 & n24488;
  assign n24629 = P1_INSTQUEUERD_ADDR_REG_0_ & ~n24529;
  assign n24630 = n24628 & n24629;
  assign n24631 = P1_INSTQUEUE_REG_0__7_ & n24630;
  assign n24632 = ~P1_INSTQUEUERD_ADDR_REG_0_ & ~n24529;
  assign n24633 = n24628 & n24632;
  assign n24634 = P1_INSTQUEUE_REG_1__7_ & n24633;
  assign n24635 = P1_INSTQUEUERD_ADDR_REG_0_ & n24529;
  assign n24636 = n24628 & n24635;
  assign n24637 = P1_INSTQUEUE_REG_2__7_ & n24636;
  assign n24638 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n24529;
  assign n24639 = n24628 & n24638;
  assign n24640 = P1_INSTQUEUE_REG_3__7_ & n24639;
  assign n24641 = ~n24631 & ~n24634;
  assign n24642 = ~n24637 & n24641;
  assign n24643 = ~n24640 & n24642;
  assign n24644 = ~n24222 & n24488;
  assign n24645 = n24629 & n24644;
  assign n24646 = P1_INSTQUEUE_REG_4__7_ & n24645;
  assign n24647 = n24632 & n24644;
  assign n24648 = P1_INSTQUEUE_REG_5__7_ & n24647;
  assign n24649 = n24635 & n24644;
  assign n24650 = P1_INSTQUEUE_REG_6__7_ & n24649;
  assign n24651 = n24638 & n24644;
  assign n24652 = P1_INSTQUEUE_REG_7__7_ & n24651;
  assign n24653 = ~n24646 & ~n24648;
  assign n24654 = ~n24650 & n24653;
  assign n24655 = ~n24652 & n24654;
  assign n24656 = n24222 & ~n24488;
  assign n24657 = n24629 & n24656;
  assign n24658 = P1_INSTQUEUE_REG_8__7_ & n24657;
  assign n24659 = n24632 & n24656;
  assign n24660 = P1_INSTQUEUE_REG_9__7_ & n24659;
  assign n24661 = n24635 & n24656;
  assign n24662 = P1_INSTQUEUE_REG_10__7_ & n24661;
  assign n24663 = n24638 & n24656;
  assign n24664 = P1_INSTQUEUE_REG_11__7_ & n24663;
  assign n24665 = ~n24658 & ~n24660;
  assign n24666 = ~n24662 & n24665;
  assign n24667 = ~n24664 & n24666;
  assign n24668 = ~n24222 & ~n24488;
  assign n24669 = n24629 & n24668;
  assign n24670 = P1_INSTQUEUE_REG_12__7_ & n24669;
  assign n24671 = n24632 & n24668;
  assign n24672 = P1_INSTQUEUE_REG_13__7_ & n24671;
  assign n24673 = n24635 & n24668;
  assign n24674 = P1_INSTQUEUE_REG_14__7_ & n24673;
  assign n24675 = n24638 & n24668;
  assign n24676 = P1_INSTQUEUE_REG_15__7_ & n24675;
  assign n24677 = ~n24670 & ~n24672;
  assign n24678 = ~n24674 & n24677;
  assign n24679 = ~n24676 & n24678;
  assign n24680 = n24643 & n24655;
  assign n24681 = n24667 & n24680;
  assign n24682 = n24679 & n24681;
  assign n24683 = n24120 & ~n24682;
  assign n24684 = ~P1_STATE2_REG_0_ & ~n24520;
  assign n24685 = n24120 & n24682;
  assign n24686 = P1_INSTQUEUE_REG_0__0_ & n24630;
  assign n24687 = P1_INSTQUEUE_REG_1__0_ & n24633;
  assign n24688 = P1_INSTQUEUE_REG_2__0_ & n24636;
  assign n24689 = P1_INSTQUEUE_REG_3__0_ & n24639;
  assign n24690 = ~n24686 & ~n24687;
  assign n24691 = ~n24688 & n24690;
  assign n24692 = ~n24689 & n24691;
  assign n24693 = P1_INSTQUEUE_REG_4__0_ & n24645;
  assign n24694 = P1_INSTQUEUE_REG_5__0_ & n24647;
  assign n24695 = P1_INSTQUEUE_REG_6__0_ & n24649;
  assign n24696 = P1_INSTQUEUE_REG_7__0_ & n24651;
  assign n24697 = ~n24693 & ~n24694;
  assign n24698 = ~n24695 & n24697;
  assign n24699 = ~n24696 & n24698;
  assign n24700 = P1_INSTQUEUE_REG_8__0_ & n24657;
  assign n24701 = P1_INSTQUEUE_REG_9__0_ & n24659;
  assign n24702 = P1_INSTQUEUE_REG_10__0_ & n24661;
  assign n24703 = P1_INSTQUEUE_REG_11__0_ & n24663;
  assign n24704 = ~n24700 & ~n24701;
  assign n24705 = ~n24702 & n24704;
  assign n24706 = ~n24703 & n24705;
  assign n24707 = P1_INSTQUEUE_REG_12__0_ & n24669;
  assign n24708 = P1_INSTQUEUE_REG_13__0_ & n24671;
  assign n24709 = P1_INSTQUEUE_REG_14__0_ & n24673;
  assign n24710 = P1_INSTQUEUE_REG_15__0_ & n24675;
  assign n24711 = ~n24707 & ~n24708;
  assign n24712 = ~n24709 & n24711;
  assign n24713 = ~n24710 & n24712;
  assign n24714 = n24692 & n24699;
  assign n24715 = n24706 & n24714;
  assign n24716 = n24713 & n24715;
  assign n24717 = n24685 & ~n24716;
  assign n24718 = n24683 & n24716;
  assign n24719 = ~n24684 & ~n24717;
  assign n24720 = ~n24718 & n24719;
  assign n24721 = ~n24683 & ~n24720;
  assign n24722 = n24683 & n24720;
  assign n24723 = P1_INSTQUEUE_REG_0__0_ & n24040;
  assign n24724 = P1_STATE2_REG_0_ & ~n24723;
  assign n24725 = n24045 & ~n24716;
  assign n24726 = n23968 & ~n24682;
  assign n24727 = n24724 & ~n24725;
  assign n24728 = ~n24726 & n24727;
  assign n24729 = ~n24721 & ~n24722;
  assign n24730 = n24728 & n24729;
  assign n24731 = n24683 & ~n24730;
  assign n24732 = ~n24728 & ~n24729;
  assign n24733 = ~n24731 & ~n24732;
  assign n24734 = ~P1_STATE2_REG_0_ & ~n24535;
  assign n24735 = P1_INSTQUEUE_REG_0__1_ & n24630;
  assign n24736 = P1_INSTQUEUE_REG_1__1_ & n24633;
  assign n24737 = P1_INSTQUEUE_REG_2__1_ & n24636;
  assign n24738 = P1_INSTQUEUE_REG_3__1_ & n24639;
  assign n24739 = ~n24735 & ~n24736;
  assign n24740 = ~n24737 & n24739;
  assign n24741 = ~n24738 & n24740;
  assign n24742 = P1_INSTQUEUE_REG_4__1_ & n24645;
  assign n24743 = P1_INSTQUEUE_REG_5__1_ & n24647;
  assign n24744 = P1_INSTQUEUE_REG_6__1_ & n24649;
  assign n24745 = P1_INSTQUEUE_REG_7__1_ & n24651;
  assign n24746 = ~n24742 & ~n24743;
  assign n24747 = ~n24744 & n24746;
  assign n24748 = ~n24745 & n24747;
  assign n24749 = P1_INSTQUEUE_REG_8__1_ & n24657;
  assign n24750 = P1_INSTQUEUE_REG_9__1_ & n24659;
  assign n24751 = P1_INSTQUEUE_REG_10__1_ & n24661;
  assign n24752 = P1_INSTQUEUE_REG_11__1_ & n24663;
  assign n24753 = ~n24749 & ~n24750;
  assign n24754 = ~n24751 & n24753;
  assign n24755 = ~n24752 & n24754;
  assign n24756 = P1_INSTQUEUE_REG_12__1_ & n24669;
  assign n24757 = P1_INSTQUEUE_REG_13__1_ & n24671;
  assign n24758 = P1_INSTQUEUE_REG_14__1_ & n24673;
  assign n24759 = P1_INSTQUEUE_REG_15__1_ & n24675;
  assign n24760 = ~n24756 & ~n24757;
  assign n24761 = ~n24758 & n24760;
  assign n24762 = ~n24759 & n24761;
  assign n24763 = n24741 & n24748;
  assign n24764 = n24755 & n24763;
  assign n24765 = n24762 & n24764;
  assign n24766 = n24685 & ~n24765;
  assign n24767 = n24683 & n24765;
  assign n24768 = ~n24734 & ~n24766;
  assign n24769 = ~n24767 & n24768;
  assign n24770 = ~n24683 & ~n24769;
  assign n24771 = n24683 & n24769;
  assign n24772 = ~n24770 & ~n24771;
  assign n24773 = P1_INSTQUEUE_REG_0__1_ & n24040;
  assign n24774 = ~n24685 & ~n24773;
  assign n24775 = n24045 & ~n24765;
  assign n24776 = n24774 & ~n24775;
  assign n24777 = ~n24772 & n24776;
  assign n24778 = n24772 & ~n24776;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 = n24733 & ~n24779;
  assign n24781 = ~n24733 & n24779;
  assign n24782 = ~n24780 & ~n24781;
  assign n24783 = ~n24730 & ~n24732;
  assign n24784 = ~n24683 & n24783;
  assign n24785 = n24683 & ~n24783;
  assign n24786 = ~n24784 & ~n24785;
  assign n24787 = ~n24782 & n24786;
  assign n24788 = n24782 & ~n24786;
  assign n24789 = ~n24787 & ~n24788;
  assign n24790 = n24786 & ~n24789;
  assign n24791 = ~n24782 & ~n24786;
  assign n24792 = P1_INSTQUEUE_REG_0__2_ & n24040;
  assign n24793 = P1_INSTQUEUE_REG_0__2_ & n24630;
  assign n24794 = P1_INSTQUEUE_REG_1__2_ & n24633;
  assign n24795 = P1_INSTQUEUE_REG_2__2_ & n24636;
  assign n24796 = P1_INSTQUEUE_REG_3__2_ & n24639;
  assign n24797 = ~n24793 & ~n24794;
  assign n24798 = ~n24795 & n24797;
  assign n24799 = ~n24796 & n24798;
  assign n24800 = P1_INSTQUEUE_REG_4__2_ & n24645;
  assign n24801 = P1_INSTQUEUE_REG_5__2_ & n24647;
  assign n24802 = P1_INSTQUEUE_REG_6__2_ & n24649;
  assign n24803 = P1_INSTQUEUE_REG_7__2_ & n24651;
  assign n24804 = ~n24800 & ~n24801;
  assign n24805 = ~n24802 & n24804;
  assign n24806 = ~n24803 & n24805;
  assign n24807 = P1_INSTQUEUE_REG_8__2_ & n24657;
  assign n24808 = P1_INSTQUEUE_REG_9__2_ & n24659;
  assign n24809 = P1_INSTQUEUE_REG_10__2_ & n24661;
  assign n24810 = P1_INSTQUEUE_REG_11__2_ & n24663;
  assign n24811 = ~n24807 & ~n24808;
  assign n24812 = ~n24809 & n24811;
  assign n24813 = ~n24810 & n24812;
  assign n24814 = P1_INSTQUEUE_REG_12__2_ & n24669;
  assign n24815 = P1_INSTQUEUE_REG_13__2_ & n24671;
  assign n24816 = P1_INSTQUEUE_REG_14__2_ & n24673;
  assign n24817 = P1_INSTQUEUE_REG_15__2_ & n24675;
  assign n24818 = ~n24814 & ~n24815;
  assign n24819 = ~n24816 & n24818;
  assign n24820 = ~n24817 & n24819;
  assign n24821 = n24799 & n24806;
  assign n24822 = n24813 & n24821;
  assign n24823 = n24820 & n24822;
  assign n24824 = n24045 & ~n24823;
  assign n24825 = ~n24792 & ~n24824;
  assign n24826 = n24683 & n24823;
  assign n24827 = n24685 & ~n24823;
  assign n24828 = ~P1_STATE2_REG_0_ & n24397;
  assign n24829 = ~n24826 & ~n24827;
  assign n24830 = ~n24828 & n24829;
  assign n24831 = ~n24683 & ~n24830;
  assign n24832 = n24683 & n24830;
  assign n24833 = ~n24831 & ~n24832;
  assign n24834 = ~n24825 & ~n24833;
  assign n24835 = n24825 & n24833;
  assign n24836 = ~n24834 & ~n24835;
  assign n24837 = ~n24772 & ~n24776;
  assign n24838 = n24772 & n24776;
  assign n24839 = ~n24733 & ~n24838;
  assign n24840 = ~n24837 & ~n24839;
  assign n24841 = n24836 & n24840;
  assign n24842 = ~n24836 & ~n24840;
  assign n24843 = ~n24841 & ~n24842;
  assign n24844 = n24791 & n24843;
  assign n24845 = ~n24791 & ~n24843;
  assign n24846 = ~n24844 & ~n24845;
  assign n24847 = ~n24835 & ~n24840;
  assign n24848 = P1_INSTQUEUE_REG_0__3_ & n24040;
  assign n24849 = P1_INSTQUEUE_REG_0__3_ & n24630;
  assign n24850 = P1_INSTQUEUE_REG_1__3_ & n24633;
  assign n24851 = P1_INSTQUEUE_REG_2__3_ & n24636;
  assign n24852 = P1_INSTQUEUE_REG_3__3_ & n24639;
  assign n24853 = ~n24849 & ~n24850;
  assign n24854 = ~n24851 & n24853;
  assign n24855 = ~n24852 & n24854;
  assign n24856 = P1_INSTQUEUE_REG_4__3_ & n24645;
  assign n24857 = P1_INSTQUEUE_REG_5__3_ & n24647;
  assign n24858 = P1_INSTQUEUE_REG_6__3_ & n24649;
  assign n24859 = P1_INSTQUEUE_REG_7__3_ & n24651;
  assign n24860 = ~n24856 & ~n24857;
  assign n24861 = ~n24858 & n24860;
  assign n24862 = ~n24859 & n24861;
  assign n24863 = P1_INSTQUEUE_REG_8__3_ & n24657;
  assign n24864 = P1_INSTQUEUE_REG_9__3_ & n24659;
  assign n24865 = P1_INSTQUEUE_REG_10__3_ & n24661;
  assign n24866 = P1_INSTQUEUE_REG_11__3_ & n24663;
  assign n24867 = ~n24863 & ~n24864;
  assign n24868 = ~n24865 & n24867;
  assign n24869 = ~n24866 & n24868;
  assign n24870 = P1_INSTQUEUE_REG_12__3_ & n24669;
  assign n24871 = P1_INSTQUEUE_REG_13__3_ & n24671;
  assign n24872 = P1_INSTQUEUE_REG_14__3_ & n24673;
  assign n24873 = P1_INSTQUEUE_REG_15__3_ & n24675;
  assign n24874 = ~n24870 & ~n24871;
  assign n24875 = ~n24872 & n24874;
  assign n24876 = ~n24873 & n24875;
  assign n24877 = n24855 & n24862;
  assign n24878 = n24869 & n24877;
  assign n24879 = n24876 & n24878;
  assign n24880 = n24045 & ~n24879;
  assign n24881 = ~n24848 & ~n24880;
  assign n24882 = n24683 & n24879;
  assign n24883 = n24685 & ~n24879;
  assign n24884 = ~P1_STATE2_REG_0_ & ~n24482;
  assign n24885 = ~n24882 & ~n24883;
  assign n24886 = ~n24884 & n24885;
  assign n24887 = ~n24683 & ~n24886;
  assign n24888 = n24683 & n24886;
  assign n24889 = ~n24887 & ~n24888;
  assign n24890 = ~n24881 & ~n24889;
  assign n24891 = n24881 & n24889;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n24834 & ~n24847;
  assign n24894 = ~n24892 & n24893;
  assign n24895 = n24892 & ~n24893;
  assign n24896 = ~n24894 & ~n24895;
  assign n24897 = n24843 & n24896;
  assign n24898 = ~n24791 & n24896;
  assign n24899 = ~n24843 & ~n24896;
  assign n24900 = n24791 & n24899;
  assign n24901 = ~n24897 & ~n24898;
  assign n24902 = ~n24900 & n24901;
  assign n24903 = ~n24846 & ~n24902;
  assign n24904 = n24790 & n24903;
  assign n24905 = ~n24843 & n24896;
  assign n24906 = n24791 & n24905;
  assign n24907 = ~n24904 & ~n24906;
  assign n24908 = P1_STATEBS16_REG & n24626;
  assign n24909 = ~P1_STATE2_REG_2_ & P1_STATE2_REG_1_;
  assign n24910 = ~n24313 & ~n24909;
  assign n24911 = ~n24590 & n24910;
  assign n24912 = ~P1_STATE2_REG_0_ & ~n24911;
  assign n24913 = n24908 & n24912;
  assign n24914 = n24907 & n24913;
  assign n24915 = ~n24627 & ~n24914;
  assign n24916 = n24625 & ~n24915;
  assign n24917 = P1_STATE2_REG_3_ & ~n24621;
  assign n24918 = ~n24384 & ~n24462;
  assign n24919 = ~P1_INSTQUEUEWR_ADDR_REG_0_ & ~n24311;
  assign n24920 = n24918 & n24919;
  assign n24921 = ~n24621 & ~n24920;
  assign n24922 = P1_STATE2_REG_2_ & n24921;
  assign n24923 = ~n24917 & ~n24922;
  assign n24924 = n24912 & n24923;
  assign n24925 = ~n24916 & n24924;
  assign n24926 = P1_INSTQUEUE_REG_15__7_ & ~n24925;
  assign n24927 = BUF1_REG_7_ & n4507;
  assign n24928 = DATAI_7_ & ~n4507;
  assign n24929 = ~n24927 & ~n24928;
  assign n24930 = n24912 & ~n24929;
  assign n24931 = P1_STATE2_REG_2_ & ~n24921;
  assign n24932 = n24907 & n24908;
  assign n24933 = ~n24627 & ~n24932;
  assign n24934 = ~n24625 & ~n24933;
  assign n24935 = ~n24931 & ~n24934;
  assign n24936 = n24930 & ~n24935;
  assign n24937 = BUF1_REG_23_ & n4507;
  assign n24938 = DATAI_23_ & ~n4507;
  assign n24939 = ~n24937 & ~n24938;
  assign n24940 = n24913 & ~n24939;
  assign n24941 = n24906 & n24940;
  assign n24942 = P1_STATE2_REG_3_ & n24912;
  assign n24943 = ~n23831 & n24942;
  assign n24944 = n24621 & n24943;
  assign n24945 = BUF1_REG_31_ & n4507;
  assign n24946 = DATAI_31_ & ~n4507;
  assign n24947 = ~n24945 & ~n24946;
  assign n24948 = n24913 & ~n24947;
  assign n24949 = n24904 & n24948;
  assign n24950 = ~n24941 & ~n24944;
  assign n24951 = ~n24949 & n24950;
  assign n24952 = ~n24926 & ~n24936;
  assign n5399 = ~n24951 | ~n24952;
  assign n24954 = P1_INSTQUEUE_REG_15__6_ & ~n24925;
  assign n24955 = BUF1_REG_6_ & n4507;
  assign n24956 = DATAI_6_ & ~n4507;
  assign n24957 = ~n24955 & ~n24956;
  assign n24958 = n24912 & ~n24957;
  assign n24959 = ~n24935 & n24958;
  assign n24960 = BUF1_REG_22_ & n4507;
  assign n24961 = DATAI_22_ & ~n4507;
  assign n24962 = ~n24960 & ~n24961;
  assign n24963 = n24913 & ~n24962;
  assign n24964 = n24906 & n24963;
  assign n24965 = ~n23800 & n24942;
  assign n24966 = n24621 & n24965;
  assign n24967 = BUF1_REG_30_ & n4507;
  assign n24968 = DATAI_30_ & ~n4507;
  assign n24969 = ~n24967 & ~n24968;
  assign n24970 = n24913 & ~n24969;
  assign n24971 = n24904 & n24970;
  assign n24972 = ~n24964 & ~n24966;
  assign n24973 = ~n24971 & n24972;
  assign n24974 = ~n24954 & ~n24959;
  assign n5404 = ~n24973 | ~n24974;
  assign n24976 = P1_INSTQUEUE_REG_15__5_ & ~n24925;
  assign n24977 = BUF1_REG_5_ & n4507;
  assign n24978 = DATAI_5_ & ~n4507;
  assign n24979 = ~n24977 & ~n24978;
  assign n24980 = n24912 & ~n24979;
  assign n24981 = ~n24935 & n24980;
  assign n24982 = BUF1_REG_21_ & n4507;
  assign n24983 = DATAI_21_ & ~n4507;
  assign n24984 = ~n24982 & ~n24983;
  assign n24985 = n24913 & ~n24984;
  assign n24986 = n24906 & n24985;
  assign n24987 = ~n23896 & n24942;
  assign n24988 = n24621 & n24987;
  assign n24989 = BUF1_REG_29_ & n4507;
  assign n24990 = DATAI_29_ & ~n4507;
  assign n24991 = ~n24989 & ~n24990;
  assign n24992 = n24913 & ~n24991;
  assign n24993 = n24904 & n24992;
  assign n24994 = ~n24986 & ~n24988;
  assign n24995 = ~n24993 & n24994;
  assign n24996 = ~n24976 & ~n24981;
  assign n5409 = ~n24995 | ~n24996;
  assign n24998 = P1_INSTQUEUE_REG_15__4_ & ~n24925;
  assign n24999 = BUF1_REG_4_ & n4507;
  assign n25000 = DATAI_4_ & ~n4507;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = n24912 & ~n25001;
  assign n25003 = ~n24935 & n25002;
  assign n25004 = BUF1_REG_20_ & n4507;
  assign n25005 = DATAI_20_ & ~n4507;
  assign n25006 = ~n25004 & ~n25005;
  assign n25007 = n24913 & ~n25006;
  assign n25008 = n24906 & n25007;
  assign n25009 = ~n23968 & n24942;
  assign n25010 = n24621 & n25009;
  assign n25011 = BUF1_REG_28_ & n4507;
  assign n25012 = DATAI_28_ & ~n4507;
  assign n25013 = ~n25011 & ~n25012;
  assign n25014 = n24913 & ~n25013;
  assign n25015 = n24904 & n25014;
  assign n25016 = ~n25008 & ~n25010;
  assign n25017 = ~n25015 & n25016;
  assign n25018 = ~n24998 & ~n25003;
  assign n5414 = ~n25017 | ~n25018;
  assign n25020 = P1_INSTQUEUE_REG_15__3_ & ~n24925;
  assign n25021 = BUF1_REG_3_ & n4507;
  assign n25022 = DATAI_3_ & ~n4507;
  assign n25023 = ~n25021 & ~n25022;
  assign n25024 = n24912 & ~n25023;
  assign n25025 = ~n24935 & n25024;
  assign n25026 = BUF1_REG_19_ & n4507;
  assign n25027 = DATAI_19_ & ~n4507;
  assign n25028 = ~n25026 & ~n25027;
  assign n25029 = n24913 & ~n25028;
  assign n25030 = n24906 & n25029;
  assign n25031 = ~n23741 & n24942;
  assign n25032 = n24621 & n25031;
  assign n25033 = BUF1_REG_27_ & n4507;
  assign n25034 = DATAI_27_ & ~n4507;
  assign n25035 = ~n25033 & ~n25034;
  assign n25036 = n24913 & ~n25035;
  assign n25037 = n24904 & n25036;
  assign n25038 = ~n25030 & ~n25032;
  assign n25039 = ~n25037 & n25038;
  assign n25040 = ~n25020 & ~n25025;
  assign n5419 = ~n25039 | ~n25040;
  assign n25042 = P1_INSTQUEUE_REG_15__2_ & ~n24925;
  assign n25043 = BUF1_REG_2_ & n4507;
  assign n25044 = DATAI_2_ & ~n4507;
  assign n25045 = ~n25043 & ~n25044;
  assign n25046 = n24912 & ~n25045;
  assign n25047 = ~n24935 & n25046;
  assign n25048 = BUF1_REG_18_ & n4507;
  assign n25049 = DATAI_18_ & ~n4507;
  assign n25050 = ~n25048 & ~n25049;
  assign n25051 = n24913 & ~n25050;
  assign n25052 = n24906 & n25051;
  assign n25053 = ~n24002 & n24942;
  assign n25054 = n24621 & n25053;
  assign n25055 = BUF1_REG_26_ & n4507;
  assign n25056 = DATAI_26_ & ~n4507;
  assign n25057 = ~n25055 & ~n25056;
  assign n25058 = n24913 & ~n25057;
  assign n25059 = n24904 & n25058;
  assign n25060 = ~n25052 & ~n25054;
  assign n25061 = ~n25059 & n25060;
  assign n25062 = ~n25042 & ~n25047;
  assign n5424 = ~n25061 | ~n25062;
  assign n25064 = P1_INSTQUEUE_REG_15__1_ & ~n24925;
  assign n25065 = BUF1_REG_1_ & n4507;
  assign n25066 = DATAI_1_ & ~n4507;
  assign n25067 = ~n25065 & ~n25066;
  assign n25068 = n24912 & ~n25067;
  assign n25069 = ~n24935 & n25068;
  assign n25070 = BUF1_REG_17_ & n4507;
  assign n25071 = DATAI_17_ & ~n4507;
  assign n25072 = ~n25070 & ~n25071;
  assign n25073 = n24913 & ~n25072;
  assign n25074 = n24906 & n25073;
  assign n25075 = ~n23709 & n24942;
  assign n25076 = n24621 & n25075;
  assign n25077 = BUF1_REG_25_ & n4507;
  assign n25078 = DATAI_25_ & ~n4507;
  assign n25079 = ~n25077 & ~n25078;
  assign n25080 = n24913 & ~n25079;
  assign n25081 = n24904 & n25080;
  assign n25082 = ~n25074 & ~n25076;
  assign n25083 = ~n25081 & n25082;
  assign n25084 = ~n25064 & ~n25069;
  assign n5429 = ~n25083 | ~n25084;
  assign n25086 = P1_INSTQUEUE_REG_15__0_ & ~n24925;
  assign n25087 = BUF1_REG_0_ & n4507;
  assign n25088 = DATAI_0_ & ~n4507;
  assign n25089 = ~n25087 & ~n25088;
  assign n25090 = n24912 & ~n25089;
  assign n25091 = ~n24935 & n25090;
  assign n25092 = BUF1_REG_16_ & n4507;
  assign n25093 = DATAI_16_ & ~n4507;
  assign n25094 = ~n25092 & ~n25093;
  assign n25095 = n24913 & ~n25094;
  assign n25096 = n24906 & n25095;
  assign n25097 = ~n23678 & n24942;
  assign n25098 = n24621 & n25097;
  assign n25099 = BUF1_REG_24_ & n4507;
  assign n25100 = DATAI_24_ & ~n4507;
  assign n25101 = ~n25099 & ~n25100;
  assign n25102 = n24913 & ~n25101;
  assign n25103 = n24904 & n25102;
  assign n25104 = ~n25096 & ~n25098;
  assign n25105 = ~n25103 & n25104;
  assign n25106 = ~n25086 & ~n25091;
  assign n5434 = ~n25105 | ~n25106;
  assign n25108 = n24310 & n24620;
  assign n25109 = n24520 & ~n24535;
  assign n25110 = n24622 & n25109;
  assign n25111 = ~n25108 & ~n25110;
  assign n25112 = ~n24786 & ~n24789;
  assign n25113 = n24903 & n25112;
  assign n25114 = n24787 & n24905;
  assign n25115 = ~n25113 & ~n25114;
  assign n25116 = n24913 & n25115;
  assign n25117 = ~n24627 & ~n25116;
  assign n25118 = n25111 & ~n25117;
  assign n25119 = P1_STATE2_REG_3_ & ~n25108;
  assign n25120 = ~n24311 & n24918;
  assign n25121 = P1_STATE2_REG_2_ & ~n25120;
  assign n25122 = ~n25119 & ~n25121;
  assign n25123 = n24912 & n25122;
  assign n25124 = ~n25118 & n25123;
  assign n25125 = P1_INSTQUEUE_REG_14__7_ & ~n25124;
  assign n25126 = P1_STATE2_REG_2_ & n25120;
  assign n25127 = n24908 & n25115;
  assign n25128 = ~n24627 & ~n25127;
  assign n25129 = ~n25111 & ~n25128;
  assign n25130 = ~n25126 & ~n25129;
  assign n25131 = n24930 & ~n25130;
  assign n25132 = n24940 & n25114;
  assign n25133 = n24943 & n25108;
  assign n25134 = n24948 & n25113;
  assign n25135 = ~n25132 & ~n25133;
  assign n25136 = ~n25134 & n25135;
  assign n25137 = ~n25125 & ~n25131;
  assign n5439 = ~n25136 | ~n25137;
  assign n25139 = P1_INSTQUEUE_REG_14__6_ & ~n25124;
  assign n25140 = n24958 & ~n25130;
  assign n25141 = n24963 & n25114;
  assign n25142 = n24965 & n25108;
  assign n25143 = n24970 & n25113;
  assign n25144 = ~n25141 & ~n25142;
  assign n25145 = ~n25143 & n25144;
  assign n25146 = ~n25139 & ~n25140;
  assign n5444 = ~n25145 | ~n25146;
  assign n25148 = P1_INSTQUEUE_REG_14__5_ & ~n25124;
  assign n25149 = n24980 & ~n25130;
  assign n25150 = n24985 & n25114;
  assign n25151 = n24987 & n25108;
  assign n25152 = n24992 & n25113;
  assign n25153 = ~n25150 & ~n25151;
  assign n25154 = ~n25152 & n25153;
  assign n25155 = ~n25148 & ~n25149;
  assign n5449 = ~n25154 | ~n25155;
  assign n25157 = P1_INSTQUEUE_REG_14__4_ & ~n25124;
  assign n25158 = n25002 & ~n25130;
  assign n25159 = n25007 & n25114;
  assign n25160 = n25009 & n25108;
  assign n25161 = n25014 & n25113;
  assign n25162 = ~n25159 & ~n25160;
  assign n25163 = ~n25161 & n25162;
  assign n25164 = ~n25157 & ~n25158;
  assign n5454 = ~n25163 | ~n25164;
  assign n25166 = P1_INSTQUEUE_REG_14__3_ & ~n25124;
  assign n25167 = n25024 & ~n25130;
  assign n25168 = n25029 & n25114;
  assign n25169 = n25031 & n25108;
  assign n25170 = n25036 & n25113;
  assign n25171 = ~n25168 & ~n25169;
  assign n25172 = ~n25170 & n25171;
  assign n25173 = ~n25166 & ~n25167;
  assign n5459 = ~n25172 | ~n25173;
  assign n25175 = P1_INSTQUEUE_REG_14__2_ & ~n25124;
  assign n25176 = n25046 & ~n25130;
  assign n25177 = n25051 & n25114;
  assign n25178 = n25053 & n25108;
  assign n25179 = n25058 & n25113;
  assign n25180 = ~n25177 & ~n25178;
  assign n25181 = ~n25179 & n25180;
  assign n25182 = ~n25175 & ~n25176;
  assign n5464 = ~n25181 | ~n25182;
  assign n25184 = P1_INSTQUEUE_REG_14__1_ & ~n25124;
  assign n25185 = n25068 & ~n25130;
  assign n25186 = n25073 & n25114;
  assign n25187 = n25075 & n25108;
  assign n25188 = n25080 & n25113;
  assign n25189 = ~n25186 & ~n25187;
  assign n25190 = ~n25188 & n25189;
  assign n25191 = ~n25184 & ~n25185;
  assign n5469 = ~n25190 | ~n25191;
  assign n25193 = P1_INSTQUEUE_REG_14__0_ & ~n25124;
  assign n25194 = n25090 & ~n25130;
  assign n25195 = n25095 & n25114;
  assign n25196 = n25097 & n25108;
  assign n25197 = n25102 & n25113;
  assign n25198 = ~n25195 & ~n25196;
  assign n25199 = ~n25197 & n25198;
  assign n25200 = ~n25193 & ~n25194;
  assign n5474 = ~n25199 | ~n25200;
  assign n25202 = n24309 & n24620;
  assign n25203 = ~n24520 & n24535;
  assign n25204 = n24622 & n25203;
  assign n25205 = ~n25202 & ~n25204;
  assign n25206 = n24786 & n24789;
  assign n25207 = n24903 & n25206;
  assign n25208 = n24788 & n24905;
  assign n25209 = ~n25207 & ~n25208;
  assign n25210 = n24913 & n25209;
  assign n25211 = ~n24627 & ~n25210;
  assign n25212 = n25205 & ~n25211;
  assign n25213 = P1_STATE2_REG_3_ & ~n25202;
  assign n25214 = ~P1_INSTQUEUEWR_ADDR_REG_0_ & n24311;
  assign n25215 = n24918 & n25214;
  assign n25216 = ~n25202 & ~n25215;
  assign n25217 = P1_STATE2_REG_2_ & n25216;
  assign n25218 = ~n25213 & ~n25217;
  assign n25219 = n24912 & n25218;
  assign n25220 = ~n25212 & n25219;
  assign n25221 = P1_INSTQUEUE_REG_13__7_ & ~n25220;
  assign n25222 = P1_STATE2_REG_2_ & ~n25216;
  assign n25223 = n24908 & n25209;
  assign n25224 = ~n24627 & ~n25223;
  assign n25225 = ~n25205 & ~n25224;
  assign n25226 = ~n25222 & ~n25225;
  assign n25227 = n24930 & ~n25226;
  assign n25228 = n24940 & n25208;
  assign n25229 = n24943 & n25202;
  assign n25230 = n24948 & n25207;
  assign n25231 = ~n25228 & ~n25229;
  assign n25232 = ~n25230 & n25231;
  assign n25233 = ~n25221 & ~n25227;
  assign n5479 = ~n25232 | ~n25233;
  assign n25235 = P1_INSTQUEUE_REG_13__6_ & ~n25220;
  assign n25236 = n24958 & ~n25226;
  assign n25237 = n24963 & n25208;
  assign n25238 = n24965 & n25202;
  assign n25239 = n24970 & n25207;
  assign n25240 = ~n25237 & ~n25238;
  assign n25241 = ~n25239 & n25240;
  assign n25242 = ~n25235 & ~n25236;
  assign n5484 = ~n25241 | ~n25242;
  assign n25244 = P1_INSTQUEUE_REG_13__5_ & ~n25220;
  assign n25245 = n24980 & ~n25226;
  assign n25246 = n24985 & n25208;
  assign n25247 = n24987 & n25202;
  assign n25248 = n24992 & n25207;
  assign n25249 = ~n25246 & ~n25247;
  assign n25250 = ~n25248 & n25249;
  assign n25251 = ~n25244 & ~n25245;
  assign n5489 = ~n25250 | ~n25251;
  assign n25253 = P1_INSTQUEUE_REG_13__4_ & ~n25220;
  assign n25254 = n25002 & ~n25226;
  assign n25255 = n25007 & n25208;
  assign n25256 = n25009 & n25202;
  assign n25257 = n25014 & n25207;
  assign n25258 = ~n25255 & ~n25256;
  assign n25259 = ~n25257 & n25258;
  assign n25260 = ~n25253 & ~n25254;
  assign n5494 = ~n25259 | ~n25260;
  assign n25262 = P1_INSTQUEUE_REG_13__3_ & ~n25220;
  assign n25263 = n25024 & ~n25226;
  assign n25264 = n25029 & n25208;
  assign n25265 = n25031 & n25202;
  assign n25266 = n25036 & n25207;
  assign n25267 = ~n25264 & ~n25265;
  assign n25268 = ~n25266 & n25267;
  assign n25269 = ~n25262 & ~n25263;
  assign n5499 = ~n25268 | ~n25269;
  assign n25271 = P1_INSTQUEUE_REG_13__2_ & ~n25220;
  assign n25272 = n25046 & ~n25226;
  assign n25273 = n25051 & n25208;
  assign n25274 = n25053 & n25202;
  assign n25275 = n25058 & n25207;
  assign n25276 = ~n25273 & ~n25274;
  assign n25277 = ~n25275 & n25276;
  assign n25278 = ~n25271 & ~n25272;
  assign n5504 = ~n25277 | ~n25278;
  assign n25280 = P1_INSTQUEUE_REG_13__1_ & ~n25220;
  assign n25281 = n25068 & ~n25226;
  assign n25282 = n25073 & n25208;
  assign n25283 = n25075 & n25202;
  assign n25284 = n25080 & n25207;
  assign n25285 = ~n25282 & ~n25283;
  assign n25286 = ~n25284 & n25285;
  assign n25287 = ~n25280 & ~n25281;
  assign n5509 = ~n25286 | ~n25287;
  assign n25289 = P1_INSTQUEUE_REG_13__0_ & ~n25220;
  assign n25290 = n25090 & ~n25226;
  assign n25291 = n25095 & n25208;
  assign n25292 = n25097 & n25202;
  assign n25293 = n25102 & n25207;
  assign n25294 = ~n25291 & ~n25292;
  assign n25295 = ~n25293 & n25294;
  assign n25296 = ~n25289 & ~n25290;
  assign n5514 = ~n25295 | ~n25296;
  assign n25298 = ~P1_INSTQUEUEWR_ADDR_REG_1_ & ~P1_INSTQUEUEWR_ADDR_REG_0_;
  assign n25299 = n24620 & n25298;
  assign n25300 = n24520 & n24535;
  assign n25301 = n24622 & n25300;
  assign n25302 = ~n25299 & ~n25301;
  assign n25303 = ~n24786 & n24789;
  assign n25304 = n24903 & n25303;
  assign n25305 = n24782 & n24786;
  assign n25306 = n24905 & n25305;
  assign n25307 = ~n25304 & ~n25306;
  assign n25308 = n24913 & n25307;
  assign n25309 = ~n24627 & ~n25308;
  assign n25310 = n25302 & ~n25309;
  assign n25311 = P1_STATE2_REG_3_ & ~n25299;
  assign n25312 = n24311 & n24918;
  assign n25313 = P1_STATE2_REG_2_ & ~n25312;
  assign n25314 = ~n25311 & ~n25313;
  assign n25315 = n24912 & n25314;
  assign n25316 = ~n25310 & n25315;
  assign n25317 = P1_INSTQUEUE_REG_12__7_ & ~n25316;
  assign n25318 = P1_STATE2_REG_2_ & n25312;
  assign n25319 = n24908 & n25307;
  assign n25320 = ~n24627 & ~n25319;
  assign n25321 = ~n25302 & ~n25320;
  assign n25322 = ~n25318 & ~n25321;
  assign n25323 = n24930 & ~n25322;
  assign n25324 = n24940 & n25306;
  assign n25325 = n24943 & n25299;
  assign n25326 = n24948 & n25304;
  assign n25327 = ~n25324 & ~n25325;
  assign n25328 = ~n25326 & n25327;
  assign n25329 = ~n25317 & ~n25323;
  assign n5519 = ~n25328 | ~n25329;
  assign n25331 = P1_INSTQUEUE_REG_12__6_ & ~n25316;
  assign n25332 = n24958 & ~n25322;
  assign n25333 = n24963 & n25306;
  assign n25334 = n24965 & n25299;
  assign n25335 = n24970 & n25304;
  assign n25336 = ~n25333 & ~n25334;
  assign n25337 = ~n25335 & n25336;
  assign n25338 = ~n25331 & ~n25332;
  assign n5524 = ~n25337 | ~n25338;
  assign n25340 = P1_INSTQUEUE_REG_12__5_ & ~n25316;
  assign n25341 = n24980 & ~n25322;
  assign n25342 = n24985 & n25306;
  assign n25343 = n24987 & n25299;
  assign n25344 = n24992 & n25304;
  assign n25345 = ~n25342 & ~n25343;
  assign n25346 = ~n25344 & n25345;
  assign n25347 = ~n25340 & ~n25341;
  assign n5529 = ~n25346 | ~n25347;
  assign n25349 = P1_INSTQUEUE_REG_12__4_ & ~n25316;
  assign n25350 = n25002 & ~n25322;
  assign n25351 = n25007 & n25306;
  assign n25352 = n25009 & n25299;
  assign n25353 = n25014 & n25304;
  assign n25354 = ~n25351 & ~n25352;
  assign n25355 = ~n25353 & n25354;
  assign n25356 = ~n25349 & ~n25350;
  assign n5534 = ~n25355 | ~n25356;
  assign n25358 = P1_INSTQUEUE_REG_12__3_ & ~n25316;
  assign n25359 = n25024 & ~n25322;
  assign n25360 = n25029 & n25306;
  assign n25361 = n25031 & n25299;
  assign n25362 = n25036 & n25304;
  assign n25363 = ~n25360 & ~n25361;
  assign n25364 = ~n25362 & n25363;
  assign n25365 = ~n25358 & ~n25359;
  assign n5539 = ~n25364 | ~n25365;
  assign n25367 = P1_INSTQUEUE_REG_12__2_ & ~n25316;
  assign n25368 = n25046 & ~n25322;
  assign n25369 = n25051 & n25306;
  assign n25370 = n25053 & n25299;
  assign n25371 = n25058 & n25304;
  assign n25372 = ~n25369 & ~n25370;
  assign n25373 = ~n25371 & n25372;
  assign n25374 = ~n25367 & ~n25368;
  assign n5544 = ~n25373 | ~n25374;
  assign n25376 = P1_INSTQUEUE_REG_12__1_ & ~n25316;
  assign n25377 = n25068 & ~n25322;
  assign n25378 = n25073 & n25306;
  assign n25379 = n25075 & n25299;
  assign n25380 = n25080 & n25304;
  assign n25381 = ~n25378 & ~n25379;
  assign n25382 = ~n25380 & n25381;
  assign n25383 = ~n25376 & ~n25377;
  assign n5549 = ~n25382 | ~n25383;
  assign n25385 = P1_INSTQUEUE_REG_12__0_ & ~n25316;
  assign n25386 = n25090 & ~n25322;
  assign n25387 = n25095 & n25306;
  assign n25388 = n25097 & n25299;
  assign n25389 = n25102 & n25304;
  assign n25390 = ~n25387 & ~n25388;
  assign n25391 = ~n25389 & n25390;
  assign n25392 = ~n25385 & ~n25386;
  assign n5554 = ~n25391 | ~n25392;
  assign n25394 = n24381 & n24457;
  assign n25395 = ~n24397 & ~n24482;
  assign n25396 = n24623 & n25395;
  assign n25397 = ~n25394 & ~n25396;
  assign n25398 = n24846 & ~n24902;
  assign n25399 = n24790 & n25398;
  assign n25400 = n24791 & n24897;
  assign n25401 = ~n25399 & ~n25400;
  assign n25402 = n24913 & n25401;
  assign n25403 = ~n24627 & ~n25402;
  assign n25404 = n25397 & ~n25403;
  assign n25405 = P1_STATE2_REG_3_ & ~n25394;
  assign n25406 = n24384 & ~n24462;
  assign n25407 = n24919 & n25406;
  assign n25408 = ~n25394 & ~n25407;
  assign n25409 = P1_STATE2_REG_2_ & n25408;
  assign n25410 = ~n25405 & ~n25409;
  assign n25411 = n24912 & n25410;
  assign n25412 = ~n25404 & n25411;
  assign n25413 = P1_INSTQUEUE_REG_11__7_ & ~n25412;
  assign n25414 = P1_STATE2_REG_2_ & ~n25408;
  assign n25415 = n24908 & n25401;
  assign n25416 = ~n24627 & ~n25415;
  assign n25417 = ~n25397 & ~n25416;
  assign n25418 = ~n25414 & ~n25417;
  assign n25419 = n24930 & ~n25418;
  assign n25420 = n24940 & n25400;
  assign n25421 = n24943 & n25394;
  assign n25422 = n24948 & n25399;
  assign n25423 = ~n25420 & ~n25421;
  assign n25424 = ~n25422 & n25423;
  assign n25425 = ~n25413 & ~n25419;
  assign n5559 = ~n25424 | ~n25425;
  assign n25427 = P1_INSTQUEUE_REG_11__6_ & ~n25412;
  assign n25428 = n24958 & ~n25418;
  assign n25429 = n24963 & n25400;
  assign n25430 = n24965 & n25394;
  assign n25431 = n24970 & n25399;
  assign n25432 = ~n25429 & ~n25430;
  assign n25433 = ~n25431 & n25432;
  assign n25434 = ~n25427 & ~n25428;
  assign n5564 = ~n25433 | ~n25434;
  assign n25436 = P1_INSTQUEUE_REG_11__5_ & ~n25412;
  assign n25437 = n24980 & ~n25418;
  assign n25438 = n24985 & n25400;
  assign n25439 = n24987 & n25394;
  assign n25440 = n24992 & n25399;
  assign n25441 = ~n25438 & ~n25439;
  assign n25442 = ~n25440 & n25441;
  assign n25443 = ~n25436 & ~n25437;
  assign n5569 = ~n25442 | ~n25443;
  assign n25445 = P1_INSTQUEUE_REG_11__4_ & ~n25412;
  assign n25446 = n25002 & ~n25418;
  assign n25447 = n25007 & n25400;
  assign n25448 = n25009 & n25394;
  assign n25449 = n25014 & n25399;
  assign n25450 = ~n25447 & ~n25448;
  assign n25451 = ~n25449 & n25450;
  assign n25452 = ~n25445 & ~n25446;
  assign n5574 = ~n25451 | ~n25452;
  assign n25454 = P1_INSTQUEUE_REG_11__3_ & ~n25412;
  assign n25455 = n25024 & ~n25418;
  assign n25456 = n25029 & n25400;
  assign n25457 = n25031 & n25394;
  assign n25458 = n25036 & n25399;
  assign n25459 = ~n25456 & ~n25457;
  assign n25460 = ~n25458 & n25459;
  assign n25461 = ~n25454 & ~n25455;
  assign n5579 = ~n25460 | ~n25461;
  assign n25463 = P1_INSTQUEUE_REG_11__2_ & ~n25412;
  assign n25464 = n25046 & ~n25418;
  assign n25465 = n25051 & n25400;
  assign n25466 = n25053 & n25394;
  assign n25467 = n25058 & n25399;
  assign n25468 = ~n25465 & ~n25466;
  assign n25469 = ~n25467 & n25468;
  assign n25470 = ~n25463 & ~n25464;
  assign n5584 = ~n25469 | ~n25470;
  assign n25472 = P1_INSTQUEUE_REG_11__1_ & ~n25412;
  assign n25473 = n25068 & ~n25418;
  assign n25474 = n25073 & n25400;
  assign n25475 = n25075 & n25394;
  assign n25476 = n25080 & n25399;
  assign n25477 = ~n25474 & ~n25475;
  assign n25478 = ~n25476 & n25477;
  assign n25479 = ~n25472 & ~n25473;
  assign n5589 = ~n25478 | ~n25479;
  assign n25481 = P1_INSTQUEUE_REG_11__0_ & ~n25412;
  assign n25482 = n25090 & ~n25418;
  assign n25483 = n25095 & n25400;
  assign n25484 = n25097 & n25394;
  assign n25485 = n25102 & n25399;
  assign n25486 = ~n25483 & ~n25484;
  assign n25487 = ~n25485 & n25486;
  assign n25488 = ~n25481 & ~n25482;
  assign n5594 = ~n25487 | ~n25488;
  assign n25490 = n24310 & n24457;
  assign n25491 = n25109 & n25395;
  assign n25492 = ~n25490 & ~n25491;
  assign n25493 = n25112 & n25398;
  assign n25494 = n24787 & n24897;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 = n24913 & n25495;
  assign n25497 = ~n24627 & ~n25496;
  assign n25498 = n25492 & ~n25497;
  assign n25499 = P1_STATE2_REG_3_ & ~n25490;
  assign n25500 = ~n24311 & n25406;
  assign n25501 = P1_STATE2_REG_2_ & ~n25500;
  assign n25502 = ~n25499 & ~n25501;
  assign n25503 = n24912 & n25502;
  assign n25504 = ~n25498 & n25503;
  assign n25505 = P1_INSTQUEUE_REG_10__7_ & ~n25504;
  assign n25506 = P1_STATE2_REG_2_ & n25500;
  assign n25507 = n24908 & n25495;
  assign n25508 = ~n24627 & ~n25507;
  assign n25509 = ~n25492 & ~n25508;
  assign n25510 = ~n25506 & ~n25509;
  assign n25511 = n24930 & ~n25510;
  assign n25512 = n24940 & n25494;
  assign n25513 = n24943 & n25490;
  assign n25514 = n24948 & n25493;
  assign n25515 = ~n25512 & ~n25513;
  assign n25516 = ~n25514 & n25515;
  assign n25517 = ~n25505 & ~n25511;
  assign n5599 = ~n25516 | ~n25517;
  assign n25519 = P1_INSTQUEUE_REG_10__6_ & ~n25504;
  assign n25520 = n24958 & ~n25510;
  assign n25521 = n24963 & n25494;
  assign n25522 = n24965 & n25490;
  assign n25523 = n24970 & n25493;
  assign n25524 = ~n25521 & ~n25522;
  assign n25525 = ~n25523 & n25524;
  assign n25526 = ~n25519 & ~n25520;
  assign n5604 = ~n25525 | ~n25526;
  assign n25528 = P1_INSTQUEUE_REG_10__5_ & ~n25504;
  assign n25529 = n24980 & ~n25510;
  assign n25530 = n24985 & n25494;
  assign n25531 = n24987 & n25490;
  assign n25532 = n24992 & n25493;
  assign n25533 = ~n25530 & ~n25531;
  assign n25534 = ~n25532 & n25533;
  assign n25535 = ~n25528 & ~n25529;
  assign n5609 = ~n25534 | ~n25535;
  assign n25537 = P1_INSTQUEUE_REG_10__4_ & ~n25504;
  assign n25538 = n25002 & ~n25510;
  assign n25539 = n25007 & n25494;
  assign n25540 = n25009 & n25490;
  assign n25541 = n25014 & n25493;
  assign n25542 = ~n25539 & ~n25540;
  assign n25543 = ~n25541 & n25542;
  assign n25544 = ~n25537 & ~n25538;
  assign n5614 = ~n25543 | ~n25544;
  assign n25546 = P1_INSTQUEUE_REG_10__3_ & ~n25504;
  assign n25547 = n25024 & ~n25510;
  assign n25548 = n25029 & n25494;
  assign n25549 = n25031 & n25490;
  assign n25550 = n25036 & n25493;
  assign n25551 = ~n25548 & ~n25549;
  assign n25552 = ~n25550 & n25551;
  assign n25553 = ~n25546 & ~n25547;
  assign n5619 = ~n25552 | ~n25553;
  assign n25555 = P1_INSTQUEUE_REG_10__2_ & ~n25504;
  assign n25556 = n25046 & ~n25510;
  assign n25557 = n25051 & n25494;
  assign n25558 = n25053 & n25490;
  assign n25559 = n25058 & n25493;
  assign n25560 = ~n25557 & ~n25558;
  assign n25561 = ~n25559 & n25560;
  assign n25562 = ~n25555 & ~n25556;
  assign n5624 = ~n25561 | ~n25562;
  assign n25564 = P1_INSTQUEUE_REG_10__1_ & ~n25504;
  assign n25565 = n25068 & ~n25510;
  assign n25566 = n25073 & n25494;
  assign n25567 = n25075 & n25490;
  assign n25568 = n25080 & n25493;
  assign n25569 = ~n25566 & ~n25567;
  assign n25570 = ~n25568 & n25569;
  assign n25571 = ~n25564 & ~n25565;
  assign n5629 = ~n25570 | ~n25571;
  assign n25573 = P1_INSTQUEUE_REG_10__0_ & ~n25504;
  assign n25574 = n25090 & ~n25510;
  assign n25575 = n25095 & n25494;
  assign n25576 = n25097 & n25490;
  assign n25577 = n25102 & n25493;
  assign n25578 = ~n25575 & ~n25576;
  assign n25579 = ~n25577 & n25578;
  assign n25580 = ~n25573 & ~n25574;
  assign n5634 = ~n25579 | ~n25580;
  assign n25582 = n24309 & n24457;
  assign n25583 = n25203 & n25395;
  assign n25584 = ~n25582 & ~n25583;
  assign n25585 = n25206 & n25398;
  assign n25586 = n24788 & n24897;
  assign n25587 = ~n25585 & ~n25586;
  assign n25588 = n24913 & n25587;
  assign n25589 = ~n24627 & ~n25588;
  assign n25590 = n25584 & ~n25589;
  assign n25591 = P1_STATE2_REG_3_ & ~n25582;
  assign n25592 = n25214 & n25406;
  assign n25593 = ~n25582 & ~n25592;
  assign n25594 = P1_STATE2_REG_2_ & n25593;
  assign n25595 = ~n25591 & ~n25594;
  assign n25596 = n24912 & n25595;
  assign n25597 = ~n25590 & n25596;
  assign n25598 = P1_INSTQUEUE_REG_9__7_ & ~n25597;
  assign n25599 = P1_STATE2_REG_2_ & ~n25593;
  assign n25600 = n24908 & n25587;
  assign n25601 = ~n24627 & ~n25600;
  assign n25602 = ~n25584 & ~n25601;
  assign n25603 = ~n25599 & ~n25602;
  assign n25604 = n24930 & ~n25603;
  assign n25605 = n24940 & n25586;
  assign n25606 = n24943 & n25582;
  assign n25607 = n24948 & n25585;
  assign n25608 = ~n25605 & ~n25606;
  assign n25609 = ~n25607 & n25608;
  assign n25610 = ~n25598 & ~n25604;
  assign n5639 = ~n25609 | ~n25610;
  assign n25612 = P1_INSTQUEUE_REG_9__6_ & ~n25597;
  assign n25613 = n24958 & ~n25603;
  assign n25614 = n24963 & n25586;
  assign n25615 = n24965 & n25582;
  assign n25616 = n24970 & n25585;
  assign n25617 = ~n25614 & ~n25615;
  assign n25618 = ~n25616 & n25617;
  assign n25619 = ~n25612 & ~n25613;
  assign n5644 = ~n25618 | ~n25619;
  assign n25621 = P1_INSTQUEUE_REG_9__5_ & ~n25597;
  assign n25622 = n24980 & ~n25603;
  assign n25623 = n24985 & n25586;
  assign n25624 = n24987 & n25582;
  assign n25625 = n24992 & n25585;
  assign n25626 = ~n25623 & ~n25624;
  assign n25627 = ~n25625 & n25626;
  assign n25628 = ~n25621 & ~n25622;
  assign n5649 = ~n25627 | ~n25628;
  assign n25630 = P1_INSTQUEUE_REG_9__4_ & ~n25597;
  assign n25631 = n25002 & ~n25603;
  assign n25632 = n25007 & n25586;
  assign n25633 = n25009 & n25582;
  assign n25634 = n25014 & n25585;
  assign n25635 = ~n25632 & ~n25633;
  assign n25636 = ~n25634 & n25635;
  assign n25637 = ~n25630 & ~n25631;
  assign n5654 = ~n25636 | ~n25637;
  assign n25639 = P1_INSTQUEUE_REG_9__3_ & ~n25597;
  assign n25640 = n25024 & ~n25603;
  assign n25641 = n25029 & n25586;
  assign n25642 = n25031 & n25582;
  assign n25643 = n25036 & n25585;
  assign n25644 = ~n25641 & ~n25642;
  assign n25645 = ~n25643 & n25644;
  assign n25646 = ~n25639 & ~n25640;
  assign n5659 = ~n25645 | ~n25646;
  assign n25648 = P1_INSTQUEUE_REG_9__2_ & ~n25597;
  assign n25649 = n25046 & ~n25603;
  assign n25650 = n25051 & n25586;
  assign n25651 = n25053 & n25582;
  assign n25652 = n25058 & n25585;
  assign n25653 = ~n25650 & ~n25651;
  assign n25654 = ~n25652 & n25653;
  assign n25655 = ~n25648 & ~n25649;
  assign n5664 = ~n25654 | ~n25655;
  assign n25657 = P1_INSTQUEUE_REG_9__1_ & ~n25597;
  assign n25658 = n25068 & ~n25603;
  assign n25659 = n25073 & n25586;
  assign n25660 = n25075 & n25582;
  assign n25661 = n25080 & n25585;
  assign n25662 = ~n25659 & ~n25660;
  assign n25663 = ~n25661 & n25662;
  assign n25664 = ~n25657 & ~n25658;
  assign n5669 = ~n25663 | ~n25664;
  assign n25666 = P1_INSTQUEUE_REG_9__0_ & ~n25597;
  assign n25667 = n25090 & ~n25603;
  assign n25668 = n25095 & n25586;
  assign n25669 = n25097 & n25582;
  assign n25670 = n25102 & n25585;
  assign n25671 = ~n25668 & ~n25669;
  assign n25672 = ~n25670 & n25671;
  assign n25673 = ~n25666 & ~n25667;
  assign n5674 = ~n25672 | ~n25673;
  assign n25675 = n24457 & n25298;
  assign n25676 = n25300 & n25395;
  assign n25677 = ~n25675 & ~n25676;
  assign n25678 = n25303 & n25398;
  assign n25679 = n24897 & n25305;
  assign n25680 = ~n25678 & ~n25679;
  assign n25681 = n24913 & n25680;
  assign n25682 = ~n24627 & ~n25681;
  assign n25683 = n25677 & ~n25682;
  assign n25684 = P1_STATE2_REG_3_ & ~n25675;
  assign n25685 = n24311 & n25406;
  assign n25686 = P1_STATE2_REG_2_ & ~n25685;
  assign n25687 = ~n25684 & ~n25686;
  assign n25688 = n24912 & n25687;
  assign n25689 = ~n25683 & n25688;
  assign n25690 = P1_INSTQUEUE_REG_8__7_ & ~n25689;
  assign n25691 = P1_STATE2_REG_2_ & n25685;
  assign n25692 = n24908 & n25680;
  assign n25693 = ~n24627 & ~n25692;
  assign n25694 = ~n25677 & ~n25693;
  assign n25695 = ~n25691 & ~n25694;
  assign n25696 = n24930 & ~n25695;
  assign n25697 = n24940 & n25679;
  assign n25698 = n24943 & n25675;
  assign n25699 = n24948 & n25678;
  assign n25700 = ~n25697 & ~n25698;
  assign n25701 = ~n25699 & n25700;
  assign n25702 = ~n25690 & ~n25696;
  assign n5679 = ~n25701 | ~n25702;
  assign n25704 = P1_INSTQUEUE_REG_8__6_ & ~n25689;
  assign n25705 = n24958 & ~n25695;
  assign n25706 = n24963 & n25679;
  assign n25707 = n24965 & n25675;
  assign n25708 = n24970 & n25678;
  assign n25709 = ~n25706 & ~n25707;
  assign n25710 = ~n25708 & n25709;
  assign n25711 = ~n25704 & ~n25705;
  assign n5684 = ~n25710 | ~n25711;
  assign n25713 = P1_INSTQUEUE_REG_8__5_ & ~n25689;
  assign n25714 = n24980 & ~n25695;
  assign n25715 = n24985 & n25679;
  assign n25716 = n24987 & n25675;
  assign n25717 = n24992 & n25678;
  assign n25718 = ~n25715 & ~n25716;
  assign n25719 = ~n25717 & n25718;
  assign n25720 = ~n25713 & ~n25714;
  assign n5689 = ~n25719 | ~n25720;
  assign n25722 = P1_INSTQUEUE_REG_8__4_ & ~n25689;
  assign n25723 = n25002 & ~n25695;
  assign n25724 = n25007 & n25679;
  assign n25725 = n25009 & n25675;
  assign n25726 = n25014 & n25678;
  assign n25727 = ~n25724 & ~n25725;
  assign n25728 = ~n25726 & n25727;
  assign n25729 = ~n25722 & ~n25723;
  assign n5694 = ~n25728 | ~n25729;
  assign n25731 = P1_INSTQUEUE_REG_8__3_ & ~n25689;
  assign n25732 = n25024 & ~n25695;
  assign n25733 = n25029 & n25679;
  assign n25734 = n25031 & n25675;
  assign n25735 = n25036 & n25678;
  assign n25736 = ~n25733 & ~n25734;
  assign n25737 = ~n25735 & n25736;
  assign n25738 = ~n25731 & ~n25732;
  assign n5699 = ~n25737 | ~n25738;
  assign n25740 = P1_INSTQUEUE_REG_8__2_ & ~n25689;
  assign n25741 = n25046 & ~n25695;
  assign n25742 = n25051 & n25679;
  assign n25743 = n25053 & n25675;
  assign n25744 = n25058 & n25678;
  assign n25745 = ~n25742 & ~n25743;
  assign n25746 = ~n25744 & n25745;
  assign n25747 = ~n25740 & ~n25741;
  assign n5704 = ~n25746 | ~n25747;
  assign n25749 = P1_INSTQUEUE_REG_8__1_ & ~n25689;
  assign n25750 = n25068 & ~n25695;
  assign n25751 = n25073 & n25679;
  assign n25752 = n25075 & n25675;
  assign n25753 = n25080 & n25678;
  assign n25754 = ~n25751 & ~n25752;
  assign n25755 = ~n25753 & n25754;
  assign n25756 = ~n25749 & ~n25750;
  assign n5709 = ~n25755 | ~n25756;
  assign n25758 = P1_INSTQUEUE_REG_8__0_ & ~n25689;
  assign n25759 = n25090 & ~n25695;
  assign n25760 = n25095 & n25679;
  assign n25761 = n25097 & n25675;
  assign n25762 = n25102 & n25678;
  assign n25763 = ~n25760 & ~n25761;
  assign n25764 = ~n25762 & n25763;
  assign n25765 = ~n25758 & ~n25759;
  assign n5714 = ~n25764 | ~n25765;
  assign n25767 = n24397 & n24482;
  assign n25768 = n24623 & n25767;
  assign n25769 = ~n24460 & ~n25768;
  assign n25770 = ~n24846 & n24902;
  assign n25771 = n24790 & n25770;
  assign n25772 = ~n24900 & ~n25771;
  assign n25773 = n24913 & n25772;
  assign n25774 = ~n24627 & ~n25773;
  assign n25775 = n25769 & ~n25774;
  assign n25776 = P1_STATE2_REG_3_ & ~n24460;
  assign n25777 = ~n24384 & n24462;
  assign n25778 = n24919 & n25777;
  assign n25779 = ~n24460 & ~n25778;
  assign n25780 = P1_STATE2_REG_2_ & n25779;
  assign n25781 = ~n25776 & ~n25780;
  assign n25782 = n24912 & n25781;
  assign n25783 = ~n25775 & n25782;
  assign n25784 = P1_INSTQUEUE_REG_7__7_ & ~n25783;
  assign n25785 = P1_STATE2_REG_2_ & ~n25779;
  assign n25786 = n24908 & n25772;
  assign n25787 = ~n24627 & ~n25786;
  assign n25788 = ~n25769 & ~n25787;
  assign n25789 = ~n25785 & ~n25788;
  assign n25790 = n24930 & ~n25789;
  assign n25791 = n24900 & n24940;
  assign n25792 = n24460 & n24943;
  assign n25793 = n24948 & n25771;
  assign n25794 = ~n25791 & ~n25792;
  assign n25795 = ~n25793 & n25794;
  assign n25796 = ~n25784 & ~n25790;
  assign n5719 = ~n25795 | ~n25796;
  assign n25798 = P1_INSTQUEUE_REG_7__6_ & ~n25783;
  assign n25799 = n24958 & ~n25789;
  assign n25800 = n24900 & n24963;
  assign n25801 = n24460 & n24965;
  assign n25802 = n24970 & n25771;
  assign n25803 = ~n25800 & ~n25801;
  assign n25804 = ~n25802 & n25803;
  assign n25805 = ~n25798 & ~n25799;
  assign n5724 = ~n25804 | ~n25805;
  assign n25807 = P1_INSTQUEUE_REG_7__5_ & ~n25783;
  assign n25808 = n24980 & ~n25789;
  assign n25809 = n24900 & n24985;
  assign n25810 = n24460 & n24987;
  assign n25811 = n24992 & n25771;
  assign n25812 = ~n25809 & ~n25810;
  assign n25813 = ~n25811 & n25812;
  assign n25814 = ~n25807 & ~n25808;
  assign n5729 = ~n25813 | ~n25814;
  assign n25816 = P1_INSTQUEUE_REG_7__4_ & ~n25783;
  assign n25817 = n25002 & ~n25789;
  assign n25818 = n24900 & n25007;
  assign n25819 = n24460 & n25009;
  assign n25820 = n25014 & n25771;
  assign n25821 = ~n25818 & ~n25819;
  assign n25822 = ~n25820 & n25821;
  assign n25823 = ~n25816 & ~n25817;
  assign n5734 = ~n25822 | ~n25823;
  assign n25825 = P1_INSTQUEUE_REG_7__3_ & ~n25783;
  assign n25826 = n25024 & ~n25789;
  assign n25827 = n24900 & n25029;
  assign n25828 = n24460 & n25031;
  assign n25829 = n25036 & n25771;
  assign n25830 = ~n25827 & ~n25828;
  assign n25831 = ~n25829 & n25830;
  assign n25832 = ~n25825 & ~n25826;
  assign n5739 = ~n25831 | ~n25832;
  assign n25834 = P1_INSTQUEUE_REG_7__2_ & ~n25783;
  assign n25835 = n25046 & ~n25789;
  assign n25836 = n24900 & n25051;
  assign n25837 = n24460 & n25053;
  assign n25838 = n25058 & n25771;
  assign n25839 = ~n25836 & ~n25837;
  assign n25840 = ~n25838 & n25839;
  assign n25841 = ~n25834 & ~n25835;
  assign n5744 = ~n25840 | ~n25841;
  assign n25843 = P1_INSTQUEUE_REG_7__1_ & ~n25783;
  assign n25844 = n25068 & ~n25789;
  assign n25845 = n24900 & n25073;
  assign n25846 = n24460 & n25075;
  assign n25847 = n25080 & n25771;
  assign n25848 = ~n25845 & ~n25846;
  assign n25849 = ~n25847 & n25848;
  assign n25850 = ~n25843 & ~n25844;
  assign n5749 = ~n25849 | ~n25850;
  assign n25852 = P1_INSTQUEUE_REG_7__0_ & ~n25783;
  assign n25853 = n25090 & ~n25789;
  assign n25854 = n24900 & n25095;
  assign n25855 = n24460 & n25097;
  assign n25856 = n25102 & n25771;
  assign n25857 = ~n25854 & ~n25855;
  assign n25858 = ~n25856 & n25857;
  assign n25859 = ~n25852 & ~n25853;
  assign n5754 = ~n25858 | ~n25859;
  assign n25861 = n24310 & n24459;
  assign n25862 = n25109 & n25767;
  assign n25863 = ~n25861 & ~n25862;
  assign n25864 = n25112 & n25770;
  assign n25865 = n24787 & n24899;
  assign n25866 = ~n25864 & ~n25865;
  assign n25867 = n24913 & n25866;
  assign n25868 = ~n24627 & ~n25867;
  assign n25869 = n25863 & ~n25868;
  assign n25870 = P1_STATE2_REG_3_ & ~n25861;
  assign n25871 = ~n24311 & n25777;
  assign n25872 = P1_STATE2_REG_2_ & ~n25871;
  assign n25873 = ~n25870 & ~n25872;
  assign n25874 = n24912 & n25873;
  assign n25875 = ~n25869 & n25874;
  assign n25876 = P1_INSTQUEUE_REG_6__7_ & ~n25875;
  assign n25877 = P1_STATE2_REG_2_ & n25871;
  assign n25878 = n24908 & n25866;
  assign n25879 = ~n24627 & ~n25878;
  assign n25880 = ~n25863 & ~n25879;
  assign n25881 = ~n25877 & ~n25880;
  assign n25882 = n24930 & ~n25881;
  assign n25883 = n24940 & n25865;
  assign n25884 = n24943 & n25861;
  assign n25885 = n24948 & n25864;
  assign n25886 = ~n25883 & ~n25884;
  assign n25887 = ~n25885 & n25886;
  assign n25888 = ~n25876 & ~n25882;
  assign n5759 = ~n25887 | ~n25888;
  assign n25890 = P1_INSTQUEUE_REG_6__6_ & ~n25875;
  assign n25891 = n24958 & ~n25881;
  assign n25892 = n24963 & n25865;
  assign n25893 = n24965 & n25861;
  assign n25894 = n24970 & n25864;
  assign n25895 = ~n25892 & ~n25893;
  assign n25896 = ~n25894 & n25895;
  assign n25897 = ~n25890 & ~n25891;
  assign n5764 = ~n25896 | ~n25897;
  assign n25899 = P1_INSTQUEUE_REG_6__5_ & ~n25875;
  assign n25900 = n24980 & ~n25881;
  assign n25901 = n24985 & n25865;
  assign n25902 = n24987 & n25861;
  assign n25903 = n24992 & n25864;
  assign n25904 = ~n25901 & ~n25902;
  assign n25905 = ~n25903 & n25904;
  assign n25906 = ~n25899 & ~n25900;
  assign n5769 = ~n25905 | ~n25906;
  assign n25908 = P1_INSTQUEUE_REG_6__4_ & ~n25875;
  assign n25909 = n25002 & ~n25881;
  assign n25910 = n25007 & n25865;
  assign n25911 = n25009 & n25861;
  assign n25912 = n25014 & n25864;
  assign n25913 = ~n25910 & ~n25911;
  assign n25914 = ~n25912 & n25913;
  assign n25915 = ~n25908 & ~n25909;
  assign n5774 = ~n25914 | ~n25915;
  assign n25917 = P1_INSTQUEUE_REG_6__3_ & ~n25875;
  assign n25918 = n25024 & ~n25881;
  assign n25919 = n25029 & n25865;
  assign n25920 = n25031 & n25861;
  assign n25921 = n25036 & n25864;
  assign n25922 = ~n25919 & ~n25920;
  assign n25923 = ~n25921 & n25922;
  assign n25924 = ~n25917 & ~n25918;
  assign n5779 = ~n25923 | ~n25924;
  assign n25926 = P1_INSTQUEUE_REG_6__2_ & ~n25875;
  assign n25927 = n25046 & ~n25881;
  assign n25928 = n25051 & n25865;
  assign n25929 = n25053 & n25861;
  assign n25930 = n25058 & n25864;
  assign n25931 = ~n25928 & ~n25929;
  assign n25932 = ~n25930 & n25931;
  assign n25933 = ~n25926 & ~n25927;
  assign n5784 = ~n25932 | ~n25933;
  assign n25935 = P1_INSTQUEUE_REG_6__1_ & ~n25875;
  assign n25936 = n25068 & ~n25881;
  assign n25937 = n25073 & n25865;
  assign n25938 = n25075 & n25861;
  assign n25939 = n25080 & n25864;
  assign n25940 = ~n25937 & ~n25938;
  assign n25941 = ~n25939 & n25940;
  assign n25942 = ~n25935 & ~n25936;
  assign n5789 = ~n25941 | ~n25942;
  assign n25944 = P1_INSTQUEUE_REG_6__0_ & ~n25875;
  assign n25945 = n25090 & ~n25881;
  assign n25946 = n25095 & n25865;
  assign n25947 = n25097 & n25861;
  assign n25948 = n25102 & n25864;
  assign n25949 = ~n25946 & ~n25947;
  assign n25950 = ~n25948 & n25949;
  assign n25951 = ~n25944 & ~n25945;
  assign n5794 = ~n25950 | ~n25951;
  assign n25953 = n24309 & n24459;
  assign n25954 = n25203 & n25767;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = n25206 & n25770;
  assign n25957 = n24788 & n24899;
  assign n25958 = ~n25956 & ~n25957;
  assign n25959 = n24913 & n25958;
  assign n25960 = ~n24627 & ~n25959;
  assign n25961 = n25955 & ~n25960;
  assign n25962 = P1_STATE2_REG_3_ & ~n25953;
  assign n25963 = n25214 & n25777;
  assign n25964 = ~n25953 & ~n25963;
  assign n25965 = P1_STATE2_REG_2_ & n25964;
  assign n25966 = ~n25962 & ~n25965;
  assign n25967 = n24912 & n25966;
  assign n25968 = ~n25961 & n25967;
  assign n25969 = P1_INSTQUEUE_REG_5__7_ & ~n25968;
  assign n25970 = P1_STATE2_REG_2_ & ~n25964;
  assign n25971 = n24908 & n25958;
  assign n25972 = ~n24627 & ~n25971;
  assign n25973 = ~n25955 & ~n25972;
  assign n25974 = ~n25970 & ~n25973;
  assign n25975 = n24930 & ~n25974;
  assign n25976 = n24940 & n25957;
  assign n25977 = n24943 & n25953;
  assign n25978 = n24948 & n25956;
  assign n25979 = ~n25976 & ~n25977;
  assign n25980 = ~n25978 & n25979;
  assign n25981 = ~n25969 & ~n25975;
  assign n5799 = ~n25980 | ~n25981;
  assign n25983 = P1_INSTQUEUE_REG_5__6_ & ~n25968;
  assign n25984 = n24958 & ~n25974;
  assign n25985 = n24963 & n25957;
  assign n25986 = n24965 & n25953;
  assign n25987 = n24970 & n25956;
  assign n25988 = ~n25985 & ~n25986;
  assign n25989 = ~n25987 & n25988;
  assign n25990 = ~n25983 & ~n25984;
  assign n5804 = ~n25989 | ~n25990;
  assign n25992 = P1_INSTQUEUE_REG_5__5_ & ~n25968;
  assign n25993 = n24980 & ~n25974;
  assign n25994 = n24985 & n25957;
  assign n25995 = n24987 & n25953;
  assign n25996 = n24992 & n25956;
  assign n25997 = ~n25994 & ~n25995;
  assign n25998 = ~n25996 & n25997;
  assign n25999 = ~n25992 & ~n25993;
  assign n5809 = ~n25998 | ~n25999;
  assign n26001 = P1_INSTQUEUE_REG_5__4_ & ~n25968;
  assign n26002 = n25002 & ~n25974;
  assign n26003 = n25007 & n25957;
  assign n26004 = n25009 & n25953;
  assign n26005 = n25014 & n25956;
  assign n26006 = ~n26003 & ~n26004;
  assign n26007 = ~n26005 & n26006;
  assign n26008 = ~n26001 & ~n26002;
  assign n5814 = ~n26007 | ~n26008;
  assign n26010 = P1_INSTQUEUE_REG_5__3_ & ~n25968;
  assign n26011 = n25024 & ~n25974;
  assign n26012 = n25029 & n25957;
  assign n26013 = n25031 & n25953;
  assign n26014 = n25036 & n25956;
  assign n26015 = ~n26012 & ~n26013;
  assign n26016 = ~n26014 & n26015;
  assign n26017 = ~n26010 & ~n26011;
  assign n5819 = ~n26016 | ~n26017;
  assign n26019 = P1_INSTQUEUE_REG_5__2_ & ~n25968;
  assign n26020 = n25046 & ~n25974;
  assign n26021 = n25051 & n25957;
  assign n26022 = n25053 & n25953;
  assign n26023 = n25058 & n25956;
  assign n26024 = ~n26021 & ~n26022;
  assign n26025 = ~n26023 & n26024;
  assign n26026 = ~n26019 & ~n26020;
  assign n5824 = ~n26025 | ~n26026;
  assign n26028 = P1_INSTQUEUE_REG_5__1_ & ~n25968;
  assign n26029 = n25068 & ~n25974;
  assign n26030 = n25073 & n25957;
  assign n26031 = n25075 & n25953;
  assign n26032 = n25080 & n25956;
  assign n26033 = ~n26030 & ~n26031;
  assign n26034 = ~n26032 & n26033;
  assign n26035 = ~n26028 & ~n26029;
  assign n5829 = ~n26034 | ~n26035;
  assign n26037 = P1_INSTQUEUE_REG_5__0_ & ~n25968;
  assign n26038 = n25090 & ~n25974;
  assign n26039 = n25095 & n25957;
  assign n26040 = n25097 & n25953;
  assign n26041 = n25102 & n25956;
  assign n26042 = ~n26039 & ~n26040;
  assign n26043 = ~n26041 & n26042;
  assign n26044 = ~n26037 & ~n26038;
  assign n5834 = ~n26043 | ~n26044;
  assign n26046 = n24459 & n25298;
  assign n26047 = n25300 & n25767;
  assign n26048 = ~n26046 & ~n26047;
  assign n26049 = n25303 & n25770;
  assign n26050 = n24899 & n25305;
  assign n26051 = ~n26049 & ~n26050;
  assign n26052 = n24913 & n26051;
  assign n26053 = ~n24627 & ~n26052;
  assign n26054 = n26048 & ~n26053;
  assign n26055 = P1_STATE2_REG_3_ & ~n26046;
  assign n26056 = n24311 & n25777;
  assign n26057 = P1_STATE2_REG_2_ & ~n26056;
  assign n26058 = ~n26055 & ~n26057;
  assign n26059 = n24912 & n26058;
  assign n26060 = ~n26054 & n26059;
  assign n26061 = P1_INSTQUEUE_REG_4__7_ & ~n26060;
  assign n26062 = P1_STATE2_REG_2_ & n26056;
  assign n26063 = n24908 & n26051;
  assign n26064 = ~n24627 & ~n26063;
  assign n26065 = ~n26048 & ~n26064;
  assign n26066 = ~n26062 & ~n26065;
  assign n26067 = n24930 & ~n26066;
  assign n26068 = n24940 & n26050;
  assign n26069 = n24943 & n26046;
  assign n26070 = n24948 & n26049;
  assign n26071 = ~n26068 & ~n26069;
  assign n26072 = ~n26070 & n26071;
  assign n26073 = ~n26061 & ~n26067;
  assign n5839 = ~n26072 | ~n26073;
  assign n26075 = P1_INSTQUEUE_REG_4__6_ & ~n26060;
  assign n26076 = n24958 & ~n26066;
  assign n26077 = n24963 & n26050;
  assign n26078 = n24965 & n26046;
  assign n26079 = n24970 & n26049;
  assign n26080 = ~n26077 & ~n26078;
  assign n26081 = ~n26079 & n26080;
  assign n26082 = ~n26075 & ~n26076;
  assign n5844 = ~n26081 | ~n26082;
  assign n26084 = P1_INSTQUEUE_REG_4__5_ & ~n26060;
  assign n26085 = n24980 & ~n26066;
  assign n26086 = n24985 & n26050;
  assign n26087 = n24987 & n26046;
  assign n26088 = n24992 & n26049;
  assign n26089 = ~n26086 & ~n26087;
  assign n26090 = ~n26088 & n26089;
  assign n26091 = ~n26084 & ~n26085;
  assign n5849 = ~n26090 | ~n26091;
  assign n26093 = P1_INSTQUEUE_REG_4__4_ & ~n26060;
  assign n26094 = n25002 & ~n26066;
  assign n26095 = n25007 & n26050;
  assign n26096 = n25009 & n26046;
  assign n26097 = n25014 & n26049;
  assign n26098 = ~n26095 & ~n26096;
  assign n26099 = ~n26097 & n26098;
  assign n26100 = ~n26093 & ~n26094;
  assign n5854 = ~n26099 | ~n26100;
  assign n26102 = P1_INSTQUEUE_REG_4__3_ & ~n26060;
  assign n26103 = n25024 & ~n26066;
  assign n26104 = n25029 & n26050;
  assign n26105 = n25031 & n26046;
  assign n26106 = n25036 & n26049;
  assign n26107 = ~n26104 & ~n26105;
  assign n26108 = ~n26106 & n26107;
  assign n26109 = ~n26102 & ~n26103;
  assign n5859 = ~n26108 | ~n26109;
  assign n26111 = P1_INSTQUEUE_REG_4__2_ & ~n26060;
  assign n26112 = n25046 & ~n26066;
  assign n26113 = n25051 & n26050;
  assign n26114 = n25053 & n26046;
  assign n26115 = n25058 & n26049;
  assign n26116 = ~n26113 & ~n26114;
  assign n26117 = ~n26115 & n26116;
  assign n26118 = ~n26111 & ~n26112;
  assign n5864 = ~n26117 | ~n26118;
  assign n26120 = P1_INSTQUEUE_REG_4__1_ & ~n26060;
  assign n26121 = n25068 & ~n26066;
  assign n26122 = n25073 & n26050;
  assign n26123 = n25075 & n26046;
  assign n26124 = n25080 & n26049;
  assign n26125 = ~n26122 & ~n26123;
  assign n26126 = ~n26124 & n26125;
  assign n26127 = ~n26120 & ~n26121;
  assign n5869 = ~n26126 | ~n26127;
  assign n26129 = P1_INSTQUEUE_REG_4__0_ & ~n26060;
  assign n26130 = n25090 & ~n26066;
  assign n26131 = n25095 & n26050;
  assign n26132 = n25097 & n26046;
  assign n26133 = n25102 & n26049;
  assign n26134 = ~n26131 & ~n26132;
  assign n26135 = ~n26133 & n26134;
  assign n26136 = ~n26129 & ~n26130;
  assign n5874 = ~n26135 | ~n26136;
  assign n26138 = ~P1_INSTQUEUEWR_ADDR_REG_3_ & ~P1_INSTQUEUEWR_ADDR_REG_2_;
  assign n26139 = n24381 & n26138;
  assign n26140 = ~n24397 & n24482;
  assign n26141 = n24623 & n26140;
  assign n26142 = ~n26139 & ~n26141;
  assign n26143 = n24846 & n24902;
  assign n26144 = n24790 & n26143;
  assign n26145 = n24843 & ~n24896;
  assign n26146 = n24791 & n26145;
  assign n26147 = ~n26144 & ~n26146;
  assign n26148 = n24913 & n26147;
  assign n26149 = ~n24627 & ~n26148;
  assign n26150 = n26142 & ~n26149;
  assign n26151 = P1_STATE2_REG_3_ & ~n26139;
  assign n26152 = n24384 & n24462;
  assign n26153 = n24919 & n26152;
  assign n26154 = ~n26139 & ~n26153;
  assign n26155 = P1_STATE2_REG_2_ & n26154;
  assign n26156 = ~n26151 & ~n26155;
  assign n26157 = n24912 & n26156;
  assign n26158 = ~n26150 & n26157;
  assign n26159 = P1_INSTQUEUE_REG_3__7_ & ~n26158;
  assign n26160 = P1_STATE2_REG_2_ & ~n26154;
  assign n26161 = n24908 & n26147;
  assign n26162 = ~n24627 & ~n26161;
  assign n26163 = ~n26142 & ~n26162;
  assign n26164 = ~n26160 & ~n26163;
  assign n26165 = n24930 & ~n26164;
  assign n26166 = n24940 & n26146;
  assign n26167 = n24943 & n26139;
  assign n26168 = n24948 & n26144;
  assign n26169 = ~n26166 & ~n26167;
  assign n26170 = ~n26168 & n26169;
  assign n26171 = ~n26159 & ~n26165;
  assign n5879 = ~n26170 | ~n26171;
  assign n26173 = P1_INSTQUEUE_REG_3__6_ & ~n26158;
  assign n26174 = n24958 & ~n26164;
  assign n26175 = n24963 & n26146;
  assign n26176 = n24965 & n26139;
  assign n26177 = n24970 & n26144;
  assign n26178 = ~n26175 & ~n26176;
  assign n26179 = ~n26177 & n26178;
  assign n26180 = ~n26173 & ~n26174;
  assign n5884 = ~n26179 | ~n26180;
  assign n26182 = P1_INSTQUEUE_REG_3__5_ & ~n26158;
  assign n26183 = n24980 & ~n26164;
  assign n26184 = n24985 & n26146;
  assign n26185 = n24987 & n26139;
  assign n26186 = n24992 & n26144;
  assign n26187 = ~n26184 & ~n26185;
  assign n26188 = ~n26186 & n26187;
  assign n26189 = ~n26182 & ~n26183;
  assign n5889 = ~n26188 | ~n26189;
  assign n26191 = P1_INSTQUEUE_REG_3__4_ & ~n26158;
  assign n26192 = n25002 & ~n26164;
  assign n26193 = n25007 & n26146;
  assign n26194 = n25009 & n26139;
  assign n26195 = n25014 & n26144;
  assign n26196 = ~n26193 & ~n26194;
  assign n26197 = ~n26195 & n26196;
  assign n26198 = ~n26191 & ~n26192;
  assign n5894 = ~n26197 | ~n26198;
  assign n26200 = P1_INSTQUEUE_REG_3__3_ & ~n26158;
  assign n26201 = n25024 & ~n26164;
  assign n26202 = n25029 & n26146;
  assign n26203 = n25031 & n26139;
  assign n26204 = n25036 & n26144;
  assign n26205 = ~n26202 & ~n26203;
  assign n26206 = ~n26204 & n26205;
  assign n26207 = ~n26200 & ~n26201;
  assign n5899 = ~n26206 | ~n26207;
  assign n26209 = P1_INSTQUEUE_REG_3__2_ & ~n26158;
  assign n26210 = n25046 & ~n26164;
  assign n26211 = n25051 & n26146;
  assign n26212 = n25053 & n26139;
  assign n26213 = n25058 & n26144;
  assign n26214 = ~n26211 & ~n26212;
  assign n26215 = ~n26213 & n26214;
  assign n26216 = ~n26209 & ~n26210;
  assign n5904 = ~n26215 | ~n26216;
  assign n26218 = P1_INSTQUEUE_REG_3__1_ & ~n26158;
  assign n26219 = n25068 & ~n26164;
  assign n26220 = n25073 & n26146;
  assign n26221 = n25075 & n26139;
  assign n26222 = n25080 & n26144;
  assign n26223 = ~n26220 & ~n26221;
  assign n26224 = ~n26222 & n26223;
  assign n26225 = ~n26218 & ~n26219;
  assign n5909 = ~n26224 | ~n26225;
  assign n26227 = P1_INSTQUEUE_REG_3__0_ & ~n26158;
  assign n26228 = n25090 & ~n26164;
  assign n26229 = n25095 & n26146;
  assign n26230 = n25097 & n26139;
  assign n26231 = n25102 & n26144;
  assign n26232 = ~n26229 & ~n26230;
  assign n26233 = ~n26231 & n26232;
  assign n26234 = ~n26227 & ~n26228;
  assign n5914 = ~n26233 | ~n26234;
  assign n26236 = n24310 & n26138;
  assign n26237 = n25109 & n26140;
  assign n26238 = ~n26236 & ~n26237;
  assign n26239 = n25112 & n26143;
  assign n26240 = n24787 & n26145;
  assign n26241 = ~n26239 & ~n26240;
  assign n26242 = n24913 & n26241;
  assign n26243 = ~n24627 & ~n26242;
  assign n26244 = n26238 & ~n26243;
  assign n26245 = P1_STATE2_REG_3_ & ~n26236;
  assign n26246 = ~n24311 & n26152;
  assign n26247 = P1_STATE2_REG_2_ & ~n26246;
  assign n26248 = ~n26245 & ~n26247;
  assign n26249 = n24912 & n26248;
  assign n26250 = ~n26244 & n26249;
  assign n26251 = P1_INSTQUEUE_REG_2__7_ & ~n26250;
  assign n26252 = P1_STATE2_REG_2_ & n26246;
  assign n26253 = n24908 & n26241;
  assign n26254 = ~n24627 & ~n26253;
  assign n26255 = ~n26238 & ~n26254;
  assign n26256 = ~n26252 & ~n26255;
  assign n26257 = n24930 & ~n26256;
  assign n26258 = n24940 & n26240;
  assign n26259 = n24943 & n26236;
  assign n26260 = n24948 & n26239;
  assign n26261 = ~n26258 & ~n26259;
  assign n26262 = ~n26260 & n26261;
  assign n26263 = ~n26251 & ~n26257;
  assign n5919 = ~n26262 | ~n26263;
  assign n26265 = P1_INSTQUEUE_REG_2__6_ & ~n26250;
  assign n26266 = n24958 & ~n26256;
  assign n26267 = n24963 & n26240;
  assign n26268 = n24965 & n26236;
  assign n26269 = n24970 & n26239;
  assign n26270 = ~n26267 & ~n26268;
  assign n26271 = ~n26269 & n26270;
  assign n26272 = ~n26265 & ~n26266;
  assign n5924 = ~n26271 | ~n26272;
  assign n26274 = P1_INSTQUEUE_REG_2__5_ & ~n26250;
  assign n26275 = n24980 & ~n26256;
  assign n26276 = n24985 & n26240;
  assign n26277 = n24987 & n26236;
  assign n26278 = n24992 & n26239;
  assign n26279 = ~n26276 & ~n26277;
  assign n26280 = ~n26278 & n26279;
  assign n26281 = ~n26274 & ~n26275;
  assign n5929 = ~n26280 | ~n26281;
  assign n26283 = P1_INSTQUEUE_REG_2__4_ & ~n26250;
  assign n26284 = n25002 & ~n26256;
  assign n26285 = n25007 & n26240;
  assign n26286 = n25009 & n26236;
  assign n26287 = n25014 & n26239;
  assign n26288 = ~n26285 & ~n26286;
  assign n26289 = ~n26287 & n26288;
  assign n26290 = ~n26283 & ~n26284;
  assign n5934 = ~n26289 | ~n26290;
  assign n26292 = P1_INSTQUEUE_REG_2__3_ & ~n26250;
  assign n26293 = n25024 & ~n26256;
  assign n26294 = n25029 & n26240;
  assign n26295 = n25031 & n26236;
  assign n26296 = n25036 & n26239;
  assign n26297 = ~n26294 & ~n26295;
  assign n26298 = ~n26296 & n26297;
  assign n26299 = ~n26292 & ~n26293;
  assign n5939 = ~n26298 | ~n26299;
  assign n26301 = P1_INSTQUEUE_REG_2__2_ & ~n26250;
  assign n26302 = n25046 & ~n26256;
  assign n26303 = n25051 & n26240;
  assign n26304 = n25053 & n26236;
  assign n26305 = n25058 & n26239;
  assign n26306 = ~n26303 & ~n26304;
  assign n26307 = ~n26305 & n26306;
  assign n26308 = ~n26301 & ~n26302;
  assign n5944 = ~n26307 | ~n26308;
  assign n26310 = P1_INSTQUEUE_REG_2__1_ & ~n26250;
  assign n26311 = n25068 & ~n26256;
  assign n26312 = n25073 & n26240;
  assign n26313 = n25075 & n26236;
  assign n26314 = n25080 & n26239;
  assign n26315 = ~n26312 & ~n26313;
  assign n26316 = ~n26314 & n26315;
  assign n26317 = ~n26310 & ~n26311;
  assign n5949 = ~n26316 | ~n26317;
  assign n26319 = P1_INSTQUEUE_REG_2__0_ & ~n26250;
  assign n26320 = n25090 & ~n26256;
  assign n26321 = n25095 & n26240;
  assign n26322 = n25097 & n26236;
  assign n26323 = n25102 & n26239;
  assign n26324 = ~n26321 & ~n26322;
  assign n26325 = ~n26323 & n26324;
  assign n26326 = ~n26319 & ~n26320;
  assign n5954 = ~n26325 | ~n26326;
  assign n26328 = n24309 & n26138;
  assign n26329 = n25203 & n26140;
  assign n26330 = ~n26328 & ~n26329;
  assign n26331 = n25206 & n26143;
  assign n26332 = n24788 & n26145;
  assign n26333 = ~n26331 & ~n26332;
  assign n26334 = n24913 & n26333;
  assign n26335 = ~n24627 & ~n26334;
  assign n26336 = n26330 & ~n26335;
  assign n26337 = P1_STATE2_REG_3_ & ~n26328;
  assign n26338 = n25214 & n26152;
  assign n26339 = ~n26328 & ~n26338;
  assign n26340 = P1_STATE2_REG_2_ & n26339;
  assign n26341 = ~n26337 & ~n26340;
  assign n26342 = n24912 & n26341;
  assign n26343 = ~n26336 & n26342;
  assign n26344 = P1_INSTQUEUE_REG_1__7_ & ~n26343;
  assign n26345 = P1_STATE2_REG_2_ & ~n26339;
  assign n26346 = n24908 & n26333;
  assign n26347 = ~n24627 & ~n26346;
  assign n26348 = ~n26330 & ~n26347;
  assign n26349 = ~n26345 & ~n26348;
  assign n26350 = n24930 & ~n26349;
  assign n26351 = n24940 & n26332;
  assign n26352 = n24943 & n26328;
  assign n26353 = n24948 & n26331;
  assign n26354 = ~n26351 & ~n26352;
  assign n26355 = ~n26353 & n26354;
  assign n26356 = ~n26344 & ~n26350;
  assign n5959 = ~n26355 | ~n26356;
  assign n26358 = P1_INSTQUEUE_REG_1__6_ & ~n26343;
  assign n26359 = n24958 & ~n26349;
  assign n26360 = n24963 & n26332;
  assign n26361 = n24965 & n26328;
  assign n26362 = n24970 & n26331;
  assign n26363 = ~n26360 & ~n26361;
  assign n26364 = ~n26362 & n26363;
  assign n26365 = ~n26358 & ~n26359;
  assign n5964 = ~n26364 | ~n26365;
  assign n26367 = P1_INSTQUEUE_REG_1__5_ & ~n26343;
  assign n26368 = n24980 & ~n26349;
  assign n26369 = n24985 & n26332;
  assign n26370 = n24987 & n26328;
  assign n26371 = n24992 & n26331;
  assign n26372 = ~n26369 & ~n26370;
  assign n26373 = ~n26371 & n26372;
  assign n26374 = ~n26367 & ~n26368;
  assign n5969 = ~n26373 | ~n26374;
  assign n26376 = P1_INSTQUEUE_REG_1__4_ & ~n26343;
  assign n26377 = n25002 & ~n26349;
  assign n26378 = n25007 & n26332;
  assign n26379 = n25009 & n26328;
  assign n26380 = n25014 & n26331;
  assign n26381 = ~n26378 & ~n26379;
  assign n26382 = ~n26380 & n26381;
  assign n26383 = ~n26376 & ~n26377;
  assign n5974 = ~n26382 | ~n26383;
  assign n26385 = P1_INSTQUEUE_REG_1__3_ & ~n26343;
  assign n26386 = n25024 & ~n26349;
  assign n26387 = n25029 & n26332;
  assign n26388 = n25031 & n26328;
  assign n26389 = n25036 & n26331;
  assign n26390 = ~n26387 & ~n26388;
  assign n26391 = ~n26389 & n26390;
  assign n26392 = ~n26385 & ~n26386;
  assign n5979 = ~n26391 | ~n26392;
  assign n26394 = P1_INSTQUEUE_REG_1__2_ & ~n26343;
  assign n26395 = n25046 & ~n26349;
  assign n26396 = n25051 & n26332;
  assign n26397 = n25053 & n26328;
  assign n26398 = n25058 & n26331;
  assign n26399 = ~n26396 & ~n26397;
  assign n26400 = ~n26398 & n26399;
  assign n26401 = ~n26394 & ~n26395;
  assign n5984 = ~n26400 | ~n26401;
  assign n26403 = P1_INSTQUEUE_REG_1__1_ & ~n26343;
  assign n26404 = n25068 & ~n26349;
  assign n26405 = n25073 & n26332;
  assign n26406 = n25075 & n26328;
  assign n26407 = n25080 & n26331;
  assign n26408 = ~n26405 & ~n26406;
  assign n26409 = ~n26407 & n26408;
  assign n26410 = ~n26403 & ~n26404;
  assign n5989 = ~n26409 | ~n26410;
  assign n26412 = P1_INSTQUEUE_REG_1__0_ & ~n26343;
  assign n26413 = n25090 & ~n26349;
  assign n26414 = n25095 & n26332;
  assign n26415 = n25097 & n26328;
  assign n26416 = n25102 & n26331;
  assign n26417 = ~n26414 & ~n26415;
  assign n26418 = ~n26416 & n26417;
  assign n26419 = ~n26412 & ~n26413;
  assign n5994 = ~n26418 | ~n26419;
  assign n26421 = n25298 & n26138;
  assign n26422 = n25300 & n26140;
  assign n26423 = ~n26421 & ~n26422;
  assign n26424 = n25303 & n26143;
  assign n26425 = n25305 & n26145;
  assign n26426 = ~n26424 & ~n26425;
  assign n26427 = n24913 & n26426;
  assign n26428 = ~n24627 & ~n26427;
  assign n26429 = n26423 & ~n26428;
  assign n26430 = P1_STATE2_REG_3_ & ~n26421;
  assign n26431 = n24311 & n26152;
  assign n26432 = P1_STATE2_REG_2_ & ~n26431;
  assign n26433 = ~n26430 & ~n26432;
  assign n26434 = n24912 & n26433;
  assign n26435 = ~n26429 & n26434;
  assign n26436 = P1_INSTQUEUE_REG_0__7_ & ~n26435;
  assign n26437 = P1_STATE2_REG_2_ & n26431;
  assign n26438 = n24908 & n26426;
  assign n26439 = ~n24627 & ~n26438;
  assign n26440 = ~n26423 & ~n26439;
  assign n26441 = ~n26437 & ~n26440;
  assign n26442 = n24930 & ~n26441;
  assign n26443 = n24940 & n26425;
  assign n26444 = n24943 & n26421;
  assign n26445 = n24948 & n26424;
  assign n26446 = ~n26443 & ~n26444;
  assign n26447 = ~n26445 & n26446;
  assign n26448 = ~n26436 & ~n26442;
  assign n5999 = ~n26447 | ~n26448;
  assign n26450 = P1_INSTQUEUE_REG_0__6_ & ~n26435;
  assign n26451 = n24958 & ~n26441;
  assign n26452 = n24963 & n26425;
  assign n26453 = n24965 & n26421;
  assign n26454 = n24970 & n26424;
  assign n26455 = ~n26452 & ~n26453;
  assign n26456 = ~n26454 & n26455;
  assign n26457 = ~n26450 & ~n26451;
  assign n6004 = ~n26456 | ~n26457;
  assign n26459 = P1_INSTQUEUE_REG_0__5_ & ~n26435;
  assign n26460 = n24980 & ~n26441;
  assign n26461 = n24985 & n26425;
  assign n26462 = n24987 & n26421;
  assign n26463 = n24992 & n26424;
  assign n26464 = ~n26461 & ~n26462;
  assign n26465 = ~n26463 & n26464;
  assign n26466 = ~n26459 & ~n26460;
  assign n6009 = ~n26465 | ~n26466;
  assign n26468 = P1_INSTQUEUE_REG_0__4_ & ~n26435;
  assign n26469 = n25002 & ~n26441;
  assign n26470 = n25007 & n26425;
  assign n26471 = n25009 & n26421;
  assign n26472 = n25014 & n26424;
  assign n26473 = ~n26470 & ~n26471;
  assign n26474 = ~n26472 & n26473;
  assign n26475 = ~n26468 & ~n26469;
  assign n6014 = ~n26474 | ~n26475;
  assign n26477 = P1_INSTQUEUE_REG_0__3_ & ~n26435;
  assign n26478 = n25024 & ~n26441;
  assign n26479 = n25029 & n26425;
  assign n26480 = n25031 & n26421;
  assign n26481 = n25036 & n26424;
  assign n26482 = ~n26479 & ~n26480;
  assign n26483 = ~n26481 & n26482;
  assign n26484 = ~n26477 & ~n26478;
  assign n6019 = ~n26483 | ~n26484;
  assign n26486 = P1_INSTQUEUE_REG_0__2_ & ~n26435;
  assign n26487 = n25046 & ~n26441;
  assign n26488 = n25051 & n26425;
  assign n26489 = n25053 & n26421;
  assign n26490 = n25058 & n26424;
  assign n26491 = ~n26488 & ~n26489;
  assign n26492 = ~n26490 & n26491;
  assign n26493 = ~n26486 & ~n26487;
  assign n6024 = ~n26492 | ~n26493;
  assign n26495 = P1_INSTQUEUE_REG_0__1_ & ~n26435;
  assign n26496 = n25068 & ~n26441;
  assign n26497 = n25073 & n26425;
  assign n26498 = n25075 & n26421;
  assign n26499 = n25080 & n26424;
  assign n26500 = ~n26497 & ~n26498;
  assign n26501 = ~n26499 & n26500;
  assign n26502 = ~n26495 & ~n26496;
  assign n6029 = ~n26501 | ~n26502;
  assign n26504 = P1_INSTQUEUE_REG_0__0_ & ~n26435;
  assign n26505 = n25090 & ~n26441;
  assign n26506 = n25095 & n26425;
  assign n26507 = n25097 & n26421;
  assign n26508 = n25102 & n26424;
  assign n26509 = ~n26506 & ~n26507;
  assign n26510 = ~n26508 & n26509;
  assign n26511 = ~n26504 & ~n26505;
  assign n6034 = ~n26510 | ~n26511;
  assign n26513 = P1_STATE2_REG_3_ & ~P1_STATE2_REG_0_;
  assign n26514 = P1_STATE2_REG_0_ & P1_FLUSH_REG;
  assign n26515 = n23609 & n26514;
  assign n26516 = ~n26513 & ~n26515;
  assign n26517 = ~n24446 & n24576;
  assign n26518 = n26516 & ~n26517;
  assign n26519 = P1_INSTQUEUERD_ADDR_REG_4_ & n26518;
  assign n26520 = n24170 & n24307;
  assign n26521 = ~n24472 & n26520;
  assign n26522 = ~n26518 & n26521;
  assign n6039 = n26519 | n26522;
  assign n26524 = n24307 & ~n24497;
  assign n26525 = ~n24488 & n24590;
  assign n26526 = ~n26524 & ~n26525;
  assign n26527 = ~n26518 & ~n26526;
  assign n26528 = P1_INSTQUEUERD_ADDR_REG_3_ & n26518;
  assign n6044 = n26527 | n26528;
  assign n26530 = n24307 & ~n24420;
  assign n26531 = n24207 & ~n24213;
  assign n26532 = ~n24222 & n24590;
  assign n26533 = ~n26530 & ~n26531;
  assign n26534 = ~n26532 & n26533;
  assign n26535 = ~n26518 & ~n26534;
  assign n26536 = P1_INSTQUEUERD_ADDR_REG_2_ & n26518;
  assign n6049 = n26535 | n26536;
  assign n26538 = n24307 & ~n24537;
  assign n26539 = n24207 & n24213;
  assign n26540 = n24529 & n24590;
  assign n26541 = ~n26538 & ~n26539;
  assign n26542 = ~n26540 & n26541;
  assign n26543 = ~n26518 & ~n26542;
  assign n26544 = P1_INSTQUEUERD_ADDR_REG_1_ & n26518;
  assign n6054 = n26543 | n26544;
  assign n26546 = n24307 & ~n24522;
  assign n26547 = P1_STATE2_REG_1_ & n24206;
  assign n26548 = ~P1_INSTQUEUERD_ADDR_REG_0_ & n24590;
  assign n26549 = ~n26546 & ~n26547;
  assign n26550 = ~n26548 & n26549;
  assign n26551 = ~n26518 & ~n26550;
  assign n26552 = P1_INSTQUEUERD_ADDR_REG_0_ & n26518;
  assign n6059 = n26551 | n26552;
  assign n26554 = P1_STATE2_REG_0_ & n23609;
  assign n26555 = ~n24609 & n26554;
  assign n26556 = ~n24912 & ~n26515;
  assign n26557 = ~n26555 & n26556;
  assign n6064 = P1_INSTQUEUEWR_ADDR_REG_4_ & n26557;
  assign n26559 = ~P1_STATE2_REG_3_ & P1_STATE2_REG_1_;
  assign n26560 = ~n24482 & ~n26559;
  assign n26561 = n24627 & n24896;
  assign n26562 = ~n26560 & ~n26561;
  assign n26563 = n24790 & ~n24846;
  assign n26564 = ~n24902 & ~n26563;
  assign n26565 = ~n25771 & ~n26564;
  assign n26566 = n24908 & ~n26565;
  assign n26567 = n26562 & ~n26566;
  assign n26568 = ~n26557 & ~n26567;
  assign n26569 = P1_INSTQUEUEWR_ADDR_REG_3_ & n26557;
  assign n6069 = n26568 | n26569;
  assign n26571 = n24397 & ~n26559;
  assign n26572 = n24627 & ~n24843;
  assign n26573 = ~n26571 & ~n26572;
  assign n26574 = ~n24790 & ~n24846;
  assign n26575 = n24790 & n24846;
  assign n26576 = ~n26574 & ~n26575;
  assign n26577 = n24908 & ~n26576;
  assign n26578 = n26573 & ~n26577;
  assign n26579 = ~n26557 & ~n26578;
  assign n26580 = P1_INSTQUEUEWR_ADDR_REG_2_ & n26557;
  assign n6074 = n26579 | n26580;
  assign n26582 = ~n24535 & ~n26559;
  assign n26583 = n24627 & ~n24782;
  assign n26584 = ~n26582 & ~n26583;
  assign n26585 = ~n25112 & ~n25206;
  assign n26586 = n24908 & ~n26585;
  assign n26587 = n26584 & ~n26586;
  assign n26588 = ~n26557 & ~n26587;
  assign n26589 = P1_INSTQUEUEWR_ADDR_REG_1_ & n26557;
  assign n6079 = n26588 | n26589;
  assign n26591 = ~n24520 & ~n26559;
  assign n26592 = n24626 & ~n24786;
  assign n26593 = ~n26591 & ~n26592;
  assign n26594 = ~n24610 & n26593;
  assign n26595 = ~n26557 & ~n26594;
  assign n26596 = P1_INSTQUEUEWR_ADDR_REG_0_ & n26557;
  assign n6084 = n26595 | n26596;
  assign n26598 = ~P1_STATE2_REG_2_ & n24308;
  assign n26599 = ~n24297 & n24313;
  assign n26600 = n24040 & n26599;
  assign n26601 = ~n26598 & ~n26600;
  assign n26602 = n24003 & n24190;
  assign n26603 = ~n23678 & ~n24240;
  assign n26604 = n23709 & ~n24195;
  assign n26605 = ~n23523 & ~n26604;
  assign n26606 = n24184 & n26605;
  assign n26607 = n26603 & ~n26606;
  assign n26608 = ~n24164 & ~n26607;
  assign n26609 = n24002 & n26608;
  assign n26610 = ~n23709 & ~n24558;
  assign n26611 = ~n24187 & ~n26610;
  assign n26612 = ~n23523 & n26611;
  assign n26613 = ~n24002 & n26612;
  assign n26614 = n24443 & ~n26602;
  assign n26615 = ~n26609 & n26614;
  assign n26616 = ~n26613 & n26615;
  assign n26617 = n24576 & ~n26616;
  assign n26618 = n26601 & ~n26617;
  assign n26619 = P1_STATE2_REG_2_ & ~n26618;
  assign n26620 = n24168 & n26619;
  assign n26621 = ~P1_INSTADDRPOINTER_REG_0_ & n26620;
  assign n26622 = n24054 & n24716;
  assign n26623 = n23678 & ~n23741;
  assign n26624 = n24136 & ~n24786;
  assign n26625 = ~n26622 & ~n26623;
  assign n26626 = ~n26624 & n26625;
  assign n26627 = ~P1_INSTADDRPOINTER_REG_0_ & ~n26626;
  assign n26628 = P1_INSTADDRPOINTER_REG_0_ & n26626;
  assign n26629 = ~n26627 & ~n26628;
  assign n26630 = n24014 & n24167;
  assign n26631 = P1_STATE2_REG_2_ & ~n23709;
  assign n26632 = ~n23678 & n26631;
  assign n26633 = n24184 & n26632;
  assign n26634 = ~n26630 & ~n26633;
  assign n26635 = n24015 & n24054;
  assign n26636 = ~n24004 & ~n24170;
  assign n26637 = ~n24291 & n26636;
  assign n26638 = n26634 & ~n26635;
  assign n26639 = n26637 & n26638;
  assign n26640 = P1_STATE2_REG_2_ & ~n26639;
  assign n26641 = ~n26618 & n26640;
  assign n26642 = ~n26629 & n26641;
  assign n26643 = ~n26621 & ~n26642;
  assign n26644 = n23678 & n24284;
  assign n26645 = n24258 & n24289;
  assign n26646 = ~n24220 & ~n24246;
  assign n26647 = ~n26645 & n26646;
  assign n26648 = n24400 & ~n26644;
  assign n26649 = n26647 & n26648;
  assign n26650 = n24417 & n26649;
  assign n26651 = n26619 & ~n26650;
  assign n26652 = ~P1_INSTADDRPOINTER_REG_0_ & n26651;
  assign n26653 = n24166 & ~n24304;
  assign n26654 = ~n24166 & n24304;
  assign n26655 = ~n26653 & ~n26654;
  assign n26656 = ~n24166 & ~n24304;
  assign n26657 = P1_EBX_REG_0_ & ~n26656;
  assign n26658 = ~n23678 & ~n24231;
  assign n26659 = P1_INSTADDRPOINTER_REG_0_ & ~n26658;
  assign n26660 = ~n26657 & ~n26659;
  assign n26661 = ~n24166 & ~n26660;
  assign n26662 = n24166 & n26660;
  assign n26663 = ~n26661 & ~n26662;
  assign n26664 = ~n26655 & n26663;
  assign n26665 = n26655 & ~n26663;
  assign n26666 = ~n26664 & ~n26665;
  assign n26667 = n24054 & n24184;
  assign n26668 = ~n24321 & ~n26667;
  assign n26669 = n26619 & ~n26668;
  assign n26670 = ~n26666 & n26669;
  assign n26671 = ~n26652 & ~n26670;
  assign n26672 = ~P1_STATE2_REG_2_ & ~n26618;
  assign n26673 = P1_REIP_REG_0_ & n26672;
  assign n26674 = P1_INSTADDRPOINTER_REG_0_ & n26618;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = n24011 & n26619;
  assign n26677 = P1_INSTADDRPOINTER_REG_0_ & n26676;
  assign n26678 = n26675 & ~n26677;
  assign n26679 = n26643 & n26671;
  assign n6089 = ~n26678 | ~n26679;
  assign n26681 = ~n24210 & n26620;
  assign n26682 = ~n23678 & n23896;
  assign n26683 = n24002 & ~n26682;
  assign n26684 = ~n23741 & n26683;
  assign n26685 = ~n24716 & n24765;
  assign n26686 = n24716 & ~n24765;
  assign n26687 = ~n26685 & ~n26686;
  assign n26688 = n24054 & ~n26687;
  assign n26689 = n24136 & ~n24782;
  assign n26690 = n26684 & ~n26688;
  assign n26691 = ~n26689 & n26690;
  assign n26692 = P1_INSTADDRPOINTER_REG_0_ & ~n26626;
  assign n26693 = ~n26691 & n26692;
  assign n26694 = P1_INSTADDRPOINTER_REG_1_ & n26693;
  assign n26695 = ~n26691 & ~n26692;
  assign n26696 = ~P1_INSTADDRPOINTER_REG_1_ & n26695;
  assign n26697 = ~n26694 & ~n26696;
  assign n26698 = ~P1_INSTADDRPOINTER_REG_1_ & n26692;
  assign n26699 = P1_INSTADDRPOINTER_REG_1_ & ~n26692;
  assign n26700 = ~n26698 & ~n26699;
  assign n26701 = n26691 & ~n26700;
  assign n26702 = n26697 & ~n26701;
  assign n26703 = n26641 & ~n26702;
  assign n26704 = ~n26681 & ~n26703;
  assign n26705 = ~n24210 & n26651;
  assign n26706 = n24166 & n24304;
  assign n26707 = ~n26656 & ~n26663;
  assign n26708 = ~n26706 & ~n26707;
  assign n26709 = P1_EBX_REG_1_ & ~n26656;
  assign n26710 = P1_INSTADDRPOINTER_REG_1_ & ~n26658;
  assign n26711 = ~n26709 & ~n26710;
  assign n26712 = ~n24166 & ~n26711;
  assign n26713 = n24166 & n26711;
  assign n26714 = ~n26712 & ~n26713;
  assign n26715 = n26658 & ~n26714;
  assign n26716 = ~n26658 & n26714;
  assign n26717 = ~n26715 & ~n26716;
  assign n26718 = n26708 & ~n26717;
  assign n26719 = ~n26708 & n26717;
  assign n26720 = ~n26718 & ~n26719;
  assign n26721 = n26669 & ~n26720;
  assign n26722 = ~n26705 & ~n26721;
  assign n26723 = P1_REIP_REG_1_ & n26672;
  assign n26724 = P1_INSTADDRPOINTER_REG_1_ & n26618;
  assign n26725 = ~n26723 & ~n26724;
  assign n26726 = ~P1_INSTADDRPOINTER_REG_1_ & n26676;
  assign n26727 = n26725 & ~n26726;
  assign n26728 = n26704 & n26722;
  assign n6094 = ~n26727 | ~n26728;
  assign n26730 = P1_INSTADDRPOINTER_REG_0_ & P1_INSTADDRPOINTER_REG_1_;
  assign n26731 = ~P1_INSTADDRPOINTER_REG_2_ & ~n26730;
  assign n26732 = P1_INSTADDRPOINTER_REG_2_ & n26730;
  assign n26733 = ~n26731 & ~n26732;
  assign n26734 = n26620 & ~n26733;
  assign n26735 = n26691 & ~n26692;
  assign n26736 = P1_INSTADDRPOINTER_REG_1_ & ~n26735;
  assign n26737 = ~n26693 & ~n26736;
  assign n26738 = ~n24716 & ~n24765;
  assign n26739 = n24823 & ~n26738;
  assign n26740 = ~n24823 & n26738;
  assign n26741 = ~n26739 & ~n26740;
  assign n26742 = n24054 & ~n26741;
  assign n26743 = n24136 & ~n24843;
  assign n26744 = ~n26623 & ~n26742;
  assign n26745 = ~n26743 & n26744;
  assign n26746 = P1_INSTADDRPOINTER_REG_2_ & n26745;
  assign n26747 = ~P1_INSTADDRPOINTER_REG_2_ & ~n26745;
  assign n26748 = ~n26746 & ~n26747;
  assign n26749 = n26737 & ~n26748;
  assign n26750 = ~n26737 & n26748;
  assign n26751 = ~n26749 & ~n26750;
  assign n26752 = n26641 & ~n26751;
  assign n26753 = ~n26734 & ~n26752;
  assign n26754 = ~P1_INSTADDRPOINTER_REG_2_ & n26730;
  assign n26755 = P1_INSTADDRPOINTER_REG_2_ & ~n26730;
  assign n26756 = ~n26754 & ~n26755;
  assign n26757 = n26651 & ~n26756;
  assign n26758 = P1_EBX_REG_2_ & ~n26656;
  assign n26759 = P1_INSTADDRPOINTER_REG_2_ & ~n26658;
  assign n26760 = ~n26758 & ~n26759;
  assign n26761 = ~n24166 & ~n26760;
  assign n26762 = n24166 & n26760;
  assign n26763 = ~n26761 & ~n26762;
  assign n26764 = ~n26658 & ~n26714;
  assign n26765 = n26658 & n26714;
  assign n26766 = ~n26708 & ~n26765;
  assign n26767 = ~n26764 & ~n26766;
  assign n26768 = ~n26763 & ~n26767;
  assign n26769 = n26763 & n26767;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = n26669 & n26770;
  assign n26772 = ~n26757 & ~n26771;
  assign n26773 = P1_REIP_REG_2_ & n26672;
  assign n26774 = P1_INSTADDRPOINTER_REG_2_ & n26618;
  assign n26775 = ~n26773 & ~n26774;
  assign n26776 = P1_INSTADDRPOINTER_REG_1_ & ~P1_INSTADDRPOINTER_REG_2_;
  assign n26777 = ~P1_INSTADDRPOINTER_REG_1_ & P1_INSTADDRPOINTER_REG_2_;
  assign n26778 = ~n26776 & ~n26777;
  assign n26779 = n26676 & ~n26778;
  assign n26780 = n26775 & ~n26779;
  assign n26781 = n26753 & n26772;
  assign n6099 = ~n26780 | ~n26781;
  assign n26783 = P1_INSTADDRPOINTER_REG_0_ & P1_INSTADDRPOINTER_REG_2_;
  assign n26784 = P1_INSTADDRPOINTER_REG_1_ & n26783;
  assign n26785 = P1_INSTADDRPOINTER_REG_3_ & ~n26784;
  assign n26786 = ~P1_INSTADDRPOINTER_REG_3_ & n26784;
  assign n26787 = ~n26785 & ~n26786;
  assign n26788 = n26651 & ~n26787;
  assign n26789 = P1_EBX_REG_3_ & ~n26656;
  assign n26790 = P1_INSTADDRPOINTER_REG_3_ & ~n26658;
  assign n26791 = ~n26789 & ~n26790;
  assign n26792 = ~n24166 & ~n26791;
  assign n26793 = n24166 & n26791;
  assign n26794 = ~n26792 & ~n26793;
  assign n26795 = ~n26768 & ~n26794;
  assign n26796 = n26768 & n26794;
  assign n26797 = ~n26795 & ~n26796;
  assign n26798 = n26669 & ~n26797;
  assign n26799 = ~P1_INSTADDRPOINTER_REG_3_ & n26731;
  assign n26800 = P1_INSTADDRPOINTER_REG_3_ & ~n26731;
  assign n26801 = ~n26799 & ~n26800;
  assign n26802 = n26620 & n26801;
  assign n26803 = ~n26788 & ~n26798;
  assign n26804 = ~n26802 & n26803;
  assign n26805 = P1_REIP_REG_3_ & n26672;
  assign n26806 = P1_INSTADDRPOINTER_REG_3_ & n26618;
  assign n26807 = ~n26805 & ~n26806;
  assign n26808 = P1_INSTADDRPOINTER_REG_1_ & P1_INSTADDRPOINTER_REG_2_;
  assign n26809 = ~P1_INSTADDRPOINTER_REG_3_ & n26808;
  assign n26810 = P1_INSTADDRPOINTER_REG_3_ & ~n26808;
  assign n26811 = ~n26809 & ~n26810;
  assign n26812 = n26676 & ~n26811;
  assign n26813 = P1_INSTADDRPOINTER_REG_2_ & ~n26745;
  assign n26814 = ~P1_INSTADDRPOINTER_REG_2_ & n26745;
  assign n26815 = ~n26737 & ~n26814;
  assign n26816 = ~n26813 & ~n26815;
  assign n26817 = n24879 & n26739;
  assign n26818 = ~n24879 & ~n26739;
  assign n26819 = ~n26817 & ~n26818;
  assign n26820 = n24054 & n26819;
  assign n26821 = n24136 & n24896;
  assign n26822 = ~n26820 & ~n26821;
  assign n26823 = P1_INSTADDRPOINTER_REG_3_ & n26822;
  assign n26824 = ~P1_INSTADDRPOINTER_REG_3_ & ~n26822;
  assign n26825 = ~n26823 & ~n26824;
  assign n26826 = n26816 & ~n26825;
  assign n26827 = ~n26816 & n26825;
  assign n26828 = ~n26826 & ~n26827;
  assign n26829 = n26641 & ~n26828;
  assign n26830 = n26807 & ~n26812;
  assign n26831 = ~n26829 & n26830;
  assign n6104 = ~n26804 | ~n26831;
  assign n26833 = P1_INSTADDRPOINTER_REG_3_ & n26784;
  assign n26834 = ~P1_INSTADDRPOINTER_REG_4_ & n26833;
  assign n26835 = P1_INSTADDRPOINTER_REG_4_ & ~n26833;
  assign n26836 = ~n26834 & ~n26835;
  assign n26837 = n26651 & ~n26836;
  assign n26838 = P1_EBX_REG_4_ & ~n26656;
  assign n26839 = P1_INSTADDRPOINTER_REG_4_ & ~n26658;
  assign n26840 = ~n26838 & ~n26839;
  assign n26841 = ~n24166 & ~n26840;
  assign n26842 = n24166 & n26840;
  assign n26843 = ~n26841 & ~n26842;
  assign n26844 = ~n26763 & ~n26794;
  assign n26845 = ~n26767 & n26844;
  assign n26846 = ~n26843 & ~n26845;
  assign n26847 = n26843 & n26845;
  assign n26848 = ~n26846 & ~n26847;
  assign n26849 = n26669 & ~n26848;
  assign n26850 = ~P1_INSTADDRPOINTER_REG_4_ & n26800;
  assign n26851 = P1_INSTADDRPOINTER_REG_4_ & ~n26800;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = n26620 & ~n26852;
  assign n26854 = ~n26837 & ~n26849;
  assign n26855 = ~n26853 & n26854;
  assign n26856 = P1_REIP_REG_4_ & n26672;
  assign n26857 = P1_INSTADDRPOINTER_REG_4_ & n26618;
  assign n26858 = ~n26856 & ~n26857;
  assign n26859 = P1_INSTADDRPOINTER_REG_3_ & n26808;
  assign n26860 = ~P1_INSTADDRPOINTER_REG_4_ & n26859;
  assign n26861 = P1_INSTADDRPOINTER_REG_4_ & ~n26859;
  assign n26862 = ~n26860 & ~n26861;
  assign n26863 = n26676 & ~n26862;
  assign n26864 = n26858 & ~n26863;
  assign n26865 = P1_INSTADDRPOINTER_REG_3_ & ~n26822;
  assign n26866 = ~P1_INSTADDRPOINTER_REG_3_ & n26822;
  assign n26867 = ~n26816 & ~n26866;
  assign n26868 = ~n26865 & ~n26867;
  assign n26869 = P1_INSTQUEUE_REG_0__4_ & n24630;
  assign n26870 = P1_INSTQUEUE_REG_1__4_ & n24633;
  assign n26871 = P1_INSTQUEUE_REG_2__4_ & n24636;
  assign n26872 = P1_INSTQUEUE_REG_3__4_ & n24639;
  assign n26873 = ~n26869 & ~n26870;
  assign n26874 = ~n26871 & n26873;
  assign n26875 = ~n26872 & n26874;
  assign n26876 = P1_INSTQUEUE_REG_4__4_ & n24645;
  assign n26877 = P1_INSTQUEUE_REG_5__4_ & n24647;
  assign n26878 = P1_INSTQUEUE_REG_6__4_ & n24649;
  assign n26879 = P1_INSTQUEUE_REG_7__4_ & n24651;
  assign n26880 = ~n26876 & ~n26877;
  assign n26881 = ~n26878 & n26880;
  assign n26882 = ~n26879 & n26881;
  assign n26883 = P1_INSTQUEUE_REG_8__4_ & n24657;
  assign n26884 = P1_INSTQUEUE_REG_9__4_ & n24659;
  assign n26885 = P1_INSTQUEUE_REG_10__4_ & n24661;
  assign n26886 = P1_INSTQUEUE_REG_11__4_ & n24663;
  assign n26887 = ~n26883 & ~n26884;
  assign n26888 = ~n26885 & n26887;
  assign n26889 = ~n26886 & n26888;
  assign n26890 = P1_INSTQUEUE_REG_12__4_ & n24669;
  assign n26891 = P1_INSTQUEUE_REG_13__4_ & n24671;
  assign n26892 = P1_INSTQUEUE_REG_14__4_ & n24673;
  assign n26893 = P1_INSTQUEUE_REG_15__4_ & n24675;
  assign n26894 = ~n26890 & ~n26891;
  assign n26895 = ~n26892 & n26894;
  assign n26896 = ~n26893 & n26895;
  assign n26897 = n26875 & n26882;
  assign n26898 = n26889 & n26897;
  assign n26899 = n26896 & n26898;
  assign n26900 = n26818 & n26899;
  assign n26901 = ~n26818 & ~n26899;
  assign n26902 = ~n26900 & ~n26901;
  assign n26903 = n24054 & ~n26902;
  assign n26904 = P1_INSTQUEUE_REG_0__4_ & n24040;
  assign n26905 = n24045 & ~n26899;
  assign n26906 = ~n26904 & ~n26905;
  assign n26907 = n24683 & n26899;
  assign n26908 = n24685 & ~n26899;
  assign n26909 = ~n26907 & ~n26908;
  assign n26910 = ~n24683 & ~n26909;
  assign n26911 = n24683 & n26909;
  assign n26912 = ~n26910 & ~n26911;
  assign n26913 = ~n26906 & ~n26912;
  assign n26914 = n26906 & n26912;
  assign n26915 = ~n26913 & ~n26914;
  assign n26916 = ~n24835 & ~n24891;
  assign n26917 = n24733 & ~n24837;
  assign n26918 = ~n24838 & ~n26917;
  assign n26919 = ~n24834 & ~n26918;
  assign n26920 = n26916 & ~n26919;
  assign n26921 = ~n24890 & ~n26920;
  assign n26922 = n26915 & n26921;
  assign n26923 = ~n26915 & ~n26921;
  assign n26924 = ~n26922 & ~n26923;
  assign n26925 = n24136 & ~n26924;
  assign n26926 = ~n26903 & ~n26925;
  assign n26927 = P1_INSTADDRPOINTER_REG_4_ & n26926;
  assign n26928 = ~P1_INSTADDRPOINTER_REG_4_ & ~n26926;
  assign n26929 = ~n26927 & ~n26928;
  assign n26930 = n26868 & ~n26929;
  assign n26931 = ~n26868 & n26929;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = n26641 & ~n26932;
  assign n26934 = n26855 & n26864;
  assign n6109 = n26933 | ~n26934;
  assign n26936 = P1_INSTADDRPOINTER_REG_3_ & P1_INSTADDRPOINTER_REG_4_;
  assign n26937 = n26784 & n26936;
  assign n26938 = P1_INSTADDRPOINTER_REG_5_ & ~n26937;
  assign n26939 = ~P1_INSTADDRPOINTER_REG_5_ & n26937;
  assign n26940 = ~n26938 & ~n26939;
  assign n26941 = n26651 & ~n26940;
  assign n26942 = P1_EBX_REG_5_ & ~n26656;
  assign n26943 = P1_INSTADDRPOINTER_REG_5_ & ~n26658;
  assign n26944 = ~n26942 & ~n26943;
  assign n26945 = ~n24166 & ~n26944;
  assign n26946 = n24166 & n26944;
  assign n26947 = ~n26945 & ~n26946;
  assign n26948 = ~n26843 & n26845;
  assign n26949 = ~n26947 & ~n26948;
  assign n26950 = n26947 & n26948;
  assign n26951 = ~n26949 & ~n26950;
  assign n26952 = n26669 & ~n26951;
  assign n26953 = P1_INSTADDRPOINTER_REG_4_ & n26800;
  assign n26954 = ~P1_INSTADDRPOINTER_REG_5_ & n26953;
  assign n26955 = P1_INSTADDRPOINTER_REG_5_ & ~n26953;
  assign n26956 = ~n26954 & ~n26955;
  assign n26957 = n26620 & ~n26956;
  assign n26958 = ~n26941 & ~n26952;
  assign n26959 = ~n26957 & n26958;
  assign n26960 = P1_REIP_REG_5_ & n26672;
  assign n26961 = P1_INSTADDRPOINTER_REG_5_ & n26618;
  assign n26962 = ~n26960 & ~n26961;
  assign n26963 = P1_INSTADDRPOINTER_REG_4_ & n26859;
  assign n26964 = ~P1_INSTADDRPOINTER_REG_5_ & n26963;
  assign n26965 = P1_INSTADDRPOINTER_REG_5_ & ~n26963;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = n26676 & ~n26966;
  assign n26968 = n26962 & ~n26967;
  assign n26969 = P1_INSTADDRPOINTER_REG_4_ & ~n26926;
  assign n26970 = ~P1_INSTADDRPOINTER_REG_4_ & n26926;
  assign n26971 = ~n26868 & ~n26970;
  assign n26972 = ~n26969 & ~n26971;
  assign n26973 = n26818 & ~n26899;
  assign n26974 = P1_INSTQUEUE_REG_0__5_ & n24630;
  assign n26975 = P1_INSTQUEUE_REG_1__5_ & n24633;
  assign n26976 = P1_INSTQUEUE_REG_2__5_ & n24636;
  assign n26977 = P1_INSTQUEUE_REG_3__5_ & n24639;
  assign n26978 = ~n26974 & ~n26975;
  assign n26979 = ~n26976 & n26978;
  assign n26980 = ~n26977 & n26979;
  assign n26981 = P1_INSTQUEUE_REG_4__5_ & n24645;
  assign n26982 = P1_INSTQUEUE_REG_5__5_ & n24647;
  assign n26983 = P1_INSTQUEUE_REG_6__5_ & n24649;
  assign n26984 = P1_INSTQUEUE_REG_7__5_ & n24651;
  assign n26985 = ~n26981 & ~n26982;
  assign n26986 = ~n26983 & n26985;
  assign n26987 = ~n26984 & n26986;
  assign n26988 = P1_INSTQUEUE_REG_8__5_ & n24657;
  assign n26989 = P1_INSTQUEUE_REG_9__5_ & n24659;
  assign n26990 = P1_INSTQUEUE_REG_10__5_ & n24661;
  assign n26991 = P1_INSTQUEUE_REG_11__5_ & n24663;
  assign n26992 = ~n26988 & ~n26989;
  assign n26993 = ~n26990 & n26992;
  assign n26994 = ~n26991 & n26993;
  assign n26995 = P1_INSTQUEUE_REG_12__5_ & n24669;
  assign n26996 = P1_INSTQUEUE_REG_13__5_ & n24671;
  assign n26997 = P1_INSTQUEUE_REG_14__5_ & n24673;
  assign n26998 = P1_INSTQUEUE_REG_15__5_ & n24675;
  assign n26999 = ~n26995 & ~n26996;
  assign n27000 = ~n26997 & n26999;
  assign n27001 = ~n26998 & n27000;
  assign n27002 = n26980 & n26987;
  assign n27003 = n26994 & n27002;
  assign n27004 = n27001 & n27003;
  assign n27005 = n26973 & n27004;
  assign n27006 = ~n26973 & ~n27004;
  assign n27007 = ~n27005 & ~n27006;
  assign n27008 = n24054 & ~n27007;
  assign n27009 = P1_INSTQUEUE_REG_0__5_ & n24040;
  assign n27010 = n24045 & ~n27004;
  assign n27011 = ~n27009 & ~n27010;
  assign n27012 = n24683 & n27004;
  assign n27013 = n24685 & ~n27004;
  assign n27014 = ~n27012 & ~n27013;
  assign n27015 = ~n24683 & ~n27014;
  assign n27016 = n24683 & n27014;
  assign n27017 = ~n27015 & ~n27016;
  assign n27018 = ~n27011 & ~n27017;
  assign n27019 = n27011 & n27017;
  assign n27020 = ~n27018 & ~n27019;
  assign n27021 = ~n24881 & ~n26914;
  assign n27022 = ~n24889 & n27021;
  assign n27023 = ~n26913 & ~n27022;
  assign n27024 = ~n24835 & ~n26914;
  assign n27025 = ~n24891 & ~n26919;
  assign n27026 = n27024 & n27025;
  assign n27027 = n27023 & ~n27026;
  assign n27028 = n27020 & n27027;
  assign n27029 = ~n27020 & ~n27027;
  assign n27030 = ~n27028 & ~n27029;
  assign n27031 = n24136 & ~n27030;
  assign n27032 = ~n27008 & ~n27031;
  assign n27033 = ~P1_INSTADDRPOINTER_REG_5_ & n27032;
  assign n27034 = ~n26972 & ~n27033;
  assign n27035 = P1_INSTADDRPOINTER_REG_5_ & ~n27032;
  assign n27036 = n27034 & ~n27035;
  assign n27037 = P1_INSTADDRPOINTER_REG_5_ & n27032;
  assign n27038 = ~P1_INSTADDRPOINTER_REG_5_ & ~n27032;
  assign n27039 = ~n27037 & ~n27038;
  assign n27040 = n26972 & n27039;
  assign n27041 = ~n27036 & ~n27040;
  assign n27042 = n26641 & n27041;
  assign n27043 = n26959 & n26968;
  assign n6114 = n27042 | ~n27043;
  assign n27045 = P1_INSTADDRPOINTER_REG_5_ & n26937;
  assign n27046 = ~P1_INSTADDRPOINTER_REG_6_ & n27045;
  assign n27047 = P1_INSTADDRPOINTER_REG_6_ & ~n27045;
  assign n27048 = ~n27046 & ~n27047;
  assign n27049 = n26651 & ~n27048;
  assign n27050 = P1_EBX_REG_6_ & ~n26656;
  assign n27051 = P1_INSTADDRPOINTER_REG_6_ & ~n26658;
  assign n27052 = ~n27050 & ~n27051;
  assign n27053 = ~n24166 & ~n27052;
  assign n27054 = n24166 & n27052;
  assign n27055 = ~n27053 & ~n27054;
  assign n27056 = ~n26843 & ~n26947;
  assign n27057 = n26845 & n27056;
  assign n27058 = ~n27055 & ~n27057;
  assign n27059 = n27055 & n27057;
  assign n27060 = ~n27058 & ~n27059;
  assign n27061 = n26669 & ~n27060;
  assign n27062 = P1_INSTADDRPOINTER_REG_5_ & n26953;
  assign n27063 = ~P1_INSTADDRPOINTER_REG_6_ & n27062;
  assign n27064 = P1_INSTADDRPOINTER_REG_6_ & ~n27062;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = n26620 & ~n27065;
  assign n27067 = ~n27049 & ~n27061;
  assign n27068 = ~n27066 & n27067;
  assign n27069 = P1_REIP_REG_6_ & n26672;
  assign n27070 = P1_INSTADDRPOINTER_REG_6_ & n26618;
  assign n27071 = ~n27069 & ~n27070;
  assign n27072 = P1_INSTADDRPOINTER_REG_5_ & n26963;
  assign n27073 = ~P1_INSTADDRPOINTER_REG_6_ & n27072;
  assign n27074 = P1_INSTADDRPOINTER_REG_6_ & ~n27072;
  assign n27075 = ~n27073 & ~n27074;
  assign n27076 = n26676 & ~n27075;
  assign n27077 = n27071 & ~n27076;
  assign n27078 = n26973 & ~n27004;
  assign n27079 = P1_INSTQUEUE_REG_0__6_ & n24630;
  assign n27080 = P1_INSTQUEUE_REG_1__6_ & n24633;
  assign n27081 = P1_INSTQUEUE_REG_2__6_ & n24636;
  assign n27082 = P1_INSTQUEUE_REG_3__6_ & n24639;
  assign n27083 = ~n27079 & ~n27080;
  assign n27084 = ~n27081 & n27083;
  assign n27085 = ~n27082 & n27084;
  assign n27086 = P1_INSTQUEUE_REG_4__6_ & n24645;
  assign n27087 = P1_INSTQUEUE_REG_5__6_ & n24647;
  assign n27088 = P1_INSTQUEUE_REG_6__6_ & n24649;
  assign n27089 = P1_INSTQUEUE_REG_7__6_ & n24651;
  assign n27090 = ~n27086 & ~n27087;
  assign n27091 = ~n27088 & n27090;
  assign n27092 = ~n27089 & n27091;
  assign n27093 = P1_INSTQUEUE_REG_8__6_ & n24657;
  assign n27094 = P1_INSTQUEUE_REG_9__6_ & n24659;
  assign n27095 = P1_INSTQUEUE_REG_10__6_ & n24661;
  assign n27096 = P1_INSTQUEUE_REG_11__6_ & n24663;
  assign n27097 = ~n27093 & ~n27094;
  assign n27098 = ~n27095 & n27097;
  assign n27099 = ~n27096 & n27098;
  assign n27100 = P1_INSTQUEUE_REG_12__6_ & n24669;
  assign n27101 = P1_INSTQUEUE_REG_13__6_ & n24671;
  assign n27102 = P1_INSTQUEUE_REG_14__6_ & n24673;
  assign n27103 = P1_INSTQUEUE_REG_15__6_ & n24675;
  assign n27104 = ~n27100 & ~n27101;
  assign n27105 = ~n27102 & n27104;
  assign n27106 = ~n27103 & n27105;
  assign n27107 = n27085 & n27092;
  assign n27108 = n27099 & n27107;
  assign n27109 = n27106 & n27108;
  assign n27110 = n27078 & n27109;
  assign n27111 = ~n27078 & ~n27109;
  assign n27112 = ~n27110 & ~n27111;
  assign n27113 = n24054 & ~n27112;
  assign n27114 = P1_INSTQUEUE_REG_0__6_ & n24040;
  assign n27115 = n24045 & ~n27109;
  assign n27116 = ~n27114 & ~n27115;
  assign n27117 = n24683 & n27109;
  assign n27118 = n24685 & ~n27109;
  assign n27119 = ~n27117 & ~n27118;
  assign n27120 = ~n24683 & ~n27119;
  assign n27121 = n24683 & n27119;
  assign n27122 = ~n27120 & ~n27121;
  assign n27123 = ~n27116 & ~n27122;
  assign n27124 = n27116 & n27122;
  assign n27125 = ~n27123 & ~n27124;
  assign n27126 = ~n27019 & ~n27027;
  assign n27127 = ~n27018 & ~n27126;
  assign n27128 = n27125 & ~n27127;
  assign n27129 = ~n27018 & ~n27125;
  assign n27130 = ~n27126 & n27129;
  assign n27131 = ~n27128 & ~n27130;
  assign n27132 = n24136 & n27131;
  assign n27133 = ~n27113 & ~n27132;
  assign n27134 = P1_INSTADDRPOINTER_REG_6_ & n27133;
  assign n27135 = ~P1_INSTADDRPOINTER_REG_6_ & ~n27133;
  assign n27136 = ~n27134 & ~n27135;
  assign n27137 = ~n27034 & ~n27035;
  assign n27138 = ~n27136 & n27137;
  assign n27139 = ~P1_INSTADDRPOINTER_REG_6_ & n27133;
  assign n27140 = P1_INSTADDRPOINTER_REG_6_ & ~n27133;
  assign n27141 = ~n27139 & ~n27140;
  assign n27142 = ~n27137 & ~n27141;
  assign n27143 = ~n27138 & ~n27142;
  assign n27144 = n26641 & ~n27143;
  assign n27145 = n27068 & n27077;
  assign n6119 = n27144 | ~n27145;
  assign n27147 = P1_INSTADDRPOINTER_REG_5_ & P1_INSTADDRPOINTER_REG_6_;
  assign n27148 = n26937 & n27147;
  assign n27149 = P1_INSTADDRPOINTER_REG_7_ & ~n27148;
  assign n27150 = ~P1_INSTADDRPOINTER_REG_7_ & n27148;
  assign n27151 = ~n27149 & ~n27150;
  assign n27152 = n26651 & ~n27151;
  assign n27153 = P1_EBX_REG_7_ & ~n26656;
  assign n27154 = P1_INSTADDRPOINTER_REG_7_ & ~n26658;
  assign n27155 = ~n27153 & ~n27154;
  assign n27156 = ~n24166 & ~n27155;
  assign n27157 = n24166 & n27155;
  assign n27158 = ~n27156 & ~n27157;
  assign n27159 = ~n27055 & n27057;
  assign n27160 = ~n27158 & ~n27159;
  assign n27161 = n27158 & n27159;
  assign n27162 = ~n27160 & ~n27161;
  assign n27163 = n26669 & ~n27162;
  assign n27164 = P1_INSTADDRPOINTER_REG_6_ & n27062;
  assign n27165 = ~P1_INSTADDRPOINTER_REG_7_ & n27164;
  assign n27166 = P1_INSTADDRPOINTER_REG_7_ & ~n27164;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = n26620 & ~n27167;
  assign n27169 = ~n27152 & ~n27163;
  assign n27170 = ~n27168 & n27169;
  assign n27171 = P1_REIP_REG_7_ & n26672;
  assign n27172 = P1_INSTADDRPOINTER_REG_7_ & n26618;
  assign n27173 = ~n27171 & ~n27172;
  assign n27174 = P1_INSTADDRPOINTER_REG_6_ & n27072;
  assign n27175 = ~P1_INSTADDRPOINTER_REG_7_ & n27174;
  assign n27176 = P1_INSTADDRPOINTER_REG_7_ & ~n27174;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = n26676 & ~n27177;
  assign n27179 = n27173 & ~n27178;
  assign n27180 = n27137 & ~n27140;
  assign n27181 = n27078 & ~n27109;
  assign n27182 = n24682 & n27181;
  assign n27183 = ~n24682 & ~n27181;
  assign n27184 = ~n27182 & ~n27183;
  assign n27185 = n24054 & ~n27184;
  assign n27186 = n24682 & n24683;
  assign n27187 = ~n24682 & n24685;
  assign n27188 = ~n27186 & ~n27187;
  assign n27189 = ~n24683 & ~n27188;
  assign n27190 = n24683 & n27188;
  assign n27191 = P1_INSTQUEUE_REG_0__7_ & n24040;
  assign n27192 = n24045 & ~n24682;
  assign n27193 = ~n27191 & ~n27192;
  assign n27194 = ~n27189 & ~n27190;
  assign n27195 = n27193 & n27194;
  assign n27196 = ~n27193 & ~n27194;
  assign n27197 = ~n27195 & ~n27196;
  assign n27198 = n27123 & n27197;
  assign n27199 = ~n27018 & ~n27197;
  assign n27200 = ~n27126 & n27199;
  assign n27201 = ~n27123 & n27200;
  assign n27202 = ~n27019 & n27197;
  assign n27203 = ~n26913 & ~n27018;
  assign n27204 = ~n27022 & n27203;
  assign n27205 = ~n27026 & n27204;
  assign n27206 = n27202 & ~n27205;
  assign n27207 = ~n27124 & n27206;
  assign n27208 = n27124 & ~n27197;
  assign n27209 = ~n27207 & ~n27208;
  assign n27210 = ~n27198 & ~n27201;
  assign n27211 = n27209 & n27210;
  assign n27212 = n24136 & n27211;
  assign n27213 = ~n27185 & ~n27212;
  assign n27214 = ~P1_INSTADDRPOINTER_REG_7_ & n27213;
  assign n27215 = ~n27139 & ~n27180;
  assign n27216 = ~n27214 & n27215;
  assign n27217 = P1_INSTADDRPOINTER_REG_7_ & ~n27213;
  assign n27218 = n27216 & ~n27217;
  assign n27219 = ~n27137 & ~n27139;
  assign n27220 = P1_INSTADDRPOINTER_REG_7_ & n27213;
  assign n27221 = ~P1_INSTADDRPOINTER_REG_7_ & ~n27213;
  assign n27222 = ~n27220 & ~n27221;
  assign n27223 = ~n27140 & ~n27219;
  assign n27224 = n27222 & n27223;
  assign n27225 = ~n27218 & ~n27224;
  assign n27226 = n26641 & n27225;
  assign n27227 = n27170 & n27179;
  assign n6124 = n27226 | ~n27227;
  assign n27229 = P1_INSTADDRPOINTER_REG_7_ & n27148;
  assign n27230 = ~P1_INSTADDRPOINTER_REG_8_ & n27229;
  assign n27231 = P1_INSTADDRPOINTER_REG_8_ & ~n27229;
  assign n27232 = ~n27230 & ~n27231;
  assign n27233 = n26651 & ~n27232;
  assign n27234 = P1_EBX_REG_8_ & ~n26656;
  assign n27235 = P1_INSTADDRPOINTER_REG_8_ & ~n26658;
  assign n27236 = ~n27234 & ~n27235;
  assign n27237 = ~n24166 & ~n27236;
  assign n27238 = n24166 & n27236;
  assign n27239 = ~n27237 & ~n27238;
  assign n27240 = ~n27055 & ~n27158;
  assign n27241 = n27057 & n27240;
  assign n27242 = ~n27239 & ~n27241;
  assign n27243 = n27239 & n27241;
  assign n27244 = ~n27242 & ~n27243;
  assign n27245 = n26669 & ~n27244;
  assign n27246 = P1_INSTADDRPOINTER_REG_7_ & n27164;
  assign n27247 = ~P1_INSTADDRPOINTER_REG_8_ & n27246;
  assign n27248 = P1_INSTADDRPOINTER_REG_8_ & ~n27246;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = n26620 & ~n27249;
  assign n27251 = ~n27233 & ~n27245;
  assign n27252 = ~n27250 & n27251;
  assign n27253 = P1_REIP_REG_8_ & n26672;
  assign n27254 = P1_INSTADDRPOINTER_REG_8_ & n26618;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = P1_INSTADDRPOINTER_REG_7_ & n27174;
  assign n27257 = ~P1_INSTADDRPOINTER_REG_8_ & n27256;
  assign n27258 = P1_INSTADDRPOINTER_REG_8_ & ~n27256;
  assign n27259 = ~n27257 & ~n27258;
  assign n27260 = n26676 & ~n27259;
  assign n27261 = n27255 & ~n27260;
  assign n27262 = ~n27216 & ~n27217;
  assign n27263 = ~n24682 & ~n27109;
  assign n27264 = n27078 & n27263;
  assign n27265 = n24054 & n27264;
  assign n27266 = n24226 & n24485;
  assign n27267 = n23662 & n27266;
  assign n27268 = P1_INSTQUEUE_REG_0__0_ & n27267;
  assign n27269 = n23655 & n27266;
  assign n27270 = P1_INSTQUEUE_REG_1__0_ & n27269;
  assign n27271 = n23624 & n27266;
  assign n27272 = P1_INSTQUEUE_REG_2__0_ & n27271;
  assign n27273 = n23665 & n27266;
  assign n27274 = P1_INSTQUEUE_REG_3__0_ & n27273;
  assign n27275 = ~n27268 & ~n27270;
  assign n27276 = ~n27272 & n27275;
  assign n27277 = ~n27274 & n27276;
  assign n27278 = ~n24226 & n24485;
  assign n27279 = n23662 & n27278;
  assign n27280 = P1_INSTQUEUE_REG_4__0_ & n27279;
  assign n27281 = n23655 & n27278;
  assign n27282 = P1_INSTQUEUE_REG_5__0_ & n27281;
  assign n27283 = n23624 & n27278;
  assign n27284 = P1_INSTQUEUE_REG_6__0_ & n27283;
  assign n27285 = n23665 & n27278;
  assign n27286 = P1_INSTQUEUE_REG_7__0_ & n27285;
  assign n27287 = ~n27280 & ~n27282;
  assign n27288 = ~n27284 & n27287;
  assign n27289 = ~n27286 & n27288;
  assign n27290 = n24226 & ~n24485;
  assign n27291 = n23662 & n27290;
  assign n27292 = P1_INSTQUEUE_REG_8__0_ & n27291;
  assign n27293 = n23655 & n27290;
  assign n27294 = P1_INSTQUEUE_REG_9__0_ & n27293;
  assign n27295 = n23624 & n27290;
  assign n27296 = P1_INSTQUEUE_REG_10__0_ & n27295;
  assign n27297 = n23665 & n27290;
  assign n27298 = P1_INSTQUEUE_REG_11__0_ & n27297;
  assign n27299 = ~n27292 & ~n27294;
  assign n27300 = ~n27296 & n27299;
  assign n27301 = ~n27298 & n27300;
  assign n27302 = ~n24226 & ~n24485;
  assign n27303 = n23662 & n27302;
  assign n27304 = P1_INSTQUEUE_REG_12__0_ & n27303;
  assign n27305 = n23655 & n27302;
  assign n27306 = P1_INSTQUEUE_REG_13__0_ & n27305;
  assign n27307 = n23624 & n27302;
  assign n27308 = P1_INSTQUEUE_REG_14__0_ & n27307;
  assign n27309 = n23665 & n27302;
  assign n27310 = P1_INSTQUEUE_REG_15__0_ & n27309;
  assign n27311 = ~n27304 & ~n27306;
  assign n27312 = ~n27308 & n27311;
  assign n27313 = ~n27310 & n27312;
  assign n27314 = n27277 & n27289;
  assign n27315 = n27301 & n27314;
  assign n27316 = n27313 & n27315;
  assign n27317 = ~n24040 & ~n24045;
  assign n27318 = ~n27316 & ~n27317;
  assign n27319 = ~n24683 & n27318;
  assign n27320 = n24683 & ~n27318;
  assign n27321 = ~n27319 & ~n27320;
  assign n27322 = ~n27124 & ~n27195;
  assign n27323 = ~n26914 & ~n27019;
  assign n27324 = n27322 & n27323;
  assign n27325 = ~n26921 & n27324;
  assign n27326 = n26913 & ~n27019;
  assign n27327 = n27322 & n27326;
  assign n27328 = n27123 & n27322;
  assign n27329 = n27018 & n27322;
  assign n27330 = ~n27196 & ~n27327;
  assign n27331 = ~n27328 & n27330;
  assign n27332 = ~n27329 & n27331;
  assign n27333 = ~n27325 & n27332;
  assign n27334 = ~n27321 & ~n27333;
  assign n27335 = n27321 & n27333;
  assign n27336 = ~n27334 & ~n27335;
  assign n27337 = n24136 & n27336;
  assign n27338 = ~n27265 & ~n27337;
  assign n27339 = P1_INSTADDRPOINTER_REG_8_ & n27338;
  assign n27340 = ~P1_INSTADDRPOINTER_REG_8_ & ~n27338;
  assign n27341 = ~n27339 & ~n27340;
  assign n27342 = n27262 & ~n27341;
  assign n27343 = ~n27262 & n27341;
  assign n27344 = ~n27342 & ~n27343;
  assign n27345 = n26641 & ~n27344;
  assign n27346 = n27252 & n27261;
  assign n6129 = n27345 | ~n27346;
  assign n27348 = P1_INSTADDRPOINTER_REG_7_ & P1_INSTADDRPOINTER_REG_8_;
  assign n27349 = n27148 & n27348;
  assign n27350 = P1_INSTADDRPOINTER_REG_9_ & ~n27349;
  assign n27351 = ~P1_INSTADDRPOINTER_REG_9_ & n27349;
  assign n27352 = ~n27350 & ~n27351;
  assign n27353 = n26651 & ~n27352;
  assign n27354 = P1_EBX_REG_9_ & ~n26656;
  assign n27355 = P1_INSTADDRPOINTER_REG_9_ & ~n26658;
  assign n27356 = ~n27354 & ~n27355;
  assign n27357 = ~n24166 & ~n27356;
  assign n27358 = n24166 & n27356;
  assign n27359 = ~n27357 & ~n27358;
  assign n27360 = ~n27239 & n27241;
  assign n27361 = ~n27359 & ~n27360;
  assign n27362 = n27359 & n27360;
  assign n27363 = ~n27361 & ~n27362;
  assign n27364 = n26669 & ~n27363;
  assign n27365 = P1_INSTADDRPOINTER_REG_8_ & n27246;
  assign n27366 = ~P1_INSTADDRPOINTER_REG_9_ & n27365;
  assign n27367 = P1_INSTADDRPOINTER_REG_9_ & ~n27365;
  assign n27368 = ~n27366 & ~n27367;
  assign n27369 = n26620 & ~n27368;
  assign n27370 = ~n27353 & ~n27364;
  assign n27371 = ~n27369 & n27370;
  assign n27372 = P1_REIP_REG_9_ & n26672;
  assign n27373 = P1_INSTADDRPOINTER_REG_9_ & n26618;
  assign n27374 = ~n27372 & ~n27373;
  assign n27375 = P1_INSTADDRPOINTER_REG_8_ & n27256;
  assign n27376 = ~P1_INSTADDRPOINTER_REG_9_ & n27375;
  assign n27377 = P1_INSTADDRPOINTER_REG_9_ & ~n27375;
  assign n27378 = ~n27376 & ~n27377;
  assign n27379 = n26676 & ~n27378;
  assign n27380 = n27374 & ~n27379;
  assign n27381 = P1_INSTQUEUE_REG_0__1_ & n27267;
  assign n27382 = P1_INSTQUEUE_REG_1__1_ & n27269;
  assign n27383 = P1_INSTQUEUE_REG_2__1_ & n27271;
  assign n27384 = P1_INSTQUEUE_REG_3__1_ & n27273;
  assign n27385 = ~n27381 & ~n27382;
  assign n27386 = ~n27383 & n27385;
  assign n27387 = ~n27384 & n27386;
  assign n27388 = P1_INSTQUEUE_REG_4__1_ & n27279;
  assign n27389 = P1_INSTQUEUE_REG_5__1_ & n27281;
  assign n27390 = P1_INSTQUEUE_REG_6__1_ & n27283;
  assign n27391 = P1_INSTQUEUE_REG_7__1_ & n27285;
  assign n27392 = ~n27388 & ~n27389;
  assign n27393 = ~n27390 & n27392;
  assign n27394 = ~n27391 & n27393;
  assign n27395 = P1_INSTQUEUE_REG_8__1_ & n27291;
  assign n27396 = P1_INSTQUEUE_REG_9__1_ & n27293;
  assign n27397 = P1_INSTQUEUE_REG_10__1_ & n27295;
  assign n27398 = P1_INSTQUEUE_REG_11__1_ & n27297;
  assign n27399 = ~n27395 & ~n27396;
  assign n27400 = ~n27397 & n27399;
  assign n27401 = ~n27398 & n27400;
  assign n27402 = P1_INSTQUEUE_REG_12__1_ & n27303;
  assign n27403 = P1_INSTQUEUE_REG_13__1_ & n27305;
  assign n27404 = P1_INSTQUEUE_REG_14__1_ & n27307;
  assign n27405 = P1_INSTQUEUE_REG_15__1_ & n27309;
  assign n27406 = ~n27402 & ~n27403;
  assign n27407 = ~n27404 & n27406;
  assign n27408 = ~n27405 & n27407;
  assign n27409 = n27387 & n27394;
  assign n27410 = n27401 & n27409;
  assign n27411 = n27408 & n27410;
  assign n27412 = ~n27317 & ~n27411;
  assign n27413 = ~n24683 & n27412;
  assign n27414 = n24683 & ~n27412;
  assign n27415 = ~n27413 & ~n27414;
  assign n27416 = ~n27334 & ~n27415;
  assign n27417 = n27334 & n27415;
  assign n27418 = ~n27416 & ~n27417;
  assign n27419 = n24136 & ~n27418;
  assign n27420 = P1_INSTADDRPOINTER_REG_9_ & n27419;
  assign n27421 = ~P1_INSTADDRPOINTER_REG_9_ & ~n27419;
  assign n27422 = ~n27420 & ~n27421;
  assign n27423 = ~P1_INSTADDRPOINTER_REG_8_ & n27338;
  assign n27424 = n27217 & ~n27423;
  assign n27425 = P1_INSTADDRPOINTER_REG_8_ & ~n27338;
  assign n27426 = ~n27424 & ~n27425;
  assign n27427 = ~n27139 & ~n27423;
  assign n27428 = ~n27180 & ~n27214;
  assign n27429 = n27427 & n27428;
  assign n27430 = n27426 & ~n27429;
  assign n27431 = n27422 & n27430;
  assign n27432 = ~n27422 & ~n27430;
  assign n27433 = ~n27431 & ~n27432;
  assign n27434 = n26641 & ~n27433;
  assign n27435 = n27371 & n27380;
  assign n6134 = n27434 | ~n27435;
  assign n27437 = P1_INSTADDRPOINTER_REG_9_ & n27349;
  assign n27438 = ~P1_INSTADDRPOINTER_REG_10_ & n27437;
  assign n27439 = P1_INSTADDRPOINTER_REG_10_ & ~n27437;
  assign n27440 = ~n27438 & ~n27439;
  assign n27441 = n26651 & ~n27440;
  assign n27442 = P1_EBX_REG_10_ & ~n26656;
  assign n27443 = P1_INSTADDRPOINTER_REG_10_ & ~n26658;
  assign n27444 = ~n27442 & ~n27443;
  assign n27445 = ~n24166 & ~n27444;
  assign n27446 = n24166 & n27444;
  assign n27447 = ~n27445 & ~n27446;
  assign n27448 = ~n27239 & ~n27359;
  assign n27449 = n27241 & n27448;
  assign n27450 = ~n27447 & ~n27449;
  assign n27451 = n27447 & n27449;
  assign n27452 = ~n27450 & ~n27451;
  assign n27453 = n26669 & ~n27452;
  assign n27454 = P1_INSTADDRPOINTER_REG_9_ & n27365;
  assign n27455 = ~P1_INSTADDRPOINTER_REG_10_ & n27454;
  assign n27456 = P1_INSTADDRPOINTER_REG_10_ & ~n27454;
  assign n27457 = ~n27455 & ~n27456;
  assign n27458 = n26620 & ~n27457;
  assign n27459 = ~n27441 & ~n27453;
  assign n27460 = ~n27458 & n27459;
  assign n27461 = P1_REIP_REG_10_ & n26672;
  assign n27462 = P1_INSTADDRPOINTER_REG_10_ & n26618;
  assign n27463 = ~n27461 & ~n27462;
  assign n27464 = P1_INSTADDRPOINTER_REG_9_ & n27375;
  assign n27465 = ~P1_INSTADDRPOINTER_REG_10_ & n27464;
  assign n27466 = P1_INSTADDRPOINTER_REG_10_ & ~n27464;
  assign n27467 = ~n27465 & ~n27466;
  assign n27468 = n26676 & ~n27467;
  assign n27469 = n27463 & ~n27468;
  assign n27470 = ~n27421 & ~n27430;
  assign n27471 = ~n27420 & ~n27470;
  assign n27472 = P1_INSTQUEUE_REG_0__2_ & n27267;
  assign n27473 = P1_INSTQUEUE_REG_1__2_ & n27269;
  assign n27474 = P1_INSTQUEUE_REG_2__2_ & n27271;
  assign n27475 = P1_INSTQUEUE_REG_3__2_ & n27273;
  assign n27476 = ~n27472 & ~n27473;
  assign n27477 = ~n27474 & n27476;
  assign n27478 = ~n27475 & n27477;
  assign n27479 = P1_INSTQUEUE_REG_4__2_ & n27279;
  assign n27480 = P1_INSTQUEUE_REG_5__2_ & n27281;
  assign n27481 = P1_INSTQUEUE_REG_6__2_ & n27283;
  assign n27482 = P1_INSTQUEUE_REG_7__2_ & n27285;
  assign n27483 = ~n27479 & ~n27480;
  assign n27484 = ~n27481 & n27483;
  assign n27485 = ~n27482 & n27484;
  assign n27486 = P1_INSTQUEUE_REG_8__2_ & n27291;
  assign n27487 = P1_INSTQUEUE_REG_9__2_ & n27293;
  assign n27488 = P1_INSTQUEUE_REG_10__2_ & n27295;
  assign n27489 = P1_INSTQUEUE_REG_11__2_ & n27297;
  assign n27490 = ~n27486 & ~n27487;
  assign n27491 = ~n27488 & n27490;
  assign n27492 = ~n27489 & n27491;
  assign n27493 = P1_INSTQUEUE_REG_12__2_ & n27303;
  assign n27494 = P1_INSTQUEUE_REG_13__2_ & n27305;
  assign n27495 = P1_INSTQUEUE_REG_14__2_ & n27307;
  assign n27496 = P1_INSTQUEUE_REG_15__2_ & n27309;
  assign n27497 = ~n27493 & ~n27494;
  assign n27498 = ~n27495 & n27497;
  assign n27499 = ~n27496 & n27498;
  assign n27500 = n27478 & n27485;
  assign n27501 = n27492 & n27500;
  assign n27502 = n27499 & n27501;
  assign n27503 = ~n27317 & ~n27502;
  assign n27504 = ~n24683 & n27503;
  assign n27505 = n24683 & ~n27503;
  assign n27506 = ~n27504 & ~n27505;
  assign n27507 = ~n27321 & ~n27415;
  assign n27508 = ~n27333 & n27507;
  assign n27509 = ~n27506 & ~n27508;
  assign n27510 = n27506 & n27508;
  assign n27511 = ~n27509 & ~n27510;
  assign n27512 = n24136 & ~n27511;
  assign n27513 = P1_INSTADDRPOINTER_REG_10_ & ~n27512;
  assign n27514 = ~P1_INSTADDRPOINTER_REG_10_ & n27512;
  assign n27515 = ~n27513 & ~n27514;
  assign n27516 = n27471 & ~n27515;
  assign n27517 = ~P1_INSTADDRPOINTER_REG_10_ & ~n27512;
  assign n27518 = P1_INSTADDRPOINTER_REG_10_ & n27512;
  assign n27519 = ~n27517 & ~n27518;
  assign n27520 = ~n27471 & ~n27519;
  assign n27521 = ~n27516 & ~n27520;
  assign n27522 = n26641 & ~n27521;
  assign n27523 = n27460 & n27469;
  assign n6139 = n27522 | ~n27523;
  assign n27525 = P1_INSTADDRPOINTER_REG_9_ & P1_INSTADDRPOINTER_REG_10_;
  assign n27526 = n27349 & n27525;
  assign n27527 = P1_INSTADDRPOINTER_REG_11_ & ~n27526;
  assign n27528 = ~P1_INSTADDRPOINTER_REG_11_ & n27526;
  assign n27529 = ~n27527 & ~n27528;
  assign n27530 = n26651 & ~n27529;
  assign n27531 = P1_EBX_REG_11_ & ~n26656;
  assign n27532 = P1_INSTADDRPOINTER_REG_11_ & ~n26658;
  assign n27533 = ~n27531 & ~n27532;
  assign n27534 = ~n24166 & ~n27533;
  assign n27535 = n24166 & n27533;
  assign n27536 = ~n27534 & ~n27535;
  assign n27537 = ~n27447 & n27449;
  assign n27538 = ~n27536 & ~n27537;
  assign n27539 = n27536 & n27537;
  assign n27540 = ~n27538 & ~n27539;
  assign n27541 = n26669 & ~n27540;
  assign n27542 = P1_INSTADDRPOINTER_REG_10_ & n27454;
  assign n27543 = ~P1_INSTADDRPOINTER_REG_11_ & n27542;
  assign n27544 = P1_INSTADDRPOINTER_REG_11_ & ~n27542;
  assign n27545 = ~n27543 & ~n27544;
  assign n27546 = n26620 & ~n27545;
  assign n27547 = ~n27530 & ~n27541;
  assign n27548 = ~n27546 & n27547;
  assign n27549 = P1_REIP_REG_11_ & n26672;
  assign n27550 = P1_INSTADDRPOINTER_REG_11_ & n26618;
  assign n27551 = ~n27549 & ~n27550;
  assign n27552 = P1_INSTADDRPOINTER_REG_10_ & n27464;
  assign n27553 = ~P1_INSTADDRPOINTER_REG_11_ & n27552;
  assign n27554 = P1_INSTADDRPOINTER_REG_11_ & ~n27552;
  assign n27555 = ~n27553 & ~n27554;
  assign n27556 = n26676 & ~n27555;
  assign n27557 = n27551 & ~n27556;
  assign n27558 = ~n27421 & ~n27517;
  assign n27559 = ~n27518 & ~n27558;
  assign n27560 = P1_INSTQUEUE_REG_0__3_ & n27267;
  assign n27561 = P1_INSTQUEUE_REG_1__3_ & n27269;
  assign n27562 = P1_INSTQUEUE_REG_2__3_ & n27271;
  assign n27563 = P1_INSTQUEUE_REG_3__3_ & n27273;
  assign n27564 = ~n27560 & ~n27561;
  assign n27565 = ~n27562 & n27564;
  assign n27566 = ~n27563 & n27565;
  assign n27567 = P1_INSTQUEUE_REG_4__3_ & n27279;
  assign n27568 = P1_INSTQUEUE_REG_5__3_ & n27281;
  assign n27569 = P1_INSTQUEUE_REG_6__3_ & n27283;
  assign n27570 = P1_INSTQUEUE_REG_7__3_ & n27285;
  assign n27571 = ~n27567 & ~n27568;
  assign n27572 = ~n27569 & n27571;
  assign n27573 = ~n27570 & n27572;
  assign n27574 = P1_INSTQUEUE_REG_8__3_ & n27291;
  assign n27575 = P1_INSTQUEUE_REG_9__3_ & n27293;
  assign n27576 = P1_INSTQUEUE_REG_10__3_ & n27295;
  assign n27577 = P1_INSTQUEUE_REG_11__3_ & n27297;
  assign n27578 = ~n27574 & ~n27575;
  assign n27579 = ~n27576 & n27578;
  assign n27580 = ~n27577 & n27579;
  assign n27581 = P1_INSTQUEUE_REG_12__3_ & n27303;
  assign n27582 = P1_INSTQUEUE_REG_13__3_ & n27305;
  assign n27583 = P1_INSTQUEUE_REG_14__3_ & n27307;
  assign n27584 = P1_INSTQUEUE_REG_15__3_ & n27309;
  assign n27585 = ~n27581 & ~n27582;
  assign n27586 = ~n27583 & n27585;
  assign n27587 = ~n27584 & n27586;
  assign n27588 = n27566 & n27573;
  assign n27589 = n27580 & n27588;
  assign n27590 = n27587 & n27589;
  assign n27591 = ~n27317 & ~n27590;
  assign n27592 = ~n24683 & n27591;
  assign n27593 = n24683 & ~n27591;
  assign n27594 = ~n27592 & ~n27593;
  assign n27595 = ~n27415 & ~n27506;
  assign n27596 = ~n27321 & n27595;
  assign n27597 = ~n27333 & n27596;
  assign n27598 = ~n27594 & ~n27597;
  assign n27599 = n27594 & n27597;
  assign n27600 = ~n27598 & ~n27599;
  assign n27601 = n24136 & ~n27600;
  assign n27602 = ~P1_INSTADDRPOINTER_REG_11_ & ~n27601;
  assign n27603 = ~n27559 & ~n27602;
  assign n27604 = ~n27425 & ~n27518;
  assign n27605 = ~n27420 & n27604;
  assign n27606 = ~n27424 & ~n27429;
  assign n27607 = n27605 & n27606;
  assign n27608 = n27603 & ~n27607;
  assign n27609 = P1_INSTADDRPOINTER_REG_11_ & n27601;
  assign n27610 = n27608 & ~n27609;
  assign n27611 = P1_INSTADDRPOINTER_REG_11_ & ~n27601;
  assign n27612 = ~P1_INSTADDRPOINTER_REG_11_ & n27601;
  assign n27613 = ~n27611 & ~n27612;
  assign n27614 = ~n27518 & n27613;
  assign n27615 = ~n27471 & ~n27517;
  assign n27616 = n27614 & ~n27615;
  assign n27617 = ~n27610 & ~n27616;
  assign n27618 = n26641 & n27617;
  assign n27619 = n27548 & n27557;
  assign n6144 = n27618 | ~n27619;
  assign n27621 = P1_INSTADDRPOINTER_REG_11_ & n27526;
  assign n27622 = ~P1_INSTADDRPOINTER_REG_12_ & n27621;
  assign n27623 = P1_INSTADDRPOINTER_REG_12_ & ~n27621;
  assign n27624 = ~n27622 & ~n27623;
  assign n27625 = n26651 & ~n27624;
  assign n27626 = P1_EBX_REG_12_ & ~n26656;
  assign n27627 = P1_INSTADDRPOINTER_REG_12_ & ~n26658;
  assign n27628 = ~n27626 & ~n27627;
  assign n27629 = ~n24166 & ~n27628;
  assign n27630 = n24166 & n27628;
  assign n27631 = ~n27629 & ~n27630;
  assign n27632 = ~n27447 & ~n27536;
  assign n27633 = n27449 & n27632;
  assign n27634 = ~n27631 & ~n27633;
  assign n27635 = n27631 & n27633;
  assign n27636 = ~n27634 & ~n27635;
  assign n27637 = n26669 & ~n27636;
  assign n27638 = P1_INSTADDRPOINTER_REG_11_ & n27542;
  assign n27639 = ~P1_INSTADDRPOINTER_REG_12_ & n27638;
  assign n27640 = P1_INSTADDRPOINTER_REG_12_ & ~n27638;
  assign n27641 = ~n27639 & ~n27640;
  assign n27642 = n26620 & ~n27641;
  assign n27643 = ~n27625 & ~n27637;
  assign n27644 = ~n27642 & n27643;
  assign n27645 = P1_REIP_REG_12_ & n26672;
  assign n27646 = P1_INSTADDRPOINTER_REG_12_ & n26618;
  assign n27647 = ~n27645 & ~n27646;
  assign n27648 = P1_INSTADDRPOINTER_REG_11_ & n27552;
  assign n27649 = ~P1_INSTADDRPOINTER_REG_12_ & n27648;
  assign n27650 = P1_INSTADDRPOINTER_REG_12_ & ~n27648;
  assign n27651 = ~n27649 & ~n27650;
  assign n27652 = n26676 & ~n27651;
  assign n27653 = n27647 & ~n27652;
  assign n27654 = P1_INSTQUEUE_REG_0__4_ & n27267;
  assign n27655 = P1_INSTQUEUE_REG_1__4_ & n27269;
  assign n27656 = P1_INSTQUEUE_REG_2__4_ & n27271;
  assign n27657 = P1_INSTQUEUE_REG_3__4_ & n27273;
  assign n27658 = ~n27654 & ~n27655;
  assign n27659 = ~n27656 & n27658;
  assign n27660 = ~n27657 & n27659;
  assign n27661 = P1_INSTQUEUE_REG_4__4_ & n27279;
  assign n27662 = P1_INSTQUEUE_REG_5__4_ & n27281;
  assign n27663 = P1_INSTQUEUE_REG_6__4_ & n27283;
  assign n27664 = P1_INSTQUEUE_REG_7__4_ & n27285;
  assign n27665 = ~n27661 & ~n27662;
  assign n27666 = ~n27663 & n27665;
  assign n27667 = ~n27664 & n27666;
  assign n27668 = P1_INSTQUEUE_REG_8__4_ & n27291;
  assign n27669 = P1_INSTQUEUE_REG_9__4_ & n27293;
  assign n27670 = P1_INSTQUEUE_REG_10__4_ & n27295;
  assign n27671 = P1_INSTQUEUE_REG_11__4_ & n27297;
  assign n27672 = ~n27668 & ~n27669;
  assign n27673 = ~n27670 & n27672;
  assign n27674 = ~n27671 & n27673;
  assign n27675 = P1_INSTQUEUE_REG_12__4_ & n27303;
  assign n27676 = P1_INSTQUEUE_REG_13__4_ & n27305;
  assign n27677 = P1_INSTQUEUE_REG_14__4_ & n27307;
  assign n27678 = P1_INSTQUEUE_REG_15__4_ & n27309;
  assign n27679 = ~n27675 & ~n27676;
  assign n27680 = ~n27677 & n27679;
  assign n27681 = ~n27678 & n27680;
  assign n27682 = n27660 & n27667;
  assign n27683 = n27674 & n27682;
  assign n27684 = n27681 & n27683;
  assign n27685 = ~n27317 & ~n27684;
  assign n27686 = ~n24683 & n27685;
  assign n27687 = n24683 & ~n27685;
  assign n27688 = ~n27686 & ~n27687;
  assign n27689 = ~n27506 & ~n27594;
  assign n27690 = ~n27415 & n27689;
  assign n27691 = ~n27321 & n27690;
  assign n27692 = ~n27333 & n27691;
  assign n27693 = ~n27688 & ~n27692;
  assign n27694 = n27688 & n27692;
  assign n27695 = ~n27693 & ~n27694;
  assign n27696 = n24136 & ~n27695;
  assign n27697 = P1_INSTADDRPOINTER_REG_12_ & n27696;
  assign n27698 = ~P1_INSTADDRPOINTER_REG_12_ & ~n27696;
  assign n27699 = ~n27697 & ~n27698;
  assign n27700 = ~n27608 & ~n27609;
  assign n27701 = n27699 & n27700;
  assign n27702 = ~n27699 & ~n27700;
  assign n27703 = ~n27701 & ~n27702;
  assign n27704 = n26641 & ~n27703;
  assign n27705 = n27644 & n27653;
  assign n6149 = n27704 | ~n27705;
  assign n27707 = P1_REIP_REG_13_ & n26672;
  assign n27708 = P1_INSTADDRPOINTER_REG_13_ & n26618;
  assign n27709 = ~n27707 & ~n27708;
  assign n27710 = P1_INSTADDRPOINTER_REG_12_ & n27648;
  assign n27711 = ~P1_INSTADDRPOINTER_REG_13_ & n27710;
  assign n27712 = P1_INSTADDRPOINTER_REG_13_ & ~n27710;
  assign n27713 = ~n27711 & ~n27712;
  assign n27714 = n26676 & ~n27713;
  assign n27715 = n27709 & ~n27714;
  assign n27716 = P1_INSTADDRPOINTER_REG_11_ & P1_INSTADDRPOINTER_REG_12_;
  assign n27717 = n27526 & n27716;
  assign n27718 = P1_INSTADDRPOINTER_REG_13_ & ~n27717;
  assign n27719 = ~P1_INSTADDRPOINTER_REG_13_ & n27717;
  assign n27720 = ~n27718 & ~n27719;
  assign n27721 = n26651 & ~n27720;
  assign n27722 = P1_INSTADDRPOINTER_REG_12_ & n27638;
  assign n27723 = ~P1_INSTADDRPOINTER_REG_13_ & n27722;
  assign n27724 = P1_INSTADDRPOINTER_REG_13_ & ~n27722;
  assign n27725 = ~n27723 & ~n27724;
  assign n27726 = n26620 & ~n27725;
  assign n27727 = ~n27721 & ~n27726;
  assign n27728 = P1_EBX_REG_13_ & ~n26656;
  assign n27729 = P1_INSTADDRPOINTER_REG_13_ & ~n26658;
  assign n27730 = ~n27728 & ~n27729;
  assign n27731 = ~n24166 & ~n27730;
  assign n27732 = n24166 & n27730;
  assign n27733 = ~n27731 & ~n27732;
  assign n27734 = ~n27631 & n27633;
  assign n27735 = ~n27733 & ~n27734;
  assign n27736 = n27733 & n27734;
  assign n27737 = ~n27735 & ~n27736;
  assign n27738 = n26669 & ~n27737;
  assign n27739 = ~n27698 & ~n27700;
  assign n27740 = ~n27697 & ~n27739;
  assign n27741 = P1_INSTQUEUE_REG_0__5_ & n27267;
  assign n27742 = P1_INSTQUEUE_REG_1__5_ & n27269;
  assign n27743 = P1_INSTQUEUE_REG_2__5_ & n27271;
  assign n27744 = P1_INSTQUEUE_REG_3__5_ & n27273;
  assign n27745 = ~n27741 & ~n27742;
  assign n27746 = ~n27743 & n27745;
  assign n27747 = ~n27744 & n27746;
  assign n27748 = P1_INSTQUEUE_REG_4__5_ & n27279;
  assign n27749 = P1_INSTQUEUE_REG_5__5_ & n27281;
  assign n27750 = P1_INSTQUEUE_REG_6__5_ & n27283;
  assign n27751 = P1_INSTQUEUE_REG_7__5_ & n27285;
  assign n27752 = ~n27748 & ~n27749;
  assign n27753 = ~n27750 & n27752;
  assign n27754 = ~n27751 & n27753;
  assign n27755 = P1_INSTQUEUE_REG_8__5_ & n27291;
  assign n27756 = P1_INSTQUEUE_REG_9__5_ & n27293;
  assign n27757 = P1_INSTQUEUE_REG_10__5_ & n27295;
  assign n27758 = P1_INSTQUEUE_REG_11__5_ & n27297;
  assign n27759 = ~n27755 & ~n27756;
  assign n27760 = ~n27757 & n27759;
  assign n27761 = ~n27758 & n27760;
  assign n27762 = P1_INSTQUEUE_REG_12__5_ & n27303;
  assign n27763 = P1_INSTQUEUE_REG_13__5_ & n27305;
  assign n27764 = P1_INSTQUEUE_REG_14__5_ & n27307;
  assign n27765 = P1_INSTQUEUE_REG_15__5_ & n27309;
  assign n27766 = ~n27762 & ~n27763;
  assign n27767 = ~n27764 & n27766;
  assign n27768 = ~n27765 & n27767;
  assign n27769 = n27747 & n27754;
  assign n27770 = n27761 & n27769;
  assign n27771 = n27768 & n27770;
  assign n27772 = ~n27317 & ~n27771;
  assign n27773 = ~n24683 & n27772;
  assign n27774 = n24683 & ~n27772;
  assign n27775 = ~n27773 & ~n27774;
  assign n27776 = ~n27688 & n27692;
  assign n27777 = ~n27775 & ~n27776;
  assign n27778 = n27775 & n27776;
  assign n27779 = ~n27777 & ~n27778;
  assign n27780 = n24136 & ~n27779;
  assign n27781 = P1_INSTADDRPOINTER_REG_13_ & ~n27780;
  assign n27782 = ~P1_INSTADDRPOINTER_REG_13_ & n27780;
  assign n27783 = ~n27781 & ~n27782;
  assign n27784 = n27740 & ~n27783;
  assign n27785 = ~P1_INSTADDRPOINTER_REG_13_ & ~n27780;
  assign n27786 = P1_INSTADDRPOINTER_REG_13_ & n27780;
  assign n27787 = ~n27785 & ~n27786;
  assign n27788 = ~n27740 & ~n27787;
  assign n27789 = ~n27784 & ~n27788;
  assign n27790 = n26641 & ~n27789;
  assign n27791 = n27715 & n27727;
  assign n27792 = ~n27738 & n27791;
  assign n6154 = n27790 | ~n27792;
  assign n27794 = P1_REIP_REG_14_ & n26672;
  assign n27795 = P1_INSTADDRPOINTER_REG_14_ & n26618;
  assign n27796 = ~n27794 & ~n27795;
  assign n27797 = P1_INSTADDRPOINTER_REG_13_ & n27710;
  assign n27798 = ~P1_INSTADDRPOINTER_REG_14_ & n27797;
  assign n27799 = P1_INSTADDRPOINTER_REG_14_ & ~n27797;
  assign n27800 = ~n27798 & ~n27799;
  assign n27801 = n26676 & ~n27800;
  assign n27802 = n27796 & ~n27801;
  assign n27803 = P1_INSTADDRPOINTER_REG_13_ & n27717;
  assign n27804 = ~P1_INSTADDRPOINTER_REG_14_ & n27803;
  assign n27805 = P1_INSTADDRPOINTER_REG_14_ & ~n27803;
  assign n27806 = ~n27804 & ~n27805;
  assign n27807 = n26651 & ~n27806;
  assign n27808 = P1_INSTADDRPOINTER_REG_13_ & n27722;
  assign n27809 = ~P1_INSTADDRPOINTER_REG_14_ & n27808;
  assign n27810 = P1_INSTADDRPOINTER_REG_14_ & ~n27808;
  assign n27811 = ~n27809 & ~n27810;
  assign n27812 = n26620 & ~n27811;
  assign n27813 = ~n27807 & ~n27812;
  assign n27814 = P1_EBX_REG_14_ & ~n26656;
  assign n27815 = P1_INSTADDRPOINTER_REG_14_ & ~n26658;
  assign n27816 = ~n27814 & ~n27815;
  assign n27817 = ~n24166 & ~n27816;
  assign n27818 = n24166 & n27816;
  assign n27819 = ~n27817 & ~n27818;
  assign n27820 = ~n27631 & ~n27733;
  assign n27821 = n27633 & n27820;
  assign n27822 = ~n27819 & ~n27821;
  assign n27823 = n27819 & n27821;
  assign n27824 = ~n27822 & ~n27823;
  assign n27825 = n26669 & ~n27824;
  assign n27826 = P1_INSTQUEUE_REG_0__6_ & n27267;
  assign n27827 = P1_INSTQUEUE_REG_1__6_ & n27269;
  assign n27828 = P1_INSTQUEUE_REG_2__6_ & n27271;
  assign n27829 = P1_INSTQUEUE_REG_3__6_ & n27273;
  assign n27830 = ~n27826 & ~n27827;
  assign n27831 = ~n27828 & n27830;
  assign n27832 = ~n27829 & n27831;
  assign n27833 = P1_INSTQUEUE_REG_4__6_ & n27279;
  assign n27834 = P1_INSTQUEUE_REG_5__6_ & n27281;
  assign n27835 = P1_INSTQUEUE_REG_6__6_ & n27283;
  assign n27836 = P1_INSTQUEUE_REG_7__6_ & n27285;
  assign n27837 = ~n27833 & ~n27834;
  assign n27838 = ~n27835 & n27837;
  assign n27839 = ~n27836 & n27838;
  assign n27840 = P1_INSTQUEUE_REG_8__6_ & n27291;
  assign n27841 = P1_INSTQUEUE_REG_9__6_ & n27293;
  assign n27842 = P1_INSTQUEUE_REG_10__6_ & n27295;
  assign n27843 = P1_INSTQUEUE_REG_11__6_ & n27297;
  assign n27844 = ~n27840 & ~n27841;
  assign n27845 = ~n27842 & n27844;
  assign n27846 = ~n27843 & n27845;
  assign n27847 = P1_INSTQUEUE_REG_12__6_ & n27303;
  assign n27848 = P1_INSTQUEUE_REG_13__6_ & n27305;
  assign n27849 = P1_INSTQUEUE_REG_14__6_ & n27307;
  assign n27850 = P1_INSTQUEUE_REG_15__6_ & n27309;
  assign n27851 = ~n27847 & ~n27848;
  assign n27852 = ~n27849 & n27851;
  assign n27853 = ~n27850 & n27852;
  assign n27854 = n27832 & n27839;
  assign n27855 = n27846 & n27854;
  assign n27856 = n27853 & n27855;
  assign n27857 = ~n27317 & ~n27856;
  assign n27858 = ~n24683 & n27857;
  assign n27859 = n24683 & ~n27857;
  assign n27860 = ~n27858 & ~n27859;
  assign n27861 = ~n27688 & ~n27775;
  assign n27862 = n27692 & n27861;
  assign n27863 = ~n27860 & ~n27862;
  assign n27864 = n27860 & n27862;
  assign n27865 = ~n27863 & ~n27864;
  assign n27866 = n24136 & ~n27865;
  assign n27867 = P1_INSTADDRPOINTER_REG_14_ & ~n27866;
  assign n27868 = ~P1_INSTADDRPOINTER_REG_14_ & n27866;
  assign n27869 = ~n27867 & ~n27868;
  assign n27870 = ~n27740 & ~n27785;
  assign n27871 = ~n27786 & ~n27870;
  assign n27872 = ~n27869 & n27871;
  assign n27873 = ~P1_INSTADDRPOINTER_REG_14_ & ~n27866;
  assign n27874 = P1_INSTADDRPOINTER_REG_14_ & n27866;
  assign n27875 = ~n27873 & ~n27874;
  assign n27876 = ~n27871 & ~n27875;
  assign n27877 = ~n27872 & ~n27876;
  assign n27878 = n26641 & ~n27877;
  assign n27879 = n27802 & n27813;
  assign n27880 = ~n27825 & n27879;
  assign n6159 = n27878 | ~n27880;
  assign n27882 = P1_REIP_REG_15_ & n26672;
  assign n27883 = P1_INSTADDRPOINTER_REG_15_ & n26618;
  assign n27884 = ~n27882 & ~n27883;
  assign n27885 = P1_INSTADDRPOINTER_REG_14_ & n27797;
  assign n27886 = ~P1_INSTADDRPOINTER_REG_15_ & n27885;
  assign n27887 = P1_INSTADDRPOINTER_REG_15_ & ~n27885;
  assign n27888 = ~n27886 & ~n27887;
  assign n27889 = n26676 & ~n27888;
  assign n27890 = n27884 & ~n27889;
  assign n27891 = P1_INSTADDRPOINTER_REG_13_ & P1_INSTADDRPOINTER_REG_14_;
  assign n27892 = n27717 & n27891;
  assign n27893 = P1_INSTADDRPOINTER_REG_15_ & ~n27892;
  assign n27894 = ~P1_INSTADDRPOINTER_REG_15_ & n27892;
  assign n27895 = ~n27893 & ~n27894;
  assign n27896 = n26651 & ~n27895;
  assign n27897 = P1_INSTADDRPOINTER_REG_14_ & n27808;
  assign n27898 = ~P1_INSTADDRPOINTER_REG_15_ & n27897;
  assign n27899 = P1_INSTADDRPOINTER_REG_15_ & ~n27897;
  assign n27900 = ~n27898 & ~n27899;
  assign n27901 = n26620 & ~n27900;
  assign n27902 = ~n27896 & ~n27901;
  assign n27903 = P1_EBX_REG_15_ & ~n26656;
  assign n27904 = P1_INSTADDRPOINTER_REG_15_ & ~n26658;
  assign n27905 = ~n27903 & ~n27904;
  assign n27906 = ~n24166 & ~n27905;
  assign n27907 = n24166 & n27905;
  assign n27908 = ~n27906 & ~n27907;
  assign n27909 = ~n27819 & n27821;
  assign n27910 = ~n27908 & ~n27909;
  assign n27911 = n27908 & n27909;
  assign n27912 = ~n27910 & ~n27911;
  assign n27913 = n26669 & ~n27912;
  assign n27914 = P1_INSTQUEUE_REG_0__7_ & n27267;
  assign n27915 = P1_INSTQUEUE_REG_1__7_ & n27269;
  assign n27916 = P1_INSTQUEUE_REG_2__7_ & n27271;
  assign n27917 = P1_INSTQUEUE_REG_3__7_ & n27273;
  assign n27918 = ~n27914 & ~n27915;
  assign n27919 = ~n27916 & n27918;
  assign n27920 = ~n27917 & n27919;
  assign n27921 = P1_INSTQUEUE_REG_4__7_ & n27279;
  assign n27922 = P1_INSTQUEUE_REG_5__7_ & n27281;
  assign n27923 = P1_INSTQUEUE_REG_6__7_ & n27283;
  assign n27924 = P1_INSTQUEUE_REG_7__7_ & n27285;
  assign n27925 = ~n27921 & ~n27922;
  assign n27926 = ~n27923 & n27925;
  assign n27927 = ~n27924 & n27926;
  assign n27928 = P1_INSTQUEUE_REG_8__7_ & n27291;
  assign n27929 = P1_INSTQUEUE_REG_9__7_ & n27293;
  assign n27930 = P1_INSTQUEUE_REG_10__7_ & n27295;
  assign n27931 = P1_INSTQUEUE_REG_11__7_ & n27297;
  assign n27932 = ~n27928 & ~n27929;
  assign n27933 = ~n27930 & n27932;
  assign n27934 = ~n27931 & n27933;
  assign n27935 = P1_INSTQUEUE_REG_12__7_ & n27303;
  assign n27936 = P1_INSTQUEUE_REG_13__7_ & n27305;
  assign n27937 = P1_INSTQUEUE_REG_14__7_ & n27307;
  assign n27938 = P1_INSTQUEUE_REG_15__7_ & n27309;
  assign n27939 = ~n27935 & ~n27936;
  assign n27940 = ~n27937 & n27939;
  assign n27941 = ~n27938 & n27940;
  assign n27942 = n27920 & n27927;
  assign n27943 = n27934 & n27942;
  assign n27944 = n27941 & n27943;
  assign n27945 = ~n27317 & ~n27944;
  assign n27946 = ~n24683 & n27945;
  assign n27947 = n24683 & ~n27945;
  assign n27948 = ~n27946 & ~n27947;
  assign n27949 = ~n27860 & n27862;
  assign n27950 = ~n27948 & ~n27949;
  assign n27951 = n27948 & n27949;
  assign n27952 = ~n27950 & ~n27951;
  assign n27953 = n24136 & ~n27952;
  assign n27954 = P1_INSTADDRPOINTER_REG_15_ & n27953;
  assign n27955 = P1_INSTADDRPOINTER_REG_15_ & ~n27873;
  assign n27956 = ~n27873 & n27953;
  assign n27957 = ~n27955 & ~n27956;
  assign n27958 = ~n27954 & ~n27957;
  assign n27959 = n27871 & ~n27874;
  assign n27960 = n27958 & ~n27959;
  assign n27961 = P1_INSTADDRPOINTER_REG_15_ & ~n27953;
  assign n27962 = ~P1_INSTADDRPOINTER_REG_15_ & n27953;
  assign n27963 = ~n27961 & ~n27962;
  assign n27964 = ~n27874 & n27963;
  assign n27965 = ~n27871 & ~n27873;
  assign n27966 = n27964 & ~n27965;
  assign n27967 = ~n27960 & ~n27966;
  assign n27968 = n26641 & n27967;
  assign n27969 = n27890 & n27902;
  assign n27970 = ~n27913 & n27969;
  assign n6164 = n27968 | ~n27970;
  assign n27972 = P1_REIP_REG_16_ & n26672;
  assign n27973 = P1_INSTADDRPOINTER_REG_16_ & n26618;
  assign n27974 = ~n27972 & ~n27973;
  assign n27975 = P1_INSTADDRPOINTER_REG_15_ & n27885;
  assign n27976 = ~P1_INSTADDRPOINTER_REG_16_ & n27975;
  assign n27977 = P1_INSTADDRPOINTER_REG_16_ & ~n27975;
  assign n27978 = ~n27976 & ~n27977;
  assign n27979 = n26676 & ~n27978;
  assign n27980 = n27974 & ~n27979;
  assign n27981 = P1_INSTADDRPOINTER_REG_15_ & n27892;
  assign n27982 = ~P1_INSTADDRPOINTER_REG_16_ & n27981;
  assign n27983 = P1_INSTADDRPOINTER_REG_16_ & ~n27981;
  assign n27984 = ~n27982 & ~n27983;
  assign n27985 = n26651 & ~n27984;
  assign n27986 = P1_INSTADDRPOINTER_REG_15_ & n27897;
  assign n27987 = ~P1_INSTADDRPOINTER_REG_16_ & n27986;
  assign n27988 = P1_INSTADDRPOINTER_REG_16_ & ~n27986;
  assign n27989 = ~n27987 & ~n27988;
  assign n27990 = n26620 & ~n27989;
  assign n27991 = ~n27985 & ~n27990;
  assign n27992 = P1_EBX_REG_16_ & ~n26656;
  assign n27993 = P1_INSTADDRPOINTER_REG_16_ & ~n26658;
  assign n27994 = ~n27992 & ~n27993;
  assign n27995 = ~n24166 & ~n27994;
  assign n27996 = n24166 & n27994;
  assign n27997 = ~n27995 & ~n27996;
  assign n27998 = ~n27819 & ~n27908;
  assign n27999 = n27821 & n27998;
  assign n28000 = ~n27997 & ~n27999;
  assign n28001 = n27997 & n27999;
  assign n28002 = ~n28000 & ~n28001;
  assign n28003 = n26669 & ~n28002;
  assign n28004 = n27697 & ~n27785;
  assign n28005 = ~n27786 & ~n28004;
  assign n28006 = ~n27874 & n28005;
  assign n28007 = ~n27957 & ~n28006;
  assign n28008 = ~n27954 & ~n28007;
  assign n28009 = ~n27953 & ~n27955;
  assign n28010 = ~n27698 & ~n27785;
  assign n28011 = ~n27873 & n28010;
  assign n28012 = ~n28009 & n28011;
  assign n28013 = ~n27700 & n28012;
  assign n28014 = n28008 & ~n28013;
  assign n28015 = n27861 & ~n27948;
  assign n28016 = ~n27860 & n28015;
  assign n28017 = n27691 & n28016;
  assign n28018 = ~n27333 & n28017;
  assign n28019 = n24683 & ~n28018;
  assign n28020 = ~n24683 & n28018;
  assign n28021 = ~n28019 & ~n28020;
  assign n28022 = n24136 & ~n28021;
  assign n28023 = P1_INSTADDRPOINTER_REG_16_ & ~n28022;
  assign n28024 = ~P1_INSTADDRPOINTER_REG_16_ & n28022;
  assign n28025 = ~n28023 & ~n28024;
  assign n28026 = n28014 & ~n28025;
  assign n28027 = ~n28014 & n28025;
  assign n28028 = ~n28026 & ~n28027;
  assign n28029 = n26641 & ~n28028;
  assign n28030 = n27980 & n27991;
  assign n28031 = ~n28003 & n28030;
  assign n6169 = n28029 | ~n28031;
  assign n28033 = P1_REIP_REG_17_ & n26672;
  assign n28034 = P1_INSTADDRPOINTER_REG_17_ & n26618;
  assign n28035 = ~n28033 & ~n28034;
  assign n28036 = P1_INSTADDRPOINTER_REG_16_ & n27975;
  assign n28037 = ~P1_INSTADDRPOINTER_REG_17_ & n28036;
  assign n28038 = P1_INSTADDRPOINTER_REG_17_ & ~n28036;
  assign n28039 = ~n28037 & ~n28038;
  assign n28040 = n26676 & ~n28039;
  assign n28041 = n28035 & ~n28040;
  assign n28042 = P1_INSTADDRPOINTER_REG_15_ & P1_INSTADDRPOINTER_REG_16_;
  assign n28043 = n27892 & n28042;
  assign n28044 = P1_INSTADDRPOINTER_REG_17_ & ~n28043;
  assign n28045 = ~P1_INSTADDRPOINTER_REG_17_ & n28043;
  assign n28046 = ~n28044 & ~n28045;
  assign n28047 = n26651 & ~n28046;
  assign n28048 = P1_INSTADDRPOINTER_REG_16_ & n27986;
  assign n28049 = ~P1_INSTADDRPOINTER_REG_17_ & n28048;
  assign n28050 = P1_INSTADDRPOINTER_REG_17_ & ~n28048;
  assign n28051 = ~n28049 & ~n28050;
  assign n28052 = n26620 & ~n28051;
  assign n28053 = ~n28047 & ~n28052;
  assign n28054 = P1_EBX_REG_17_ & ~n26656;
  assign n28055 = P1_INSTADDRPOINTER_REG_17_ & ~n26658;
  assign n28056 = ~n28054 & ~n28055;
  assign n28057 = ~n24166 & ~n28056;
  assign n28058 = n24166 & n28056;
  assign n28059 = ~n28057 & ~n28058;
  assign n28060 = ~n27997 & n27999;
  assign n28061 = ~n28059 & ~n28060;
  assign n28062 = n28059 & n28060;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = n26669 & ~n28063;
  assign n28065 = P1_INSTADDRPOINTER_REG_16_ & n28022;
  assign n28066 = ~P1_INSTADDRPOINTER_REG_16_ & ~n28022;
  assign n28067 = ~n28014 & ~n28066;
  assign n28068 = ~n28065 & ~n28067;
  assign n28069 = n24136 & n28019;
  assign n28070 = P1_INSTADDRPOINTER_REG_17_ & ~n28069;
  assign n28071 = ~P1_INSTADDRPOINTER_REG_17_ & n28069;
  assign n28072 = ~n28070 & ~n28071;
  assign n28073 = n28068 & ~n28072;
  assign n28074 = ~n28068 & n28072;
  assign n28075 = ~n28073 & ~n28074;
  assign n28076 = n26641 & ~n28075;
  assign n28077 = n28041 & n28053;
  assign n28078 = ~n28064 & n28077;
  assign n6174 = n28076 | ~n28078;
  assign n28080 = P1_REIP_REG_18_ & n26672;
  assign n28081 = P1_INSTADDRPOINTER_REG_18_ & n26618;
  assign n28082 = ~n28080 & ~n28081;
  assign n28083 = P1_INSTADDRPOINTER_REG_17_ & n28036;
  assign n28084 = ~P1_INSTADDRPOINTER_REG_18_ & n28083;
  assign n28085 = P1_INSTADDRPOINTER_REG_18_ & ~n28083;
  assign n28086 = ~n28084 & ~n28085;
  assign n28087 = n26676 & ~n28086;
  assign n28088 = n28082 & ~n28087;
  assign n28089 = P1_INSTADDRPOINTER_REG_17_ & n28043;
  assign n28090 = ~P1_INSTADDRPOINTER_REG_18_ & n28089;
  assign n28091 = P1_INSTADDRPOINTER_REG_18_ & ~n28089;
  assign n28092 = ~n28090 & ~n28091;
  assign n28093 = n26651 & ~n28092;
  assign n28094 = P1_INSTADDRPOINTER_REG_17_ & n28048;
  assign n28095 = ~P1_INSTADDRPOINTER_REG_18_ & n28094;
  assign n28096 = P1_INSTADDRPOINTER_REG_18_ & ~n28094;
  assign n28097 = ~n28095 & ~n28096;
  assign n28098 = n26620 & ~n28097;
  assign n28099 = ~n28093 & ~n28098;
  assign n28100 = P1_EBX_REG_18_ & ~n26656;
  assign n28101 = P1_INSTADDRPOINTER_REG_18_ & ~n26658;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = ~n24166 & ~n28102;
  assign n28104 = n24166 & n28102;
  assign n28105 = ~n28103 & ~n28104;
  assign n28106 = ~n27997 & ~n28059;
  assign n28107 = n27999 & n28106;
  assign n28108 = ~n28105 & ~n28107;
  assign n28109 = n28105 & n28107;
  assign n28110 = ~n28108 & ~n28109;
  assign n28111 = n26669 & ~n28110;
  assign n28112 = P1_INSTADDRPOINTER_REG_17_ & n28069;
  assign n28113 = ~n28065 & ~n28112;
  assign n28114 = ~P1_INSTADDRPOINTER_REG_17_ & ~n28069;
  assign n28115 = ~n28113 & ~n28114;
  assign n28116 = ~n28066 & ~n28114;
  assign n28117 = ~n28014 & n28116;
  assign n28118 = ~n28115 & ~n28117;
  assign n28119 = P1_INSTADDRPOINTER_REG_18_ & ~n28069;
  assign n28120 = ~P1_INSTADDRPOINTER_REG_18_ & n28069;
  assign n28121 = ~n28119 & ~n28120;
  assign n28122 = n28118 & ~n28121;
  assign n28123 = ~n28118 & n28121;
  assign n28124 = ~n28122 & ~n28123;
  assign n28125 = n26641 & ~n28124;
  assign n28126 = n28088 & n28099;
  assign n28127 = ~n28111 & n28126;
  assign n6179 = n28125 | ~n28127;
  assign n28129 = P1_REIP_REG_19_ & n26672;
  assign n28130 = P1_INSTADDRPOINTER_REG_19_ & n26618;
  assign n28131 = ~n28129 & ~n28130;
  assign n28132 = P1_INSTADDRPOINTER_REG_18_ & n28083;
  assign n28133 = ~P1_INSTADDRPOINTER_REG_19_ & n28132;
  assign n28134 = P1_INSTADDRPOINTER_REG_19_ & ~n28132;
  assign n28135 = ~n28133 & ~n28134;
  assign n28136 = n26676 & ~n28135;
  assign n28137 = n28131 & ~n28136;
  assign n28138 = P1_INSTADDRPOINTER_REG_17_ & P1_INSTADDRPOINTER_REG_18_;
  assign n28139 = n28043 & n28138;
  assign n28140 = P1_INSTADDRPOINTER_REG_19_ & ~n28139;
  assign n28141 = ~P1_INSTADDRPOINTER_REG_19_ & n28139;
  assign n28142 = ~n28140 & ~n28141;
  assign n28143 = n26651 & ~n28142;
  assign n28144 = P1_INSTADDRPOINTER_REG_18_ & n28094;
  assign n28145 = ~P1_INSTADDRPOINTER_REG_19_ & n28144;
  assign n28146 = P1_INSTADDRPOINTER_REG_19_ & ~n28144;
  assign n28147 = ~n28145 & ~n28146;
  assign n28148 = n26620 & ~n28147;
  assign n28149 = ~n28143 & ~n28148;
  assign n28150 = P1_EBX_REG_19_ & ~n26656;
  assign n28151 = P1_INSTADDRPOINTER_REG_19_ & ~n26658;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = ~n24166 & ~n28152;
  assign n28154 = n24166 & n28152;
  assign n28155 = ~n28153 & ~n28154;
  assign n28156 = ~n28105 & n28107;
  assign n28157 = ~n28155 & ~n28156;
  assign n28158 = n28155 & n28156;
  assign n28159 = ~n28157 & ~n28158;
  assign n28160 = n26669 & ~n28159;
  assign n28161 = ~P1_INSTADDRPOINTER_REG_18_ & ~n28069;
  assign n28162 = ~n28114 & ~n28161;
  assign n28163 = ~n28113 & n28162;
  assign n28164 = P1_INSTADDRPOINTER_REG_18_ & n28069;
  assign n28165 = ~n28163 & ~n28164;
  assign n28166 = n28116 & ~n28161;
  assign n28167 = ~n28014 & n28166;
  assign n28168 = n28165 & ~n28167;
  assign n28169 = P1_INSTADDRPOINTER_REG_19_ & ~n28069;
  assign n28170 = ~P1_INSTADDRPOINTER_REG_19_ & n28069;
  assign n28171 = ~n28169 & ~n28170;
  assign n28172 = n28168 & ~n28171;
  assign n28173 = ~n28168 & n28171;
  assign n28174 = ~n28172 & ~n28173;
  assign n28175 = n26641 & ~n28174;
  assign n28176 = n28137 & n28149;
  assign n28177 = ~n28160 & n28176;
  assign n6184 = n28175 | ~n28177;
  assign n28179 = P1_REIP_REG_20_ & n26672;
  assign n28180 = P1_INSTADDRPOINTER_REG_20_ & n26618;
  assign n28181 = ~n28179 & ~n28180;
  assign n28182 = P1_INSTADDRPOINTER_REG_19_ & n28132;
  assign n28183 = ~P1_INSTADDRPOINTER_REG_20_ & n28182;
  assign n28184 = P1_INSTADDRPOINTER_REG_20_ & ~n28182;
  assign n28185 = ~n28183 & ~n28184;
  assign n28186 = n26676 & ~n28185;
  assign n28187 = n28181 & ~n28186;
  assign n28188 = P1_INSTADDRPOINTER_REG_19_ & n28139;
  assign n28189 = ~P1_INSTADDRPOINTER_REG_20_ & n28188;
  assign n28190 = P1_INSTADDRPOINTER_REG_20_ & ~n28188;
  assign n28191 = ~n28189 & ~n28190;
  assign n28192 = n26651 & ~n28191;
  assign n28193 = P1_INSTADDRPOINTER_REG_19_ & n28144;
  assign n28194 = ~P1_INSTADDRPOINTER_REG_20_ & n28193;
  assign n28195 = P1_INSTADDRPOINTER_REG_20_ & ~n28193;
  assign n28196 = ~n28194 & ~n28195;
  assign n28197 = n26620 & ~n28196;
  assign n28198 = ~n28192 & ~n28197;
  assign n28199 = P1_EBX_REG_20_ & ~n26656;
  assign n28200 = P1_INSTADDRPOINTER_REG_20_ & ~n26658;
  assign n28201 = ~n28199 & ~n28200;
  assign n28202 = ~n24166 & ~n28201;
  assign n28203 = n24166 & n28201;
  assign n28204 = ~n28202 & ~n28203;
  assign n28205 = ~n28155 & n28156;
  assign n28206 = ~n28204 & ~n28205;
  assign n28207 = n28204 & n28205;
  assign n28208 = ~n28206 & ~n28207;
  assign n28209 = n26669 & ~n28208;
  assign n28210 = P1_INSTADDRPOINTER_REG_19_ & n28069;
  assign n28211 = ~P1_INSTADDRPOINTER_REG_19_ & ~n28069;
  assign n28212 = ~n28168 & ~n28211;
  assign n28213 = ~n28210 & ~n28212;
  assign n28214 = P1_INSTADDRPOINTER_REG_20_ & ~n28069;
  assign n28215 = ~P1_INSTADDRPOINTER_REG_20_ & n28069;
  assign n28216 = ~n28214 & ~n28215;
  assign n28217 = n28213 & ~n28216;
  assign n28218 = ~n28213 & n28216;
  assign n28219 = ~n28217 & ~n28218;
  assign n28220 = n26641 & ~n28219;
  assign n28221 = n28187 & n28198;
  assign n28222 = ~n28209 & n28221;
  assign n6189 = n28220 | ~n28222;
  assign n28224 = P1_REIP_REG_21_ & n26672;
  assign n28225 = P1_INSTADDRPOINTER_REG_21_ & n26618;
  assign n28226 = ~n28224 & ~n28225;
  assign n28227 = P1_INSTADDRPOINTER_REG_20_ & n28182;
  assign n28228 = ~P1_INSTADDRPOINTER_REG_21_ & n28227;
  assign n28229 = P1_INSTADDRPOINTER_REG_21_ & ~n28227;
  assign n28230 = ~n28228 & ~n28229;
  assign n28231 = n26676 & ~n28230;
  assign n28232 = n28226 & ~n28231;
  assign n28233 = P1_INSTADDRPOINTER_REG_19_ & P1_INSTADDRPOINTER_REG_20_;
  assign n28234 = n28139 & n28233;
  assign n28235 = P1_INSTADDRPOINTER_REG_21_ & ~n28234;
  assign n28236 = ~P1_INSTADDRPOINTER_REG_21_ & n28234;
  assign n28237 = ~n28235 & ~n28236;
  assign n28238 = n26651 & ~n28237;
  assign n28239 = P1_INSTADDRPOINTER_REG_20_ & n28193;
  assign n28240 = ~P1_INSTADDRPOINTER_REG_21_ & n28239;
  assign n28241 = P1_INSTADDRPOINTER_REG_21_ & ~n28239;
  assign n28242 = ~n28240 & ~n28241;
  assign n28243 = n26620 & ~n28242;
  assign n28244 = ~n28238 & ~n28243;
  assign n28245 = P1_EBX_REG_21_ & ~n26656;
  assign n28246 = P1_INSTADDRPOINTER_REG_21_ & ~n26658;
  assign n28247 = ~n28245 & ~n28246;
  assign n28248 = ~n24166 & ~n28247;
  assign n28249 = n24166 & n28247;
  assign n28250 = ~n28248 & ~n28249;
  assign n28251 = ~n28204 & n28205;
  assign n28252 = ~n28250 & ~n28251;
  assign n28253 = n28250 & n28251;
  assign n28254 = ~n28252 & ~n28253;
  assign n28255 = n26669 & ~n28254;
  assign n28256 = ~P1_INSTADDRPOINTER_REG_20_ & ~n28069;
  assign n28257 = n28210 & ~n28256;
  assign n28258 = P1_INSTADDRPOINTER_REG_20_ & n28069;
  assign n28259 = ~n28257 & ~n28258;
  assign n28260 = ~n28211 & ~n28256;
  assign n28261 = ~n28168 & n28260;
  assign n28262 = n28259 & ~n28261;
  assign n28263 = P1_INSTADDRPOINTER_REG_21_ & ~n28069;
  assign n28264 = ~P1_INSTADDRPOINTER_REG_21_ & n28069;
  assign n28265 = ~n28263 & ~n28264;
  assign n28266 = n28262 & ~n28265;
  assign n28267 = ~n28262 & n28265;
  assign n28268 = ~n28266 & ~n28267;
  assign n28269 = n26641 & ~n28268;
  assign n28270 = n28232 & n28244;
  assign n28271 = ~n28255 & n28270;
  assign n6194 = n28269 | ~n28271;
  assign n28273 = P1_REIP_REG_22_ & n26672;
  assign n28274 = P1_INSTADDRPOINTER_REG_22_ & n26618;
  assign n28275 = ~n28273 & ~n28274;
  assign n28276 = P1_INSTADDRPOINTER_REG_21_ & n28227;
  assign n28277 = ~P1_INSTADDRPOINTER_REG_22_ & n28276;
  assign n28278 = P1_INSTADDRPOINTER_REG_22_ & ~n28276;
  assign n28279 = ~n28277 & ~n28278;
  assign n28280 = n26676 & ~n28279;
  assign n28281 = n28275 & ~n28280;
  assign n28282 = P1_INSTADDRPOINTER_REG_21_ & n28234;
  assign n28283 = ~P1_INSTADDRPOINTER_REG_22_ & n28282;
  assign n28284 = P1_INSTADDRPOINTER_REG_22_ & ~n28282;
  assign n28285 = ~n28283 & ~n28284;
  assign n28286 = n26651 & ~n28285;
  assign n28287 = P1_INSTADDRPOINTER_REG_21_ & n28239;
  assign n28288 = ~P1_INSTADDRPOINTER_REG_22_ & n28287;
  assign n28289 = P1_INSTADDRPOINTER_REG_22_ & ~n28287;
  assign n28290 = ~n28288 & ~n28289;
  assign n28291 = n26620 & ~n28290;
  assign n28292 = ~n28286 & ~n28291;
  assign n28293 = P1_EBX_REG_22_ & ~n26656;
  assign n28294 = P1_INSTADDRPOINTER_REG_22_ & ~n26658;
  assign n28295 = ~n28293 & ~n28294;
  assign n28296 = ~n24166 & ~n28295;
  assign n28297 = n24166 & n28295;
  assign n28298 = ~n28296 & ~n28297;
  assign n28299 = ~n28250 & n28251;
  assign n28300 = ~n28298 & ~n28299;
  assign n28301 = n28298 & n28299;
  assign n28302 = ~n28300 & ~n28301;
  assign n28303 = n26669 & ~n28302;
  assign n28304 = ~P1_INSTADDRPOINTER_REG_21_ & ~n28069;
  assign n28305 = ~n28259 & ~n28304;
  assign n28306 = P1_INSTADDRPOINTER_REG_21_ & n28069;
  assign n28307 = ~n28305 & ~n28306;
  assign n28308 = n28260 & ~n28304;
  assign n28309 = ~n28168 & n28308;
  assign n28310 = n28307 & ~n28309;
  assign n28311 = P1_INSTADDRPOINTER_REG_22_ & ~n28069;
  assign n28312 = ~P1_INSTADDRPOINTER_REG_22_ & n28069;
  assign n28313 = ~n28311 & ~n28312;
  assign n28314 = n28310 & ~n28313;
  assign n28315 = ~n28310 & n28313;
  assign n28316 = ~n28314 & ~n28315;
  assign n28317 = n26641 & ~n28316;
  assign n28318 = n28281 & n28292;
  assign n28319 = ~n28303 & n28318;
  assign n6199 = n28317 | ~n28319;
  assign n28321 = P1_REIP_REG_23_ & n26672;
  assign n28322 = P1_INSTADDRPOINTER_REG_23_ & n26618;
  assign n28323 = ~n28321 & ~n28322;
  assign n28324 = P1_INSTADDRPOINTER_REG_22_ & n28276;
  assign n28325 = ~P1_INSTADDRPOINTER_REG_23_ & n28324;
  assign n28326 = P1_INSTADDRPOINTER_REG_23_ & ~n28324;
  assign n28327 = ~n28325 & ~n28326;
  assign n28328 = n26676 & ~n28327;
  assign n28329 = n28323 & ~n28328;
  assign n28330 = P1_INSTADDRPOINTER_REG_21_ & P1_INSTADDRPOINTER_REG_22_;
  assign n28331 = n28234 & n28330;
  assign n28332 = P1_INSTADDRPOINTER_REG_23_ & ~n28331;
  assign n28333 = ~P1_INSTADDRPOINTER_REG_23_ & n28331;
  assign n28334 = ~n28332 & ~n28333;
  assign n28335 = n26651 & ~n28334;
  assign n28336 = P1_INSTADDRPOINTER_REG_22_ & n28287;
  assign n28337 = ~P1_INSTADDRPOINTER_REG_23_ & n28336;
  assign n28338 = P1_INSTADDRPOINTER_REG_23_ & ~n28336;
  assign n28339 = ~n28337 & ~n28338;
  assign n28340 = n26620 & ~n28339;
  assign n28341 = ~n28335 & ~n28340;
  assign n28342 = P1_EBX_REG_23_ & ~n26656;
  assign n28343 = P1_INSTADDRPOINTER_REG_23_ & ~n26658;
  assign n28344 = ~n28342 & ~n28343;
  assign n28345 = ~n24166 & ~n28344;
  assign n28346 = n24166 & n28344;
  assign n28347 = ~n28345 & ~n28346;
  assign n28348 = ~n28298 & n28299;
  assign n28349 = ~n28347 & ~n28348;
  assign n28350 = n28347 & n28348;
  assign n28351 = ~n28349 & ~n28350;
  assign n28352 = n26669 & ~n28351;
  assign n28353 = ~P1_INSTADDRPOINTER_REG_22_ & ~n28069;
  assign n28354 = n28162 & n28308;
  assign n28355 = ~n28113 & n28354;
  assign n28356 = ~n28353 & n28355;
  assign n28357 = n28164 & ~n28353;
  assign n28358 = n28308 & n28357;
  assign n28359 = ~n28356 & ~n28358;
  assign n28360 = n28308 & ~n28353;
  assign n28361 = n28166 & n28360;
  assign n28362 = ~n28014 & n28361;
  assign n28363 = ~n28307 & ~n28353;
  assign n28364 = P1_INSTADDRPOINTER_REG_22_ & n28069;
  assign n28365 = ~n28363 & ~n28364;
  assign n28366 = n28359 & ~n28362;
  assign n28367 = n28365 & n28366;
  assign n28368 = P1_INSTADDRPOINTER_REG_23_ & ~n28069;
  assign n28369 = ~P1_INSTADDRPOINTER_REG_23_ & n28069;
  assign n28370 = ~n28368 & ~n28369;
  assign n28371 = n28367 & ~n28370;
  assign n28372 = ~n28367 & n28370;
  assign n28373 = ~n28371 & ~n28372;
  assign n28374 = n26641 & ~n28373;
  assign n28375 = n28329 & n28341;
  assign n28376 = ~n28352 & n28375;
  assign n6204 = n28374 | ~n28376;
  assign n28378 = P1_REIP_REG_24_ & n26672;
  assign n28379 = P1_INSTADDRPOINTER_REG_24_ & n26618;
  assign n28380 = ~n28378 & ~n28379;
  assign n28381 = P1_INSTADDRPOINTER_REG_23_ & n28324;
  assign n28382 = ~P1_INSTADDRPOINTER_REG_24_ & n28381;
  assign n28383 = P1_INSTADDRPOINTER_REG_24_ & ~n28381;
  assign n28384 = ~n28382 & ~n28383;
  assign n28385 = n26676 & ~n28384;
  assign n28386 = n28380 & ~n28385;
  assign n28387 = P1_INSTADDRPOINTER_REG_23_ & n28331;
  assign n28388 = ~P1_INSTADDRPOINTER_REG_24_ & n28387;
  assign n28389 = P1_INSTADDRPOINTER_REG_24_ & ~n28387;
  assign n28390 = ~n28388 & ~n28389;
  assign n28391 = n26651 & ~n28390;
  assign n28392 = P1_INSTADDRPOINTER_REG_23_ & n28336;
  assign n28393 = ~P1_INSTADDRPOINTER_REG_24_ & n28392;
  assign n28394 = P1_INSTADDRPOINTER_REG_24_ & ~n28392;
  assign n28395 = ~n28393 & ~n28394;
  assign n28396 = n26620 & ~n28395;
  assign n28397 = ~n28391 & ~n28396;
  assign n28398 = P1_EBX_REG_24_ & ~n26656;
  assign n28399 = P1_INSTADDRPOINTER_REG_24_ & ~n26658;
  assign n28400 = ~n28398 & ~n28399;
  assign n28401 = ~n24166 & ~n28400;
  assign n28402 = n24166 & n28400;
  assign n28403 = ~n28401 & ~n28402;
  assign n28404 = ~n28347 & n28348;
  assign n28405 = ~n28403 & ~n28404;
  assign n28406 = n28403 & n28404;
  assign n28407 = ~n28405 & ~n28406;
  assign n28408 = n26669 & ~n28407;
  assign n28409 = ~P1_INSTADDRPOINTER_REG_23_ & ~n28069;
  assign n28410 = ~n28367 & ~n28409;
  assign n28411 = P1_INSTADDRPOINTER_REG_23_ & n28069;
  assign n28412 = ~n28410 & ~n28411;
  assign n28413 = P1_INSTADDRPOINTER_REG_24_ & ~n28069;
  assign n28414 = ~P1_INSTADDRPOINTER_REG_24_ & n28069;
  assign n28415 = ~n28413 & ~n28414;
  assign n28416 = n28412 & ~n28415;
  assign n28417 = ~n28412 & n28415;
  assign n28418 = ~n28416 & ~n28417;
  assign n28419 = n26641 & ~n28418;
  assign n28420 = n28386 & n28397;
  assign n28421 = ~n28408 & n28420;
  assign n6209 = n28419 | ~n28421;
  assign n28423 = P1_REIP_REG_25_ & n26672;
  assign n28424 = P1_INSTADDRPOINTER_REG_25_ & n26618;
  assign n28425 = ~n28423 & ~n28424;
  assign n28426 = P1_INSTADDRPOINTER_REG_24_ & n28381;
  assign n28427 = ~P1_INSTADDRPOINTER_REG_25_ & n28426;
  assign n28428 = P1_INSTADDRPOINTER_REG_25_ & ~n28426;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 = n26676 & ~n28429;
  assign n28431 = n28425 & ~n28430;
  assign n28432 = P1_INSTADDRPOINTER_REG_23_ & P1_INSTADDRPOINTER_REG_24_;
  assign n28433 = n28331 & n28432;
  assign n28434 = P1_INSTADDRPOINTER_REG_25_ & ~n28433;
  assign n28435 = ~P1_INSTADDRPOINTER_REG_25_ & n28433;
  assign n28436 = ~n28434 & ~n28435;
  assign n28437 = n26651 & ~n28436;
  assign n28438 = P1_INSTADDRPOINTER_REG_24_ & n28392;
  assign n28439 = ~P1_INSTADDRPOINTER_REG_25_ & n28438;
  assign n28440 = P1_INSTADDRPOINTER_REG_25_ & ~n28438;
  assign n28441 = ~n28439 & ~n28440;
  assign n28442 = n26620 & ~n28441;
  assign n28443 = ~n28437 & ~n28442;
  assign n28444 = P1_EBX_REG_25_ & ~n26656;
  assign n28445 = P1_INSTADDRPOINTER_REG_25_ & ~n26658;
  assign n28446 = ~n28444 & ~n28445;
  assign n28447 = ~n24166 & ~n28446;
  assign n28448 = n24166 & n28446;
  assign n28449 = ~n28447 & ~n28448;
  assign n28450 = ~n28403 & n28404;
  assign n28451 = ~n28449 & ~n28450;
  assign n28452 = n28449 & n28450;
  assign n28453 = ~n28451 & ~n28452;
  assign n28454 = n26669 & ~n28453;
  assign n28455 = ~P1_INSTADDRPOINTER_REG_24_ & ~n28069;
  assign n28456 = n28411 & ~n28455;
  assign n28457 = P1_INSTADDRPOINTER_REG_24_ & n28069;
  assign n28458 = ~n28456 & ~n28457;
  assign n28459 = ~n28409 & ~n28455;
  assign n28460 = ~n28367 & n28459;
  assign n28461 = n28458 & ~n28460;
  assign n28462 = P1_INSTADDRPOINTER_REG_25_ & ~n28069;
  assign n28463 = ~P1_INSTADDRPOINTER_REG_25_ & n28069;
  assign n28464 = ~n28462 & ~n28463;
  assign n28465 = n28461 & ~n28464;
  assign n28466 = ~n28461 & n28464;
  assign n28467 = ~n28465 & ~n28466;
  assign n28468 = n26641 & ~n28467;
  assign n28469 = n28431 & n28443;
  assign n28470 = ~n28454 & n28469;
  assign n6214 = n28468 | ~n28470;
  assign n28472 = P1_REIP_REG_26_ & n26672;
  assign n28473 = P1_INSTADDRPOINTER_REG_26_ & n26618;
  assign n28474 = ~n28472 & ~n28473;
  assign n28475 = P1_INSTADDRPOINTER_REG_25_ & n28426;
  assign n28476 = ~P1_INSTADDRPOINTER_REG_26_ & n28475;
  assign n28477 = P1_INSTADDRPOINTER_REG_26_ & ~n28475;
  assign n28478 = ~n28476 & ~n28477;
  assign n28479 = n26676 & ~n28478;
  assign n28480 = n28474 & ~n28479;
  assign n28481 = P1_INSTADDRPOINTER_REG_25_ & n28433;
  assign n28482 = ~P1_INSTADDRPOINTER_REG_26_ & n28481;
  assign n28483 = P1_INSTADDRPOINTER_REG_26_ & ~n28481;
  assign n28484 = ~n28482 & ~n28483;
  assign n28485 = n26651 & ~n28484;
  assign n28486 = P1_INSTADDRPOINTER_REG_25_ & n28438;
  assign n28487 = ~P1_INSTADDRPOINTER_REG_26_ & n28486;
  assign n28488 = P1_INSTADDRPOINTER_REG_26_ & ~n28486;
  assign n28489 = ~n28487 & ~n28488;
  assign n28490 = n26620 & ~n28489;
  assign n28491 = ~n28485 & ~n28490;
  assign n28492 = P1_EBX_REG_26_ & ~n26656;
  assign n28493 = P1_INSTADDRPOINTER_REG_26_ & ~n26658;
  assign n28494 = ~n28492 & ~n28493;
  assign n28495 = ~n24166 & ~n28494;
  assign n28496 = n24166 & n28494;
  assign n28497 = ~n28495 & ~n28496;
  assign n28498 = ~n28449 & n28450;
  assign n28499 = ~n28497 & ~n28498;
  assign n28500 = n28497 & n28498;
  assign n28501 = ~n28499 & ~n28500;
  assign n28502 = n26669 & ~n28501;
  assign n28503 = ~P1_INSTADDRPOINTER_REG_25_ & ~n28069;
  assign n28504 = ~n28458 & ~n28503;
  assign n28505 = P1_INSTADDRPOINTER_REG_25_ & n28069;
  assign n28506 = ~n28504 & ~n28505;
  assign n28507 = n28459 & ~n28503;
  assign n28508 = ~n28367 & n28507;
  assign n28509 = n28506 & ~n28508;
  assign n28510 = P1_INSTADDRPOINTER_REG_26_ & ~n28069;
  assign n28511 = ~P1_INSTADDRPOINTER_REG_26_ & n28069;
  assign n28512 = ~n28510 & ~n28511;
  assign n28513 = n28509 & ~n28512;
  assign n28514 = ~n28509 & n28512;
  assign n28515 = ~n28513 & ~n28514;
  assign n28516 = n26641 & ~n28515;
  assign n28517 = n28480 & n28491;
  assign n28518 = ~n28502 & n28517;
  assign n6219 = n28516 | ~n28518;
  assign n28520 = P1_REIP_REG_27_ & n26672;
  assign n28521 = P1_INSTADDRPOINTER_REG_27_ & n26618;
  assign n28522 = ~n28520 & ~n28521;
  assign n28523 = P1_INSTADDRPOINTER_REG_26_ & n28475;
  assign n28524 = ~P1_INSTADDRPOINTER_REG_27_ & n28523;
  assign n28525 = P1_INSTADDRPOINTER_REG_27_ & ~n28523;
  assign n28526 = ~n28524 & ~n28525;
  assign n28527 = n26676 & ~n28526;
  assign n28528 = n28522 & ~n28527;
  assign n28529 = P1_INSTADDRPOINTER_REG_25_ & P1_INSTADDRPOINTER_REG_26_;
  assign n28530 = n28433 & n28529;
  assign n28531 = P1_INSTADDRPOINTER_REG_27_ & ~n28530;
  assign n28532 = ~P1_INSTADDRPOINTER_REG_27_ & n28530;
  assign n28533 = ~n28531 & ~n28532;
  assign n28534 = n26651 & ~n28533;
  assign n28535 = P1_INSTADDRPOINTER_REG_26_ & n28486;
  assign n28536 = ~P1_INSTADDRPOINTER_REG_27_ & n28535;
  assign n28537 = P1_INSTADDRPOINTER_REG_27_ & ~n28535;
  assign n28538 = ~n28536 & ~n28537;
  assign n28539 = n26620 & ~n28538;
  assign n28540 = ~n28534 & ~n28539;
  assign n28541 = P1_EBX_REG_27_ & ~n26656;
  assign n28542 = P1_INSTADDRPOINTER_REG_27_ & ~n26658;
  assign n28543 = ~n28541 & ~n28542;
  assign n28544 = ~n24166 & ~n28543;
  assign n28545 = n24166 & n28543;
  assign n28546 = ~n28544 & ~n28545;
  assign n28547 = ~n28497 & n28498;
  assign n28548 = ~n28546 & ~n28547;
  assign n28549 = n28546 & n28547;
  assign n28550 = ~n28548 & ~n28549;
  assign n28551 = n26669 & ~n28550;
  assign n28552 = ~P1_INSTADDRPOINTER_REG_26_ & ~n28069;
  assign n28553 = n28507 & ~n28552;
  assign n28554 = ~n28367 & n28553;
  assign n28555 = P1_INSTADDRPOINTER_REG_26_ & n28069;
  assign n28556 = ~n28505 & ~n28555;
  assign n28557 = ~n28504 & n28556;
  assign n28558 = ~n28552 & ~n28557;
  assign n28559 = ~n28554 & ~n28558;
  assign n28560 = P1_INSTADDRPOINTER_REG_27_ & ~n28069;
  assign n28561 = ~P1_INSTADDRPOINTER_REG_27_ & n28069;
  assign n28562 = ~n28560 & ~n28561;
  assign n28563 = n28559 & ~n28562;
  assign n28564 = ~n28559 & n28562;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = n26641 & ~n28565;
  assign n28567 = n28528 & n28540;
  assign n28568 = ~n28551 & n28567;
  assign n6224 = n28566 | ~n28568;
  assign n28570 = P1_REIP_REG_28_ & n26672;
  assign n28571 = P1_INSTADDRPOINTER_REG_28_ & n26618;
  assign n28572 = ~n28570 & ~n28571;
  assign n28573 = P1_INSTADDRPOINTER_REG_27_ & n28523;
  assign n28574 = ~P1_INSTADDRPOINTER_REG_28_ & n28573;
  assign n28575 = P1_INSTADDRPOINTER_REG_28_ & ~n28573;
  assign n28576 = ~n28574 & ~n28575;
  assign n28577 = n26676 & ~n28576;
  assign n28578 = n28572 & ~n28577;
  assign n28579 = P1_INSTADDRPOINTER_REG_27_ & n28530;
  assign n28580 = ~P1_INSTADDRPOINTER_REG_28_ & n28579;
  assign n28581 = P1_INSTADDRPOINTER_REG_28_ & ~n28579;
  assign n28582 = ~n28580 & ~n28581;
  assign n28583 = n26651 & ~n28582;
  assign n28584 = P1_INSTADDRPOINTER_REG_27_ & n28535;
  assign n28585 = ~P1_INSTADDRPOINTER_REG_28_ & n28584;
  assign n28586 = P1_INSTADDRPOINTER_REG_28_ & ~n28584;
  assign n28587 = ~n28585 & ~n28586;
  assign n28588 = n26620 & ~n28587;
  assign n28589 = ~n28583 & ~n28588;
  assign n28590 = P1_EBX_REG_28_ & ~n26656;
  assign n28591 = P1_INSTADDRPOINTER_REG_28_ & ~n26658;
  assign n28592 = ~n28590 & ~n28591;
  assign n28593 = ~n24166 & ~n28592;
  assign n28594 = n24166 & n28592;
  assign n28595 = ~n28593 & ~n28594;
  assign n28596 = ~n28546 & n28547;
  assign n28597 = ~n28595 & ~n28596;
  assign n28598 = n28595 & n28596;
  assign n28599 = ~n28597 & ~n28598;
  assign n28600 = n26669 & ~n28599;
  assign n28601 = ~P1_INSTADDRPOINTER_REG_27_ & ~n28069;
  assign n28602 = ~n28552 & ~n28601;
  assign n28603 = n28507 & n28602;
  assign n28604 = ~n28367 & n28603;
  assign n28605 = P1_INSTADDRPOINTER_REG_27_ & n28069;
  assign n28606 = ~n28558 & ~n28605;
  assign n28607 = ~n28601 & ~n28606;
  assign n28608 = ~n28604 & ~n28607;
  assign n28609 = ~P1_INSTADDRPOINTER_REG_28_ & n28069;
  assign n28610 = P1_INSTADDRPOINTER_REG_28_ & ~n28069;
  assign n28611 = ~n28609 & ~n28610;
  assign n28612 = n28608 & ~n28611;
  assign n28613 = ~n28608 & n28611;
  assign n28614 = ~n28612 & ~n28613;
  assign n28615 = n26641 & ~n28614;
  assign n28616 = n28578 & n28589;
  assign n28617 = ~n28600 & n28616;
  assign n6229 = n28615 | ~n28617;
  assign n28619 = P1_REIP_REG_29_ & n26672;
  assign n28620 = P1_INSTADDRPOINTER_REG_29_ & n26618;
  assign n28621 = ~n28619 & ~n28620;
  assign n28622 = P1_INSTADDRPOINTER_REG_28_ & n28573;
  assign n28623 = ~P1_INSTADDRPOINTER_REG_29_ & n28622;
  assign n28624 = P1_INSTADDRPOINTER_REG_29_ & ~n28622;
  assign n28625 = ~n28623 & ~n28624;
  assign n28626 = n26676 & ~n28625;
  assign n28627 = n28621 & ~n28626;
  assign n28628 = P1_INSTADDRPOINTER_REG_27_ & P1_INSTADDRPOINTER_REG_28_;
  assign n28629 = n28530 & n28628;
  assign n28630 = P1_INSTADDRPOINTER_REG_29_ & ~n28629;
  assign n28631 = ~P1_INSTADDRPOINTER_REG_29_ & n28629;
  assign n28632 = ~n28630 & ~n28631;
  assign n28633 = n26651 & ~n28632;
  assign n28634 = P1_INSTADDRPOINTER_REG_28_ & n28584;
  assign n28635 = ~P1_INSTADDRPOINTER_REG_29_ & n28634;
  assign n28636 = P1_INSTADDRPOINTER_REG_29_ & ~n28634;
  assign n28637 = ~n28635 & ~n28636;
  assign n28638 = n26620 & ~n28637;
  assign n28639 = ~n28633 & ~n28638;
  assign n28640 = P1_EBX_REG_29_ & ~n26656;
  assign n28641 = P1_INSTADDRPOINTER_REG_29_ & ~n26658;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = ~n24166 & ~n28642;
  assign n28644 = n24166 & n28642;
  assign n28645 = ~n28643 & ~n28644;
  assign n28646 = ~n28595 & n28596;
  assign n28647 = ~n28645 & ~n28646;
  assign n28648 = n28645 & n28646;
  assign n28649 = ~n28647 & ~n28648;
  assign n28650 = n26669 & ~n28649;
  assign n28651 = ~P1_INSTADDRPOINTER_REG_28_ & ~n28069;
  assign n28652 = ~n28353 & ~n28651;
  assign n28653 = n28603 & n28652;
  assign n28654 = ~n28307 & n28653;
  assign n28655 = n28602 & ~n28651;
  assign n28656 = ~n28557 & n28655;
  assign n28657 = ~n28654 & ~n28656;
  assign n28658 = n28360 & ~n28651;
  assign n28659 = n28166 & n28658;
  assign n28660 = ~n28014 & n28603;
  assign n28661 = n28659 & n28660;
  assign n28662 = n28605 & ~n28651;
  assign n28663 = P1_INSTADDRPOINTER_REG_28_ & n28069;
  assign n28664 = ~n28662 & ~n28663;
  assign n28665 = n28364 & ~n28651;
  assign n28666 = n28603 & n28665;
  assign n28667 = n28603 & ~n28651;
  assign n28668 = n28358 & n28667;
  assign n28669 = n28664 & ~n28666;
  assign n28670 = ~n28668 & n28669;
  assign n28671 = n28356 & n28667;
  assign n28672 = n28670 & ~n28671;
  assign n28673 = n28657 & ~n28661;
  assign n28674 = n28672 & n28673;
  assign n28675 = ~P1_INSTADDRPOINTER_REG_29_ & n28069;
  assign n28676 = P1_INSTADDRPOINTER_REG_29_ & ~n28069;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = n28674 & ~n28677;
  assign n28679 = ~n28674 & n28677;
  assign n28680 = ~n28678 & ~n28679;
  assign n28681 = n26641 & ~n28680;
  assign n28682 = n28627 & n28639;
  assign n28683 = ~n28650 & n28682;
  assign n6234 = n28681 | ~n28683;
  assign n28685 = P1_REIP_REG_30_ & n26672;
  assign n28686 = P1_INSTADDRPOINTER_REG_30_ & n26618;
  assign n28687 = ~n28685 & ~n28686;
  assign n28688 = P1_INSTADDRPOINTER_REG_29_ & n28622;
  assign n28689 = ~P1_INSTADDRPOINTER_REG_30_ & n28688;
  assign n28690 = P1_INSTADDRPOINTER_REG_30_ & ~n28688;
  assign n28691 = ~n28689 & ~n28690;
  assign n28692 = n26676 & ~n28691;
  assign n28693 = n28687 & ~n28692;
  assign n28694 = P1_INSTADDRPOINTER_REG_29_ & n28629;
  assign n28695 = ~P1_INSTADDRPOINTER_REG_30_ & n28694;
  assign n28696 = P1_INSTADDRPOINTER_REG_30_ & ~n28694;
  assign n28697 = ~n28695 & ~n28696;
  assign n28698 = n26651 & ~n28697;
  assign n28699 = P1_INSTADDRPOINTER_REG_29_ & n28634;
  assign n28700 = ~P1_INSTADDRPOINTER_REG_30_ & n28699;
  assign n28701 = P1_INSTADDRPOINTER_REG_30_ & ~n28699;
  assign n28702 = ~n28700 & ~n28701;
  assign n28703 = n26620 & ~n28702;
  assign n28704 = ~n28698 & ~n28703;
  assign n28705 = P1_EBX_REG_30_ & ~n26656;
  assign n28706 = P1_INSTADDRPOINTER_REG_30_ & ~n26658;
  assign n28707 = ~n28705 & ~n28706;
  assign n28708 = ~n24166 & ~n28707;
  assign n28709 = n24166 & n28707;
  assign n28710 = ~n28708 & ~n28709;
  assign n28711 = ~n28645 & n28646;
  assign n28712 = ~n28710 & ~n28711;
  assign n28713 = n28710 & n28711;
  assign n28714 = ~n28712 & ~n28713;
  assign n28715 = n26669 & ~n28714;
  assign n28716 = ~P1_INSTADDRPOINTER_REG_29_ & ~n28069;
  assign n28717 = n28671 & ~n28716;
  assign n28718 = n28603 & ~n28716;
  assign n28719 = ~n28014 & n28718;
  assign n28720 = n28659 & n28719;
  assign n28721 = ~n28670 & ~n28716;
  assign n28722 = n28656 & ~n28716;
  assign n28723 = P1_INSTADDRPOINTER_REG_29_ & n28069;
  assign n28724 = n28654 & ~n28716;
  assign n28725 = ~n28722 & ~n28723;
  assign n28726 = ~n28724 & n28725;
  assign n28727 = ~n28717 & ~n28720;
  assign n28728 = ~n28721 & n28727;
  assign n28729 = n28726 & n28728;
  assign n28730 = ~P1_INSTADDRPOINTER_REG_30_ & n28069;
  assign n28731 = P1_INSTADDRPOINTER_REG_30_ & ~n28069;
  assign n28732 = ~n28730 & ~n28731;
  assign n28733 = n28729 & ~n28732;
  assign n28734 = ~n28729 & n28732;
  assign n28735 = ~n28733 & ~n28734;
  assign n28736 = n26641 & ~n28735;
  assign n28737 = n28693 & n28704;
  assign n28738 = ~n28715 & n28737;
  assign n6239 = n28736 | ~n28738;
  assign n28740 = P1_REIP_REG_31_ & n26672;
  assign n28741 = P1_INSTADDRPOINTER_REG_31_ & n26618;
  assign n28742 = ~n28740 & ~n28741;
  assign n28743 = P1_INSTADDRPOINTER_REG_30_ & n28688;
  assign n28744 = ~P1_INSTADDRPOINTER_REG_31_ & n28743;
  assign n28745 = P1_INSTADDRPOINTER_REG_31_ & ~n28743;
  assign n28746 = ~n28744 & ~n28745;
  assign n28747 = n26676 & ~n28746;
  assign n28748 = n28742 & ~n28747;
  assign n28749 = P1_INSTADDRPOINTER_REG_30_ & n28694;
  assign n28750 = ~P1_INSTADDRPOINTER_REG_31_ & n28749;
  assign n28751 = P1_INSTADDRPOINTER_REG_31_ & ~n28749;
  assign n28752 = ~n28750 & ~n28751;
  assign n28753 = n26651 & ~n28752;
  assign n28754 = P1_INSTADDRPOINTER_REG_30_ & n28699;
  assign n28755 = ~P1_INSTADDRPOINTER_REG_31_ & n28754;
  assign n28756 = P1_INSTADDRPOINTER_REG_31_ & ~n28754;
  assign n28757 = ~n28755 & ~n28756;
  assign n28758 = n26620 & ~n28757;
  assign n28759 = ~n28753 & ~n28758;
  assign n28760 = P1_EBX_REG_31_ & ~n26656;
  assign n28761 = P1_INSTADDRPOINTER_REG_31_ & ~n26658;
  assign n28762 = ~n28760 & ~n28761;
  assign n28763 = ~n24166 & ~n28762;
  assign n28764 = n24166 & n28762;
  assign n28765 = ~n28763 & ~n28764;
  assign n28766 = ~n28645 & ~n28710;
  assign n28767 = n28646 & n28766;
  assign n28768 = ~n28765 & ~n28767;
  assign n28769 = n28765 & n28767;
  assign n28770 = ~n28768 & ~n28769;
  assign n28771 = n26669 & ~n28770;
  assign n28772 = ~P1_INSTADDRPOINTER_REG_31_ & n28069;
  assign n28773 = P1_INSTADDRPOINTER_REG_31_ & ~n28069;
  assign n28774 = ~n28772 & ~n28773;
  assign n28775 = n28069 & ~n28774;
  assign n28776 = P1_INSTADDRPOINTER_REG_30_ & n28775;
  assign n28777 = ~n28069 & n28774;
  assign n28778 = ~P1_INSTADDRPOINTER_REG_30_ & n28777;
  assign n28779 = ~n28776 & ~n28778;
  assign n28780 = ~P1_INSTADDRPOINTER_REG_30_ & ~n28069;
  assign n28781 = ~n28774 & ~n28780;
  assign n28782 = ~n28716 & n28781;
  assign n28783 = ~n28674 & n28782;
  assign n28784 = n28723 & n28781;
  assign n28785 = n28652 & ~n28716;
  assign n28786 = n28603 & n28785;
  assign n28787 = ~n28307 & n28786;
  assign n28788 = ~n28651 & ~n28716;
  assign n28789 = ~n28601 & n28788;
  assign n28790 = ~n28552 & n28789;
  assign n28791 = ~n28557 & n28790;
  assign n28792 = P1_INSTADDRPOINTER_REG_30_ & n28069;
  assign n28793 = n28666 & ~n28716;
  assign n28794 = n28668 & ~n28716;
  assign n28795 = ~n28664 & ~n28716;
  assign n28796 = n28603 & n28788;
  assign n28797 = n28356 & n28796;
  assign n28798 = n28774 & ~n28795;
  assign n28799 = ~n28797 & n28798;
  assign n28800 = ~n28791 & ~n28792;
  assign n28801 = ~n28793 & n28800;
  assign n28802 = ~n28794 & n28801;
  assign n28803 = n28799 & n28802;
  assign n28804 = ~n28720 & ~n28787;
  assign n28805 = n28803 & n28804;
  assign n28806 = ~n28723 & n28805;
  assign n28807 = n28779 & ~n28783;
  assign n28808 = ~n28784 & n28807;
  assign n28809 = ~n28806 & n28808;
  assign n28810 = n26641 & n28809;
  assign n28811 = n28748 & n28759;
  assign n28812 = ~n28771 & n28811;
  assign n6244 = n28810 | ~n28812;
  assign n28814 = ~P1_STATE2_REG_0_ & n24626;
  assign n28815 = ~n24308 & ~n28814;
  assign n28816 = P1_STATE2_REG_2_ & n24240;
  assign n28817 = ~P1_STATE2_REG_1_ & ~n23741;
  assign n28818 = n24002 & n28817;
  assign n28819 = n24050 & n28816;
  assign n28820 = n28818 & n28819;
  assign n28821 = n24179 & n28820;
  assign n28822 = n28815 & ~n28821;
  assign n28823 = P1_STATE2_REG_0_ & ~n28822;
  assign n28824 = ~n26629 & n28823;
  assign n28825 = P1_STATE2_REG_1_ & ~P1_STATEBS16_REG;
  assign n28826 = P1_STATE2_REG_2_ & ~P1_STATE2_REG_0_;
  assign n28827 = ~n28825 & ~n28826;
  assign n28828 = ~n28822 & ~n28827;
  assign n28829 = P1_PHYADDRPOINTER_REG_0_ & n28828;
  assign n28830 = n24591 & ~n28822;
  assign n28831 = P1_REIP_REG_0_ & n28830;
  assign n28832 = P1_PHYADDRPOINTER_REG_0_ & n28822;
  assign n28833 = P1_STATE2_REG_2_ & n23831;
  assign n28834 = n23800 & ~n28833;
  assign n28835 = n24786 & n28834;
  assign n28836 = P1_STATE2_REG_2_ & ~n28835;
  assign n28837 = ~P1_STATE2_REG_2_ & P1_STATEBS16_REG;
  assign n28838 = P1_PHYADDRPOINTER_REG_0_ & n28837;
  assign n28839 = P1_STATE2_REG_2_ & n23800;
  assign n28840 = ~n26631 & ~n28839;
  assign n28841 = ~n24520 & ~n28840;
  assign n28842 = P1_EAX_REG_0_ & n28833;
  assign n28843 = P1_INSTQUEUERD_ADDR_REG_0_ & n28816;
  assign n28844 = P1_PHYADDRPOINTER_REG_0_ & n24584;
  assign n28845 = ~n28838 & ~n28841;
  assign n28846 = ~n28842 & n28845;
  assign n28847 = ~n28843 & n28846;
  assign n28848 = ~n28844 & n28847;
  assign n28849 = ~n24584 & ~n28848;
  assign n28850 = n24584 & n28848;
  assign n28851 = ~n28849 & ~n28850;
  assign n28852 = n28836 & ~n28851;
  assign n28853 = ~n28836 & n28851;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = ~n24584 & n28854;
  assign n28856 = n24584 & ~n28854;
  assign n28857 = ~n28855 & ~n28856;
  assign n28858 = P1_STATE2_REG_1_ & P1_STATEBS16_REG;
  assign n28859 = ~n28822 & n28858;
  assign n28860 = ~n28857 & n28859;
  assign n28861 = ~n28824 & ~n28829;
  assign n28862 = ~n28831 & n28861;
  assign n28863 = ~n28832 & n28862;
  assign n6249 = n28860 | ~n28863;
  assign n28865 = ~n26702 & n28823;
  assign n28866 = ~P1_PHYADDRPOINTER_REG_1_ & n28828;
  assign n28867 = P1_REIP_REG_1_ & n28830;
  assign n28868 = P1_PHYADDRPOINTER_REG_1_ & n28822;
  assign n28869 = ~n24782 & ~n28840;
  assign n28870 = P1_INSTQUEUERD_ADDR_REG_1_ & n28816;
  assign n28871 = ~P1_PHYADDRPOINTER_REG_1_ & n24584;
  assign n28872 = P1_EAX_REG_1_ & n28833;
  assign n28873 = P1_PHYADDRPOINTER_REG_1_ & n28837;
  assign n28874 = ~n28872 & ~n28873;
  assign n28875 = ~n24535 & ~n28840;
  assign n28876 = ~n28870 & ~n28871;
  assign n28877 = n28874 & n28876;
  assign n28878 = ~n28875 & n28877;
  assign n28879 = ~n24584 & ~n28878;
  assign n28880 = n24584 & n28878;
  assign n28881 = ~n28879 & ~n28880;
  assign n28882 = n28869 & ~n28881;
  assign n28883 = ~n28869 & n28881;
  assign n28884 = ~n28882 & ~n28883;
  assign n28885 = n24584 & ~n28853;
  assign n28886 = ~n28852 & ~n28885;
  assign n28887 = n28884 & n28886;
  assign n28888 = ~n28884 & ~n28886;
  assign n28889 = ~n28887 & ~n28888;
  assign n28890 = n28859 & ~n28889;
  assign n28891 = ~n28865 & ~n28866;
  assign n28892 = ~n28867 & n28891;
  assign n28893 = ~n28868 & n28892;
  assign n6254 = n28890 | ~n28893;
  assign n28895 = P1_REIP_REG_2_ & n28830;
  assign n28896 = P1_PHYADDRPOINTER_REG_1_ & ~P1_PHYADDRPOINTER_REG_2_;
  assign n28897 = ~P1_PHYADDRPOINTER_REG_1_ & P1_PHYADDRPOINTER_REG_2_;
  assign n28898 = ~n28896 & ~n28897;
  assign n28899 = n28828 & ~n28898;
  assign n28900 = ~n26751 & n28823;
  assign n28901 = P1_PHYADDRPOINTER_REG_2_ & n28822;
  assign n28902 = ~n28883 & ~n28886;
  assign n28903 = ~n28882 & ~n28902;
  assign n28904 = P1_INSTQUEUERD_ADDR_REG_2_ & n28816;
  assign n28905 = n24584 & ~n28898;
  assign n28906 = P1_EAX_REG_2_ & n28833;
  assign n28907 = P1_PHYADDRPOINTER_REG_2_ & n28837;
  assign n28908 = ~n28906 & ~n28907;
  assign n28909 = n24397 & ~n28840;
  assign n28910 = ~n28904 & ~n28905;
  assign n28911 = n28908 & n28910;
  assign n28912 = ~n28909 & n28911;
  assign n28913 = ~n24584 & ~n28912;
  assign n28914 = n24584 & n28912;
  assign n28915 = ~n24843 & ~n28840;
  assign n28916 = ~n28837 & ~n28915;
  assign n28917 = ~n28913 & ~n28914;
  assign n28918 = n28916 & n28917;
  assign n28919 = ~n28903 & ~n28918;
  assign n28920 = ~n28916 & ~n28917;
  assign n28921 = n28919 & ~n28920;
  assign n28922 = ~n28918 & ~n28920;
  assign n28923 = n28903 & ~n28922;
  assign n28924 = ~n28921 & ~n28923;
  assign n28925 = n28859 & n28924;
  assign n28926 = ~n28895 & ~n28899;
  assign n28927 = ~n28900 & n28926;
  assign n28928 = ~n28901 & n28927;
  assign n6259 = n28925 | ~n28928;
  assign n28930 = P1_REIP_REG_3_ & n28830;
  assign n28931 = P1_PHYADDRPOINTER_REG_1_ & P1_PHYADDRPOINTER_REG_2_;
  assign n28932 = ~P1_PHYADDRPOINTER_REG_3_ & n28931;
  assign n28933 = P1_PHYADDRPOINTER_REG_3_ & ~n28931;
  assign n28934 = ~n28932 & ~n28933;
  assign n28935 = n28828 & ~n28934;
  assign n28936 = ~n26828 & n28823;
  assign n28937 = P1_PHYADDRPOINTER_REG_3_ & n28822;
  assign n28938 = P1_INSTQUEUERD_ADDR_REG_3_ & n28816;
  assign n28939 = n24584 & ~n28934;
  assign n28940 = P1_EAX_REG_3_ & n28833;
  assign n28941 = P1_PHYADDRPOINTER_REG_3_ & n28837;
  assign n28942 = ~n28940 & ~n28941;
  assign n28943 = ~n24482 & ~n28840;
  assign n28944 = ~n28938 & ~n28939;
  assign n28945 = n28942 & n28944;
  assign n28946 = ~n28943 & n28945;
  assign n28947 = ~n24584 & ~n28946;
  assign n28948 = n24584 & n28946;
  assign n28949 = n24896 & ~n28840;
  assign n28950 = ~n28947 & ~n28948;
  assign n28951 = ~n28949 & n28950;
  assign n28952 = n28949 & ~n28950;
  assign n28953 = ~n28951 & ~n28952;
  assign n28954 = ~n28919 & ~n28920;
  assign n28955 = ~n28953 & n28954;
  assign n28956 = n28953 & ~n28954;
  assign n28957 = ~n28955 & ~n28956;
  assign n28958 = n28859 & n28957;
  assign n28959 = ~n28930 & ~n28935;
  assign n28960 = ~n28936 & n28959;
  assign n28961 = ~n28937 & n28960;
  assign n6264 = n28958 | ~n28961;
  assign n28963 = P1_REIP_REG_4_ & n28830;
  assign n28964 = P1_PHYADDRPOINTER_REG_3_ & n28931;
  assign n28965 = ~P1_PHYADDRPOINTER_REG_4_ & n28964;
  assign n28966 = P1_PHYADDRPOINTER_REG_4_ & ~n28964;
  assign n28967 = ~n28965 & ~n28966;
  assign n28968 = n28828 & ~n28967;
  assign n28969 = ~n26932 & n28823;
  assign n28970 = P1_PHYADDRPOINTER_REG_4_ & n28822;
  assign n28971 = P1_INSTQUEUERD_ADDR_REG_4_ & n28816;
  assign n28972 = n24584 & ~n28967;
  assign n28973 = P1_EAX_REG_4_ & n28833;
  assign n28974 = P1_PHYADDRPOINTER_REG_4_ & n28837;
  assign n28975 = ~n28973 & ~n28974;
  assign n28976 = ~n24472 & ~n28840;
  assign n28977 = ~n28971 & ~n28972;
  assign n28978 = n28975 & n28977;
  assign n28979 = ~n28976 & n28978;
  assign n28980 = ~n24584 & ~n28979;
  assign n28981 = n24584 & n28979;
  assign n28982 = ~n26924 & ~n28840;
  assign n28983 = ~n28980 & ~n28981;
  assign n28984 = ~n28982 & n28983;
  assign n28985 = n28982 & ~n28983;
  assign n28986 = ~n28984 & ~n28985;
  assign n28987 = ~n28918 & ~n28951;
  assign n28988 = ~n28853 & ~n28883;
  assign n28989 = ~n24584 & ~n28852;
  assign n28990 = n28988 & ~n28989;
  assign n28991 = ~n28882 & ~n28990;
  assign n28992 = ~n28920 & n28991;
  assign n28993 = n28987 & ~n28992;
  assign n28994 = ~n28952 & ~n28993;
  assign n28995 = n28986 & n28994;
  assign n28996 = ~n28986 & ~n28994;
  assign n28997 = ~n28995 & ~n28996;
  assign n28998 = n28859 & ~n28997;
  assign n28999 = ~n28963 & ~n28968;
  assign n29000 = ~n28969 & n28999;
  assign n29001 = ~n28970 & n29000;
  assign n6269 = n28998 | ~n29001;
  assign n29003 = P1_REIP_REG_5_ & n28830;
  assign n29004 = P1_PHYADDRPOINTER_REG_4_ & n28964;
  assign n29005 = ~P1_PHYADDRPOINTER_REG_5_ & n29004;
  assign n29006 = P1_PHYADDRPOINTER_REG_5_ & ~n29004;
  assign n29007 = ~n29005 & ~n29006;
  assign n29008 = n28828 & ~n29007;
  assign n29009 = n27041 & n28823;
  assign n29010 = P1_PHYADDRPOINTER_REG_5_ & n28822;
  assign n29011 = ~n27030 & ~n28840;
  assign n29012 = n24456 & n24469;
  assign n29013 = ~n28840 & n29012;
  assign n29014 = P1_EAX_REG_5_ & n28833;
  assign n29015 = n24584 & ~n29007;
  assign n29016 = P1_PHYADDRPOINTER_REG_5_ & n28837;
  assign n29017 = ~n29015 & ~n29016;
  assign n29018 = ~n29014 & n29017;
  assign n29019 = ~n29013 & n29018;
  assign n29020 = ~n24584 & ~n29019;
  assign n29021 = n24584 & n29019;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = n29011 & ~n29022;
  assign n29024 = ~n29011 & n29022;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = ~n28984 & ~n28994;
  assign n29027 = ~n28985 & ~n29026;
  assign n29028 = n29025 & n29027;
  assign n29029 = ~n29025 & ~n29027;
  assign n29030 = ~n29028 & ~n29029;
  assign n29031 = n28859 & ~n29030;
  assign n29032 = ~n29003 & ~n29008;
  assign n29033 = ~n29009 & n29032;
  assign n29034 = ~n29010 & n29033;
  assign n6274 = n29031 | ~n29034;
  assign n29036 = P1_REIP_REG_6_ & n28830;
  assign n29037 = P1_PHYADDRPOINTER_REG_5_ & n29004;
  assign n29038 = ~P1_PHYADDRPOINTER_REG_6_ & n29037;
  assign n29039 = P1_PHYADDRPOINTER_REG_6_ & ~n29037;
  assign n29040 = ~n29038 & ~n29039;
  assign n29041 = n28828 & ~n29040;
  assign n29042 = ~n27143 & n28823;
  assign n29043 = P1_PHYADDRPOINTER_REG_6_ & n28822;
  assign n29044 = ~n29024 & ~n29027;
  assign n29045 = ~n29023 & ~n29044;
  assign n29046 = P1_EAX_REG_6_ & n28833;
  assign n29047 = n24584 & ~n29040;
  assign n29048 = P1_PHYADDRPOINTER_REG_6_ & n28837;
  assign n29049 = ~n29047 & ~n29048;
  assign n29050 = ~n29046 & n29049;
  assign n29051 = ~n24584 & ~n29050;
  assign n29052 = n24584 & n29050;
  assign n29053 = n27131 & ~n28840;
  assign n29054 = ~n29051 & ~n29052;
  assign n29055 = ~n29053 & n29054;
  assign n29056 = ~n29045 & ~n29055;
  assign n29057 = n29053 & ~n29054;
  assign n29058 = n29056 & ~n29057;
  assign n29059 = ~n29055 & ~n29057;
  assign n29060 = n29045 & ~n29059;
  assign n29061 = ~n29058 & ~n29060;
  assign n29062 = n28859 & n29061;
  assign n29063 = ~n29036 & ~n29041;
  assign n29064 = ~n29042 & n29063;
  assign n29065 = ~n29043 & n29064;
  assign n6279 = n29062 | ~n29065;
  assign n29067 = P1_REIP_REG_7_ & n28830;
  assign n29068 = P1_PHYADDRPOINTER_REG_6_ & n29037;
  assign n29069 = ~P1_PHYADDRPOINTER_REG_7_ & n29068;
  assign n29070 = P1_PHYADDRPOINTER_REG_7_ & ~n29068;
  assign n29071 = ~n29069 & ~n29070;
  assign n29072 = n28828 & ~n29071;
  assign n29073 = n27225 & n28823;
  assign n29074 = P1_PHYADDRPOINTER_REG_7_ & n28822;
  assign n29075 = P1_EAX_REG_7_ & n28833;
  assign n29076 = n24584 & ~n29071;
  assign n29077 = P1_PHYADDRPOINTER_REG_7_ & n28837;
  assign n29078 = ~n29076 & ~n29077;
  assign n29079 = ~n29075 & n29078;
  assign n29080 = ~n24584 & ~n29079;
  assign n29081 = n24584 & n29079;
  assign n29082 = n27211 & ~n28840;
  assign n29083 = ~n29080 & ~n29081;
  assign n29084 = ~n29082 & n29083;
  assign n29085 = n29082 & ~n29083;
  assign n29086 = ~n29084 & ~n29085;
  assign n29087 = ~n29056 & ~n29057;
  assign n29088 = ~n29086 & n29087;
  assign n29089 = n29086 & ~n29087;
  assign n29090 = ~n29088 & ~n29089;
  assign n29091 = n28859 & n29090;
  assign n29092 = ~n29067 & ~n29072;
  assign n29093 = ~n29073 & n29092;
  assign n29094 = ~n29074 & n29093;
  assign n6284 = n29091 | ~n29094;
  assign n29096 = P1_REIP_REG_8_ & n28830;
  assign n29097 = P1_PHYADDRPOINTER_REG_7_ & n29068;
  assign n29098 = ~P1_PHYADDRPOINTER_REG_8_ & n29097;
  assign n29099 = P1_PHYADDRPOINTER_REG_8_ & ~n29097;
  assign n29100 = ~n29098 & ~n29099;
  assign n29101 = n28828 & ~n29100;
  assign n29102 = P1_PHYADDRPOINTER_REG_8_ & n28822;
  assign n29103 = ~n27344 & n28823;
  assign n29104 = P1_EAX_REG_8_ & n28833;
  assign n29105 = n24584 & ~n29100;
  assign n29106 = P1_PHYADDRPOINTER_REG_8_ & n28837;
  assign n29107 = ~n29105 & ~n29106;
  assign n29108 = ~n29104 & n29107;
  assign n29109 = ~n24584 & ~n29108;
  assign n29110 = n24584 & n29108;
  assign n29111 = n27336 & ~n28840;
  assign n29112 = ~n29109 & ~n29110;
  assign n29113 = ~n29111 & n29112;
  assign n29114 = n29111 & ~n29112;
  assign n29115 = ~n29113 & ~n29114;
  assign n29116 = ~n29024 & n29026;
  assign n29117 = ~n29055 & n29116;
  assign n29118 = ~n29084 & n29117;
  assign n29119 = n28985 & ~n29024;
  assign n29120 = ~n29023 & ~n29119;
  assign n29121 = ~n29057 & n29120;
  assign n29122 = ~n29055 & ~n29121;
  assign n29123 = ~n29084 & n29122;
  assign n29124 = ~n29085 & ~n29118;
  assign n29125 = ~n29123 & n29124;
  assign n29126 = n29115 & n29125;
  assign n29127 = ~n29115 & ~n29125;
  assign n29128 = ~n29126 & ~n29127;
  assign n29129 = n28859 & ~n29128;
  assign n29130 = ~n29096 & ~n29101;
  assign n29131 = ~n29102 & n29130;
  assign n29132 = ~n29103 & n29131;
  assign n6289 = n29129 | ~n29132;
  assign n29134 = P1_REIP_REG_9_ & n28830;
  assign n29135 = P1_PHYADDRPOINTER_REG_8_ & n29097;
  assign n29136 = ~P1_PHYADDRPOINTER_REG_9_ & n29135;
  assign n29137 = P1_PHYADDRPOINTER_REG_9_ & ~n29135;
  assign n29138 = ~n29136 & ~n29137;
  assign n29139 = n28828 & ~n29138;
  assign n29140 = P1_PHYADDRPOINTER_REG_9_ & n28822;
  assign n29141 = ~n27433 & n28823;
  assign n29142 = ~n27418 & ~n28840;
  assign n29143 = P1_EAX_REG_9_ & n28833;
  assign n29144 = n24584 & ~n29138;
  assign n29145 = P1_PHYADDRPOINTER_REG_9_ & n28837;
  assign n29146 = ~n29144 & ~n29145;
  assign n29147 = ~n29143 & n29146;
  assign n29148 = ~n24584 & ~n29147;
  assign n29149 = n24584 & n29147;
  assign n29150 = ~n29148 & ~n29149;
  assign n29151 = n29142 & ~n29150;
  assign n29152 = ~n29142 & n29150;
  assign n29153 = ~n29151 & ~n29152;
  assign n29154 = ~n29113 & ~n29125;
  assign n29155 = ~n29114 & ~n29154;
  assign n29156 = n29153 & n29155;
  assign n29157 = ~n29153 & ~n29155;
  assign n29158 = ~n29156 & ~n29157;
  assign n29159 = n28859 & ~n29158;
  assign n29160 = ~n29134 & ~n29139;
  assign n29161 = ~n29140 & n29160;
  assign n29162 = ~n29141 & n29161;
  assign n6294 = n29159 | ~n29162;
  assign n29164 = P1_REIP_REG_10_ & n28830;
  assign n29165 = P1_PHYADDRPOINTER_REG_9_ & n29135;
  assign n29166 = ~P1_PHYADDRPOINTER_REG_10_ & n29165;
  assign n29167 = P1_PHYADDRPOINTER_REG_10_ & ~n29165;
  assign n29168 = ~n29166 & ~n29167;
  assign n29169 = n28828 & ~n29168;
  assign n29170 = P1_PHYADDRPOINTER_REG_10_ & n28822;
  assign n29171 = ~n27521 & n28823;
  assign n29172 = ~n29152 & ~n29155;
  assign n29173 = ~n29151 & ~n29172;
  assign n29174 = P1_EAX_REG_10_ & n28833;
  assign n29175 = n24584 & ~n29168;
  assign n29176 = P1_PHYADDRPOINTER_REG_10_ & n28837;
  assign n29177 = ~n29175 & ~n29176;
  assign n29178 = ~n29174 & n29177;
  assign n29179 = ~n24584 & ~n29178;
  assign n29180 = n24584 & n29178;
  assign n29181 = ~n27511 & ~n28840;
  assign n29182 = ~n29179 & ~n29180;
  assign n29183 = ~n29181 & n29182;
  assign n29184 = ~n29173 & ~n29183;
  assign n29185 = n29181 & ~n29182;
  assign n29186 = n29184 & ~n29185;
  assign n29187 = ~n29183 & ~n29185;
  assign n29188 = n29173 & ~n29187;
  assign n29189 = ~n29186 & ~n29188;
  assign n29190 = n28859 & n29189;
  assign n29191 = ~n29164 & ~n29169;
  assign n29192 = ~n29170 & n29191;
  assign n29193 = ~n29171 & n29192;
  assign n6299 = n29190 | ~n29193;
  assign n29195 = P1_REIP_REG_11_ & n28830;
  assign n29196 = P1_PHYADDRPOINTER_REG_10_ & n29165;
  assign n29197 = ~P1_PHYADDRPOINTER_REG_11_ & n29196;
  assign n29198 = P1_PHYADDRPOINTER_REG_11_ & ~n29196;
  assign n29199 = ~n29197 & ~n29198;
  assign n29200 = n28828 & ~n29199;
  assign n29201 = P1_PHYADDRPOINTER_REG_11_ & n28822;
  assign n29202 = n27617 & n28823;
  assign n29203 = P1_EAX_REG_11_ & n28833;
  assign n29204 = P1_PHYADDRPOINTER_REG_11_ & n28837;
  assign n29205 = n24584 & ~n29199;
  assign n29206 = ~n29203 & ~n29204;
  assign n29207 = ~n29205 & n29206;
  assign n29208 = ~n24584 & ~n29207;
  assign n29209 = n24584 & n29207;
  assign n29210 = ~n29208 & ~n29209;
  assign n29211 = ~n27600 & ~n28840;
  assign n29212 = n29210 & ~n29211;
  assign n29213 = ~n29210 & n29211;
  assign n29214 = ~n29212 & ~n29213;
  assign n29215 = ~n29185 & ~n29214;
  assign n29216 = ~n29184 & n29215;
  assign n29217 = ~n29184 & ~n29185;
  assign n29218 = n29214 & ~n29217;
  assign n29219 = ~n29216 & ~n29218;
  assign n29220 = n28859 & n29219;
  assign n29221 = ~n29195 & ~n29200;
  assign n29222 = ~n29201 & n29221;
  assign n29223 = ~n29202 & n29222;
  assign n6304 = n29220 | ~n29223;
  assign n29225 = P1_REIP_REG_12_ & n28830;
  assign n29226 = P1_PHYADDRPOINTER_REG_11_ & n29196;
  assign n29227 = ~P1_PHYADDRPOINTER_REG_12_ & n29226;
  assign n29228 = P1_PHYADDRPOINTER_REG_12_ & ~n29226;
  assign n29229 = ~n29227 & ~n29228;
  assign n29230 = n28828 & ~n29229;
  assign n29231 = P1_PHYADDRPOINTER_REG_12_ & n28822;
  assign n29232 = ~n27703 & n28823;
  assign n29233 = ~n27695 & ~n28840;
  assign n29234 = P1_EAX_REG_12_ & n28833;
  assign n29235 = P1_PHYADDRPOINTER_REG_12_ & n28837;
  assign n29236 = n24584 & ~n29229;
  assign n29237 = ~n29234 & ~n29235;
  assign n29238 = ~n29236 & n29237;
  assign n29239 = ~n24584 & ~n29238;
  assign n29240 = n24584 & n29238;
  assign n29241 = ~n29239 & ~n29240;
  assign n29242 = n29233 & ~n29241;
  assign n29243 = ~n29233 & n29241;
  assign n29244 = ~n29242 & ~n29243;
  assign n29245 = ~n29113 & ~n29152;
  assign n29246 = ~n29183 & ~n29212;
  assign n29247 = ~n29125 & n29245;
  assign n29248 = n29246 & n29247;
  assign n29249 = n29152 & ~n29185;
  assign n29250 = ~n29114 & ~n29151;
  assign n29251 = ~n29185 & n29250;
  assign n29252 = ~n29212 & ~n29249;
  assign n29253 = ~n29251 & n29252;
  assign n29254 = ~n29183 & n29253;
  assign n29255 = ~n29213 & ~n29248;
  assign n29256 = ~n29254 & n29255;
  assign n29257 = n29244 & n29256;
  assign n29258 = ~n29244 & ~n29256;
  assign n29259 = ~n29257 & ~n29258;
  assign n29260 = n28859 & ~n29259;
  assign n29261 = ~n29225 & ~n29230;
  assign n29262 = ~n29231 & n29261;
  assign n29263 = ~n29232 & n29262;
  assign n6309 = n29260 | ~n29263;
  assign n29265 = P1_REIP_REG_13_ & n28830;
  assign n29266 = P1_PHYADDRPOINTER_REG_12_ & n29226;
  assign n29267 = ~P1_PHYADDRPOINTER_REG_13_ & n29266;
  assign n29268 = P1_PHYADDRPOINTER_REG_13_ & ~n29266;
  assign n29269 = ~n29267 & ~n29268;
  assign n29270 = n28828 & ~n29269;
  assign n29271 = P1_PHYADDRPOINTER_REG_13_ & n28822;
  assign n29272 = ~n27789 & n28823;
  assign n29273 = ~n27779 & ~n28840;
  assign n29274 = P1_EAX_REG_13_ & n28833;
  assign n29275 = P1_PHYADDRPOINTER_REG_13_ & n28837;
  assign n29276 = n24584 & ~n29269;
  assign n29277 = ~n29274 & ~n29275;
  assign n29278 = ~n29276 & n29277;
  assign n29279 = ~n24584 & ~n29278;
  assign n29280 = n24584 & n29278;
  assign n29281 = ~n29279 & ~n29280;
  assign n29282 = n29273 & ~n29281;
  assign n29283 = ~n29273 & n29281;
  assign n29284 = ~n29282 & ~n29283;
  assign n29285 = ~n29243 & ~n29256;
  assign n29286 = ~n29242 & ~n29285;
  assign n29287 = n29284 & n29286;
  assign n29288 = ~n29284 & ~n29286;
  assign n29289 = ~n29287 & ~n29288;
  assign n29290 = n28859 & ~n29289;
  assign n29291 = ~n29265 & ~n29270;
  assign n29292 = ~n29271 & n29291;
  assign n29293 = ~n29272 & n29292;
  assign n6314 = n29290 | ~n29293;
  assign n29295 = P1_REIP_REG_14_ & n28830;
  assign n29296 = P1_PHYADDRPOINTER_REG_13_ & n29266;
  assign n29297 = ~P1_PHYADDRPOINTER_REG_14_ & n29296;
  assign n29298 = P1_PHYADDRPOINTER_REG_14_ & ~n29296;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = n28828 & ~n29299;
  assign n29301 = P1_PHYADDRPOINTER_REG_14_ & n28822;
  assign n29302 = ~n27877 & n28823;
  assign n29303 = ~n29283 & ~n29286;
  assign n29304 = ~n29282 & ~n29303;
  assign n29305 = P1_EAX_REG_14_ & n28833;
  assign n29306 = P1_PHYADDRPOINTER_REG_14_ & n28837;
  assign n29307 = n24584 & ~n29299;
  assign n29308 = ~n29305 & ~n29306;
  assign n29309 = ~n29307 & n29308;
  assign n29310 = ~n24584 & ~n29309;
  assign n29311 = n24584 & n29309;
  assign n29312 = ~n27865 & ~n28840;
  assign n29313 = ~n29310 & ~n29311;
  assign n29314 = ~n29312 & n29313;
  assign n29315 = ~n29304 & ~n29314;
  assign n29316 = n29312 & ~n29313;
  assign n29317 = n29315 & ~n29316;
  assign n29318 = ~n29314 & ~n29316;
  assign n29319 = n29304 & ~n29318;
  assign n29320 = ~n29317 & ~n29319;
  assign n29321 = n28859 & n29320;
  assign n29322 = ~n29295 & ~n29300;
  assign n29323 = ~n29301 & n29322;
  assign n29324 = ~n29302 & n29323;
  assign n6319 = n29321 | ~n29324;
  assign n29326 = P1_REIP_REG_15_ & n28830;
  assign n29327 = P1_PHYADDRPOINTER_REG_14_ & n29296;
  assign n29328 = ~P1_PHYADDRPOINTER_REG_15_ & n29327;
  assign n29329 = P1_PHYADDRPOINTER_REG_15_ & ~n29327;
  assign n29330 = ~n29328 & ~n29329;
  assign n29331 = n28828 & ~n29330;
  assign n29332 = P1_PHYADDRPOINTER_REG_15_ & n28822;
  assign n29333 = n27967 & n28823;
  assign n29334 = P1_EAX_REG_15_ & n28833;
  assign n29335 = P1_PHYADDRPOINTER_REG_15_ & n28837;
  assign n29336 = n24584 & ~n29330;
  assign n29337 = ~n29334 & ~n29335;
  assign n29338 = ~n29336 & n29337;
  assign n29339 = ~n24584 & ~n29338;
  assign n29340 = n24584 & n29338;
  assign n29341 = ~n29339 & ~n29340;
  assign n29342 = ~n27952 & ~n28840;
  assign n29343 = n29341 & ~n29342;
  assign n29344 = ~n29341 & n29342;
  assign n29345 = ~n29343 & ~n29344;
  assign n29346 = ~n29316 & ~n29345;
  assign n29347 = ~n29315 & n29346;
  assign n29348 = ~n29315 & ~n29316;
  assign n29349 = n29345 & ~n29348;
  assign n29350 = ~n29347 & ~n29349;
  assign n29351 = n28859 & n29350;
  assign n29352 = ~n29326 & ~n29331;
  assign n29353 = ~n29332 & n29352;
  assign n29354 = ~n29333 & n29353;
  assign n6324 = n29351 | ~n29354;
  assign n29356 = P1_REIP_REG_16_ & n28830;
  assign n29357 = P1_PHYADDRPOINTER_REG_15_ & n29327;
  assign n29358 = ~P1_PHYADDRPOINTER_REG_16_ & n29357;
  assign n29359 = P1_PHYADDRPOINTER_REG_16_ & ~n29357;
  assign n29360 = ~n29358 & ~n29359;
  assign n29361 = n28828 & ~n29360;
  assign n29362 = P1_PHYADDRPOINTER_REG_16_ & n28822;
  assign n29363 = ~n28028 & n28823;
  assign n29364 = ~n28021 & ~n28840;
  assign n29365 = P1_INSTQUEUERD_ADDR_REG_2_ & ~n23624;
  assign n29366 = ~P1_INSTQUEUERD_ADDR_REG_3_ & n29365;
  assign n29367 = P1_INSTQUEUERD_ADDR_REG_3_ & ~n29365;
  assign n29368 = ~n29366 & ~n29367;
  assign n29369 = ~n23638 & ~n29365;
  assign n29370 = n29368 & n29369;
  assign n29371 = n24632 & n29370;
  assign n29372 = P1_INSTQUEUE_REG_7__0_ & n29371;
  assign n29373 = n24629 & n29370;
  assign n29374 = P1_INSTQUEUE_REG_6__0_ & n29373;
  assign n29375 = n24638 & n29370;
  assign n29376 = P1_INSTQUEUE_REG_5__0_ & n29375;
  assign n29377 = n24635 & n29370;
  assign n29378 = P1_INSTQUEUE_REG_4__0_ & n29377;
  assign n29379 = ~n29372 & ~n29374;
  assign n29380 = ~n29376 & n29379;
  assign n29381 = ~n29378 & n29380;
  assign n29382 = n29368 & ~n29369;
  assign n29383 = n24632 & n29382;
  assign n29384 = P1_INSTQUEUE_REG_3__0_ & n29383;
  assign n29385 = n24629 & n29382;
  assign n29386 = P1_INSTQUEUE_REG_2__0_ & n29385;
  assign n29387 = n24638 & n29382;
  assign n29388 = P1_INSTQUEUE_REG_1__0_ & n29387;
  assign n29389 = n24635 & n29382;
  assign n29390 = P1_INSTQUEUE_REG_0__0_ & n29389;
  assign n29391 = ~n29384 & ~n29386;
  assign n29392 = ~n29388 & n29391;
  assign n29393 = ~n29390 & n29392;
  assign n29394 = ~n29368 & n29369;
  assign n29395 = n24632 & n29394;
  assign n29396 = P1_INSTQUEUE_REG_15__0_ & n29395;
  assign n29397 = n24629 & n29394;
  assign n29398 = P1_INSTQUEUE_REG_14__0_ & n29397;
  assign n29399 = n24638 & n29394;
  assign n29400 = P1_INSTQUEUE_REG_13__0_ & n29399;
  assign n29401 = n24635 & n29394;
  assign n29402 = P1_INSTQUEUE_REG_12__0_ & n29401;
  assign n29403 = ~n29396 & ~n29398;
  assign n29404 = ~n29400 & n29403;
  assign n29405 = ~n29402 & n29404;
  assign n29406 = ~n29368 & ~n29369;
  assign n29407 = n24632 & n29406;
  assign n29408 = P1_INSTQUEUE_REG_11__0_ & n29407;
  assign n29409 = n24629 & n29406;
  assign n29410 = P1_INSTQUEUE_REG_10__0_ & n29409;
  assign n29411 = n24638 & n29406;
  assign n29412 = P1_INSTQUEUE_REG_9__0_ & n29411;
  assign n29413 = n24635 & n29406;
  assign n29414 = P1_INSTQUEUE_REG_8__0_ & n29413;
  assign n29415 = ~n29408 & ~n29410;
  assign n29416 = ~n29412 & n29415;
  assign n29417 = ~n29414 & n29416;
  assign n29418 = n29381 & n29393;
  assign n29419 = n29405 & n29418;
  assign n29420 = n29417 & n29419;
  assign n29421 = P1_STATE2_REG_0_ & n24168;
  assign n29422 = n24003 & n24046;
  assign n29423 = ~n29421 & ~n29422;
  assign n29424 = ~n29420 & ~n29423;
  assign n29425 = ~n28840 & n29424;
  assign n29426 = P1_EAX_REG_16_ & n28833;
  assign n29427 = P1_PHYADDRPOINTER_REG_16_ & n28837;
  assign n29428 = n24584 & ~n29360;
  assign n29429 = ~n29426 & ~n29427;
  assign n29430 = ~n29428 & n29429;
  assign n29431 = ~n29425 & n29430;
  assign n29432 = ~n24584 & ~n29431;
  assign n29433 = n24584 & n29431;
  assign n29434 = ~n29432 & ~n29433;
  assign n29435 = n29364 & ~n29434;
  assign n29436 = ~n29364 & n29434;
  assign n29437 = ~n29435 & ~n29436;
  assign n29438 = ~n29243 & ~n29283;
  assign n29439 = ~n29314 & n29438;
  assign n29440 = ~n29343 & n29439;
  assign n29441 = ~n29256 & n29440;
  assign n29442 = n29242 & ~n29283;
  assign n29443 = ~n29314 & n29442;
  assign n29444 = ~n29343 & n29443;
  assign n29445 = n29316 & ~n29343;
  assign n29446 = n29282 & ~n29314;
  assign n29447 = ~n29343 & n29446;
  assign n29448 = ~n29344 & ~n29444;
  assign n29449 = ~n29445 & n29448;
  assign n29450 = ~n29447 & n29449;
  assign n29451 = ~n29441 & n29450;
  assign n29452 = n29437 & n29451;
  assign n29453 = ~n29437 & ~n29451;
  assign n29454 = ~n29452 & ~n29453;
  assign n29455 = n28859 & ~n29454;
  assign n29456 = ~n29356 & ~n29361;
  assign n29457 = ~n29362 & n29456;
  assign n29458 = ~n29363 & n29457;
  assign n6329 = n29455 | ~n29458;
  assign n29460 = P1_REIP_REG_17_ & n28830;
  assign n29461 = P1_PHYADDRPOINTER_REG_16_ & n29357;
  assign n29462 = ~P1_PHYADDRPOINTER_REG_17_ & n29461;
  assign n29463 = P1_PHYADDRPOINTER_REG_17_ & ~n29461;
  assign n29464 = ~n29462 & ~n29463;
  assign n29465 = n28828 & ~n29464;
  assign n29466 = P1_PHYADDRPOINTER_REG_17_ & n28822;
  assign n29467 = ~n28075 & n28823;
  assign n29468 = n28019 & ~n28840;
  assign n29469 = P1_INSTQUEUE_REG_7__1_ & n29371;
  assign n29470 = P1_INSTQUEUE_REG_6__1_ & n29373;
  assign n29471 = P1_INSTQUEUE_REG_5__1_ & n29375;
  assign n29472 = P1_INSTQUEUE_REG_4__1_ & n29377;
  assign n29473 = ~n29469 & ~n29470;
  assign n29474 = ~n29471 & n29473;
  assign n29475 = ~n29472 & n29474;
  assign n29476 = P1_INSTQUEUE_REG_3__1_ & n29383;
  assign n29477 = P1_INSTQUEUE_REG_2__1_ & n29385;
  assign n29478 = P1_INSTQUEUE_REG_1__1_ & n29387;
  assign n29479 = P1_INSTQUEUE_REG_0__1_ & n29389;
  assign n29480 = ~n29476 & ~n29477;
  assign n29481 = ~n29478 & n29480;
  assign n29482 = ~n29479 & n29481;
  assign n29483 = P1_INSTQUEUE_REG_15__1_ & n29395;
  assign n29484 = P1_INSTQUEUE_REG_14__1_ & n29397;
  assign n29485 = P1_INSTQUEUE_REG_13__1_ & n29399;
  assign n29486 = P1_INSTQUEUE_REG_12__1_ & n29401;
  assign n29487 = ~n29483 & ~n29484;
  assign n29488 = ~n29485 & n29487;
  assign n29489 = ~n29486 & n29488;
  assign n29490 = P1_INSTQUEUE_REG_11__1_ & n29407;
  assign n29491 = P1_INSTQUEUE_REG_10__1_ & n29409;
  assign n29492 = P1_INSTQUEUE_REG_9__1_ & n29411;
  assign n29493 = P1_INSTQUEUE_REG_8__1_ & n29413;
  assign n29494 = ~n29490 & ~n29491;
  assign n29495 = ~n29492 & n29494;
  assign n29496 = ~n29493 & n29495;
  assign n29497 = n29475 & n29482;
  assign n29498 = n29489 & n29497;
  assign n29499 = n29496 & n29498;
  assign n29500 = ~n29423 & ~n29499;
  assign n29501 = ~n28840 & n29500;
  assign n29502 = P1_EAX_REG_17_ & n28833;
  assign n29503 = P1_PHYADDRPOINTER_REG_17_ & n28837;
  assign n29504 = n24584 & ~n29464;
  assign n29505 = ~n29502 & ~n29503;
  assign n29506 = ~n29504 & n29505;
  assign n29507 = ~n29501 & n29506;
  assign n29508 = ~n24584 & ~n29507;
  assign n29509 = n24584 & n29507;
  assign n29510 = ~n29508 & ~n29509;
  assign n29511 = n29468 & ~n29510;
  assign n29512 = ~n29468 & n29510;
  assign n29513 = ~n29511 & ~n29512;
  assign n29514 = ~n29436 & ~n29451;
  assign n29515 = ~n29435 & ~n29514;
  assign n29516 = n29513 & n29515;
  assign n29517 = ~n29513 & ~n29515;
  assign n29518 = ~n29516 & ~n29517;
  assign n29519 = n28859 & ~n29518;
  assign n29520 = ~n29460 & ~n29465;
  assign n29521 = ~n29466 & n29520;
  assign n29522 = ~n29467 & n29521;
  assign n6334 = n29519 | ~n29522;
  assign n29524 = P1_REIP_REG_18_ & n28830;
  assign n29525 = P1_PHYADDRPOINTER_REG_17_ & n29461;
  assign n29526 = ~P1_PHYADDRPOINTER_REG_18_ & n29525;
  assign n29527 = P1_PHYADDRPOINTER_REG_18_ & ~n29525;
  assign n29528 = ~n29526 & ~n29527;
  assign n29529 = n28828 & ~n29528;
  assign n29530 = P1_PHYADDRPOINTER_REG_18_ & n28822;
  assign n29531 = ~n28124 & n28823;
  assign n29532 = P1_INSTQUEUE_REG_7__2_ & n29371;
  assign n29533 = P1_INSTQUEUE_REG_6__2_ & n29373;
  assign n29534 = P1_INSTQUEUE_REG_5__2_ & n29375;
  assign n29535 = P1_INSTQUEUE_REG_4__2_ & n29377;
  assign n29536 = ~n29532 & ~n29533;
  assign n29537 = ~n29534 & n29536;
  assign n29538 = ~n29535 & n29537;
  assign n29539 = P1_INSTQUEUE_REG_3__2_ & n29383;
  assign n29540 = P1_INSTQUEUE_REG_2__2_ & n29385;
  assign n29541 = P1_INSTQUEUE_REG_1__2_ & n29387;
  assign n29542 = P1_INSTQUEUE_REG_0__2_ & n29389;
  assign n29543 = ~n29539 & ~n29540;
  assign n29544 = ~n29541 & n29543;
  assign n29545 = ~n29542 & n29544;
  assign n29546 = P1_INSTQUEUE_REG_15__2_ & n29395;
  assign n29547 = P1_INSTQUEUE_REG_14__2_ & n29397;
  assign n29548 = P1_INSTQUEUE_REG_13__2_ & n29399;
  assign n29549 = P1_INSTQUEUE_REG_12__2_ & n29401;
  assign n29550 = ~n29546 & ~n29547;
  assign n29551 = ~n29548 & n29550;
  assign n29552 = ~n29549 & n29551;
  assign n29553 = P1_INSTQUEUE_REG_11__2_ & n29407;
  assign n29554 = P1_INSTQUEUE_REG_10__2_ & n29409;
  assign n29555 = P1_INSTQUEUE_REG_9__2_ & n29411;
  assign n29556 = P1_INSTQUEUE_REG_8__2_ & n29413;
  assign n29557 = ~n29553 & ~n29554;
  assign n29558 = ~n29555 & n29557;
  assign n29559 = ~n29556 & n29558;
  assign n29560 = n29538 & n29545;
  assign n29561 = n29552 & n29560;
  assign n29562 = n29559 & n29561;
  assign n29563 = ~n29423 & ~n29562;
  assign n29564 = ~n28840 & n29563;
  assign n29565 = P1_EAX_REG_18_ & n28833;
  assign n29566 = P1_PHYADDRPOINTER_REG_18_ & n28837;
  assign n29567 = n24584 & ~n29528;
  assign n29568 = ~n29565 & ~n29566;
  assign n29569 = ~n29567 & n29568;
  assign n29570 = ~n29564 & n29569;
  assign n29571 = ~n24584 & ~n29570;
  assign n29572 = n24584 & n29570;
  assign n29573 = ~n29571 & ~n29572;
  assign n29574 = n29468 & ~n29573;
  assign n29575 = ~n29468 & n29573;
  assign n29576 = ~n29574 & ~n29575;
  assign n29577 = n29435 & ~n29512;
  assign n29578 = ~n29511 & ~n29577;
  assign n29579 = ~n29436 & ~n29512;
  assign n29580 = ~n29451 & n29579;
  assign n29581 = n29578 & ~n29580;
  assign n29582 = n29576 & n29581;
  assign n29583 = ~n29576 & ~n29581;
  assign n29584 = ~n29582 & ~n29583;
  assign n29585 = n28859 & ~n29584;
  assign n29586 = ~n29524 & ~n29529;
  assign n29587 = ~n29530 & n29586;
  assign n29588 = ~n29531 & n29587;
  assign n6339 = n29585 | ~n29588;
  assign n29590 = P1_REIP_REG_19_ & n28830;
  assign n29591 = P1_PHYADDRPOINTER_REG_18_ & n29525;
  assign n29592 = ~P1_PHYADDRPOINTER_REG_19_ & n29591;
  assign n29593 = P1_PHYADDRPOINTER_REG_19_ & ~n29591;
  assign n29594 = ~n29592 & ~n29593;
  assign n29595 = n28828 & ~n29594;
  assign n29596 = P1_PHYADDRPOINTER_REG_19_ & n28822;
  assign n29597 = ~n28174 & n28823;
  assign n29598 = P1_INSTQUEUE_REG_7__3_ & n29371;
  assign n29599 = P1_INSTQUEUE_REG_6__3_ & n29373;
  assign n29600 = P1_INSTQUEUE_REG_5__3_ & n29375;
  assign n29601 = P1_INSTQUEUE_REG_4__3_ & n29377;
  assign n29602 = ~n29598 & ~n29599;
  assign n29603 = ~n29600 & n29602;
  assign n29604 = ~n29601 & n29603;
  assign n29605 = P1_INSTQUEUE_REG_3__3_ & n29383;
  assign n29606 = P1_INSTQUEUE_REG_2__3_ & n29385;
  assign n29607 = P1_INSTQUEUE_REG_1__3_ & n29387;
  assign n29608 = P1_INSTQUEUE_REG_0__3_ & n29389;
  assign n29609 = ~n29605 & ~n29606;
  assign n29610 = ~n29607 & n29609;
  assign n29611 = ~n29608 & n29610;
  assign n29612 = P1_INSTQUEUE_REG_15__3_ & n29395;
  assign n29613 = P1_INSTQUEUE_REG_14__3_ & n29397;
  assign n29614 = P1_INSTQUEUE_REG_13__3_ & n29399;
  assign n29615 = P1_INSTQUEUE_REG_12__3_ & n29401;
  assign n29616 = ~n29612 & ~n29613;
  assign n29617 = ~n29614 & n29616;
  assign n29618 = ~n29615 & n29617;
  assign n29619 = P1_INSTQUEUE_REG_11__3_ & n29407;
  assign n29620 = P1_INSTQUEUE_REG_10__3_ & n29409;
  assign n29621 = P1_INSTQUEUE_REG_9__3_ & n29411;
  assign n29622 = P1_INSTQUEUE_REG_8__3_ & n29413;
  assign n29623 = ~n29619 & ~n29620;
  assign n29624 = ~n29621 & n29623;
  assign n29625 = ~n29622 & n29624;
  assign n29626 = n29604 & n29611;
  assign n29627 = n29618 & n29626;
  assign n29628 = n29625 & n29627;
  assign n29629 = ~n29423 & ~n29628;
  assign n29630 = ~n28840 & n29629;
  assign n29631 = P1_EAX_REG_19_ & n28833;
  assign n29632 = P1_PHYADDRPOINTER_REG_19_ & n28837;
  assign n29633 = n24584 & ~n29594;
  assign n29634 = ~n29631 & ~n29632;
  assign n29635 = ~n29633 & n29634;
  assign n29636 = ~n29630 & n29635;
  assign n29637 = ~n24584 & ~n29636;
  assign n29638 = n24584 & n29636;
  assign n29639 = ~n29637 & ~n29638;
  assign n29640 = n29468 & ~n29639;
  assign n29641 = ~n29468 & n29639;
  assign n29642 = ~n29640 & ~n29641;
  assign n29643 = ~n29575 & ~n29578;
  assign n29644 = ~n29574 & ~n29643;
  assign n29645 = ~n29575 & n29579;
  assign n29646 = ~n29451 & n29645;
  assign n29647 = n29644 & ~n29646;
  assign n29648 = n29642 & n29647;
  assign n29649 = ~n29642 & ~n29647;
  assign n29650 = ~n29648 & ~n29649;
  assign n29651 = n28859 & ~n29650;
  assign n29652 = ~n29590 & ~n29595;
  assign n29653 = ~n29596 & n29652;
  assign n29654 = ~n29597 & n29653;
  assign n6344 = n29651 | ~n29654;
  assign n29656 = P1_REIP_REG_20_ & n28830;
  assign n29657 = P1_PHYADDRPOINTER_REG_19_ & n29591;
  assign n29658 = ~P1_PHYADDRPOINTER_REG_20_ & n29657;
  assign n29659 = P1_PHYADDRPOINTER_REG_20_ & ~n29657;
  assign n29660 = ~n29658 & ~n29659;
  assign n29661 = n28828 & ~n29660;
  assign n29662 = P1_PHYADDRPOINTER_REG_20_ & n28822;
  assign n29663 = ~n28219 & n28823;
  assign n29664 = P1_INSTQUEUE_REG_0__4_ & n29389;
  assign n29665 = P1_INSTQUEUE_REG_7__4_ & n29371;
  assign n29666 = P1_INSTQUEUE_REG_6__4_ & n29373;
  assign n29667 = P1_INSTQUEUE_REG_5__4_ & n29375;
  assign n29668 = ~n29664 & ~n29665;
  assign n29669 = ~n29666 & n29668;
  assign n29670 = ~n29667 & n29669;
  assign n29671 = P1_INSTQUEUE_REG_4__4_ & n29377;
  assign n29672 = P1_INSTQUEUE_REG_3__4_ & n29383;
  assign n29673 = P1_INSTQUEUE_REG_2__4_ & n29385;
  assign n29674 = P1_INSTQUEUE_REG_1__4_ & n29387;
  assign n29675 = ~n29671 & ~n29672;
  assign n29676 = ~n29673 & n29675;
  assign n29677 = ~n29674 & n29676;
  assign n29678 = P1_INSTQUEUE_REG_15__4_ & n29395;
  assign n29679 = P1_INSTQUEUE_REG_14__4_ & n29397;
  assign n29680 = P1_INSTQUEUE_REG_13__4_ & n29399;
  assign n29681 = P1_INSTQUEUE_REG_12__4_ & n29401;
  assign n29682 = ~n29678 & ~n29679;
  assign n29683 = ~n29680 & n29682;
  assign n29684 = ~n29681 & n29683;
  assign n29685 = P1_INSTQUEUE_REG_11__4_ & n29407;
  assign n29686 = P1_INSTQUEUE_REG_10__4_ & n29409;
  assign n29687 = P1_INSTQUEUE_REG_9__4_ & n29411;
  assign n29688 = P1_INSTQUEUE_REG_8__4_ & n29413;
  assign n29689 = ~n29685 & ~n29686;
  assign n29690 = ~n29687 & n29689;
  assign n29691 = ~n29688 & n29690;
  assign n29692 = n29670 & n29677;
  assign n29693 = n29684 & n29692;
  assign n29694 = n29691 & n29693;
  assign n29695 = ~n29423 & ~n29694;
  assign n29696 = ~n28840 & n29695;
  assign n29697 = P1_EAX_REG_20_ & n28833;
  assign n29698 = P1_PHYADDRPOINTER_REG_20_ & n28837;
  assign n29699 = n24584 & ~n29660;
  assign n29700 = ~n29697 & ~n29698;
  assign n29701 = ~n29699 & n29700;
  assign n29702 = ~n29696 & n29701;
  assign n29703 = ~n24584 & ~n29702;
  assign n29704 = n24584 & n29702;
  assign n29705 = ~n29703 & ~n29704;
  assign n29706 = n29468 & ~n29705;
  assign n29707 = ~n29468 & n29705;
  assign n29708 = ~n29706 & ~n29707;
  assign n29709 = ~n29641 & ~n29647;
  assign n29710 = ~n29640 & ~n29709;
  assign n29711 = n29708 & n29710;
  assign n29712 = ~n29708 & ~n29710;
  assign n29713 = ~n29711 & ~n29712;
  assign n29714 = n28859 & ~n29713;
  assign n29715 = ~n29656 & ~n29661;
  assign n29716 = ~n29662 & n29715;
  assign n29717 = ~n29663 & n29716;
  assign n6349 = n29714 | ~n29717;
  assign n29719 = P1_REIP_REG_21_ & n28830;
  assign n29720 = P1_PHYADDRPOINTER_REG_20_ & n29657;
  assign n29721 = ~P1_PHYADDRPOINTER_REG_21_ & n29720;
  assign n29722 = P1_PHYADDRPOINTER_REG_21_ & ~n29720;
  assign n29723 = ~n29721 & ~n29722;
  assign n29724 = n28828 & ~n29723;
  assign n29725 = P1_PHYADDRPOINTER_REG_21_ & n28822;
  assign n29726 = ~n28268 & n28823;
  assign n29727 = P1_INSTQUEUE_REG_7__5_ & n29371;
  assign n29728 = P1_INSTQUEUE_REG_6__5_ & n29373;
  assign n29729 = P1_INSTQUEUE_REG_5__5_ & n29375;
  assign n29730 = P1_INSTQUEUE_REG_4__5_ & n29377;
  assign n29731 = ~n29727 & ~n29728;
  assign n29732 = ~n29729 & n29731;
  assign n29733 = ~n29730 & n29732;
  assign n29734 = P1_INSTQUEUE_REG_3__5_ & n29383;
  assign n29735 = P1_INSTQUEUE_REG_2__5_ & n29385;
  assign n29736 = P1_INSTQUEUE_REG_1__5_ & n29387;
  assign n29737 = P1_INSTQUEUE_REG_0__5_ & n29389;
  assign n29738 = ~n29734 & ~n29735;
  assign n29739 = ~n29736 & n29738;
  assign n29740 = ~n29737 & n29739;
  assign n29741 = P1_INSTQUEUE_REG_15__5_ & n29395;
  assign n29742 = P1_INSTQUEUE_REG_14__5_ & n29397;
  assign n29743 = P1_INSTQUEUE_REG_13__5_ & n29399;
  assign n29744 = P1_INSTQUEUE_REG_12__5_ & n29401;
  assign n29745 = ~n29741 & ~n29742;
  assign n29746 = ~n29743 & n29745;
  assign n29747 = ~n29744 & n29746;
  assign n29748 = P1_INSTQUEUE_REG_11__5_ & n29407;
  assign n29749 = P1_INSTQUEUE_REG_10__5_ & n29409;
  assign n29750 = P1_INSTQUEUE_REG_9__5_ & n29411;
  assign n29751 = P1_INSTQUEUE_REG_8__5_ & n29413;
  assign n29752 = ~n29748 & ~n29749;
  assign n29753 = ~n29750 & n29752;
  assign n29754 = ~n29751 & n29753;
  assign n29755 = n29733 & n29740;
  assign n29756 = n29747 & n29755;
  assign n29757 = n29754 & n29756;
  assign n29758 = ~n29423 & ~n29757;
  assign n29759 = ~n28840 & n29758;
  assign n29760 = P1_EAX_REG_21_ & n28833;
  assign n29761 = P1_PHYADDRPOINTER_REG_21_ & n28837;
  assign n29762 = n24584 & ~n29723;
  assign n29763 = ~n29760 & ~n29761;
  assign n29764 = ~n29762 & n29763;
  assign n29765 = ~n29759 & n29764;
  assign n29766 = ~n24584 & ~n29765;
  assign n29767 = n24584 & n29765;
  assign n29768 = ~n29766 & ~n29767;
  assign n29769 = n29468 & ~n29768;
  assign n29770 = ~n29468 & n29768;
  assign n29771 = ~n29769 & ~n29770;
  assign n29772 = n29640 & ~n29707;
  assign n29773 = ~n29706 & ~n29772;
  assign n29774 = ~n29641 & ~n29707;
  assign n29775 = ~n29647 & n29774;
  assign n29776 = n29773 & ~n29775;
  assign n29777 = n29771 & n29776;
  assign n29778 = ~n29771 & ~n29776;
  assign n29779 = ~n29777 & ~n29778;
  assign n29780 = n28859 & ~n29779;
  assign n29781 = ~n29719 & ~n29724;
  assign n29782 = ~n29725 & n29781;
  assign n29783 = ~n29726 & n29782;
  assign n6354 = n29780 | ~n29783;
  assign n29785 = P1_REIP_REG_22_ & n28830;
  assign n29786 = P1_PHYADDRPOINTER_REG_21_ & n29720;
  assign n29787 = ~P1_PHYADDRPOINTER_REG_22_ & n29786;
  assign n29788 = P1_PHYADDRPOINTER_REG_22_ & ~n29786;
  assign n29789 = ~n29787 & ~n29788;
  assign n29790 = n28828 & ~n29789;
  assign n29791 = P1_PHYADDRPOINTER_REG_22_ & n28822;
  assign n29792 = ~n28316 & n28823;
  assign n29793 = P1_INSTQUEUE_REG_7__6_ & n29371;
  assign n29794 = P1_INSTQUEUE_REG_6__6_ & n29373;
  assign n29795 = P1_INSTQUEUE_REG_5__6_ & n29375;
  assign n29796 = P1_INSTQUEUE_REG_4__6_ & n29377;
  assign n29797 = ~n29793 & ~n29794;
  assign n29798 = ~n29795 & n29797;
  assign n29799 = ~n29796 & n29798;
  assign n29800 = P1_INSTQUEUE_REG_3__6_ & n29383;
  assign n29801 = P1_INSTQUEUE_REG_2__6_ & n29385;
  assign n29802 = P1_INSTQUEUE_REG_1__6_ & n29387;
  assign n29803 = P1_INSTQUEUE_REG_0__6_ & n29389;
  assign n29804 = ~n29800 & ~n29801;
  assign n29805 = ~n29802 & n29804;
  assign n29806 = ~n29803 & n29805;
  assign n29807 = P1_INSTQUEUE_REG_15__6_ & n29395;
  assign n29808 = P1_INSTQUEUE_REG_14__6_ & n29397;
  assign n29809 = P1_INSTQUEUE_REG_13__6_ & n29399;
  assign n29810 = P1_INSTQUEUE_REG_12__6_ & n29401;
  assign n29811 = ~n29807 & ~n29808;
  assign n29812 = ~n29809 & n29811;
  assign n29813 = ~n29810 & n29812;
  assign n29814 = P1_INSTQUEUE_REG_11__6_ & n29407;
  assign n29815 = P1_INSTQUEUE_REG_10__6_ & n29409;
  assign n29816 = P1_INSTQUEUE_REG_9__6_ & n29411;
  assign n29817 = P1_INSTQUEUE_REG_8__6_ & n29413;
  assign n29818 = ~n29814 & ~n29815;
  assign n29819 = ~n29816 & n29818;
  assign n29820 = ~n29817 & n29819;
  assign n29821 = n29799 & n29806;
  assign n29822 = n29813 & n29821;
  assign n29823 = n29820 & n29822;
  assign n29824 = ~n29423 & ~n29823;
  assign n29825 = ~n28840 & n29824;
  assign n29826 = P1_EAX_REG_22_ & n28833;
  assign n29827 = P1_PHYADDRPOINTER_REG_22_ & n28837;
  assign n29828 = n24584 & ~n29789;
  assign n29829 = ~n29826 & ~n29827;
  assign n29830 = ~n29828 & n29829;
  assign n29831 = ~n29825 & n29830;
  assign n29832 = ~n24584 & ~n29831;
  assign n29833 = n24584 & n29831;
  assign n29834 = ~n29832 & ~n29833;
  assign n29835 = n29468 & ~n29834;
  assign n29836 = ~n29468 & n29834;
  assign n29837 = ~n29835 & ~n29836;
  assign n29838 = ~n29770 & ~n29773;
  assign n29839 = ~n29769 & ~n29838;
  assign n29840 = ~n29770 & n29774;
  assign n29841 = ~n29647 & n29840;
  assign n29842 = n29839 & ~n29841;
  assign n29843 = n29837 & n29842;
  assign n29844 = ~n29837 & ~n29842;
  assign n29845 = ~n29843 & ~n29844;
  assign n29846 = n28859 & ~n29845;
  assign n29847 = ~n29785 & ~n29790;
  assign n29848 = ~n29791 & n29847;
  assign n29849 = ~n29792 & n29848;
  assign n6359 = n29846 | ~n29849;
  assign n29851 = P1_REIP_REG_23_ & n28830;
  assign n29852 = P1_PHYADDRPOINTER_REG_22_ & n29786;
  assign n29853 = ~P1_PHYADDRPOINTER_REG_23_ & n29852;
  assign n29854 = P1_PHYADDRPOINTER_REG_23_ & ~n29852;
  assign n29855 = ~n29853 & ~n29854;
  assign n29856 = n28828 & ~n29855;
  assign n29857 = P1_PHYADDRPOINTER_REG_23_ & n28822;
  assign n29858 = ~n28373 & n28823;
  assign n29859 = P1_INSTQUEUERD_ADDR_REG_3_ & ~P1_INSTQUEUERD_ADDR_REG_2_;
  assign n29860 = ~n23652 & ~n29859;
  assign n29861 = n23856 & n29860;
  assign n29862 = P1_INSTQUEUE_REG_7__0_ & n29861;
  assign n29863 = n23860 & n29860;
  assign n29864 = P1_INSTQUEUE_REG_6__0_ & n29863;
  assign n29865 = P1_INSTQUEUERD_ADDR_REG_0_ & n23635;
  assign n29866 = n29860 & n29865;
  assign n29867 = P1_INSTQUEUE_REG_5__0_ & n29866;
  assign n29868 = n23638 & n29860;
  assign n29869 = P1_INSTQUEUE_REG_4__0_ & n29868;
  assign n29870 = ~n29862 & ~n29864;
  assign n29871 = ~n29867 & n29870;
  assign n29872 = ~n29869 & n29871;
  assign n29873 = P1_INSTQUEUERD_ADDR_REG_2_ & n29860;
  assign n29874 = n23655 & n29873;
  assign n29875 = P1_INSTQUEUE_REG_3__0_ & n29874;
  assign n29876 = n23662 & n29873;
  assign n29877 = P1_INSTQUEUE_REG_2__0_ & n29876;
  assign n29878 = n23665 & n29873;
  assign n29879 = P1_INSTQUEUE_REG_1__0_ & n29878;
  assign n29880 = n23624 & n29873;
  assign n29881 = P1_INSTQUEUE_REG_0__0_ & n29880;
  assign n29882 = ~n29875 & ~n29877;
  assign n29883 = ~n29879 & n29882;
  assign n29884 = ~n29881 & n29883;
  assign n29885 = n23856 & ~n29860;
  assign n29886 = P1_INSTQUEUE_REG_15__0_ & n29885;
  assign n29887 = n23860 & ~n29860;
  assign n29888 = P1_INSTQUEUE_REG_14__0_ & n29887;
  assign n29889 = ~n29860 & n29865;
  assign n29890 = P1_INSTQUEUE_REG_13__0_ & n29889;
  assign n29891 = n23638 & ~n29860;
  assign n29892 = P1_INSTQUEUE_REG_12__0_ & n29891;
  assign n29893 = ~n29886 & ~n29888;
  assign n29894 = ~n29890 & n29893;
  assign n29895 = ~n29892 & n29894;
  assign n29896 = P1_INSTQUEUERD_ADDR_REG_2_ & ~n29860;
  assign n29897 = n23655 & n29896;
  assign n29898 = P1_INSTQUEUE_REG_11__0_ & n29897;
  assign n29899 = n23662 & n29896;
  assign n29900 = P1_INSTQUEUE_REG_10__0_ & n29899;
  assign n29901 = n23665 & n29896;
  assign n29902 = P1_INSTQUEUE_REG_9__0_ & n29901;
  assign n29903 = n23624 & n29896;
  assign n29904 = P1_INSTQUEUE_REG_8__0_ & n29903;
  assign n29905 = ~n29898 & ~n29900;
  assign n29906 = ~n29902 & n29905;
  assign n29907 = ~n29904 & n29906;
  assign n29908 = n29872 & n29884;
  assign n29909 = n29895 & n29908;
  assign n29910 = n29907 & n29909;
  assign n29911 = ~n29423 & ~n29910;
  assign n29912 = P1_INSTQUEUE_REG_7__7_ & n29371;
  assign n29913 = P1_INSTQUEUE_REG_6__7_ & n29373;
  assign n29914 = P1_INSTQUEUE_REG_5__7_ & n29375;
  assign n29915 = P1_INSTQUEUE_REG_4__7_ & n29377;
  assign n29916 = ~n29912 & ~n29913;
  assign n29917 = ~n29914 & n29916;
  assign n29918 = ~n29915 & n29917;
  assign n29919 = P1_INSTQUEUE_REG_3__7_ & n29383;
  assign n29920 = P1_INSTQUEUE_REG_2__7_ & n29385;
  assign n29921 = P1_INSTQUEUE_REG_1__7_ & n29387;
  assign n29922 = P1_INSTQUEUE_REG_0__7_ & n29389;
  assign n29923 = ~n29919 & ~n29920;
  assign n29924 = ~n29921 & n29923;
  assign n29925 = ~n29922 & n29924;
  assign n29926 = P1_INSTQUEUE_REG_15__7_ & n29395;
  assign n29927 = P1_INSTQUEUE_REG_14__7_ & n29397;
  assign n29928 = P1_INSTQUEUE_REG_13__7_ & n29399;
  assign n29929 = P1_INSTQUEUE_REG_12__7_ & n29401;
  assign n29930 = ~n29926 & ~n29927;
  assign n29931 = ~n29928 & n29930;
  assign n29932 = ~n29929 & n29931;
  assign n29933 = P1_INSTQUEUE_REG_11__7_ & n29407;
  assign n29934 = P1_INSTQUEUE_REG_10__7_ & n29409;
  assign n29935 = P1_INSTQUEUE_REG_9__7_ & n29411;
  assign n29936 = P1_INSTQUEUE_REG_8__7_ & n29413;
  assign n29937 = ~n29933 & ~n29934;
  assign n29938 = ~n29935 & n29937;
  assign n29939 = ~n29936 & n29938;
  assign n29940 = n29918 & n29925;
  assign n29941 = n29932 & n29940;
  assign n29942 = n29939 & n29941;
  assign n29943 = ~n29423 & ~n29942;
  assign n29944 = ~n29911 & ~n29943;
  assign n29945 = n29911 & n29943;
  assign n29946 = ~n29944 & ~n29945;
  assign n29947 = ~n28840 & n29946;
  assign n29948 = P1_EAX_REG_23_ & n28833;
  assign n29949 = P1_PHYADDRPOINTER_REG_23_ & n28837;
  assign n29950 = n24584 & ~n29855;
  assign n29951 = ~n29948 & ~n29949;
  assign n29952 = ~n29950 & n29951;
  assign n29953 = ~n29947 & n29952;
  assign n29954 = ~n24584 & ~n29953;
  assign n29955 = n24584 & n29953;
  assign n29956 = ~n29954 & ~n29955;
  assign n29957 = n29468 & ~n29956;
  assign n29958 = ~n29468 & n29956;
  assign n29959 = ~n29957 & ~n29958;
  assign n29960 = ~n29836 & ~n29839;
  assign n29961 = ~n29835 & ~n29960;
  assign n29962 = ~n29836 & n29840;
  assign n29963 = ~n29647 & n29962;
  assign n29964 = n29961 & ~n29963;
  assign n29965 = n29959 & n29964;
  assign n29966 = ~n29959 & ~n29964;
  assign n29967 = ~n29965 & ~n29966;
  assign n29968 = n28859 & ~n29967;
  assign n29969 = ~n29851 & ~n29856;
  assign n29970 = ~n29857 & n29969;
  assign n29971 = ~n29858 & n29970;
  assign n6364 = n29968 | ~n29971;
  assign n29973 = P1_REIP_REG_24_ & n28830;
  assign n29974 = P1_PHYADDRPOINTER_REG_23_ & n29852;
  assign n29975 = ~P1_PHYADDRPOINTER_REG_24_ & n29974;
  assign n29976 = P1_PHYADDRPOINTER_REG_24_ & ~n29974;
  assign n29977 = ~n29975 & ~n29976;
  assign n29978 = n28828 & ~n29977;
  assign n29979 = P1_PHYADDRPOINTER_REG_24_ & n28822;
  assign n29980 = ~n28418 & n28823;
  assign n29981 = P1_INSTQUEUE_REG_7__1_ & n29861;
  assign n29982 = P1_INSTQUEUE_REG_6__1_ & n29863;
  assign n29983 = P1_INSTQUEUE_REG_5__1_ & n29866;
  assign n29984 = P1_INSTQUEUE_REG_4__1_ & n29868;
  assign n29985 = ~n29981 & ~n29982;
  assign n29986 = ~n29983 & n29985;
  assign n29987 = ~n29984 & n29986;
  assign n29988 = P1_INSTQUEUE_REG_3__1_ & n29874;
  assign n29989 = P1_INSTQUEUE_REG_2__1_ & n29876;
  assign n29990 = P1_INSTQUEUE_REG_1__1_ & n29878;
  assign n29991 = P1_INSTQUEUE_REG_0__1_ & n29880;
  assign n29992 = ~n29988 & ~n29989;
  assign n29993 = ~n29990 & n29992;
  assign n29994 = ~n29991 & n29993;
  assign n29995 = P1_INSTQUEUE_REG_15__1_ & n29885;
  assign n29996 = P1_INSTQUEUE_REG_14__1_ & n29887;
  assign n29997 = P1_INSTQUEUE_REG_13__1_ & n29889;
  assign n29998 = P1_INSTQUEUE_REG_12__1_ & n29891;
  assign n29999 = ~n29995 & ~n29996;
  assign n30000 = ~n29997 & n29999;
  assign n30001 = ~n29998 & n30000;
  assign n30002 = P1_INSTQUEUE_REG_11__1_ & n29897;
  assign n30003 = P1_INSTQUEUE_REG_10__1_ & n29899;
  assign n30004 = P1_INSTQUEUE_REG_9__1_ & n29901;
  assign n30005 = P1_INSTQUEUE_REG_8__1_ & n29903;
  assign n30006 = ~n30002 & ~n30003;
  assign n30007 = ~n30004 & n30006;
  assign n30008 = ~n30005 & n30007;
  assign n30009 = n29987 & n29994;
  assign n30010 = n30001 & n30009;
  assign n30011 = n30008 & n30010;
  assign n30012 = ~n29423 & ~n30011;
  assign n30013 = ~n29945 & n30012;
  assign n30014 = n29945 & ~n30012;
  assign n30015 = ~n30013 & ~n30014;
  assign n30016 = ~n28840 & ~n30015;
  assign n30017 = P1_EAX_REG_24_ & n28833;
  assign n30018 = P1_PHYADDRPOINTER_REG_24_ & n28837;
  assign n30019 = n24584 & ~n29977;
  assign n30020 = ~n30017 & ~n30018;
  assign n30021 = ~n30019 & n30020;
  assign n30022 = ~n30016 & n30021;
  assign n30023 = ~n24584 & ~n30022;
  assign n30024 = n24584 & n30022;
  assign n30025 = ~n30023 & ~n30024;
  assign n30026 = n29468 & ~n30025;
  assign n30027 = ~n29468 & n30025;
  assign n30028 = ~n30026 & ~n30027;
  assign n30029 = ~n29958 & ~n29964;
  assign n30030 = ~n29957 & ~n30029;
  assign n30031 = n30028 & n30030;
  assign n30032 = ~n30028 & ~n30030;
  assign n30033 = ~n30031 & ~n30032;
  assign n30034 = n28859 & ~n30033;
  assign n30035 = ~n29973 & ~n29978;
  assign n30036 = ~n29979 & n30035;
  assign n30037 = ~n29980 & n30036;
  assign n6369 = n30034 | ~n30037;
  assign n30039 = P1_REIP_REG_25_ & n28830;
  assign n30040 = P1_PHYADDRPOINTER_REG_24_ & n29974;
  assign n30041 = ~P1_PHYADDRPOINTER_REG_25_ & n30040;
  assign n30042 = P1_PHYADDRPOINTER_REG_25_ & ~n30040;
  assign n30043 = ~n30041 & ~n30042;
  assign n30044 = n28828 & ~n30043;
  assign n30045 = P1_PHYADDRPOINTER_REG_25_ & n28822;
  assign n30046 = ~n28467 & n28823;
  assign n30047 = n29945 & n30012;
  assign n30048 = P1_INSTQUEUE_REG_7__2_ & n29861;
  assign n30049 = P1_INSTQUEUE_REG_6__2_ & n29863;
  assign n30050 = P1_INSTQUEUE_REG_5__2_ & n29866;
  assign n30051 = P1_INSTQUEUE_REG_4__2_ & n29868;
  assign n30052 = ~n30048 & ~n30049;
  assign n30053 = ~n30050 & n30052;
  assign n30054 = ~n30051 & n30053;
  assign n30055 = P1_INSTQUEUE_REG_3__2_ & n29874;
  assign n30056 = P1_INSTQUEUE_REG_2__2_ & n29876;
  assign n30057 = P1_INSTQUEUE_REG_1__2_ & n29878;
  assign n30058 = P1_INSTQUEUE_REG_0__2_ & n29880;
  assign n30059 = ~n30055 & ~n30056;
  assign n30060 = ~n30057 & n30059;
  assign n30061 = ~n30058 & n30060;
  assign n30062 = P1_INSTQUEUE_REG_15__2_ & n29885;
  assign n30063 = P1_INSTQUEUE_REG_14__2_ & n29887;
  assign n30064 = P1_INSTQUEUE_REG_13__2_ & n29889;
  assign n30065 = P1_INSTQUEUE_REG_12__2_ & n29891;
  assign n30066 = ~n30062 & ~n30063;
  assign n30067 = ~n30064 & n30066;
  assign n30068 = ~n30065 & n30067;
  assign n30069 = P1_INSTQUEUE_REG_11__2_ & n29897;
  assign n30070 = P1_INSTQUEUE_REG_10__2_ & n29899;
  assign n30071 = P1_INSTQUEUE_REG_9__2_ & n29901;
  assign n30072 = P1_INSTQUEUE_REG_8__2_ & n29903;
  assign n30073 = ~n30069 & ~n30070;
  assign n30074 = ~n30071 & n30073;
  assign n30075 = ~n30072 & n30074;
  assign n30076 = n30054 & n30061;
  assign n30077 = n30068 & n30076;
  assign n30078 = n30075 & n30077;
  assign n30079 = ~n29423 & ~n30078;
  assign n30080 = n30047 & ~n30079;
  assign n30081 = ~n30047 & n30079;
  assign n30082 = ~n30080 & ~n30081;
  assign n30083 = ~n28840 & ~n30082;
  assign n30084 = P1_EAX_REG_25_ & n28833;
  assign n30085 = P1_PHYADDRPOINTER_REG_25_ & n28837;
  assign n30086 = n24584 & ~n30043;
  assign n30087 = ~n30084 & ~n30085;
  assign n30088 = ~n30086 & n30087;
  assign n30089 = ~n30083 & n30088;
  assign n30090 = ~n24584 & ~n30089;
  assign n30091 = n24584 & n30089;
  assign n30092 = ~n30090 & ~n30091;
  assign n30093 = n29468 & ~n30092;
  assign n30094 = ~n29468 & n30092;
  assign n30095 = ~n30093 & ~n30094;
  assign n30096 = n29957 & ~n30027;
  assign n30097 = ~n30026 & ~n30096;
  assign n30098 = ~n29958 & ~n30027;
  assign n30099 = ~n29964 & n30098;
  assign n30100 = n30097 & ~n30099;
  assign n30101 = n30095 & n30100;
  assign n30102 = ~n30095 & ~n30100;
  assign n30103 = ~n30101 & ~n30102;
  assign n30104 = n28859 & ~n30103;
  assign n30105 = ~n30039 & ~n30044;
  assign n30106 = ~n30045 & n30105;
  assign n30107 = ~n30046 & n30106;
  assign n6374 = n30104 | ~n30107;
  assign n30109 = P1_REIP_REG_26_ & n28830;
  assign n30110 = P1_PHYADDRPOINTER_REG_25_ & n30040;
  assign n30111 = ~P1_PHYADDRPOINTER_REG_26_ & n30110;
  assign n30112 = P1_PHYADDRPOINTER_REG_26_ & ~n30110;
  assign n30113 = ~n30111 & ~n30112;
  assign n30114 = n28828 & ~n30113;
  assign n30115 = P1_PHYADDRPOINTER_REG_26_ & n28822;
  assign n30116 = ~n28515 & n28823;
  assign n30117 = P1_INSTQUEUE_REG_7__3_ & n29861;
  assign n30118 = P1_INSTQUEUE_REG_6__3_ & n29863;
  assign n30119 = P1_INSTQUEUE_REG_5__3_ & n29866;
  assign n30120 = P1_INSTQUEUE_REG_4__3_ & n29868;
  assign n30121 = ~n30117 & ~n30118;
  assign n30122 = ~n30119 & n30121;
  assign n30123 = ~n30120 & n30122;
  assign n30124 = P1_INSTQUEUE_REG_3__3_ & n29874;
  assign n30125 = P1_INSTQUEUE_REG_2__3_ & n29876;
  assign n30126 = P1_INSTQUEUE_REG_1__3_ & n29878;
  assign n30127 = P1_INSTQUEUE_REG_0__3_ & n29880;
  assign n30128 = ~n30124 & ~n30125;
  assign n30129 = ~n30126 & n30128;
  assign n30130 = ~n30127 & n30129;
  assign n30131 = P1_INSTQUEUE_REG_15__3_ & n29885;
  assign n30132 = P1_INSTQUEUE_REG_14__3_ & n29887;
  assign n30133 = P1_INSTQUEUE_REG_13__3_ & n29889;
  assign n30134 = P1_INSTQUEUE_REG_12__3_ & n29891;
  assign n30135 = ~n30131 & ~n30132;
  assign n30136 = ~n30133 & n30135;
  assign n30137 = ~n30134 & n30136;
  assign n30138 = P1_INSTQUEUE_REG_11__3_ & n29897;
  assign n30139 = P1_INSTQUEUE_REG_10__3_ & n29899;
  assign n30140 = P1_INSTQUEUE_REG_9__3_ & n29901;
  assign n30141 = P1_INSTQUEUE_REG_8__3_ & n29903;
  assign n30142 = ~n30138 & ~n30139;
  assign n30143 = ~n30140 & n30142;
  assign n30144 = ~n30141 & n30143;
  assign n30145 = n30123 & n30130;
  assign n30146 = n30137 & n30145;
  assign n30147 = n30144 & n30146;
  assign n30148 = ~n29423 & ~n30147;
  assign n30149 = n30012 & n30079;
  assign n30150 = n29945 & n30149;
  assign n30151 = n30148 & ~n30150;
  assign n30152 = ~n30148 & n30150;
  assign n30153 = ~n30151 & ~n30152;
  assign n30154 = ~n28840 & ~n30153;
  assign n30155 = P1_EAX_REG_26_ & n28833;
  assign n30156 = P1_PHYADDRPOINTER_REG_26_ & n28837;
  assign n30157 = n24584 & ~n30113;
  assign n30158 = ~n30155 & ~n30156;
  assign n30159 = ~n30157 & n30158;
  assign n30160 = ~n30154 & n30159;
  assign n30161 = ~n24584 & ~n30160;
  assign n30162 = n24584 & n30160;
  assign n30163 = ~n30161 & ~n30162;
  assign n30164 = n29468 & ~n30163;
  assign n30165 = ~n29468 & n30163;
  assign n30166 = ~n30164 & ~n30165;
  assign n30167 = ~n30094 & ~n30097;
  assign n30168 = ~n30093 & ~n30167;
  assign n30169 = ~n30094 & n30098;
  assign n30170 = ~n29964 & n30169;
  assign n30171 = n30168 & ~n30170;
  assign n30172 = n30166 & n30171;
  assign n30173 = ~n30166 & ~n30171;
  assign n30174 = ~n30172 & ~n30173;
  assign n30175 = n28859 & ~n30174;
  assign n30176 = ~n30109 & ~n30114;
  assign n30177 = ~n30115 & n30176;
  assign n30178 = ~n30116 & n30177;
  assign n6379 = n30175 | ~n30178;
  assign n30180 = P1_REIP_REG_27_ & n28830;
  assign n30181 = P1_PHYADDRPOINTER_REG_26_ & n30110;
  assign n30182 = ~P1_PHYADDRPOINTER_REG_27_ & n30181;
  assign n30183 = P1_PHYADDRPOINTER_REG_27_ & ~n30181;
  assign n30184 = ~n30182 & ~n30183;
  assign n30185 = n28828 & ~n30184;
  assign n30186 = P1_PHYADDRPOINTER_REG_27_ & n28822;
  assign n30187 = ~n28565 & n28823;
  assign n30188 = n30148 & n30150;
  assign n30189 = P1_INSTQUEUE_REG_0__4_ & n29880;
  assign n30190 = P1_INSTQUEUE_REG_7__4_ & n29861;
  assign n30191 = P1_INSTQUEUE_REG_6__4_ & n29863;
  assign n30192 = P1_INSTQUEUE_REG_5__4_ & n29866;
  assign n30193 = ~n30191 & ~n30192;
  assign n30194 = ~n30189 & ~n30190;
  assign n30195 = n30193 & n30194;
  assign n30196 = P1_INSTQUEUE_REG_4__4_ & n29868;
  assign n30197 = P1_INSTQUEUE_REG_3__4_ & n29874;
  assign n30198 = P1_INSTQUEUE_REG_2__4_ & n29876;
  assign n30199 = P1_INSTQUEUE_REG_1__4_ & n29878;
  assign n30200 = ~n30196 & ~n30197;
  assign n30201 = ~n30198 & n30200;
  assign n30202 = ~n30199 & n30201;
  assign n30203 = P1_INSTQUEUE_REG_15__4_ & n29885;
  assign n30204 = P1_INSTQUEUE_REG_14__4_ & n29887;
  assign n30205 = P1_INSTQUEUE_REG_13__4_ & n29889;
  assign n30206 = P1_INSTQUEUE_REG_12__4_ & n29891;
  assign n30207 = ~n30203 & ~n30204;
  assign n30208 = ~n30205 & n30207;
  assign n30209 = ~n30206 & n30208;
  assign n30210 = P1_INSTQUEUE_REG_11__4_ & n29897;
  assign n30211 = P1_INSTQUEUE_REG_10__4_ & n29899;
  assign n30212 = P1_INSTQUEUE_REG_9__4_ & n29901;
  assign n30213 = P1_INSTQUEUE_REG_8__4_ & n29903;
  assign n30214 = ~n30210 & ~n30211;
  assign n30215 = ~n30212 & n30214;
  assign n30216 = ~n30213 & n30215;
  assign n30217 = n30195 & n30202;
  assign n30218 = n30209 & n30217;
  assign n30219 = n30216 & n30218;
  assign n30220 = ~n29423 & ~n30219;
  assign n30221 = n30188 & ~n30220;
  assign n30222 = ~n30188 & n30220;
  assign n30223 = ~n30221 & ~n30222;
  assign n30224 = ~n28840 & ~n30223;
  assign n30225 = P1_EAX_REG_27_ & n28833;
  assign n30226 = P1_PHYADDRPOINTER_REG_27_ & n28837;
  assign n30227 = n24584 & ~n30184;
  assign n30228 = ~n30225 & ~n30226;
  assign n30229 = ~n30227 & n30228;
  assign n30230 = ~n30224 & n30229;
  assign n30231 = ~n24584 & ~n30230;
  assign n30232 = n24584 & n30230;
  assign n30233 = ~n30231 & ~n30232;
  assign n30234 = n29468 & ~n30233;
  assign n30235 = ~n29468 & n30233;
  assign n30236 = ~n30234 & ~n30235;
  assign n30237 = ~n30165 & ~n30168;
  assign n30238 = ~n30164 & ~n30237;
  assign n30239 = ~n30165 & n30169;
  assign n30240 = ~n29964 & n30239;
  assign n30241 = n30238 & ~n30240;
  assign n30242 = n30236 & n30241;
  assign n30243 = ~n30236 & ~n30241;
  assign n30244 = ~n30242 & ~n30243;
  assign n30245 = n28859 & ~n30244;
  assign n30246 = ~n30180 & ~n30185;
  assign n30247 = ~n30186 & n30246;
  assign n30248 = ~n30187 & n30247;
  assign n6384 = n30245 | ~n30248;
  assign n30250 = P1_REIP_REG_28_ & n28830;
  assign n30251 = P1_PHYADDRPOINTER_REG_27_ & n30181;
  assign n30252 = ~P1_PHYADDRPOINTER_REG_28_ & n30251;
  assign n30253 = P1_PHYADDRPOINTER_REG_28_ & ~n30251;
  assign n30254 = ~n30252 & ~n30253;
  assign n30255 = n28828 & ~n30254;
  assign n30256 = P1_PHYADDRPOINTER_REG_28_ & n28822;
  assign n30257 = ~n28614 & n28823;
  assign n30258 = P1_INSTQUEUE_REG_7__5_ & n29861;
  assign n30259 = P1_INSTQUEUE_REG_6__5_ & n29863;
  assign n30260 = P1_INSTQUEUE_REG_5__5_ & n29866;
  assign n30261 = P1_INSTQUEUE_REG_4__5_ & n29868;
  assign n30262 = ~n30258 & ~n30259;
  assign n30263 = ~n30260 & n30262;
  assign n30264 = ~n30261 & n30263;
  assign n30265 = P1_INSTQUEUE_REG_3__5_ & n29874;
  assign n30266 = P1_INSTQUEUE_REG_2__5_ & n29876;
  assign n30267 = P1_INSTQUEUE_REG_1__5_ & n29878;
  assign n30268 = P1_INSTQUEUE_REG_0__5_ & n29880;
  assign n30269 = ~n30265 & ~n30266;
  assign n30270 = ~n30267 & n30269;
  assign n30271 = ~n30268 & n30270;
  assign n30272 = P1_INSTQUEUE_REG_15__5_ & n29885;
  assign n30273 = P1_INSTQUEUE_REG_14__5_ & n29887;
  assign n30274 = P1_INSTQUEUE_REG_13__5_ & n29889;
  assign n30275 = P1_INSTQUEUE_REG_12__5_ & n29891;
  assign n30276 = ~n30272 & ~n30273;
  assign n30277 = ~n30274 & n30276;
  assign n30278 = ~n30275 & n30277;
  assign n30279 = P1_INSTQUEUE_REG_11__5_ & n29897;
  assign n30280 = P1_INSTQUEUE_REG_10__5_ & n29899;
  assign n30281 = P1_INSTQUEUE_REG_9__5_ & n29901;
  assign n30282 = P1_INSTQUEUE_REG_8__5_ & n29903;
  assign n30283 = ~n30279 & ~n30280;
  assign n30284 = ~n30281 & n30283;
  assign n30285 = ~n30282 & n30284;
  assign n30286 = n30264 & n30271;
  assign n30287 = n30278 & n30286;
  assign n30288 = n30285 & n30287;
  assign n30289 = ~n29423 & ~n30288;
  assign n30290 = n30148 & n30220;
  assign n30291 = n30150 & n30290;
  assign n30292 = n30289 & ~n30291;
  assign n30293 = ~n30289 & n30291;
  assign n30294 = ~n30292 & ~n30293;
  assign n30295 = ~n28840 & ~n30294;
  assign n30296 = P1_EAX_REG_28_ & n28833;
  assign n30297 = P1_PHYADDRPOINTER_REG_28_ & n28837;
  assign n30298 = n24584 & ~n30254;
  assign n30299 = ~n30296 & ~n30297;
  assign n30300 = ~n30298 & n30299;
  assign n30301 = ~n30295 & n30300;
  assign n30302 = ~n24584 & ~n30301;
  assign n30303 = n24584 & n30301;
  assign n30304 = ~n30302 & ~n30303;
  assign n30305 = n29468 & ~n30304;
  assign n30306 = ~n29468 & n30304;
  assign n30307 = ~n30305 & ~n30306;
  assign n30308 = ~n30235 & ~n30238;
  assign n30309 = ~n30234 & ~n30308;
  assign n30310 = ~n30235 & n30239;
  assign n30311 = ~n29964 & n30310;
  assign n30312 = n30309 & ~n30311;
  assign n30313 = n30307 & n30312;
  assign n30314 = ~n30307 & ~n30312;
  assign n30315 = ~n30313 & ~n30314;
  assign n30316 = n28859 & ~n30315;
  assign n30317 = ~n30250 & ~n30255;
  assign n30318 = ~n30256 & n30317;
  assign n30319 = ~n30257 & n30318;
  assign n6389 = n30316 | ~n30319;
  assign n30321 = P1_REIP_REG_29_ & n28830;
  assign n30322 = P1_PHYADDRPOINTER_REG_28_ & n30251;
  assign n30323 = ~P1_PHYADDRPOINTER_REG_29_ & n30322;
  assign n30324 = P1_PHYADDRPOINTER_REG_29_ & ~n30322;
  assign n30325 = ~n30323 & ~n30324;
  assign n30326 = n28828 & ~n30325;
  assign n30327 = P1_PHYADDRPOINTER_REG_29_ & n28822;
  assign n30328 = ~n28680 & n28823;
  assign n30329 = n30289 & n30291;
  assign n30330 = P1_INSTQUEUE_REG_7__6_ & n29861;
  assign n30331 = P1_INSTQUEUE_REG_6__6_ & n29863;
  assign n30332 = P1_INSTQUEUE_REG_5__6_ & n29866;
  assign n30333 = P1_INSTQUEUE_REG_4__6_ & n29868;
  assign n30334 = ~n30330 & ~n30331;
  assign n30335 = ~n30332 & n30334;
  assign n30336 = ~n30333 & n30335;
  assign n30337 = P1_INSTQUEUE_REG_3__6_ & n29874;
  assign n30338 = P1_INSTQUEUE_REG_2__6_ & n29876;
  assign n30339 = P1_INSTQUEUE_REG_1__6_ & n29878;
  assign n30340 = P1_INSTQUEUE_REG_0__6_ & n29880;
  assign n30341 = ~n30337 & ~n30338;
  assign n30342 = ~n30339 & n30341;
  assign n30343 = ~n30340 & n30342;
  assign n30344 = P1_INSTQUEUE_REG_15__6_ & n29885;
  assign n30345 = P1_INSTQUEUE_REG_14__6_ & n29887;
  assign n30346 = P1_INSTQUEUE_REG_13__6_ & n29889;
  assign n30347 = P1_INSTQUEUE_REG_12__6_ & n29891;
  assign n30348 = ~n30344 & ~n30345;
  assign n30349 = ~n30346 & n30348;
  assign n30350 = ~n30347 & n30349;
  assign n30351 = P1_INSTQUEUE_REG_11__6_ & n29897;
  assign n30352 = P1_INSTQUEUE_REG_10__6_ & n29899;
  assign n30353 = P1_INSTQUEUE_REG_9__6_ & n29901;
  assign n30354 = P1_INSTQUEUE_REG_8__6_ & n29903;
  assign n30355 = ~n30351 & ~n30352;
  assign n30356 = ~n30353 & n30355;
  assign n30357 = ~n30354 & n30356;
  assign n30358 = n30336 & n30343;
  assign n30359 = n30350 & n30358;
  assign n30360 = n30357 & n30359;
  assign n30361 = ~n29423 & ~n30360;
  assign n30362 = n30329 & ~n30361;
  assign n30363 = ~n30329 & n30361;
  assign n30364 = ~n30362 & ~n30363;
  assign n30365 = ~n28840 & ~n30364;
  assign n30366 = P1_EAX_REG_29_ & n28833;
  assign n30367 = P1_PHYADDRPOINTER_REG_29_ & n28837;
  assign n30368 = n24584 & ~n30325;
  assign n30369 = ~n30366 & ~n30367;
  assign n30370 = ~n30368 & n30369;
  assign n30371 = ~n30365 & n30370;
  assign n30372 = ~n24584 & ~n30371;
  assign n30373 = n24584 & n30371;
  assign n30374 = ~n30372 & ~n30373;
  assign n30375 = n29468 & ~n30374;
  assign n30376 = ~n29468 & n30374;
  assign n30377 = ~n30375 & ~n30376;
  assign n30378 = ~n30306 & ~n30312;
  assign n30379 = ~n30305 & ~n30378;
  assign n30380 = n30377 & n30379;
  assign n30381 = ~n30377 & ~n30379;
  assign n30382 = ~n30380 & ~n30381;
  assign n30383 = n28859 & ~n30382;
  assign n30384 = ~n30321 & ~n30326;
  assign n30385 = ~n30327 & n30384;
  assign n30386 = ~n30328 & n30385;
  assign n6394 = n30383 | ~n30386;
  assign n30388 = P1_REIP_REG_30_ & n28830;
  assign n30389 = P1_PHYADDRPOINTER_REG_29_ & n30322;
  assign n30390 = ~P1_PHYADDRPOINTER_REG_30_ & n30389;
  assign n30391 = P1_PHYADDRPOINTER_REG_30_ & ~n30389;
  assign n30392 = ~n30390 & ~n30391;
  assign n30393 = n28828 & ~n30392;
  assign n30394 = P1_PHYADDRPOINTER_REG_30_ & n28822;
  assign n30395 = ~n28735 & n28823;
  assign n30396 = ~n30376 & ~n30379;
  assign n30397 = ~n30375 & ~n30396;
  assign n30398 = n30329 & n30361;
  assign n30399 = P1_INSTQUEUE_REG_7__7_ & n29861;
  assign n30400 = P1_INSTQUEUE_REG_6__7_ & n29863;
  assign n30401 = P1_INSTQUEUE_REG_5__7_ & n29866;
  assign n30402 = P1_INSTQUEUE_REG_4__7_ & n29868;
  assign n30403 = ~n30399 & ~n30400;
  assign n30404 = ~n30401 & n30403;
  assign n30405 = ~n30402 & n30404;
  assign n30406 = P1_INSTQUEUE_REG_3__7_ & n29874;
  assign n30407 = P1_INSTQUEUE_REG_2__7_ & n29876;
  assign n30408 = P1_INSTQUEUE_REG_1__7_ & n29878;
  assign n30409 = P1_INSTQUEUE_REG_0__7_ & n29880;
  assign n30410 = ~n30406 & ~n30407;
  assign n30411 = ~n30408 & n30410;
  assign n30412 = ~n30409 & n30411;
  assign n30413 = P1_INSTQUEUE_REG_15__7_ & n29885;
  assign n30414 = P1_INSTQUEUE_REG_14__7_ & n29887;
  assign n30415 = P1_INSTQUEUE_REG_13__7_ & n29889;
  assign n30416 = P1_INSTQUEUE_REG_12__7_ & n29891;
  assign n30417 = ~n30413 & ~n30414;
  assign n30418 = ~n30415 & n30417;
  assign n30419 = ~n30416 & n30418;
  assign n30420 = P1_INSTQUEUE_REG_11__7_ & n29897;
  assign n30421 = P1_INSTQUEUE_REG_10__7_ & n29899;
  assign n30422 = P1_INSTQUEUE_REG_9__7_ & n29901;
  assign n30423 = P1_INSTQUEUE_REG_8__7_ & n29903;
  assign n30424 = ~n30420 & ~n30421;
  assign n30425 = ~n30422 & n30424;
  assign n30426 = ~n30423 & n30425;
  assign n30427 = n30405 & n30412;
  assign n30428 = n30419 & n30427;
  assign n30429 = n30426 & n30428;
  assign n30430 = ~n29423 & ~n30429;
  assign n30431 = n30398 & ~n30430;
  assign n30432 = ~n30398 & n30430;
  assign n30433 = ~n30431 & ~n30432;
  assign n30434 = ~n28840 & ~n30433;
  assign n30435 = P1_EAX_REG_30_ & n28833;
  assign n30436 = P1_PHYADDRPOINTER_REG_30_ & n28837;
  assign n30437 = n24584 & ~n30392;
  assign n30438 = ~n30435 & ~n30436;
  assign n30439 = ~n30437 & n30438;
  assign n30440 = ~n30434 & n30439;
  assign n30441 = ~n24584 & ~n30440;
  assign n30442 = n24584 & n30440;
  assign n30443 = ~n30441 & ~n30442;
  assign n30444 = ~n29468 & ~n30443;
  assign n30445 = n29468 & n30443;
  assign n30446 = ~n30444 & ~n30445;
  assign n30447 = n30397 & ~n30446;
  assign n30448 = ~n30397 & n30446;
  assign n30449 = ~n30447 & ~n30448;
  assign n30450 = n28859 & ~n30449;
  assign n30451 = ~n30388 & ~n30393;
  assign n30452 = ~n30394 & n30451;
  assign n30453 = ~n30395 & n30452;
  assign n6399 = n30450 | ~n30453;
  assign n30455 = P1_REIP_REG_31_ & n28830;
  assign n30456 = P1_PHYADDRPOINTER_REG_30_ & n30389;
  assign n30457 = ~P1_PHYADDRPOINTER_REG_31_ & n30456;
  assign n30458 = P1_PHYADDRPOINTER_REG_31_ & ~n30456;
  assign n30459 = ~n30457 & ~n30458;
  assign n30460 = n28828 & ~n30459;
  assign n30461 = P1_PHYADDRPOINTER_REG_31_ & n28822;
  assign n30462 = n28809 & n28823;
  assign n30463 = P1_PHYADDRPOINTER_REG_31_ & n28837;
  assign n30464 = P1_EAX_REG_31_ & n28833;
  assign n30465 = n24584 & ~n30459;
  assign n30466 = ~n30463 & ~n30464;
  assign n30467 = ~n30465 & n30466;
  assign n30468 = ~n24584 & ~n30467;
  assign n30469 = n24584 & n30467;
  assign n30470 = ~n30468 & ~n30469;
  assign n30471 = ~n29468 & n30443;
  assign n30472 = ~n30470 & ~n30471;
  assign n30473 = n30375 & n30472;
  assign n30474 = n29468 & ~n30443;
  assign n30475 = n30470 & ~n30474;
  assign n30476 = ~n30396 & n30475;
  assign n30477 = ~n30375 & n30476;
  assign n30478 = ~n30443 & ~n30470;
  assign n30479 = n29468 & n30478;
  assign n30480 = n30443 & n30470;
  assign n30481 = ~n29468 & n30480;
  assign n30482 = ~n30479 & ~n30481;
  assign n30483 = n30396 & n30472;
  assign n30484 = n30482 & ~n30483;
  assign n30485 = ~n30473 & ~n30477;
  assign n30486 = n30484 & n30485;
  assign n30487 = n28859 & n30486;
  assign n30488 = ~n30455 & ~n30460;
  assign n30489 = ~n30461 & n30488;
  assign n30490 = ~n30462 & n30489;
  assign n6404 = n30487 | ~n30490;
  assign n30492 = BUF1_REG_15_ & n4507;
  assign n30493 = DATAI_15_ & ~n4507;
  assign n30494 = ~n30492 & ~n30493;
  assign n30495 = n23523 & ~n24054;
  assign n30496 = ~n23678 & n24576;
  assign n30497 = ~n30495 & n30496;
  assign n30498 = ~n24164 & n30497;
  assign n30499 = ~n23709 & n30498;
  assign n30500 = ~n30494 & n30499;
  assign n30501 = n23709 & n30498;
  assign n30502 = P1_EAX_REG_15_ & n30501;
  assign n30503 = ~n30500 & ~n30502;
  assign n30504 = n24184 & ~n30503;
  assign n30505 = n24184 & n30498;
  assign n30506 = P1_LWORD_REG_15_ & ~n30505;
  assign n6409 = n30504 | n30506;
  assign n30508 = BUF1_REG_14_ & n4507;
  assign n30509 = DATAI_14_ & ~n4507;
  assign n30510 = ~n30508 & ~n30509;
  assign n30511 = n30499 & ~n30510;
  assign n30512 = P1_EAX_REG_14_ & n30501;
  assign n30513 = ~n30511 & ~n30512;
  assign n30514 = n24184 & ~n30513;
  assign n30515 = P1_LWORD_REG_14_ & ~n30505;
  assign n6414 = n30514 | n30515;
  assign n30517 = BUF1_REG_13_ & n4507;
  assign n30518 = DATAI_13_ & ~n4507;
  assign n30519 = ~n30517 & ~n30518;
  assign n30520 = n30499 & ~n30519;
  assign n30521 = P1_EAX_REG_13_ & n30501;
  assign n30522 = ~n30520 & ~n30521;
  assign n30523 = n24184 & ~n30522;
  assign n30524 = P1_LWORD_REG_13_ & ~n30505;
  assign n6419 = n30523 | n30524;
  assign n30526 = BUF1_REG_12_ & n4507;
  assign n30527 = DATAI_12_ & ~n4507;
  assign n30528 = ~n30526 & ~n30527;
  assign n30529 = n30499 & ~n30528;
  assign n30530 = P1_EAX_REG_12_ & n30501;
  assign n30531 = ~n30529 & ~n30530;
  assign n30532 = n24184 & ~n30531;
  assign n30533 = P1_LWORD_REG_12_ & ~n30505;
  assign n6424 = n30532 | n30533;
  assign n30535 = BUF1_REG_11_ & n4507;
  assign n30536 = DATAI_11_ & ~n4507;
  assign n30537 = ~n30535 & ~n30536;
  assign n30538 = n30499 & ~n30537;
  assign n30539 = P1_EAX_REG_11_ & n30501;
  assign n30540 = ~n30538 & ~n30539;
  assign n30541 = n24184 & ~n30540;
  assign n30542 = P1_LWORD_REG_11_ & ~n30505;
  assign n6429 = n30541 | n30542;
  assign n30544 = BUF1_REG_10_ & n4507;
  assign n30545 = DATAI_10_ & ~n4507;
  assign n30546 = ~n30544 & ~n30545;
  assign n30547 = n30499 & ~n30546;
  assign n30548 = P1_EAX_REG_10_ & n30501;
  assign n30549 = ~n30547 & ~n30548;
  assign n30550 = n24184 & ~n30549;
  assign n30551 = P1_LWORD_REG_10_ & ~n30505;
  assign n6434 = n30550 | n30551;
  assign n30553 = BUF1_REG_9_ & n4507;
  assign n30554 = DATAI_9_ & ~n4507;
  assign n30555 = ~n30553 & ~n30554;
  assign n30556 = n30499 & ~n30555;
  assign n30557 = P1_EAX_REG_9_ & n30501;
  assign n30558 = ~n30556 & ~n30557;
  assign n30559 = n24184 & ~n30558;
  assign n30560 = P1_LWORD_REG_9_ & ~n30505;
  assign n6439 = n30559 | n30560;
  assign n30562 = BUF1_REG_8_ & n4507;
  assign n30563 = DATAI_8_ & ~n4507;
  assign n30564 = ~n30562 & ~n30563;
  assign n30565 = n30499 & ~n30564;
  assign n30566 = P1_EAX_REG_8_ & n30501;
  assign n30567 = ~n30565 & ~n30566;
  assign n30568 = n24184 & ~n30567;
  assign n30569 = P1_LWORD_REG_8_ & ~n30505;
  assign n6444 = n30568 | n30569;
  assign n30571 = ~n24929 & n30499;
  assign n30572 = P1_EAX_REG_7_ & n30501;
  assign n30573 = ~n30571 & ~n30572;
  assign n30574 = n24184 & ~n30573;
  assign n30575 = P1_LWORD_REG_7_ & ~n30505;
  assign n6449 = n30574 | n30575;
  assign n30577 = ~n24957 & n30499;
  assign n30578 = P1_EAX_REG_6_ & n30501;
  assign n30579 = ~n30577 & ~n30578;
  assign n30580 = n24184 & ~n30579;
  assign n30581 = P1_LWORD_REG_6_ & ~n30505;
  assign n6454 = n30580 | n30581;
  assign n30583 = ~n24979 & n30499;
  assign n30584 = P1_EAX_REG_5_ & n30501;
  assign n30585 = ~n30583 & ~n30584;
  assign n30586 = n24184 & ~n30585;
  assign n30587 = P1_LWORD_REG_5_ & ~n30505;
  assign n6459 = n30586 | n30587;
  assign n30589 = ~n25001 & n30499;
  assign n30590 = P1_EAX_REG_4_ & n30501;
  assign n30591 = ~n30589 & ~n30590;
  assign n30592 = n24184 & ~n30591;
  assign n30593 = P1_LWORD_REG_4_ & ~n30505;
  assign n6464 = n30592 | n30593;
  assign n30595 = ~n25023 & n30499;
  assign n30596 = P1_EAX_REG_3_ & n30501;
  assign n30597 = ~n30595 & ~n30596;
  assign n30598 = n24184 & ~n30597;
  assign n30599 = P1_LWORD_REG_3_ & ~n30505;
  assign n6469 = n30598 | n30599;
  assign n30601 = ~n25045 & n30499;
  assign n30602 = P1_EAX_REG_2_ & n30501;
  assign n30603 = ~n30601 & ~n30602;
  assign n30604 = n24184 & ~n30603;
  assign n30605 = P1_LWORD_REG_2_ & ~n30505;
  assign n6474 = n30604 | n30605;
  assign n30607 = ~n25067 & n30499;
  assign n30608 = P1_EAX_REG_1_ & n30501;
  assign n30609 = ~n30607 & ~n30608;
  assign n30610 = n24184 & ~n30609;
  assign n30611 = P1_LWORD_REG_1_ & ~n30505;
  assign n6479 = n30610 | n30611;
  assign n30613 = ~n25089 & n30499;
  assign n30614 = P1_EAX_REG_0_ & n30501;
  assign n30615 = ~n30613 & ~n30614;
  assign n30616 = n24184 & ~n30615;
  assign n30617 = P1_LWORD_REG_0_ & ~n30505;
  assign n6484 = n30616 | n30617;
  assign n30619 = P1_EAX_REG_30_ & n30501;
  assign n30620 = ~n30511 & ~n30619;
  assign n30621 = n24184 & ~n30620;
  assign n30622 = P1_UWORD_REG_14_ & ~n30505;
  assign n6489 = n30621 | n30622;
  assign n30624 = P1_EAX_REG_29_ & n30501;
  assign n30625 = ~n30520 & ~n30624;
  assign n30626 = n24184 & ~n30625;
  assign n30627 = P1_UWORD_REG_13_ & ~n30505;
  assign n6494 = n30626 | n30627;
  assign n30629 = P1_EAX_REG_28_ & n30501;
  assign n30630 = ~n30529 & ~n30629;
  assign n30631 = n24184 & ~n30630;
  assign n30632 = P1_UWORD_REG_12_ & ~n30505;
  assign n6499 = n30631 | n30632;
  assign n30634 = P1_EAX_REG_27_ & n30501;
  assign n30635 = ~n30538 & ~n30634;
  assign n30636 = n24184 & ~n30635;
  assign n30637 = P1_UWORD_REG_11_ & ~n30505;
  assign n6504 = n30636 | n30637;
  assign n30639 = P1_EAX_REG_26_ & n30501;
  assign n30640 = ~n30547 & ~n30639;
  assign n30641 = n24184 & ~n30640;
  assign n30642 = P1_UWORD_REG_10_ & ~n30505;
  assign n6509 = n30641 | n30642;
  assign n30644 = P1_EAX_REG_25_ & n30501;
  assign n30645 = ~n30556 & ~n30644;
  assign n30646 = n24184 & ~n30645;
  assign n30647 = P1_UWORD_REG_9_ & ~n30505;
  assign n6514 = n30646 | n30647;
  assign n30649 = P1_EAX_REG_24_ & n30501;
  assign n30650 = ~n30565 & ~n30649;
  assign n30651 = n24184 & ~n30650;
  assign n30652 = P1_UWORD_REG_8_ & ~n30505;
  assign n6519 = n30651 | n30652;
  assign n30654 = P1_EAX_REG_23_ & n30501;
  assign n30655 = ~n30571 & ~n30654;
  assign n30656 = n24184 & ~n30655;
  assign n30657 = P1_UWORD_REG_7_ & ~n30505;
  assign n6524 = n30656 | n30657;
  assign n30659 = P1_EAX_REG_22_ & n30501;
  assign n30660 = ~n30577 & ~n30659;
  assign n30661 = n24184 & ~n30660;
  assign n30662 = P1_UWORD_REG_6_ & ~n30505;
  assign n6529 = n30661 | n30662;
  assign n30664 = P1_EAX_REG_21_ & n30501;
  assign n30665 = ~n30583 & ~n30664;
  assign n30666 = n24184 & ~n30665;
  assign n30667 = P1_UWORD_REG_5_ & ~n30505;
  assign n6534 = n30666 | n30667;
  assign n30669 = P1_EAX_REG_20_ & n30501;
  assign n30670 = ~n30589 & ~n30669;
  assign n30671 = n24184 & ~n30670;
  assign n30672 = P1_UWORD_REG_4_ & ~n30505;
  assign n6539 = n30671 | n30672;
  assign n30674 = P1_EAX_REG_19_ & n30501;
  assign n30675 = ~n30595 & ~n30674;
  assign n30676 = n24184 & ~n30675;
  assign n30677 = P1_UWORD_REG_3_ & ~n30505;
  assign n6544 = n30676 | n30677;
  assign n30679 = P1_EAX_REG_18_ & n30501;
  assign n30680 = ~n30601 & ~n30679;
  assign n30681 = n24184 & ~n30680;
  assign n30682 = P1_UWORD_REG_2_ & ~n30505;
  assign n6549 = n30681 | n30682;
  assign n30684 = P1_EAX_REG_17_ & n30501;
  assign n30685 = ~n30607 & ~n30684;
  assign n30686 = n24184 & ~n30685;
  assign n30687 = P1_UWORD_REG_1_ & ~n30505;
  assign n6554 = n30686 | n30687;
  assign n30689 = P1_EAX_REG_16_ & n30501;
  assign n30690 = ~n30613 & ~n30689;
  assign n30691 = n24184 & ~n30690;
  assign n30692 = P1_UWORD_REG_0_ & ~n30505;
  assign n6559 = n30691 | n30692;
  assign n30694 = ~P1_STATE2_REG_0_ & n23609;
  assign n30695 = n24054 & n24576;
  assign n30696 = n24184 & n30695;
  assign n30697 = ~n24454 & ~n30696;
  assign n30698 = n24313 & ~n30697;
  assign n30699 = n24558 & n30698;
  assign n30700 = ~n30694 & ~n30699;
  assign n30701 = P1_STATE2_REG_0_ & ~n30700;
  assign n30702 = P1_EAX_REG_0_ & n30701;
  assign n30703 = ~P1_STATE2_REG_0_ & ~n30700;
  assign n30704 = P1_LWORD_REG_0_ & n30703;
  assign n30705 = P1_DATAO_REG_0_ & n30700;
  assign n30706 = ~n30702 & ~n30704;
  assign n6564 = n30705 | ~n30706;
  assign n30708 = P1_EAX_REG_1_ & n30701;
  assign n30709 = P1_LWORD_REG_1_ & n30703;
  assign n30710 = P1_DATAO_REG_1_ & n30700;
  assign n30711 = ~n30708 & ~n30709;
  assign n6569 = n30710 | ~n30711;
  assign n30713 = P1_EAX_REG_2_ & n30701;
  assign n30714 = P1_LWORD_REG_2_ & n30703;
  assign n30715 = P1_DATAO_REG_2_ & n30700;
  assign n30716 = ~n30713 & ~n30714;
  assign n6574 = n30715 | ~n30716;
  assign n30718 = P1_EAX_REG_3_ & n30701;
  assign n30719 = P1_LWORD_REG_3_ & n30703;
  assign n30720 = P1_DATAO_REG_3_ & n30700;
  assign n30721 = ~n30718 & ~n30719;
  assign n6579 = n30720 | ~n30721;
  assign n30723 = P1_EAX_REG_4_ & n30701;
  assign n30724 = P1_LWORD_REG_4_ & n30703;
  assign n30725 = P1_DATAO_REG_4_ & n30700;
  assign n30726 = ~n30723 & ~n30724;
  assign n6584 = n30725 | ~n30726;
  assign n30728 = P1_EAX_REG_5_ & n30701;
  assign n30729 = P1_LWORD_REG_5_ & n30703;
  assign n30730 = P1_DATAO_REG_5_ & n30700;
  assign n30731 = ~n30728 & ~n30729;
  assign n6589 = n30730 | ~n30731;
  assign n30733 = P1_EAX_REG_6_ & n30701;
  assign n30734 = P1_LWORD_REG_6_ & n30703;
  assign n30735 = P1_DATAO_REG_6_ & n30700;
  assign n30736 = ~n30733 & ~n30734;
  assign n6594 = n30735 | ~n30736;
  assign n30738 = P1_EAX_REG_7_ & n30701;
  assign n30739 = P1_LWORD_REG_7_ & n30703;
  assign n30740 = P1_DATAO_REG_7_ & n30700;
  assign n30741 = ~n30738 & ~n30739;
  assign n6599 = n30740 | ~n30741;
  assign n30743 = P1_EAX_REG_8_ & n30701;
  assign n30744 = P1_LWORD_REG_8_ & n30703;
  assign n30745 = P1_DATAO_REG_8_ & n30700;
  assign n30746 = ~n30743 & ~n30744;
  assign n6604 = n30745 | ~n30746;
  assign n30748 = P1_EAX_REG_9_ & n30701;
  assign n30749 = P1_LWORD_REG_9_ & n30703;
  assign n30750 = P1_DATAO_REG_9_ & n30700;
  assign n30751 = ~n30748 & ~n30749;
  assign n6609 = n30750 | ~n30751;
  assign n30753 = P1_EAX_REG_10_ & n30701;
  assign n30754 = P1_LWORD_REG_10_ & n30703;
  assign n30755 = P1_DATAO_REG_10_ & n30700;
  assign n30756 = ~n30753 & ~n30754;
  assign n6614 = n30755 | ~n30756;
  assign n30758 = P1_EAX_REG_11_ & n30701;
  assign n30759 = P1_LWORD_REG_11_ & n30703;
  assign n30760 = P1_DATAO_REG_11_ & n30700;
  assign n30761 = ~n30758 & ~n30759;
  assign n6619 = n30760 | ~n30761;
  assign n30763 = P1_EAX_REG_12_ & n30701;
  assign n30764 = P1_LWORD_REG_12_ & n30703;
  assign n30765 = P1_DATAO_REG_12_ & n30700;
  assign n30766 = ~n30763 & ~n30764;
  assign n6624 = n30765 | ~n30766;
  assign n30768 = P1_EAX_REG_13_ & n30701;
  assign n30769 = P1_LWORD_REG_13_ & n30703;
  assign n30770 = P1_DATAO_REG_13_ & n30700;
  assign n30771 = ~n30768 & ~n30769;
  assign n6629 = n30770 | ~n30771;
  assign n30773 = P1_EAX_REG_14_ & n30701;
  assign n30774 = P1_LWORD_REG_14_ & n30703;
  assign n30775 = P1_DATAO_REG_14_ & n30700;
  assign n30776 = ~n30773 & ~n30774;
  assign n6634 = n30775 | ~n30776;
  assign n30778 = P1_EAX_REG_15_ & n30701;
  assign n30779 = P1_LWORD_REG_15_ & n30703;
  assign n30780 = P1_DATAO_REG_15_ & n30700;
  assign n30781 = ~n30778 & ~n30779;
  assign n6639 = n30780 | ~n30781;
  assign n30783 = P1_UWORD_REG_0_ & n30703;
  assign n30784 = P1_DATAO_REG_16_ & n30700;
  assign n30785 = ~n30783 & ~n30784;
  assign n30786 = ~n23678 & n30701;
  assign n30787 = P1_EAX_REG_16_ & n30786;
  assign n6644 = ~n30785 | n30787;
  assign n30789 = P1_UWORD_REG_1_ & n30703;
  assign n30790 = P1_DATAO_REG_17_ & n30700;
  assign n30791 = ~n30789 & ~n30790;
  assign n30792 = P1_EAX_REG_17_ & n30786;
  assign n6649 = ~n30791 | n30792;
  assign n30794 = P1_UWORD_REG_2_ & n30703;
  assign n30795 = P1_DATAO_REG_18_ & n30700;
  assign n30796 = ~n30794 & ~n30795;
  assign n30797 = P1_EAX_REG_18_ & n30786;
  assign n6654 = ~n30796 | n30797;
  assign n30799 = P1_UWORD_REG_3_ & n30703;
  assign n30800 = P1_DATAO_REG_19_ & n30700;
  assign n30801 = ~n30799 & ~n30800;
  assign n30802 = P1_EAX_REG_19_ & n30786;
  assign n6659 = ~n30801 | n30802;
  assign n30804 = P1_UWORD_REG_4_ & n30703;
  assign n30805 = P1_DATAO_REG_20_ & n30700;
  assign n30806 = ~n30804 & ~n30805;
  assign n30807 = P1_EAX_REG_20_ & n30786;
  assign n6664 = ~n30806 | n30807;
  assign n30809 = P1_UWORD_REG_5_ & n30703;
  assign n30810 = P1_DATAO_REG_21_ & n30700;
  assign n30811 = ~n30809 & ~n30810;
  assign n30812 = P1_EAX_REG_21_ & n30786;
  assign n6669 = ~n30811 | n30812;
  assign n30814 = P1_UWORD_REG_6_ & n30703;
  assign n30815 = P1_DATAO_REG_22_ & n30700;
  assign n30816 = ~n30814 & ~n30815;
  assign n30817 = P1_EAX_REG_22_ & n30786;
  assign n6674 = ~n30816 | n30817;
  assign n30819 = P1_UWORD_REG_7_ & n30703;
  assign n30820 = P1_DATAO_REG_23_ & n30700;
  assign n30821 = ~n30819 & ~n30820;
  assign n30822 = P1_EAX_REG_23_ & n30786;
  assign n6679 = ~n30821 | n30822;
  assign n30824 = P1_UWORD_REG_8_ & n30703;
  assign n30825 = P1_DATAO_REG_24_ & n30700;
  assign n30826 = ~n30824 & ~n30825;
  assign n30827 = P1_EAX_REG_24_ & n30786;
  assign n6684 = ~n30826 | n30827;
  assign n30829 = P1_UWORD_REG_9_ & n30703;
  assign n30830 = P1_DATAO_REG_25_ & n30700;
  assign n30831 = ~n30829 & ~n30830;
  assign n30832 = P1_EAX_REG_25_ & n30786;
  assign n6689 = ~n30831 | n30832;
  assign n30834 = P1_UWORD_REG_10_ & n30703;
  assign n30835 = P1_DATAO_REG_26_ & n30700;
  assign n30836 = ~n30834 & ~n30835;
  assign n30837 = P1_EAX_REG_26_ & n30786;
  assign n6694 = ~n30836 | n30837;
  assign n30839 = P1_UWORD_REG_11_ & n30703;
  assign n30840 = P1_DATAO_REG_27_ & n30700;
  assign n30841 = ~n30839 & ~n30840;
  assign n30842 = P1_EAX_REG_27_ & n30786;
  assign n6699 = ~n30841 | n30842;
  assign n30844 = P1_UWORD_REG_12_ & n30703;
  assign n30845 = P1_DATAO_REG_28_ & n30700;
  assign n30846 = ~n30844 & ~n30845;
  assign n30847 = P1_EAX_REG_28_ & n30786;
  assign n6704 = ~n30846 | n30847;
  assign n30849 = P1_UWORD_REG_13_ & n30703;
  assign n30850 = P1_DATAO_REG_29_ & n30700;
  assign n30851 = ~n30849 & ~n30850;
  assign n30852 = P1_EAX_REG_29_ & n30786;
  assign n6709 = ~n30851 | n30852;
  assign n30854 = P1_UWORD_REG_14_ & n30703;
  assign n30855 = P1_DATAO_REG_30_ & n30700;
  assign n30856 = ~n30854 & ~n30855;
  assign n30857 = P1_EAX_REG_30_ & n30786;
  assign n6714 = ~n30856 | n30857;
  assign n6719 = P1_DATAO_REG_31_ & n30700;
  assign n30860 = ~n23741 & n29422;
  assign n30861 = ~n24164 & n30860;
  assign n30862 = n24217 & n24317;
  assign n30863 = n24046 & n30862;
  assign n30864 = ~n30861 & ~n30863;
  assign n30865 = n24184 & n24233;
  assign n30866 = ~n24164 & n30865;
  assign n30867 = n24010 & n24046;
  assign n30868 = n24174 & n30867;
  assign n30869 = ~n30866 & ~n30868;
  assign n30870 = ~n23523 & ~n30869;
  assign n30871 = n30864 & ~n30870;
  assign n30872 = n24313 & ~n30871;
  assign n30873 = ~n23831 & ~n24297;
  assign n30874 = n30872 & ~n30873;
  assign n30875 = ~n28857 & n30874;
  assign n30876 = n30872 & n30873;
  assign n30877 = ~n25089 & n30876;
  assign n30878 = P1_EAX_REG_0_ & ~n30872;
  assign n30879 = ~n30875 & ~n30877;
  assign n6724 = n30878 | ~n30879;
  assign n30881 = ~n28889 & n30874;
  assign n30882 = ~n25067 & n30876;
  assign n30883 = P1_EAX_REG_1_ & ~n30872;
  assign n30884 = ~n30881 & ~n30882;
  assign n6729 = n30883 | ~n30884;
  assign n30886 = P1_EAX_REG_2_ & ~n30872;
  assign n30887 = ~n25045 & n30876;
  assign n30888 = n28924 & n30874;
  assign n30889 = ~n30886 & ~n30887;
  assign n6734 = n30888 | ~n30889;
  assign n30891 = P1_EAX_REG_3_ & ~n30872;
  assign n30892 = ~n25023 & n30876;
  assign n30893 = n28957 & n30874;
  assign n30894 = ~n30891 & ~n30892;
  assign n6739 = n30893 | ~n30894;
  assign n30896 = P1_EAX_REG_4_ & ~n30872;
  assign n30897 = ~n25001 & n30876;
  assign n30898 = ~n28997 & n30874;
  assign n30899 = ~n30896 & ~n30897;
  assign n6744 = n30898 | ~n30899;
  assign n30901 = P1_EAX_REG_5_ & ~n30872;
  assign n30902 = ~n24979 & n30876;
  assign n30903 = ~n29030 & n30874;
  assign n30904 = ~n30901 & ~n30902;
  assign n6749 = n30903 | ~n30904;
  assign n30906 = P1_EAX_REG_6_ & ~n30872;
  assign n30907 = ~n24957 & n30876;
  assign n30908 = n29061 & n30874;
  assign n30909 = ~n30906 & ~n30907;
  assign n6754 = n30908 | ~n30909;
  assign n30911 = P1_EAX_REG_7_ & ~n30872;
  assign n30912 = ~n24929 & n30876;
  assign n30913 = n29090 & n30874;
  assign n30914 = ~n30911 & ~n30912;
  assign n6759 = n30913 | ~n30914;
  assign n30916 = P1_EAX_REG_8_ & ~n30872;
  assign n30917 = ~n30564 & n30876;
  assign n30918 = ~n29128 & n30874;
  assign n30919 = ~n30916 & ~n30917;
  assign n6764 = n30918 | ~n30919;
  assign n30921 = P1_EAX_REG_9_ & ~n30872;
  assign n30922 = ~n30555 & n30876;
  assign n30923 = ~n29158 & n30874;
  assign n30924 = ~n30921 & ~n30922;
  assign n6769 = n30923 | ~n30924;
  assign n30926 = P1_EAX_REG_10_ & ~n30872;
  assign n30927 = ~n30546 & n30876;
  assign n30928 = n29189 & n30874;
  assign n30929 = ~n30926 & ~n30927;
  assign n6774 = n30928 | ~n30929;
  assign n30931 = P1_EAX_REG_11_ & ~n30872;
  assign n30932 = ~n30537 & n30876;
  assign n30933 = n29219 & n30874;
  assign n30934 = ~n30931 & ~n30932;
  assign n6779 = n30933 | ~n30934;
  assign n30936 = P1_EAX_REG_12_ & ~n30872;
  assign n30937 = ~n30528 & n30876;
  assign n30938 = ~n29259 & n30874;
  assign n30939 = ~n30936 & ~n30937;
  assign n6784 = n30938 | ~n30939;
  assign n30941 = P1_EAX_REG_13_ & ~n30872;
  assign n30942 = ~n30519 & n30876;
  assign n30943 = ~n29289 & n30874;
  assign n30944 = ~n30941 & ~n30942;
  assign n6789 = n30943 | ~n30944;
  assign n30946 = P1_EAX_REG_14_ & ~n30872;
  assign n30947 = ~n30510 & n30876;
  assign n30948 = n29320 & n30874;
  assign n30949 = ~n30946 & ~n30947;
  assign n6794 = n30948 | ~n30949;
  assign n30951 = P1_EAX_REG_15_ & ~n30872;
  assign n30952 = ~n30494 & n30876;
  assign n30953 = n29350 & n30874;
  assign n30954 = ~n30951 & ~n30952;
  assign n6799 = n30953 | ~n30954;
  assign n30956 = ~n23831 & n23896;
  assign n30957 = n30872 & n30956;
  assign n30958 = ~n25089 & n30957;
  assign n30959 = n24240 & n30872;
  assign n30960 = ~n25094 & n30959;
  assign n30961 = P1_EAX_REG_16_ & ~n30872;
  assign n30962 = ~n29454 & n30874;
  assign n30963 = ~n30958 & ~n30960;
  assign n30964 = ~n30961 & n30963;
  assign n6804 = n30962 | ~n30964;
  assign n30966 = ~n25067 & n30957;
  assign n30967 = ~n25072 & n30959;
  assign n30968 = P1_EAX_REG_17_ & ~n30872;
  assign n30969 = ~n29518 & n30874;
  assign n30970 = ~n30966 & ~n30967;
  assign n30971 = ~n30968 & n30970;
  assign n6809 = n30969 | ~n30971;
  assign n30973 = ~n25045 & n30957;
  assign n30974 = ~n25050 & n30959;
  assign n30975 = P1_EAX_REG_18_ & ~n30872;
  assign n30976 = ~n29584 & n30874;
  assign n30977 = ~n30973 & ~n30974;
  assign n30978 = ~n30975 & n30977;
  assign n6814 = n30976 | ~n30978;
  assign n30980 = ~n25023 & n30957;
  assign n30981 = ~n25028 & n30959;
  assign n30982 = P1_EAX_REG_19_ & ~n30872;
  assign n30983 = ~n29650 & n30874;
  assign n30984 = ~n30980 & ~n30981;
  assign n30985 = ~n30982 & n30984;
  assign n6819 = n30983 | ~n30985;
  assign n30987 = ~n25001 & n30957;
  assign n30988 = ~n25006 & n30959;
  assign n30989 = P1_EAX_REG_20_ & ~n30872;
  assign n30990 = ~n29713 & n30874;
  assign n30991 = ~n30987 & ~n30988;
  assign n30992 = ~n30989 & n30991;
  assign n6824 = n30990 | ~n30992;
  assign n30994 = ~n24979 & n30957;
  assign n30995 = ~n24984 & n30959;
  assign n30996 = P1_EAX_REG_21_ & ~n30872;
  assign n30997 = ~n29779 & n30874;
  assign n30998 = ~n30994 & ~n30995;
  assign n30999 = ~n30996 & n30998;
  assign n6829 = n30997 | ~n30999;
  assign n31001 = ~n24957 & n30957;
  assign n31002 = ~n24962 & n30959;
  assign n31003 = P1_EAX_REG_22_ & ~n30872;
  assign n31004 = ~n29845 & n30874;
  assign n31005 = ~n31001 & ~n31002;
  assign n31006 = ~n31003 & n31005;
  assign n6834 = n31004 | ~n31006;
  assign n31008 = ~n24929 & n30957;
  assign n31009 = ~n24939 & n30959;
  assign n31010 = P1_EAX_REG_23_ & ~n30872;
  assign n31011 = ~n29967 & n30874;
  assign n31012 = ~n31008 & ~n31009;
  assign n31013 = ~n31010 & n31012;
  assign n6839 = n31011 | ~n31013;
  assign n31015 = ~n30564 & n30957;
  assign n31016 = ~n25101 & n30959;
  assign n31017 = P1_EAX_REG_24_ & ~n30872;
  assign n31018 = ~n30033 & n30874;
  assign n31019 = ~n31015 & ~n31016;
  assign n31020 = ~n31017 & n31019;
  assign n6844 = n31018 | ~n31020;
  assign n31022 = ~n30555 & n30957;
  assign n31023 = ~n25079 & n30959;
  assign n31024 = P1_EAX_REG_25_ & ~n30872;
  assign n31025 = ~n30103 & n30874;
  assign n31026 = ~n31022 & ~n31023;
  assign n31027 = ~n31024 & n31026;
  assign n6849 = n31025 | ~n31027;
  assign n31029 = ~n30546 & n30957;
  assign n31030 = ~n25057 & n30959;
  assign n31031 = P1_EAX_REG_26_ & ~n30872;
  assign n31032 = ~n30174 & n30874;
  assign n31033 = ~n31029 & ~n31030;
  assign n31034 = ~n31031 & n31033;
  assign n6854 = n31032 | ~n31034;
  assign n31036 = ~n30537 & n30957;
  assign n31037 = ~n25035 & n30959;
  assign n31038 = P1_EAX_REG_27_ & ~n30872;
  assign n31039 = ~n30244 & n30874;
  assign n31040 = ~n31036 & ~n31037;
  assign n31041 = ~n31038 & n31040;
  assign n6859 = n31039 | ~n31041;
  assign n31043 = ~n30528 & n30957;
  assign n31044 = ~n25013 & n30959;
  assign n31045 = P1_EAX_REG_28_ & ~n30872;
  assign n31046 = ~n30315 & n30874;
  assign n31047 = ~n31043 & ~n31044;
  assign n31048 = ~n31045 & n31047;
  assign n6864 = n31046 | ~n31048;
  assign n31050 = ~n30519 & n30957;
  assign n31051 = ~n24991 & n30959;
  assign n31052 = P1_EAX_REG_29_ & ~n30872;
  assign n31053 = ~n30382 & n30874;
  assign n31054 = ~n31050 & ~n31051;
  assign n31055 = ~n31052 & n31054;
  assign n6869 = n31053 | ~n31055;
  assign n31057 = ~n30510 & n30957;
  assign n31058 = ~n24969 & n30959;
  assign n31059 = P1_EAX_REG_30_ & ~n30872;
  assign n31060 = ~n30449 & n30874;
  assign n31061 = ~n31057 & ~n31058;
  assign n31062 = ~n31059 & n31061;
  assign n6874 = n31060 | ~n31062;
  assign n31064 = n23831 & n30486;
  assign n31065 = n30872 & n31064;
  assign n31066 = P1_EAX_REG_31_ & ~n30872;
  assign n31067 = ~n31065 & ~n31066;
  assign n31068 = ~n24947 & n30959;
  assign n6879 = ~n31067 | n31068;
  assign n31070 = P1_STATE2_REG_0_ & ~n23709;
  assign n31071 = n24002 & n31070;
  assign n31072 = n24304 & n31071;
  assign n31073 = n24317 & n31072;
  assign n31074 = n24164 & n29421;
  assign n31075 = ~n31073 & ~n31074;
  assign n31076 = n24313 & ~n31075;
  assign n31077 = n23831 & n31076;
  assign n31078 = ~n26666 & n31077;
  assign n31079 = ~n23831 & n31076;
  assign n31080 = ~n28857 & n31079;
  assign n31081 = P1_EBX_REG_0_ & ~n31076;
  assign n31082 = ~n31078 & ~n31080;
  assign n6884 = n31081 | ~n31082;
  assign n31084 = ~n26720 & n31077;
  assign n31085 = P1_EBX_REG_1_ & ~n31076;
  assign n31086 = ~n28889 & n31079;
  assign n31087 = ~n31084 & ~n31085;
  assign n6889 = n31086 | ~n31087;
  assign n31089 = n26770 & n31077;
  assign n31090 = P1_EBX_REG_2_ & ~n31076;
  assign n31091 = n28924 & n31079;
  assign n31092 = ~n31089 & ~n31090;
  assign n6894 = n31091 | ~n31092;
  assign n31094 = ~n26797 & n31077;
  assign n31095 = P1_EBX_REG_3_ & ~n31076;
  assign n31096 = n28957 & n31079;
  assign n31097 = ~n31094 & ~n31095;
  assign n6899 = n31096 | ~n31097;
  assign n31099 = ~n26848 & n31077;
  assign n31100 = P1_EBX_REG_4_ & ~n31076;
  assign n31101 = ~n28997 & n31079;
  assign n31102 = ~n31099 & ~n31100;
  assign n6904 = n31101 | ~n31102;
  assign n31104 = ~n26951 & n31077;
  assign n31105 = P1_EBX_REG_5_ & ~n31076;
  assign n31106 = ~n29030 & n31079;
  assign n31107 = ~n31104 & ~n31105;
  assign n6909 = n31106 | ~n31107;
  assign n31109 = ~n27060 & n31077;
  assign n31110 = P1_EBX_REG_6_ & ~n31076;
  assign n31111 = n29061 & n31079;
  assign n31112 = ~n31109 & ~n31110;
  assign n6914 = n31111 | ~n31112;
  assign n31114 = ~n27162 & n31077;
  assign n31115 = P1_EBX_REG_7_ & ~n31076;
  assign n31116 = n29090 & n31079;
  assign n31117 = ~n31114 & ~n31115;
  assign n6919 = n31116 | ~n31117;
  assign n31119 = ~n27244 & n31077;
  assign n31120 = P1_EBX_REG_8_ & ~n31076;
  assign n31121 = ~n29128 & n31079;
  assign n31122 = ~n31119 & ~n31120;
  assign n6924 = n31121 | ~n31122;
  assign n31124 = ~n27363 & n31077;
  assign n31125 = P1_EBX_REG_9_ & ~n31076;
  assign n31126 = ~n29158 & n31079;
  assign n31127 = ~n31124 & ~n31125;
  assign n6929 = n31126 | ~n31127;
  assign n31129 = ~n27452 & n31077;
  assign n31130 = P1_EBX_REG_10_ & ~n31076;
  assign n31131 = n29189 & n31079;
  assign n31132 = ~n31129 & ~n31130;
  assign n6934 = n31131 | ~n31132;
  assign n31134 = ~n27540 & n31077;
  assign n31135 = P1_EBX_REG_11_ & ~n31076;
  assign n31136 = n29219 & n31079;
  assign n31137 = ~n31134 & ~n31135;
  assign n6939 = n31136 | ~n31137;
  assign n31139 = ~n27636 & n31077;
  assign n31140 = P1_EBX_REG_12_ & ~n31076;
  assign n31141 = ~n29259 & n31079;
  assign n31142 = ~n31139 & ~n31140;
  assign n6944 = n31141 | ~n31142;
  assign n31144 = ~n27737 & n31077;
  assign n31145 = P1_EBX_REG_13_ & ~n31076;
  assign n31146 = ~n29289 & n31079;
  assign n31147 = ~n31144 & ~n31145;
  assign n6949 = n31146 | ~n31147;
  assign n31149 = ~n27824 & n31077;
  assign n31150 = P1_EBX_REG_14_ & ~n31076;
  assign n31151 = n29320 & n31079;
  assign n31152 = ~n31149 & ~n31150;
  assign n6954 = n31151 | ~n31152;
  assign n31154 = ~n27912 & n31077;
  assign n31155 = P1_EBX_REG_15_ & ~n31076;
  assign n31156 = n29350 & n31079;
  assign n31157 = ~n31154 & ~n31155;
  assign n6959 = n31156 | ~n31157;
  assign n31159 = ~n28002 & n31077;
  assign n31160 = P1_EBX_REG_16_ & ~n31076;
  assign n31161 = ~n29454 & n31079;
  assign n31162 = ~n31159 & ~n31160;
  assign n6964 = n31161 | ~n31162;
  assign n31164 = ~n28063 & n31077;
  assign n31165 = P1_EBX_REG_17_ & ~n31076;
  assign n31166 = ~n29518 & n31079;
  assign n31167 = ~n31164 & ~n31165;
  assign n6969 = n31166 | ~n31167;
  assign n31169 = ~n28110 & n31077;
  assign n31170 = P1_EBX_REG_18_ & ~n31076;
  assign n31171 = ~n29584 & n31079;
  assign n31172 = ~n31169 & ~n31170;
  assign n6974 = n31171 | ~n31172;
  assign n31174 = ~n28159 & n31077;
  assign n31175 = P1_EBX_REG_19_ & ~n31076;
  assign n31176 = ~n29650 & n31079;
  assign n31177 = ~n31174 & ~n31175;
  assign n6979 = n31176 | ~n31177;
  assign n31179 = ~n28208 & n31077;
  assign n31180 = P1_EBX_REG_20_ & ~n31076;
  assign n31181 = ~n29713 & n31079;
  assign n31182 = ~n31179 & ~n31180;
  assign n6984 = n31181 | ~n31182;
  assign n31184 = ~n28254 & n31077;
  assign n31185 = P1_EBX_REG_21_ & ~n31076;
  assign n31186 = ~n29779 & n31079;
  assign n31187 = ~n31184 & ~n31185;
  assign n6989 = n31186 | ~n31187;
  assign n31189 = ~n28302 & n31077;
  assign n31190 = P1_EBX_REG_22_ & ~n31076;
  assign n31191 = ~n29845 & n31079;
  assign n31192 = ~n31189 & ~n31190;
  assign n6994 = n31191 | ~n31192;
  assign n31194 = ~n28351 & n31077;
  assign n31195 = P1_EBX_REG_23_ & ~n31076;
  assign n31196 = ~n29967 & n31079;
  assign n31197 = ~n31194 & ~n31195;
  assign n6999 = n31196 | ~n31197;
  assign n31199 = ~n28407 & n31077;
  assign n31200 = P1_EBX_REG_24_ & ~n31076;
  assign n31201 = ~n30033 & n31079;
  assign n31202 = ~n31199 & ~n31200;
  assign n7004 = n31201 | ~n31202;
  assign n31204 = ~n28453 & n31077;
  assign n31205 = P1_EBX_REG_25_ & ~n31076;
  assign n31206 = ~n30103 & n31079;
  assign n31207 = ~n31204 & ~n31205;
  assign n7009 = n31206 | ~n31207;
  assign n31209 = ~n28501 & n31077;
  assign n31210 = P1_EBX_REG_26_ & ~n31076;
  assign n31211 = ~n30174 & n31079;
  assign n31212 = ~n31209 & ~n31210;
  assign n7014 = n31211 | ~n31212;
  assign n31214 = ~n28550 & n31077;
  assign n31215 = P1_EBX_REG_27_ & ~n31076;
  assign n31216 = ~n30244 & n31079;
  assign n31217 = ~n31214 & ~n31215;
  assign n7019 = n31216 | ~n31217;
  assign n31219 = ~n28599 & n31077;
  assign n31220 = P1_EBX_REG_28_ & ~n31076;
  assign n31221 = ~n30315 & n31079;
  assign n31222 = ~n31219 & ~n31220;
  assign n7024 = n31221 | ~n31222;
  assign n31224 = ~n28649 & n31077;
  assign n31225 = P1_EBX_REG_29_ & ~n31076;
  assign n31226 = ~n30382 & n31079;
  assign n31227 = ~n31224 & ~n31225;
  assign n7029 = n31226 | ~n31227;
  assign n31229 = ~n28714 & n31077;
  assign n31230 = P1_EBX_REG_30_ & ~n31076;
  assign n31231 = ~n30449 & n31079;
  assign n31232 = ~n31229 & ~n31230;
  assign n7034 = n31231 | ~n31232;
  assign n31234 = P1_EBX_REG_31_ & ~n31076;
  assign n31235 = ~n28770 & n31077;
  assign n7039 = n31234 | n31235;
  assign n31237 = ~n24164 & n24454;
  assign n31238 = n24174 & n24238;
  assign n31239 = n24179 & n24576;
  assign n31240 = n24184 & n31239;
  assign n31241 = ~n31237 & ~n31238;
  assign n31242 = ~n31240 & n31241;
  assign n31243 = n24313 & ~n31242;
  assign n31244 = ~n24586 & ~n24614;
  assign n31245 = ~n26598 & n31244;
  assign n31246 = ~n31243 & n31245;
  assign n31247 = P1_STATE2_REG_2_ & ~n31246;
  assign n31248 = n24054 & n31247;
  assign n31249 = n24195 & n31248;
  assign n31250 = n24556 & n31249;
  assign n31251 = n24051 & n31247;
  assign n31252 = n24556 & n31251;
  assign n31253 = ~n31250 & ~n31252;
  assign n31254 = P1_REIP_REG_0_ & ~n31253;
  assign n31255 = ~n24556 & n31251;
  assign n31256 = P1_EBX_REG_31_ & n31255;
  assign n31257 = ~n26666 & n31256;
  assign n31258 = ~P1_EBX_REG_31_ & n31255;
  assign n31259 = ~n24195 & n31248;
  assign n31260 = ~n24556 & n31249;
  assign n31261 = ~n31258 & ~n31259;
  assign n31262 = ~n31260 & n31261;
  assign n31263 = P1_EBX_REG_0_ & ~n31262;
  assign n31264 = P1_STATE2_REG_3_ & ~n31246;
  assign n31265 = P1_PHYADDRPOINTER_REG_0_ & n31264;
  assign n31266 = n23678 & n26631;
  assign n31267 = ~n31246 & n31266;
  assign n31268 = ~n24520 & n31267;
  assign n31269 = P1_REIP_REG_0_ & n31246;
  assign n31270 = P1_STATE2_REG_1_ & ~n31246;
  assign n31271 = n30459 & n31270;
  assign n31272 = P1_PHYADDRPOINTER_REG_0_ & n31271;
  assign n31273 = P1_STATE2_REG_1_ & ~n30459;
  assign n31274 = P1_STATE2_REG_2_ & n23710;
  assign n31275 = ~n31273 & ~n31274;
  assign n31276 = ~n31246 & ~n31275;
  assign n31277 = ~n28857 & n31276;
  assign n31278 = ~n31265 & ~n31268;
  assign n31279 = ~n31269 & n31278;
  assign n31280 = ~n31272 & n31279;
  assign n31281 = ~n31277 & n31280;
  assign n31282 = ~n31254 & ~n31257;
  assign n31283 = ~n31263 & n31282;
  assign n7044 = ~n31281 | ~n31283;
  assign n31285 = ~P1_REIP_REG_1_ & ~n31253;
  assign n31286 = ~n26720 & n31256;
  assign n31287 = P1_EBX_REG_1_ & ~n31262;
  assign n31288 = P1_PHYADDRPOINTER_REG_1_ & n31264;
  assign n31289 = ~n24535 & n31267;
  assign n31290 = P1_REIP_REG_1_ & n31246;
  assign n31291 = ~P1_PHYADDRPOINTER_REG_1_ & n31271;
  assign n31292 = ~n28889 & n31276;
  assign n31293 = ~n31288 & ~n31289;
  assign n31294 = ~n31290 & n31293;
  assign n31295 = ~n31291 & n31294;
  assign n31296 = ~n31292 & n31295;
  assign n31297 = ~n31285 & ~n31286;
  assign n31298 = ~n31287 & n31297;
  assign n7049 = ~n31296 | ~n31298;
  assign n31300 = P1_REIP_REG_1_ & ~P1_REIP_REG_2_;
  assign n31301 = ~P1_REIP_REG_1_ & P1_REIP_REG_2_;
  assign n31302 = ~n31300 & ~n31301;
  assign n31303 = ~n31253 & ~n31302;
  assign n31304 = n26770 & n31256;
  assign n31305 = P1_EBX_REG_2_ & ~n31262;
  assign n31306 = P1_PHYADDRPOINTER_REG_2_ & n31264;
  assign n31307 = n24397 & n31267;
  assign n31308 = P1_REIP_REG_2_ & n31246;
  assign n31309 = ~n28898 & n31271;
  assign n31310 = n28924 & n31276;
  assign n31311 = ~n31306 & ~n31307;
  assign n31312 = ~n31308 & n31311;
  assign n31313 = ~n31309 & n31312;
  assign n31314 = ~n31310 & n31313;
  assign n31315 = ~n31303 & ~n31304;
  assign n31316 = ~n31305 & n31315;
  assign n7054 = ~n31314 | ~n31316;
  assign n31318 = P1_REIP_REG_1_ & P1_REIP_REG_2_;
  assign n31319 = ~P1_REIP_REG_3_ & n31318;
  assign n31320 = P1_REIP_REG_3_ & ~n31318;
  assign n31321 = ~n31319 & ~n31320;
  assign n31322 = ~n31253 & ~n31321;
  assign n31323 = ~n26797 & n31256;
  assign n31324 = P1_EBX_REG_3_ & ~n31262;
  assign n31325 = P1_PHYADDRPOINTER_REG_3_ & n31264;
  assign n31326 = ~n24482 & n31267;
  assign n31327 = P1_REIP_REG_3_ & n31246;
  assign n31328 = ~n28934 & n31271;
  assign n31329 = n28957 & n31276;
  assign n31330 = ~n31325 & ~n31326;
  assign n31331 = ~n31327 & n31330;
  assign n31332 = ~n31328 & n31331;
  assign n31333 = ~n31329 & n31332;
  assign n31334 = ~n31322 & ~n31323;
  assign n31335 = ~n31324 & n31334;
  assign n7059 = ~n31333 | ~n31335;
  assign n31337 = ~n26848 & n31256;
  assign n31338 = ~P1_STATE2_REG_1_ & n24626;
  assign n31339 = ~n31246 & n31338;
  assign n31340 = ~n31337 & ~n31339;
  assign n31341 = P1_REIP_REG_3_ & n31318;
  assign n31342 = ~P1_REIP_REG_4_ & n31341;
  assign n31343 = P1_REIP_REG_4_ & ~n31341;
  assign n31344 = ~n31342 & ~n31343;
  assign n31345 = ~n31253 & ~n31344;
  assign n31346 = P1_PHYADDRPOINTER_REG_4_ & n31264;
  assign n31347 = ~n24472 & n31267;
  assign n31348 = P1_REIP_REG_4_ & n31246;
  assign n31349 = ~n28967 & n31271;
  assign n31350 = ~n31346 & ~n31347;
  assign n31351 = ~n31348 & n31350;
  assign n31352 = ~n31349 & n31351;
  assign n31353 = ~n28997 & n31276;
  assign n31354 = P1_EBX_REG_4_ & ~n31262;
  assign n31355 = n31340 & ~n31345;
  assign n31356 = n31352 & n31355;
  assign n31357 = ~n31353 & n31356;
  assign n7064 = n31354 | ~n31357;
  assign n31359 = ~n26951 & n31256;
  assign n31360 = ~n31339 & ~n31359;
  assign n31361 = P1_REIP_REG_4_ & n31341;
  assign n31362 = ~P1_REIP_REG_5_ & n31361;
  assign n31363 = P1_REIP_REG_5_ & ~n31361;
  assign n31364 = ~n31362 & ~n31363;
  assign n31365 = ~n31253 & ~n31364;
  assign n31366 = P1_EBX_REG_5_ & ~n31262;
  assign n31367 = P1_PHYADDRPOINTER_REG_5_ & n31264;
  assign n31368 = n29012 & n31267;
  assign n31369 = P1_REIP_REG_5_ & n31246;
  assign n31370 = ~n29007 & n31271;
  assign n31371 = ~n29030 & n31276;
  assign n31372 = ~n31367 & ~n31368;
  assign n31373 = ~n31369 & n31372;
  assign n31374 = ~n31370 & n31373;
  assign n31375 = ~n31371 & n31374;
  assign n31376 = n31360 & ~n31365;
  assign n31377 = ~n31366 & n31376;
  assign n7069 = ~n31375 | ~n31377;
  assign n31379 = P1_REIP_REG_6_ & n31246;
  assign n31380 = P1_PHYADDRPOINTER_REG_6_ & n31264;
  assign n31381 = ~n29040 & n31271;
  assign n31382 = ~n31379 & ~n31380;
  assign n31383 = ~n31381 & n31382;
  assign n31384 = P1_EBX_REG_6_ & ~n31262;
  assign n31385 = ~n27060 & n31256;
  assign n31386 = ~n31339 & ~n31385;
  assign n31387 = P1_REIP_REG_5_ & n31361;
  assign n31388 = ~P1_REIP_REG_6_ & n31387;
  assign n31389 = P1_REIP_REG_6_ & ~n31387;
  assign n31390 = ~n31388 & ~n31389;
  assign n31391 = ~n31253 & ~n31390;
  assign n31392 = ~n30459 & n31270;
  assign n31393 = n29061 & n31392;
  assign n31394 = n31383 & ~n31384;
  assign n31395 = n31386 & n31394;
  assign n31396 = ~n31391 & n31395;
  assign n7074 = n31393 | ~n31396;
  assign n31398 = P1_REIP_REG_7_ & n31246;
  assign n31399 = P1_PHYADDRPOINTER_REG_7_ & n31264;
  assign n31400 = ~n29071 & n31271;
  assign n31401 = ~n31398 & ~n31399;
  assign n31402 = ~n31400 & n31401;
  assign n31403 = P1_EBX_REG_7_ & ~n31262;
  assign n31404 = ~n27162 & n31256;
  assign n31405 = ~n31339 & ~n31404;
  assign n31406 = P1_REIP_REG_6_ & n31387;
  assign n31407 = ~P1_REIP_REG_7_ & n31406;
  assign n31408 = P1_REIP_REG_7_ & ~n31406;
  assign n31409 = ~n31407 & ~n31408;
  assign n31410 = ~n31253 & ~n31409;
  assign n31411 = n29090 & n31392;
  assign n31412 = n31402 & ~n31403;
  assign n31413 = n31405 & n31412;
  assign n31414 = ~n31410 & n31413;
  assign n7079 = n31411 | ~n31414;
  assign n31416 = P1_REIP_REG_8_ & n31246;
  assign n31417 = P1_PHYADDRPOINTER_REG_8_ & n31264;
  assign n31418 = ~n29100 & n31271;
  assign n31419 = ~n31416 & ~n31417;
  assign n31420 = ~n31418 & n31419;
  assign n31421 = P1_EBX_REG_8_ & ~n31262;
  assign n31422 = ~n27244 & n31256;
  assign n31423 = ~n31339 & ~n31422;
  assign n31424 = P1_REIP_REG_7_ & n31406;
  assign n31425 = ~P1_REIP_REG_8_ & n31424;
  assign n31426 = P1_REIP_REG_8_ & ~n31424;
  assign n31427 = ~n31425 & ~n31426;
  assign n31428 = ~n31253 & ~n31427;
  assign n31429 = ~n29128 & n31392;
  assign n31430 = n31420 & ~n31421;
  assign n31431 = n31423 & n31430;
  assign n31432 = ~n31428 & n31431;
  assign n7084 = n31429 | ~n31432;
  assign n31434 = P1_REIP_REG_9_ & n31246;
  assign n31435 = P1_PHYADDRPOINTER_REG_9_ & n31264;
  assign n31436 = ~n29138 & n31271;
  assign n31437 = ~n31434 & ~n31435;
  assign n31438 = ~n31436 & n31437;
  assign n31439 = P1_EBX_REG_9_ & ~n31262;
  assign n31440 = ~n27363 & n31256;
  assign n31441 = ~n31339 & ~n31440;
  assign n31442 = P1_REIP_REG_8_ & n31424;
  assign n31443 = ~P1_REIP_REG_9_ & n31442;
  assign n31444 = P1_REIP_REG_9_ & ~n31442;
  assign n31445 = ~n31443 & ~n31444;
  assign n31446 = ~n31253 & ~n31445;
  assign n31447 = ~n29158 & n31392;
  assign n31448 = n31438 & ~n31439;
  assign n31449 = n31441 & n31448;
  assign n31450 = ~n31446 & n31449;
  assign n7089 = n31447 | ~n31450;
  assign n31452 = P1_REIP_REG_10_ & n31246;
  assign n31453 = P1_PHYADDRPOINTER_REG_10_ & n31264;
  assign n31454 = ~n29168 & n31271;
  assign n31455 = ~n31452 & ~n31453;
  assign n31456 = ~n31454 & n31455;
  assign n31457 = P1_EBX_REG_10_ & ~n31262;
  assign n31458 = ~n27452 & n31256;
  assign n31459 = ~n31339 & ~n31458;
  assign n31460 = P1_REIP_REG_9_ & n31442;
  assign n31461 = ~P1_REIP_REG_10_ & n31460;
  assign n31462 = P1_REIP_REG_10_ & ~n31460;
  assign n31463 = ~n31461 & ~n31462;
  assign n31464 = ~n31253 & ~n31463;
  assign n31465 = n29189 & n31392;
  assign n31466 = n31456 & ~n31457;
  assign n31467 = n31459 & n31466;
  assign n31468 = ~n31464 & n31467;
  assign n7094 = n31465 | ~n31468;
  assign n31470 = P1_REIP_REG_11_ & n31246;
  assign n31471 = P1_PHYADDRPOINTER_REG_11_ & n31264;
  assign n31472 = ~n29199 & n31271;
  assign n31473 = ~n31470 & ~n31471;
  assign n31474 = ~n31472 & n31473;
  assign n31475 = P1_EBX_REG_11_ & ~n31262;
  assign n31476 = ~n27540 & n31256;
  assign n31477 = ~n31339 & ~n31476;
  assign n31478 = P1_REIP_REG_10_ & n31460;
  assign n31479 = ~P1_REIP_REG_11_ & n31478;
  assign n31480 = P1_REIP_REG_11_ & ~n31478;
  assign n31481 = ~n31479 & ~n31480;
  assign n31482 = ~n31253 & ~n31481;
  assign n31483 = n29219 & n31392;
  assign n31484 = n31474 & ~n31475;
  assign n31485 = n31477 & n31484;
  assign n31486 = ~n31482 & n31485;
  assign n7099 = n31483 | ~n31486;
  assign n31488 = P1_REIP_REG_12_ & n31246;
  assign n31489 = P1_PHYADDRPOINTER_REG_12_ & n31264;
  assign n31490 = ~n29229 & n31271;
  assign n31491 = ~n31488 & ~n31489;
  assign n31492 = ~n31490 & n31491;
  assign n31493 = P1_EBX_REG_12_ & ~n31262;
  assign n31494 = ~n27636 & n31256;
  assign n31495 = ~n31339 & ~n31494;
  assign n31496 = P1_REIP_REG_11_ & n31478;
  assign n31497 = ~P1_REIP_REG_12_ & n31496;
  assign n31498 = P1_REIP_REG_12_ & ~n31496;
  assign n31499 = ~n31497 & ~n31498;
  assign n31500 = ~n31253 & ~n31499;
  assign n31501 = ~n29259 & n31392;
  assign n31502 = n31492 & ~n31493;
  assign n31503 = n31495 & n31502;
  assign n31504 = ~n31500 & n31503;
  assign n7104 = n31501 | ~n31504;
  assign n31506 = P1_REIP_REG_13_ & n31246;
  assign n31507 = P1_PHYADDRPOINTER_REG_13_ & n31264;
  assign n31508 = ~n29269 & n31271;
  assign n31509 = ~n31506 & ~n31507;
  assign n31510 = ~n31508 & n31509;
  assign n31511 = P1_EBX_REG_13_ & ~n31262;
  assign n31512 = ~n27737 & n31256;
  assign n31513 = ~n31339 & ~n31512;
  assign n31514 = P1_REIP_REG_12_ & n31496;
  assign n31515 = ~P1_REIP_REG_13_ & n31514;
  assign n31516 = P1_REIP_REG_13_ & ~n31514;
  assign n31517 = ~n31515 & ~n31516;
  assign n31518 = ~n31253 & ~n31517;
  assign n31519 = ~n29289 & n31392;
  assign n31520 = n31510 & ~n31511;
  assign n31521 = n31513 & n31520;
  assign n31522 = ~n31518 & n31521;
  assign n7109 = n31519 | ~n31522;
  assign n31524 = P1_REIP_REG_14_ & n31246;
  assign n31525 = P1_PHYADDRPOINTER_REG_14_ & n31264;
  assign n31526 = ~n29299 & n31271;
  assign n31527 = ~n31524 & ~n31525;
  assign n31528 = ~n31526 & n31527;
  assign n31529 = P1_EBX_REG_14_ & ~n31262;
  assign n31530 = ~n27824 & n31256;
  assign n31531 = ~n31339 & ~n31530;
  assign n31532 = P1_REIP_REG_13_ & n31514;
  assign n31533 = ~P1_REIP_REG_14_ & n31532;
  assign n31534 = P1_REIP_REG_14_ & ~n31532;
  assign n31535 = ~n31533 & ~n31534;
  assign n31536 = ~n31253 & ~n31535;
  assign n31537 = n29320 & n31392;
  assign n31538 = n31528 & ~n31529;
  assign n31539 = n31531 & n31538;
  assign n31540 = ~n31536 & n31539;
  assign n7114 = n31537 | ~n31540;
  assign n31542 = P1_EBX_REG_15_ & ~n31262;
  assign n31543 = P1_REIP_REG_14_ & n31532;
  assign n31544 = ~P1_REIP_REG_15_ & n31543;
  assign n31545 = P1_REIP_REG_15_ & ~n31543;
  assign n31546 = ~n31544 & ~n31545;
  assign n31547 = ~n31253 & ~n31546;
  assign n31548 = P1_REIP_REG_15_ & n31246;
  assign n31549 = P1_PHYADDRPOINTER_REG_15_ & n31264;
  assign n31550 = ~n29330 & n31271;
  assign n31551 = ~n31548 & ~n31549;
  assign n31552 = ~n31550 & n31551;
  assign n31553 = ~n27912 & n31256;
  assign n31554 = ~n31339 & ~n31553;
  assign n31555 = n29350 & n31392;
  assign n31556 = ~n31542 & ~n31547;
  assign n31557 = n31552 & n31556;
  assign n31558 = n31554 & n31557;
  assign n7119 = n31555 | ~n31558;
  assign n31560 = P1_EBX_REG_16_ & ~n31262;
  assign n31561 = P1_REIP_REG_15_ & n31543;
  assign n31562 = ~P1_REIP_REG_16_ & n31561;
  assign n31563 = P1_REIP_REG_16_ & ~n31561;
  assign n31564 = ~n31562 & ~n31563;
  assign n31565 = ~n31253 & ~n31564;
  assign n31566 = P1_REIP_REG_16_ & n31246;
  assign n31567 = P1_PHYADDRPOINTER_REG_16_ & n31264;
  assign n31568 = ~n29360 & n31271;
  assign n31569 = ~n31566 & ~n31567;
  assign n31570 = ~n31568 & n31569;
  assign n31571 = ~n28002 & n31256;
  assign n31572 = ~n31339 & ~n31571;
  assign n31573 = ~n29454 & n31392;
  assign n31574 = ~n31560 & ~n31565;
  assign n31575 = n31570 & n31574;
  assign n31576 = n31572 & n31575;
  assign n7124 = n31573 | ~n31576;
  assign n31578 = P1_REIP_REG_16_ & n31561;
  assign n31579 = ~P1_REIP_REG_17_ & n31578;
  assign n31580 = P1_REIP_REG_17_ & ~n31578;
  assign n31581 = ~n31579 & ~n31580;
  assign n31582 = ~n31253 & ~n31581;
  assign n31583 = ~n31339 & ~n31582;
  assign n31584 = P1_EBX_REG_17_ & ~n31262;
  assign n31585 = P1_REIP_REG_17_ & n31246;
  assign n31586 = P1_PHYADDRPOINTER_REG_17_ & n31264;
  assign n31587 = ~n29464 & n31271;
  assign n31588 = ~n31585 & ~n31586;
  assign n31589 = ~n31587 & n31588;
  assign n31590 = ~n28063 & n31256;
  assign n31591 = ~n29518 & n31392;
  assign n31592 = n31583 & ~n31584;
  assign n31593 = n31589 & n31592;
  assign n31594 = ~n31590 & n31593;
  assign n7129 = n31591 | ~n31594;
  assign n31596 = P1_REIP_REG_17_ & n31578;
  assign n31597 = ~P1_REIP_REG_18_ & n31596;
  assign n31598 = P1_REIP_REG_18_ & ~n31596;
  assign n31599 = ~n31597 & ~n31598;
  assign n31600 = ~n31253 & ~n31599;
  assign n31601 = ~n31339 & ~n31600;
  assign n31602 = P1_EBX_REG_18_ & ~n31262;
  assign n31603 = P1_REIP_REG_18_ & n31246;
  assign n31604 = P1_PHYADDRPOINTER_REG_18_ & n31264;
  assign n31605 = ~n29528 & n31271;
  assign n31606 = ~n31603 & ~n31604;
  assign n31607 = ~n31605 & n31606;
  assign n31608 = ~n28110 & n31256;
  assign n31609 = ~n29584 & n31392;
  assign n31610 = n31601 & ~n31602;
  assign n31611 = n31607 & n31610;
  assign n31612 = ~n31608 & n31611;
  assign n7134 = n31609 | ~n31612;
  assign n31614 = P1_REIP_REG_18_ & n31596;
  assign n31615 = ~P1_REIP_REG_19_ & n31614;
  assign n31616 = P1_REIP_REG_19_ & ~n31614;
  assign n31617 = ~n31615 & ~n31616;
  assign n31618 = ~n31253 & ~n31617;
  assign n31619 = ~n31339 & ~n31618;
  assign n31620 = P1_EBX_REG_19_ & ~n31262;
  assign n31621 = P1_REIP_REG_19_ & n31246;
  assign n31622 = P1_PHYADDRPOINTER_REG_19_ & n31264;
  assign n31623 = ~n29594 & n31271;
  assign n31624 = ~n31621 & ~n31622;
  assign n31625 = ~n31623 & n31624;
  assign n31626 = ~n28159 & n31256;
  assign n31627 = ~n29650 & n31392;
  assign n31628 = n31619 & ~n31620;
  assign n31629 = n31625 & n31628;
  assign n31630 = ~n31626 & n31629;
  assign n7139 = n31627 | ~n31630;
  assign n31632 = P1_EBX_REG_20_ & ~n31262;
  assign n31633 = P1_PHYADDRPOINTER_REG_20_ & n31264;
  assign n31634 = P1_REIP_REG_19_ & n31614;
  assign n31635 = ~P1_REIP_REG_20_ & n31634;
  assign n31636 = P1_REIP_REG_20_ & ~n31634;
  assign n31637 = ~n31635 & ~n31636;
  assign n31638 = ~n31253 & ~n31637;
  assign n31639 = ~n31633 & ~n31638;
  assign n31640 = ~n29660 & n31271;
  assign n31641 = P1_REIP_REG_20_ & n31246;
  assign n31642 = ~n31640 & ~n31641;
  assign n31643 = ~n28208 & n31256;
  assign n31644 = ~n29713 & n31392;
  assign n31645 = ~n31632 & n31639;
  assign n31646 = n31642 & n31645;
  assign n31647 = ~n31643 & n31646;
  assign n7144 = n31644 | ~n31647;
  assign n31649 = P1_EBX_REG_21_ & ~n31262;
  assign n31650 = P1_PHYADDRPOINTER_REG_21_ & n31264;
  assign n31651 = P1_REIP_REG_20_ & n31634;
  assign n31652 = ~P1_REIP_REG_21_ & n31651;
  assign n31653 = P1_REIP_REG_21_ & ~n31651;
  assign n31654 = ~n31652 & ~n31653;
  assign n31655 = ~n31253 & ~n31654;
  assign n31656 = ~n31650 & ~n31655;
  assign n31657 = ~n29723 & n31271;
  assign n31658 = P1_REIP_REG_21_ & n31246;
  assign n31659 = ~n31657 & ~n31658;
  assign n31660 = ~n28254 & n31256;
  assign n31661 = ~n29779 & n31392;
  assign n31662 = ~n31649 & n31656;
  assign n31663 = n31659 & n31662;
  assign n31664 = ~n31660 & n31663;
  assign n7149 = n31661 | ~n31664;
  assign n31666 = P1_EBX_REG_22_ & ~n31262;
  assign n31667 = P1_PHYADDRPOINTER_REG_22_ & n31264;
  assign n31668 = P1_REIP_REG_21_ & n31651;
  assign n31669 = ~P1_REIP_REG_22_ & n31668;
  assign n31670 = P1_REIP_REG_22_ & ~n31668;
  assign n31671 = ~n31669 & ~n31670;
  assign n31672 = ~n31253 & ~n31671;
  assign n31673 = ~n31667 & ~n31672;
  assign n31674 = ~n29789 & n31271;
  assign n31675 = P1_REIP_REG_22_ & n31246;
  assign n31676 = ~n31674 & ~n31675;
  assign n31677 = ~n28302 & n31256;
  assign n31678 = ~n29845 & n31392;
  assign n31679 = ~n31666 & n31673;
  assign n31680 = n31676 & n31679;
  assign n31681 = ~n31677 & n31680;
  assign n7154 = n31678 | ~n31681;
  assign n31683 = P1_EBX_REG_23_ & ~n31262;
  assign n31684 = P1_PHYADDRPOINTER_REG_23_ & n31264;
  assign n31685 = P1_REIP_REG_22_ & n31668;
  assign n31686 = ~P1_REIP_REG_23_ & n31685;
  assign n31687 = P1_REIP_REG_23_ & ~n31685;
  assign n31688 = ~n31686 & ~n31687;
  assign n31689 = ~n31253 & ~n31688;
  assign n31690 = ~n31684 & ~n31689;
  assign n31691 = ~n29855 & n31271;
  assign n31692 = P1_REIP_REG_23_ & n31246;
  assign n31693 = ~n31691 & ~n31692;
  assign n31694 = ~n28351 & n31256;
  assign n31695 = ~n29967 & n31392;
  assign n31696 = ~n31683 & n31690;
  assign n31697 = n31693 & n31696;
  assign n31698 = ~n31694 & n31697;
  assign n7159 = n31695 | ~n31698;
  assign n31700 = P1_EBX_REG_24_ & ~n31262;
  assign n31701 = P1_PHYADDRPOINTER_REG_24_ & n31264;
  assign n31702 = P1_REIP_REG_23_ & n31685;
  assign n31703 = ~P1_REIP_REG_24_ & n31702;
  assign n31704 = P1_REIP_REG_24_ & ~n31702;
  assign n31705 = ~n31703 & ~n31704;
  assign n31706 = ~n31253 & ~n31705;
  assign n31707 = ~n31701 & ~n31706;
  assign n31708 = ~n29977 & n31271;
  assign n31709 = P1_REIP_REG_24_ & n31246;
  assign n31710 = ~n31708 & ~n31709;
  assign n31711 = ~n28407 & n31256;
  assign n31712 = ~n30033 & n31392;
  assign n31713 = ~n31700 & n31707;
  assign n31714 = n31710 & n31713;
  assign n31715 = ~n31711 & n31714;
  assign n7164 = n31712 | ~n31715;
  assign n31717 = P1_EBX_REG_25_ & ~n31262;
  assign n31718 = P1_PHYADDRPOINTER_REG_25_ & n31264;
  assign n31719 = P1_REIP_REG_24_ & n31702;
  assign n31720 = ~P1_REIP_REG_25_ & n31719;
  assign n31721 = P1_REIP_REG_25_ & ~n31719;
  assign n31722 = ~n31720 & ~n31721;
  assign n31723 = ~n31253 & ~n31722;
  assign n31724 = ~n31718 & ~n31723;
  assign n31725 = ~n30043 & n31271;
  assign n31726 = P1_REIP_REG_25_ & n31246;
  assign n31727 = ~n31725 & ~n31726;
  assign n31728 = ~n28453 & n31256;
  assign n31729 = ~n30103 & n31392;
  assign n31730 = ~n31717 & n31724;
  assign n31731 = n31727 & n31730;
  assign n31732 = ~n31728 & n31731;
  assign n7169 = n31729 | ~n31732;
  assign n31734 = P1_EBX_REG_26_ & ~n31262;
  assign n31735 = P1_PHYADDRPOINTER_REG_26_ & n31264;
  assign n31736 = P1_REIP_REG_25_ & n31719;
  assign n31737 = ~P1_REIP_REG_26_ & n31736;
  assign n31738 = P1_REIP_REG_26_ & ~n31736;
  assign n31739 = ~n31737 & ~n31738;
  assign n31740 = ~n31253 & ~n31739;
  assign n31741 = ~n31735 & ~n31740;
  assign n31742 = ~n30113 & n31271;
  assign n31743 = P1_REIP_REG_26_ & n31246;
  assign n31744 = ~n31742 & ~n31743;
  assign n31745 = ~n28501 & n31256;
  assign n31746 = ~n30174 & n31392;
  assign n31747 = ~n31734 & n31741;
  assign n31748 = n31744 & n31747;
  assign n31749 = ~n31745 & n31748;
  assign n7174 = n31746 | ~n31749;
  assign n31751 = P1_EBX_REG_27_ & ~n31262;
  assign n31752 = P1_PHYADDRPOINTER_REG_27_ & n31264;
  assign n31753 = P1_REIP_REG_26_ & n31736;
  assign n31754 = ~P1_REIP_REG_27_ & n31753;
  assign n31755 = P1_REIP_REG_27_ & ~n31753;
  assign n31756 = ~n31754 & ~n31755;
  assign n31757 = ~n31253 & ~n31756;
  assign n31758 = ~n31752 & ~n31757;
  assign n31759 = ~n30184 & n31271;
  assign n31760 = P1_REIP_REG_27_ & n31246;
  assign n31761 = ~n31759 & ~n31760;
  assign n31762 = ~n28550 & n31256;
  assign n31763 = ~n30244 & n31392;
  assign n31764 = ~n31751 & n31758;
  assign n31765 = n31761 & n31764;
  assign n31766 = ~n31762 & n31765;
  assign n7179 = n31763 | ~n31766;
  assign n31768 = P1_EBX_REG_28_ & ~n31262;
  assign n31769 = P1_PHYADDRPOINTER_REG_28_ & n31264;
  assign n31770 = P1_REIP_REG_27_ & n31753;
  assign n31771 = ~P1_REIP_REG_28_ & n31770;
  assign n31772 = P1_REIP_REG_28_ & ~n31770;
  assign n31773 = ~n31771 & ~n31772;
  assign n31774 = ~n31253 & ~n31773;
  assign n31775 = ~n31769 & ~n31774;
  assign n31776 = ~n30254 & n31271;
  assign n31777 = P1_REIP_REG_28_ & n31246;
  assign n31778 = ~n31776 & ~n31777;
  assign n31779 = ~n28599 & n31256;
  assign n31780 = ~n30315 & n31392;
  assign n31781 = ~n31768 & n31775;
  assign n31782 = n31778 & n31781;
  assign n31783 = ~n31779 & n31782;
  assign n7184 = n31780 | ~n31783;
  assign n31785 = P1_EBX_REG_29_ & ~n31262;
  assign n31786 = P1_PHYADDRPOINTER_REG_29_ & n31264;
  assign n31787 = P1_REIP_REG_28_ & n31770;
  assign n31788 = ~P1_REIP_REG_29_ & n31787;
  assign n31789 = P1_REIP_REG_29_ & ~n31787;
  assign n31790 = ~n31788 & ~n31789;
  assign n31791 = ~n31253 & ~n31790;
  assign n31792 = ~n31786 & ~n31791;
  assign n31793 = ~n30325 & n31271;
  assign n31794 = P1_REIP_REG_29_ & n31246;
  assign n31795 = ~n31793 & ~n31794;
  assign n31796 = ~n28649 & n31256;
  assign n31797 = ~n30382 & n31392;
  assign n31798 = ~n31785 & n31792;
  assign n31799 = n31795 & n31798;
  assign n31800 = ~n31796 & n31799;
  assign n7189 = n31797 | ~n31800;
  assign n31802 = P1_EBX_REG_30_ & ~n31262;
  assign n31803 = P1_PHYADDRPOINTER_REG_30_ & n31264;
  assign n31804 = P1_REIP_REG_29_ & n31787;
  assign n31805 = ~P1_REIP_REG_30_ & n31804;
  assign n31806 = P1_REIP_REG_30_ & ~n31804;
  assign n31807 = ~n31805 & ~n31806;
  assign n31808 = ~n31253 & ~n31807;
  assign n31809 = ~n31803 & ~n31808;
  assign n31810 = ~n30392 & n31271;
  assign n31811 = P1_REIP_REG_30_ & n31246;
  assign n31812 = ~n31810 & ~n31811;
  assign n31813 = ~n28714 & n31256;
  assign n31814 = ~n30449 & n31392;
  assign n31815 = ~n31802 & n31809;
  assign n31816 = n31812 & n31815;
  assign n31817 = ~n31813 & n31816;
  assign n7194 = n31814 | ~n31817;
  assign n31819 = P1_EBX_REG_31_ & ~n31262;
  assign n31820 = P1_PHYADDRPOINTER_REG_31_ & n31264;
  assign n31821 = P1_REIP_REG_30_ & n31804;
  assign n31822 = ~P1_REIP_REG_31_ & n31821;
  assign n31823 = P1_REIP_REG_31_ & ~n31821;
  assign n31824 = ~n31822 & ~n31823;
  assign n31825 = ~n31253 & ~n31824;
  assign n31826 = ~n31820 & ~n31825;
  assign n31827 = ~n30459 & n31271;
  assign n31828 = P1_REIP_REG_31_ & n31246;
  assign n31829 = ~n31827 & ~n31828;
  assign n31830 = ~n28770 & n31256;
  assign n31831 = n30486 & n31392;
  assign n31832 = ~n31819 & n31826;
  assign n31833 = n31829 & n31832;
  assign n31834 = ~n31830 & n31833;
  assign n7199 = n31831 | ~n31834;
  assign n31836 = ~P1_DATAWIDTH_REG_1_ & ~P1_REIP_REG_1_;
  assign n31837 = ~P1_DATAWIDTH_REG_30_ & ~P1_DATAWIDTH_REG_31_;
  assign n31838 = P1_DATAWIDTH_REG_0_ & P1_DATAWIDTH_REG_1_;
  assign n31839 = ~P1_DATAWIDTH_REG_28_ & ~P1_DATAWIDTH_REG_29_;
  assign n31840 = ~P1_DATAWIDTH_REG_26_ & ~P1_DATAWIDTH_REG_27_;
  assign n31841 = n31837 & ~n31838;
  assign n31842 = n31839 & n31841;
  assign n31843 = n31840 & n31842;
  assign n31844 = ~P1_DATAWIDTH_REG_22_ & ~P1_DATAWIDTH_REG_23_;
  assign n31845 = ~P1_DATAWIDTH_REG_24_ & n31844;
  assign n31846 = ~P1_DATAWIDTH_REG_25_ & n31845;
  assign n31847 = ~P1_DATAWIDTH_REG_18_ & ~P1_DATAWIDTH_REG_19_;
  assign n31848 = ~P1_DATAWIDTH_REG_20_ & n31847;
  assign n31849 = ~P1_DATAWIDTH_REG_21_ & n31848;
  assign n31850 = n31846 & n31849;
  assign n31851 = ~P1_DATAWIDTH_REG_14_ & ~P1_DATAWIDTH_REG_15_;
  assign n31852 = ~P1_DATAWIDTH_REG_16_ & n31851;
  assign n31853 = ~P1_DATAWIDTH_REG_17_ & n31852;
  assign n31854 = ~P1_DATAWIDTH_REG_10_ & ~P1_DATAWIDTH_REG_11_;
  assign n31855 = ~P1_DATAWIDTH_REG_12_ & n31854;
  assign n31856 = ~P1_DATAWIDTH_REG_13_ & n31855;
  assign n31857 = n31853 & n31856;
  assign n31858 = ~P1_DATAWIDTH_REG_6_ & ~P1_DATAWIDTH_REG_7_;
  assign n31859 = ~P1_DATAWIDTH_REG_8_ & n31858;
  assign n31860 = ~P1_DATAWIDTH_REG_9_ & n31859;
  assign n31861 = ~P1_DATAWIDTH_REG_2_ & ~P1_DATAWIDTH_REG_3_;
  assign n31862 = ~P1_DATAWIDTH_REG_4_ & n31861;
  assign n31863 = ~P1_DATAWIDTH_REG_5_ & n31862;
  assign n31864 = n31860 & n31863;
  assign n31865 = n31843 & n31850;
  assign n31866 = n31857 & n31865;
  assign n31867 = n31864 & n31866;
  assign n31868 = n31836 & n31867;
  assign n31869 = P1_BYTEENABLE_REG_3_ & ~n31867;
  assign n31870 = ~P1_DATAWIDTH_REG_0_ & ~P1_REIP_REG_0_;
  assign n31871 = ~P1_DATAWIDTH_REG_1_ & n31870;
  assign n31872 = n31867 & n31871;
  assign n31873 = ~n31868 & ~n31869;
  assign n7204 = n31872 | ~n31873;
  assign n31875 = P1_REIP_REG_0_ & P1_REIP_REG_1_;
  assign n31876 = P1_DATAWIDTH_REG_0_ & ~P1_REIP_REG_0_;
  assign n31877 = ~P1_DATAWIDTH_REG_0_ & ~P1_DATAWIDTH_REG_1_;
  assign n31878 = ~n31876 & ~n31877;
  assign n31879 = ~P1_REIP_REG_1_ & ~n31878;
  assign n31880 = ~n31875 & ~n31879;
  assign n31881 = n31867 & ~n31880;
  assign n31882 = P1_BYTEENABLE_REG_2_ & ~n31867;
  assign n7209 = n31881 | n31882;
  assign n31884 = P1_REIP_REG_1_ & n31867;
  assign n31885 = P1_BYTEENABLE_REG_1_ & ~n31867;
  assign n31886 = ~n31884 & ~n31885;
  assign n7214 = n31872 | ~n31886;
  assign n31888 = ~P1_REIP_REG_0_ & ~P1_REIP_REG_1_;
  assign n31889 = n31867 & ~n31888;
  assign n31890 = P1_BYTEENABLE_REG_0_ & ~n31867;
  assign n7219 = n31889 | n31890;
  assign n31892 = P1_W_R_N_REG & ~n23355;
  assign n31893 = ~P1_READREQUEST_REG & n23355;
  assign n7224 = n31892 | n31893;
  assign n31895 = ~n24199 & n24576;
  assign n31896 = P1_FLUSH_REG & ~n31895;
  assign n7229 = n28821 | n31896;
  assign n31898 = n24178 & n31895;
  assign n31899 = P1_MORE_REG & ~n31895;
  assign n7234 = n31898 | n31899;
  assign n31901 = BS16 & ~n23572;
  assign n31902 = P1_STATEBS16_REG & n23572;
  assign n31903 = ~P1_STATE_REG_0_ & n23526;
  assign n31904 = ~n31901 & ~n31902;
  assign n7239 = n31903 | ~n31904;
  assign n31906 = n24047 & ~n24195;
  assign n31907 = ~n24591 & ~n31906;
  assign n31908 = P1_STATE2_REG_2_ & ~n23523;
  assign n31909 = P1_STATEBS16_REG & n24195;
  assign n31910 = n24054 & ~n31909;
  assign n31911 = n31908 & ~n31910;
  assign n31912 = P1_STATE2_REG_0_ & ~n31911;
  assign n31913 = n31907 & ~n31912;
  assign n31914 = ~P1_STATE2_REG_0_ & ~n23523;
  assign n31915 = n23609 & n31914;
  assign n31916 = ~n24308 & ~n24626;
  assign n31917 = ~n31915 & n31916;
  assign n31918 = ~n31243 & n31917;
  assign n31919 = ~n31913 & ~n31918;
  assign n31920 = P1_REQUESTPENDING_REG & n31918;
  assign n7244 = n31919 | n31920;
  assign n31922 = P1_D_C_N_REG & ~n23355;
  assign n31923 = ~P1_CODEFETCH_REG & n23355;
  assign n31924 = ~n31922 & ~n31923;
  assign n7249 = n31903 | ~n31924;
  assign n31926 = P1_MEMORYFETCH_REG & n23355;
  assign n31927 = P1_M_IO_N_REG & ~n23355;
  assign n7254 = n31926 | n31927;
  assign n31929 = P1_STATE2_REG_0_ & n31338;
  assign n31930 = n24192 & n24576;
  assign n31931 = P1_CODEFETCH_REG & ~n31930;
  assign n7259 = n31929 | n31931;
  assign n31933 = P1_STATE_REG_0_ & P1_ADS_N_REG;
  assign n7264 = ~n23572 | n31933;
  assign n31935 = P1_STATE2_REG_2_ & ~n23710;
  assign n31936 = ~n24167 & n31935;
  assign n31937 = ~n31243 & ~n31338;
  assign n31938 = ~n31936 & ~n31937;
  assign n31939 = P1_READREQUEST_REG & n31937;
  assign n7268 = n31938 | n31939;
  assign n31941 = n24045 & n24313;
  assign n31942 = n24188 & n31941;
  assign n31943 = ~n24190 & n31942;
  assign n31944 = P1_MEMORYFETCH_REG & ~n31943;
  assign n31945 = ~n31338 & ~n31944;
  assign n7273 = n31240 | ~n31945;
  always @ (posedge clock) begin
    BUF1_REG_0_ <= n270;
    BUF1_REG_1_ <= n275;
    BUF1_REG_2_ <= n280;
    BUF1_REG_3_ <= n285;
    BUF1_REG_4_ <= n290;
    BUF1_REG_5_ <= n295;
    BUF1_REG_6_ <= n300;
    BUF1_REG_7_ <= n305;
    BUF1_REG_8_ <= n310;
    BUF1_REG_9_ <= n315;
    BUF1_REG_10_ <= n320;
    BUF1_REG_11_ <= n325;
    BUF1_REG_12_ <= n330;
    BUF1_REG_13_ <= n335;
    BUF1_REG_14_ <= n340;
    BUF1_REG_15_ <= n345;
    BUF1_REG_16_ <= n350;
    BUF1_REG_17_ <= n355;
    BUF1_REG_18_ <= n360;
    BUF1_REG_19_ <= n365;
    BUF1_REG_20_ <= n370;
    BUF1_REG_21_ <= n375;
    BUF1_REG_22_ <= n380;
    BUF1_REG_23_ <= n385;
    BUF1_REG_24_ <= n390;
    BUF1_REG_25_ <= n395;
    BUF1_REG_26_ <= n400;
    BUF1_REG_27_ <= n405;
    BUF1_REG_28_ <= n410;
    BUF1_REG_29_ <= n415;
    BUF1_REG_30_ <= n420;
    BUF1_REG_31_ <= n425;
    BUF2_REG_0_ <= n430;
    BUF2_REG_1_ <= n435;
    BUF2_REG_2_ <= n440;
    BUF2_REG_3_ <= n445;
    BUF2_REG_4_ <= n450;
    BUF2_REG_5_ <= n455;
    BUF2_REG_6_ <= n460;
    BUF2_REG_7_ <= n465;
    BUF2_REG_8_ <= n470;
    BUF2_REG_9_ <= n475;
    BUF2_REG_10_ <= n480;
    BUF2_REG_11_ <= n485;
    BUF2_REG_12_ <= n490;
    BUF2_REG_13_ <= n495;
    BUF2_REG_14_ <= n500;
    BUF2_REG_15_ <= n505;
    BUF2_REG_16_ <= n510;
    BUF2_REG_17_ <= n515;
    BUF2_REG_18_ <= n520;
    BUF2_REG_19_ <= n525;
    BUF2_REG_20_ <= n530;
    BUF2_REG_21_ <= n535;
    BUF2_REG_22_ <= n540;
    BUF2_REG_23_ <= n545;
    BUF2_REG_24_ <= n550;
    BUF2_REG_25_ <= n555;
    BUF2_REG_26_ <= n560;
    BUF2_REG_27_ <= n565;
    BUF2_REG_28_ <= n570;
    BUF2_REG_29_ <= n575;
    BUF2_REG_30_ <= n580;
    BUF2_REG_31_ <= n585;
    READY12_REG <= n590;
    READY21_REG <= n595;
    READY22_REG <= n600;
    READY11_REG <= n605;
    P3_BE_N_REG_3_ <= n610;
    P3_BE_N_REG_2_ <= n615;
    P3_BE_N_REG_1_ <= n620;
    P3_BE_N_REG_0_ <= n625;
    P3_ADDRESS_REG_29_ <= n630;
    P3_ADDRESS_REG_28_ <= n635;
    P3_ADDRESS_REG_27_ <= n640;
    P3_ADDRESS_REG_26_ <= n645;
    P3_ADDRESS_REG_25_ <= n650;
    P3_ADDRESS_REG_24_ <= n655;
    P3_ADDRESS_REG_23_ <= n660;
    P3_ADDRESS_REG_22_ <= n665;
    P3_ADDRESS_REG_21_ <= n670;
    P3_ADDRESS_REG_20_ <= n675;
    P3_ADDRESS_REG_19_ <= n680;
    P3_ADDRESS_REG_18_ <= n685;
    P3_ADDRESS_REG_17_ <= n690;
    P3_ADDRESS_REG_16_ <= n695;
    P3_ADDRESS_REG_15_ <= n700;
    P3_ADDRESS_REG_14_ <= n705;
    P3_ADDRESS_REG_13_ <= n710;
    P3_ADDRESS_REG_12_ <= n715;
    P3_ADDRESS_REG_11_ <= n720;
    P3_ADDRESS_REG_10_ <= n725;
    P3_ADDRESS_REG_9_ <= n730;
    P3_ADDRESS_REG_8_ <= n735;
    P3_ADDRESS_REG_7_ <= n740;
    P3_ADDRESS_REG_6_ <= n745;
    P3_ADDRESS_REG_5_ <= n750;
    P3_ADDRESS_REG_4_ <= n755;
    P3_ADDRESS_REG_3_ <= n760;
    P3_ADDRESS_REG_2_ <= n765;
    P3_ADDRESS_REG_1_ <= n770;
    P3_ADDRESS_REG_0_ <= n775;
    P3_STATE_REG_2_ <= n780;
    P3_STATE_REG_1_ <= n785;
    P3_STATE_REG_0_ <= n790;
    P3_DATAWIDTH_REG_0_ <= n795;
    P3_DATAWIDTH_REG_1_ <= n800;
    P3_DATAWIDTH_REG_2_ <= n805;
    P3_DATAWIDTH_REG_3_ <= n810;
    P3_DATAWIDTH_REG_4_ <= n815;
    P3_DATAWIDTH_REG_5_ <= n820;
    P3_DATAWIDTH_REG_6_ <= n825;
    P3_DATAWIDTH_REG_7_ <= n830;
    P3_DATAWIDTH_REG_8_ <= n835;
    P3_DATAWIDTH_REG_9_ <= n840;
    P3_DATAWIDTH_REG_10_ <= n845;
    P3_DATAWIDTH_REG_11_ <= n850;
    P3_DATAWIDTH_REG_12_ <= n855;
    P3_DATAWIDTH_REG_13_ <= n860;
    P3_DATAWIDTH_REG_14_ <= n865;
    P3_DATAWIDTH_REG_15_ <= n870;
    P3_DATAWIDTH_REG_16_ <= n875;
    P3_DATAWIDTH_REG_17_ <= n880;
    P3_DATAWIDTH_REG_18_ <= n885;
    P3_DATAWIDTH_REG_19_ <= n890;
    P3_DATAWIDTH_REG_20_ <= n895;
    P3_DATAWIDTH_REG_21_ <= n900;
    P3_DATAWIDTH_REG_22_ <= n905;
    P3_DATAWIDTH_REG_23_ <= n910;
    P3_DATAWIDTH_REG_24_ <= n915;
    P3_DATAWIDTH_REG_25_ <= n920;
    P3_DATAWIDTH_REG_26_ <= n925;
    P3_DATAWIDTH_REG_27_ <= n930;
    P3_DATAWIDTH_REG_28_ <= n935;
    P3_DATAWIDTH_REG_29_ <= n940;
    P3_DATAWIDTH_REG_30_ <= n945;
    P3_DATAWIDTH_REG_31_ <= n950;
    P3_STATE2_REG_3_ <= n955;
    P3_STATE2_REG_2_ <= n960;
    P3_STATE2_REG_1_ <= n965;
    P3_STATE2_REG_0_ <= n970;
    P3_INSTQUEUE_REG_15__7_ <= n975;
    P3_INSTQUEUE_REG_15__6_ <= n980;
    P3_INSTQUEUE_REG_15__5_ <= n985;
    P3_INSTQUEUE_REG_15__4_ <= n990;
    P3_INSTQUEUE_REG_15__3_ <= n995;
    P3_INSTQUEUE_REG_15__2_ <= n1000;
    P3_INSTQUEUE_REG_15__1_ <= n1005;
    P3_INSTQUEUE_REG_15__0_ <= n1010;
    P3_INSTQUEUE_REG_14__7_ <= n1015;
    P3_INSTQUEUE_REG_14__6_ <= n1020;
    P3_INSTQUEUE_REG_14__5_ <= n1025;
    P3_INSTQUEUE_REG_14__4_ <= n1030;
    P3_INSTQUEUE_REG_14__3_ <= n1035;
    P3_INSTQUEUE_REG_14__2_ <= n1040;
    P3_INSTQUEUE_REG_14__1_ <= n1045;
    P3_INSTQUEUE_REG_14__0_ <= n1050;
    P3_INSTQUEUE_REG_13__7_ <= n1055;
    P3_INSTQUEUE_REG_13__6_ <= n1060;
    P3_INSTQUEUE_REG_13__5_ <= n1065;
    P3_INSTQUEUE_REG_13__4_ <= n1070;
    P3_INSTQUEUE_REG_13__3_ <= n1075;
    P3_INSTQUEUE_REG_13__2_ <= n1080;
    P3_INSTQUEUE_REG_13__1_ <= n1085;
    P3_INSTQUEUE_REG_13__0_ <= n1090;
    P3_INSTQUEUE_REG_12__7_ <= n1095;
    P3_INSTQUEUE_REG_12__6_ <= n1100;
    P3_INSTQUEUE_REG_12__5_ <= n1105;
    P3_INSTQUEUE_REG_12__4_ <= n1110;
    P3_INSTQUEUE_REG_12__3_ <= n1115;
    P3_INSTQUEUE_REG_12__2_ <= n1120;
    P3_INSTQUEUE_REG_12__1_ <= n1125;
    P3_INSTQUEUE_REG_12__0_ <= n1130;
    P3_INSTQUEUE_REG_11__7_ <= n1135;
    P3_INSTQUEUE_REG_11__6_ <= n1140;
    P3_INSTQUEUE_REG_11__5_ <= n1145;
    P3_INSTQUEUE_REG_11__4_ <= n1150;
    P3_INSTQUEUE_REG_11__3_ <= n1155;
    P3_INSTQUEUE_REG_11__2_ <= n1160;
    P3_INSTQUEUE_REG_11__1_ <= n1165;
    P3_INSTQUEUE_REG_11__0_ <= n1170;
    P3_INSTQUEUE_REG_10__7_ <= n1175;
    P3_INSTQUEUE_REG_10__6_ <= n1180;
    P3_INSTQUEUE_REG_10__5_ <= n1185;
    P3_INSTQUEUE_REG_10__4_ <= n1190;
    P3_INSTQUEUE_REG_10__3_ <= n1195;
    P3_INSTQUEUE_REG_10__2_ <= n1200;
    P3_INSTQUEUE_REG_10__1_ <= n1205;
    P3_INSTQUEUE_REG_10__0_ <= n1210;
    P3_INSTQUEUE_REG_9__7_ <= n1215;
    P3_INSTQUEUE_REG_9__6_ <= n1220;
    P3_INSTQUEUE_REG_9__5_ <= n1225;
    P3_INSTQUEUE_REG_9__4_ <= n1230;
    P3_INSTQUEUE_REG_9__3_ <= n1235;
    P3_INSTQUEUE_REG_9__2_ <= n1240;
    P3_INSTQUEUE_REG_9__1_ <= n1245;
    P3_INSTQUEUE_REG_9__0_ <= n1250;
    P3_INSTQUEUE_REG_8__7_ <= n1255;
    P3_INSTQUEUE_REG_8__6_ <= n1260;
    P3_INSTQUEUE_REG_8__5_ <= n1265;
    P3_INSTQUEUE_REG_8__4_ <= n1270;
    P3_INSTQUEUE_REG_8__3_ <= n1275;
    P3_INSTQUEUE_REG_8__2_ <= n1280;
    P3_INSTQUEUE_REG_8__1_ <= n1285;
    P3_INSTQUEUE_REG_8__0_ <= n1290;
    P3_INSTQUEUE_REG_7__7_ <= n1295;
    P3_INSTQUEUE_REG_7__6_ <= n1300;
    P3_INSTQUEUE_REG_7__5_ <= n1305;
    P3_INSTQUEUE_REG_7__4_ <= n1310;
    P3_INSTQUEUE_REG_7__3_ <= n1315;
    P3_INSTQUEUE_REG_7__2_ <= n1320;
    P3_INSTQUEUE_REG_7__1_ <= n1325;
    P3_INSTQUEUE_REG_7__0_ <= n1330;
    P3_INSTQUEUE_REG_6__7_ <= n1335;
    P3_INSTQUEUE_REG_6__6_ <= n1340;
    P3_INSTQUEUE_REG_6__5_ <= n1345;
    P3_INSTQUEUE_REG_6__4_ <= n1350;
    P3_INSTQUEUE_REG_6__3_ <= n1355;
    P3_INSTQUEUE_REG_6__2_ <= n1360;
    P3_INSTQUEUE_REG_6__1_ <= n1365;
    P3_INSTQUEUE_REG_6__0_ <= n1370;
    P3_INSTQUEUE_REG_5__7_ <= n1375;
    P3_INSTQUEUE_REG_5__6_ <= n1380;
    P3_INSTQUEUE_REG_5__5_ <= n1385;
    P3_INSTQUEUE_REG_5__4_ <= n1390;
    P3_INSTQUEUE_REG_5__3_ <= n1395;
    P3_INSTQUEUE_REG_5__2_ <= n1400;
    P3_INSTQUEUE_REG_5__1_ <= n1405;
    P3_INSTQUEUE_REG_5__0_ <= n1410;
    P3_INSTQUEUE_REG_4__7_ <= n1415;
    P3_INSTQUEUE_REG_4__6_ <= n1420;
    P3_INSTQUEUE_REG_4__5_ <= n1425;
    P3_INSTQUEUE_REG_4__4_ <= n1430;
    P3_INSTQUEUE_REG_4__3_ <= n1435;
    P3_INSTQUEUE_REG_4__2_ <= n1440;
    P3_INSTQUEUE_REG_4__1_ <= n1445;
    P3_INSTQUEUE_REG_4__0_ <= n1450;
    P3_INSTQUEUE_REG_3__7_ <= n1455;
    P3_INSTQUEUE_REG_3__6_ <= n1460;
    P3_INSTQUEUE_REG_3__5_ <= n1465;
    P3_INSTQUEUE_REG_3__4_ <= n1470;
    P3_INSTQUEUE_REG_3__3_ <= n1475;
    P3_INSTQUEUE_REG_3__2_ <= n1480;
    P3_INSTQUEUE_REG_3__1_ <= n1485;
    P3_INSTQUEUE_REG_3__0_ <= n1490;
    P3_INSTQUEUE_REG_2__7_ <= n1495;
    P3_INSTQUEUE_REG_2__6_ <= n1500;
    P3_INSTQUEUE_REG_2__5_ <= n1505;
    P3_INSTQUEUE_REG_2__4_ <= n1510;
    P3_INSTQUEUE_REG_2__3_ <= n1515;
    P3_INSTQUEUE_REG_2__2_ <= n1520;
    P3_INSTQUEUE_REG_2__1_ <= n1525;
    P3_INSTQUEUE_REG_2__0_ <= n1530;
    P3_INSTQUEUE_REG_1__7_ <= n1535;
    P3_INSTQUEUE_REG_1__6_ <= n1540;
    P3_INSTQUEUE_REG_1__5_ <= n1545;
    P3_INSTQUEUE_REG_1__4_ <= n1550;
    P3_INSTQUEUE_REG_1__3_ <= n1555;
    P3_INSTQUEUE_REG_1__2_ <= n1560;
    P3_INSTQUEUE_REG_1__1_ <= n1565;
    P3_INSTQUEUE_REG_1__0_ <= n1570;
    P3_INSTQUEUE_REG_0__7_ <= n1575;
    P3_INSTQUEUE_REG_0__6_ <= n1580;
    P3_INSTQUEUE_REG_0__5_ <= n1585;
    P3_INSTQUEUE_REG_0__4_ <= n1590;
    P3_INSTQUEUE_REG_0__3_ <= n1595;
    P3_INSTQUEUE_REG_0__2_ <= n1600;
    P3_INSTQUEUE_REG_0__1_ <= n1605;
    P3_INSTQUEUE_REG_0__0_ <= n1610;
    P3_INSTQUEUERD_ADDR_REG_4_ <= n1615;
    P3_INSTQUEUERD_ADDR_REG_3_ <= n1620;
    P3_INSTQUEUERD_ADDR_REG_2_ <= n1625;
    P3_INSTQUEUERD_ADDR_REG_1_ <= n1630;
    P3_INSTQUEUERD_ADDR_REG_0_ <= n1635;
    P3_INSTQUEUEWR_ADDR_REG_4_ <= n1640;
    P3_INSTQUEUEWR_ADDR_REG_3_ <= n1645;
    P3_INSTQUEUEWR_ADDR_REG_2_ <= n1650;
    P3_INSTQUEUEWR_ADDR_REG_1_ <= n1655;
    P3_INSTQUEUEWR_ADDR_REG_0_ <= n1660;
    P3_INSTADDRPOINTER_REG_0_ <= n1665;
    P3_INSTADDRPOINTER_REG_1_ <= n1670;
    P3_INSTADDRPOINTER_REG_2_ <= n1675;
    P3_INSTADDRPOINTER_REG_3_ <= n1680;
    P3_INSTADDRPOINTER_REG_4_ <= n1685;
    P3_INSTADDRPOINTER_REG_5_ <= n1690;
    P3_INSTADDRPOINTER_REG_6_ <= n1695;
    P3_INSTADDRPOINTER_REG_7_ <= n1700;
    P3_INSTADDRPOINTER_REG_8_ <= n1705;
    P3_INSTADDRPOINTER_REG_9_ <= n1710;
    P3_INSTADDRPOINTER_REG_10_ <= n1715;
    P3_INSTADDRPOINTER_REG_11_ <= n1720;
    P3_INSTADDRPOINTER_REG_12_ <= n1725;
    P3_INSTADDRPOINTER_REG_13_ <= n1730;
    P3_INSTADDRPOINTER_REG_14_ <= n1735;
    P3_INSTADDRPOINTER_REG_15_ <= n1740;
    P3_INSTADDRPOINTER_REG_16_ <= n1745;
    P3_INSTADDRPOINTER_REG_17_ <= n1750;
    P3_INSTADDRPOINTER_REG_18_ <= n1755;
    P3_INSTADDRPOINTER_REG_19_ <= n1760;
    P3_INSTADDRPOINTER_REG_20_ <= n1765;
    P3_INSTADDRPOINTER_REG_21_ <= n1770;
    P3_INSTADDRPOINTER_REG_22_ <= n1775;
    P3_INSTADDRPOINTER_REG_23_ <= n1780;
    P3_INSTADDRPOINTER_REG_24_ <= n1785;
    P3_INSTADDRPOINTER_REG_25_ <= n1790;
    P3_INSTADDRPOINTER_REG_26_ <= n1795;
    P3_INSTADDRPOINTER_REG_27_ <= n1800;
    P3_INSTADDRPOINTER_REG_28_ <= n1805;
    P3_INSTADDRPOINTER_REG_29_ <= n1810;
    P3_INSTADDRPOINTER_REG_30_ <= n1815;
    P3_INSTADDRPOINTER_REG_31_ <= n1820;
    P3_PHYADDRPOINTER_REG_0_ <= n1825;
    P3_PHYADDRPOINTER_REG_1_ <= n1830;
    P3_PHYADDRPOINTER_REG_2_ <= n1835;
    P3_PHYADDRPOINTER_REG_3_ <= n1840;
    P3_PHYADDRPOINTER_REG_4_ <= n1845;
    P3_PHYADDRPOINTER_REG_5_ <= n1850;
    P3_PHYADDRPOINTER_REG_6_ <= n1855;
    P3_PHYADDRPOINTER_REG_7_ <= n1860;
    P3_PHYADDRPOINTER_REG_8_ <= n1865;
    P3_PHYADDRPOINTER_REG_9_ <= n1870;
    P3_PHYADDRPOINTER_REG_10_ <= n1875;
    P3_PHYADDRPOINTER_REG_11_ <= n1880;
    P3_PHYADDRPOINTER_REG_12_ <= n1885;
    P3_PHYADDRPOINTER_REG_13_ <= n1890;
    P3_PHYADDRPOINTER_REG_14_ <= n1895;
    P3_PHYADDRPOINTER_REG_15_ <= n1900;
    P3_PHYADDRPOINTER_REG_16_ <= n1905;
    P3_PHYADDRPOINTER_REG_17_ <= n1910;
    P3_PHYADDRPOINTER_REG_18_ <= n1915;
    P3_PHYADDRPOINTER_REG_19_ <= n1920;
    P3_PHYADDRPOINTER_REG_20_ <= n1925;
    P3_PHYADDRPOINTER_REG_21_ <= n1930;
    P3_PHYADDRPOINTER_REG_22_ <= n1935;
    P3_PHYADDRPOINTER_REG_23_ <= n1940;
    P3_PHYADDRPOINTER_REG_24_ <= n1945;
    P3_PHYADDRPOINTER_REG_25_ <= n1950;
    P3_PHYADDRPOINTER_REG_26_ <= n1955;
    P3_PHYADDRPOINTER_REG_27_ <= n1960;
    P3_PHYADDRPOINTER_REG_28_ <= n1965;
    P3_PHYADDRPOINTER_REG_29_ <= n1970;
    P3_PHYADDRPOINTER_REG_30_ <= n1975;
    P3_PHYADDRPOINTER_REG_31_ <= n1980;
    P3_LWORD_REG_15_ <= n1985;
    P3_LWORD_REG_14_ <= n1990;
    P3_LWORD_REG_13_ <= n1995;
    P3_LWORD_REG_12_ <= n2000;
    P3_LWORD_REG_11_ <= n2005;
    P3_LWORD_REG_10_ <= n2010;
    P3_LWORD_REG_9_ <= n2015;
    P3_LWORD_REG_8_ <= n2020;
    P3_LWORD_REG_7_ <= n2025;
    P3_LWORD_REG_6_ <= n2030;
    P3_LWORD_REG_5_ <= n2035;
    P3_LWORD_REG_4_ <= n2040;
    P3_LWORD_REG_3_ <= n2045;
    P3_LWORD_REG_2_ <= n2050;
    P3_LWORD_REG_1_ <= n2055;
    P3_LWORD_REG_0_ <= n2060;
    P3_UWORD_REG_14_ <= n2065;
    P3_UWORD_REG_13_ <= n2070;
    P3_UWORD_REG_12_ <= n2075;
    P3_UWORD_REG_11_ <= n2080;
    P3_UWORD_REG_10_ <= n2085;
    P3_UWORD_REG_9_ <= n2090;
    P3_UWORD_REG_8_ <= n2095;
    P3_UWORD_REG_7_ <= n2100;
    P3_UWORD_REG_6_ <= n2105;
    P3_UWORD_REG_5_ <= n2110;
    P3_UWORD_REG_4_ <= n2115;
    P3_UWORD_REG_3_ <= n2120;
    P3_UWORD_REG_2_ <= n2125;
    P3_UWORD_REG_1_ <= n2130;
    P3_UWORD_REG_0_ <= n2135;
    P3_DATAO_REG_0_ <= n2140;
    P3_DATAO_REG_1_ <= n2144;
    P3_DATAO_REG_2_ <= n2148;
    P3_DATAO_REG_3_ <= n2152;
    P3_DATAO_REG_4_ <= n2156;
    P3_DATAO_REG_5_ <= n2160;
    P3_DATAO_REG_6_ <= n2164;
    P3_DATAO_REG_7_ <= n2168;
    P3_DATAO_REG_8_ <= n2172;
    P3_DATAO_REG_9_ <= n2176;
    P3_DATAO_REG_10_ <= n2180;
    P3_DATAO_REG_11_ <= n2184;
    P3_DATAO_REG_12_ <= n2188;
    P3_DATAO_REG_13_ <= n2192;
    P3_DATAO_REG_14_ <= n2196;
    P3_DATAO_REG_15_ <= n2200;
    P3_DATAO_REG_16_ <= n2204;
    P3_DATAO_REG_17_ <= n2208;
    P3_DATAO_REG_18_ <= n2212;
    P3_DATAO_REG_19_ <= n2216;
    P3_DATAO_REG_20_ <= n2220;
    P3_DATAO_REG_21_ <= n2224;
    P3_DATAO_REG_22_ <= n2228;
    P3_DATAO_REG_23_ <= n2232;
    P3_DATAO_REG_24_ <= n2236;
    P3_DATAO_REG_25_ <= n2240;
    P3_DATAO_REG_26_ <= n2244;
    P3_DATAO_REG_27_ <= n2248;
    P3_DATAO_REG_28_ <= n2252;
    P3_DATAO_REG_29_ <= n2256;
    P3_DATAO_REG_30_ <= n2260;
    P3_DATAO_REG_31_ <= n2264;
    P3_EAX_REG_0_ <= n2268;
    P3_EAX_REG_1_ <= n2273;
    P3_EAX_REG_2_ <= n2278;
    P3_EAX_REG_3_ <= n2283;
    P3_EAX_REG_4_ <= n2288;
    P3_EAX_REG_5_ <= n2293;
    P3_EAX_REG_6_ <= n2298;
    P3_EAX_REG_7_ <= n2303;
    P3_EAX_REG_8_ <= n2308;
    P3_EAX_REG_9_ <= n2313;
    P3_EAX_REG_10_ <= n2318;
    P3_EAX_REG_11_ <= n2323;
    P3_EAX_REG_12_ <= n2328;
    P3_EAX_REG_13_ <= n2333;
    P3_EAX_REG_14_ <= n2338;
    P3_EAX_REG_15_ <= n2343;
    P3_EAX_REG_16_ <= n2348;
    P3_EAX_REG_17_ <= n2353;
    P3_EAX_REG_18_ <= n2358;
    P3_EAX_REG_19_ <= n2363;
    P3_EAX_REG_20_ <= n2368;
    P3_EAX_REG_21_ <= n2373;
    P3_EAX_REG_22_ <= n2378;
    P3_EAX_REG_23_ <= n2383;
    P3_EAX_REG_24_ <= n2388;
    P3_EAX_REG_25_ <= n2393;
    P3_EAX_REG_26_ <= n2398;
    P3_EAX_REG_27_ <= n2403;
    P3_EAX_REG_28_ <= n2408;
    P3_EAX_REG_29_ <= n2413;
    P3_EAX_REG_30_ <= n2418;
    P3_EAX_REG_31_ <= n2423;
    P3_EBX_REG_0_ <= n2428;
    P3_EBX_REG_1_ <= n2433;
    P3_EBX_REG_2_ <= n2438;
    P3_EBX_REG_3_ <= n2443;
    P3_EBX_REG_4_ <= n2448;
    P3_EBX_REG_5_ <= n2453;
    P3_EBX_REG_6_ <= n2458;
    P3_EBX_REG_7_ <= n2463;
    P3_EBX_REG_8_ <= n2468;
    P3_EBX_REG_9_ <= n2473;
    P3_EBX_REG_10_ <= n2478;
    P3_EBX_REG_11_ <= n2483;
    P3_EBX_REG_12_ <= n2488;
    P3_EBX_REG_13_ <= n2493;
    P3_EBX_REG_14_ <= n2498;
    P3_EBX_REG_15_ <= n2503;
    P3_EBX_REG_16_ <= n2508;
    P3_EBX_REG_17_ <= n2513;
    P3_EBX_REG_18_ <= n2518;
    P3_EBX_REG_19_ <= n2523;
    P3_EBX_REG_20_ <= n2528;
    P3_EBX_REG_21_ <= n2533;
    P3_EBX_REG_22_ <= n2538;
    P3_EBX_REG_23_ <= n2543;
    P3_EBX_REG_24_ <= n2548;
    P3_EBX_REG_25_ <= n2553;
    P3_EBX_REG_26_ <= n2558;
    P3_EBX_REG_27_ <= n2563;
    P3_EBX_REG_28_ <= n2568;
    P3_EBX_REG_29_ <= n2573;
    P3_EBX_REG_30_ <= n2578;
    P3_EBX_REG_31_ <= n2583;
    P3_REIP_REG_0_ <= n2588;
    P3_REIP_REG_1_ <= n2593;
    P3_REIP_REG_2_ <= n2598;
    P3_REIP_REG_3_ <= n2603;
    P3_REIP_REG_4_ <= n2608;
    P3_REIP_REG_5_ <= n2613;
    P3_REIP_REG_6_ <= n2618;
    P3_REIP_REG_7_ <= n2623;
    P3_REIP_REG_8_ <= n2628;
    P3_REIP_REG_9_ <= n2633;
    P3_REIP_REG_10_ <= n2638;
    P3_REIP_REG_11_ <= n2643;
    P3_REIP_REG_12_ <= n2648;
    P3_REIP_REG_13_ <= n2653;
    P3_REIP_REG_14_ <= n2658;
    P3_REIP_REG_15_ <= n2663;
    P3_REIP_REG_16_ <= n2668;
    P3_REIP_REG_17_ <= n2673;
    P3_REIP_REG_18_ <= n2678;
    P3_REIP_REG_19_ <= n2683;
    P3_REIP_REG_20_ <= n2688;
    P3_REIP_REG_21_ <= n2693;
    P3_REIP_REG_22_ <= n2698;
    P3_REIP_REG_23_ <= n2703;
    P3_REIP_REG_24_ <= n2708;
    P3_REIP_REG_25_ <= n2713;
    P3_REIP_REG_26_ <= n2718;
    P3_REIP_REG_27_ <= n2723;
    P3_REIP_REG_28_ <= n2728;
    P3_REIP_REG_29_ <= n2733;
    P3_REIP_REG_30_ <= n2738;
    P3_REIP_REG_31_ <= n2743;
    P3_BYTEENABLE_REG_3_ <= n2748;
    P3_BYTEENABLE_REG_2_ <= n2753;
    P3_BYTEENABLE_REG_1_ <= n2758;
    P3_BYTEENABLE_REG_0_ <= n2763;
    P3_W_R_N_REG <= n2768;
    P3_FLUSH_REG <= n2772;
    P3_MORE_REG <= n2777;
    P3_STATEBS16_REG <= n2782;
    P3_REQUESTPENDING_REG <= n2787;
    P3_D_C_N_REG <= n2792;
    P3_M_IO_N_REG <= n2796;
    P3_CODEFETCH_REG <= n2800;
    P3_ADS_N_REG <= n2805;
    P3_READREQUEST_REG <= n2809;
    P3_MEMORYFETCH_REG <= n2814;
    P2_BE_N_REG_3_ <= n2819;
    P2_BE_N_REG_2_ <= n2824;
    P2_BE_N_REG_1_ <= n2829;
    P2_BE_N_REG_0_ <= n2834;
    P2_ADDRESS_REG_29_ <= n2839;
    P2_ADDRESS_REG_28_ <= n2844;
    P2_ADDRESS_REG_27_ <= n2849;
    P2_ADDRESS_REG_26_ <= n2854;
    P2_ADDRESS_REG_25_ <= n2859;
    P2_ADDRESS_REG_24_ <= n2864;
    P2_ADDRESS_REG_23_ <= n2869;
    P2_ADDRESS_REG_22_ <= n2874;
    P2_ADDRESS_REG_21_ <= n2879;
    P2_ADDRESS_REG_20_ <= n2884;
    P2_ADDRESS_REG_19_ <= n2889;
    P2_ADDRESS_REG_18_ <= n2894;
    P2_ADDRESS_REG_17_ <= n2899;
    P2_ADDRESS_REG_16_ <= n2904;
    P2_ADDRESS_REG_15_ <= n2909;
    P2_ADDRESS_REG_14_ <= n2914;
    P2_ADDRESS_REG_13_ <= n2919;
    P2_ADDRESS_REG_12_ <= n2924;
    P2_ADDRESS_REG_11_ <= n2929;
    P2_ADDRESS_REG_10_ <= n2934;
    P2_ADDRESS_REG_9_ <= n2939;
    P2_ADDRESS_REG_8_ <= n2944;
    P2_ADDRESS_REG_7_ <= n2949;
    P2_ADDRESS_REG_6_ <= n2954;
    P2_ADDRESS_REG_5_ <= n2959;
    P2_ADDRESS_REG_4_ <= n2964;
    P2_ADDRESS_REG_3_ <= n2969;
    P2_ADDRESS_REG_2_ <= n2974;
    P2_ADDRESS_REG_1_ <= n2979;
    P2_ADDRESS_REG_0_ <= n2984;
    P2_STATE_REG_2_ <= n2989;
    P2_STATE_REG_1_ <= n2994;
    P2_STATE_REG_0_ <= n2999;
    P2_DATAWIDTH_REG_0_ <= n3004;
    P2_DATAWIDTH_REG_1_ <= n3009;
    P2_DATAWIDTH_REG_2_ <= n3014;
    P2_DATAWIDTH_REG_3_ <= n3019;
    P2_DATAWIDTH_REG_4_ <= n3024;
    P2_DATAWIDTH_REG_5_ <= n3029;
    P2_DATAWIDTH_REG_6_ <= n3034;
    P2_DATAWIDTH_REG_7_ <= n3039;
    P2_DATAWIDTH_REG_8_ <= n3044;
    P2_DATAWIDTH_REG_9_ <= n3049;
    P2_DATAWIDTH_REG_10_ <= n3054;
    P2_DATAWIDTH_REG_11_ <= n3059;
    P2_DATAWIDTH_REG_12_ <= n3064;
    P2_DATAWIDTH_REG_13_ <= n3069;
    P2_DATAWIDTH_REG_14_ <= n3074;
    P2_DATAWIDTH_REG_15_ <= n3079;
    P2_DATAWIDTH_REG_16_ <= n3084;
    P2_DATAWIDTH_REG_17_ <= n3089;
    P2_DATAWIDTH_REG_18_ <= n3094;
    P2_DATAWIDTH_REG_19_ <= n3099;
    P2_DATAWIDTH_REG_20_ <= n3104;
    P2_DATAWIDTH_REG_21_ <= n3109;
    P2_DATAWIDTH_REG_22_ <= n3114;
    P2_DATAWIDTH_REG_23_ <= n3119;
    P2_DATAWIDTH_REG_24_ <= n3124;
    P2_DATAWIDTH_REG_25_ <= n3129;
    P2_DATAWIDTH_REG_26_ <= n3134;
    P2_DATAWIDTH_REG_27_ <= n3139;
    P2_DATAWIDTH_REG_28_ <= n3144;
    P2_DATAWIDTH_REG_29_ <= n3149;
    P2_DATAWIDTH_REG_30_ <= n3154;
    P2_DATAWIDTH_REG_31_ <= n3159;
    P2_STATE2_REG_3_ <= n3164;
    P2_STATE2_REG_2_ <= n3169;
    P2_STATE2_REG_1_ <= n3174;
    P2_STATE2_REG_0_ <= n3179;
    P2_INSTQUEUE_REG_15__7_ <= n3184;
    P2_INSTQUEUE_REG_15__6_ <= n3189;
    P2_INSTQUEUE_REG_15__5_ <= n3194;
    P2_INSTQUEUE_REG_15__4_ <= n3199;
    P2_INSTQUEUE_REG_15__3_ <= n3204;
    P2_INSTQUEUE_REG_15__2_ <= n3209;
    P2_INSTQUEUE_REG_15__1_ <= n3214;
    P2_INSTQUEUE_REG_15__0_ <= n3219;
    P2_INSTQUEUE_REG_14__7_ <= n3224;
    P2_INSTQUEUE_REG_14__6_ <= n3229;
    P2_INSTQUEUE_REG_14__5_ <= n3234;
    P2_INSTQUEUE_REG_14__4_ <= n3239;
    P2_INSTQUEUE_REG_14__3_ <= n3244;
    P2_INSTQUEUE_REG_14__2_ <= n3249;
    P2_INSTQUEUE_REG_14__1_ <= n3254;
    P2_INSTQUEUE_REG_14__0_ <= n3259;
    P2_INSTQUEUE_REG_13__7_ <= n3264;
    P2_INSTQUEUE_REG_13__6_ <= n3269;
    P2_INSTQUEUE_REG_13__5_ <= n3274;
    P2_INSTQUEUE_REG_13__4_ <= n3279;
    P2_INSTQUEUE_REG_13__3_ <= n3284;
    P2_INSTQUEUE_REG_13__2_ <= n3289;
    P2_INSTQUEUE_REG_13__1_ <= n3294;
    P2_INSTQUEUE_REG_13__0_ <= n3299;
    P2_INSTQUEUE_REG_12__7_ <= n3304;
    P2_INSTQUEUE_REG_12__6_ <= n3309;
    P2_INSTQUEUE_REG_12__5_ <= n3314;
    P2_INSTQUEUE_REG_12__4_ <= n3319;
    P2_INSTQUEUE_REG_12__3_ <= n3324;
    P2_INSTQUEUE_REG_12__2_ <= n3329;
    P2_INSTQUEUE_REG_12__1_ <= n3334;
    P2_INSTQUEUE_REG_12__0_ <= n3339;
    P2_INSTQUEUE_REG_11__7_ <= n3344;
    P2_INSTQUEUE_REG_11__6_ <= n3349;
    P2_INSTQUEUE_REG_11__5_ <= n3354;
    P2_INSTQUEUE_REG_11__4_ <= n3359;
    P2_INSTQUEUE_REG_11__3_ <= n3364;
    P2_INSTQUEUE_REG_11__2_ <= n3369;
    P2_INSTQUEUE_REG_11__1_ <= n3374;
    P2_INSTQUEUE_REG_11__0_ <= n3379;
    P2_INSTQUEUE_REG_10__7_ <= n3384;
    P2_INSTQUEUE_REG_10__6_ <= n3389;
    P2_INSTQUEUE_REG_10__5_ <= n3394;
    P2_INSTQUEUE_REG_10__4_ <= n3399;
    P2_INSTQUEUE_REG_10__3_ <= n3404;
    P2_INSTQUEUE_REG_10__2_ <= n3409;
    P2_INSTQUEUE_REG_10__1_ <= n3414;
    P2_INSTQUEUE_REG_10__0_ <= n3419;
    P2_INSTQUEUE_REG_9__7_ <= n3424;
    P2_INSTQUEUE_REG_9__6_ <= n3429;
    P2_INSTQUEUE_REG_9__5_ <= n3434;
    P2_INSTQUEUE_REG_9__4_ <= n3439;
    P2_INSTQUEUE_REG_9__3_ <= n3444;
    P2_INSTQUEUE_REG_9__2_ <= n3449;
    P2_INSTQUEUE_REG_9__1_ <= n3454;
    P2_INSTQUEUE_REG_9__0_ <= n3459;
    P2_INSTQUEUE_REG_8__7_ <= n3464;
    P2_INSTQUEUE_REG_8__6_ <= n3469;
    P2_INSTQUEUE_REG_8__5_ <= n3474;
    P2_INSTQUEUE_REG_8__4_ <= n3479;
    P2_INSTQUEUE_REG_8__3_ <= n3484;
    P2_INSTQUEUE_REG_8__2_ <= n3489;
    P2_INSTQUEUE_REG_8__1_ <= n3494;
    P2_INSTQUEUE_REG_8__0_ <= n3499;
    P2_INSTQUEUE_REG_7__7_ <= n3504;
    P2_INSTQUEUE_REG_7__6_ <= n3509;
    P2_INSTQUEUE_REG_7__5_ <= n3514;
    P2_INSTQUEUE_REG_7__4_ <= n3519;
    P2_INSTQUEUE_REG_7__3_ <= n3524;
    P2_INSTQUEUE_REG_7__2_ <= n3529;
    P2_INSTQUEUE_REG_7__1_ <= n3534;
    P2_INSTQUEUE_REG_7__0_ <= n3539;
    P2_INSTQUEUE_REG_6__7_ <= n3544;
    P2_INSTQUEUE_REG_6__6_ <= n3549;
    P2_INSTQUEUE_REG_6__5_ <= n3554;
    P2_INSTQUEUE_REG_6__4_ <= n3559;
    P2_INSTQUEUE_REG_6__3_ <= n3564;
    P2_INSTQUEUE_REG_6__2_ <= n3569;
    P2_INSTQUEUE_REG_6__1_ <= n3574;
    P2_INSTQUEUE_REG_6__0_ <= n3579;
    P2_INSTQUEUE_REG_5__7_ <= n3584;
    P2_INSTQUEUE_REG_5__6_ <= n3589;
    P2_INSTQUEUE_REG_5__5_ <= n3594;
    P2_INSTQUEUE_REG_5__4_ <= n3599;
    P2_INSTQUEUE_REG_5__3_ <= n3604;
    P2_INSTQUEUE_REG_5__2_ <= n3609;
    P2_INSTQUEUE_REG_5__1_ <= n3614;
    P2_INSTQUEUE_REG_5__0_ <= n3619;
    P2_INSTQUEUE_REG_4__7_ <= n3624;
    P2_INSTQUEUE_REG_4__6_ <= n3629;
    P2_INSTQUEUE_REG_4__5_ <= n3634;
    P2_INSTQUEUE_REG_4__4_ <= n3639;
    P2_INSTQUEUE_REG_4__3_ <= n3644;
    P2_INSTQUEUE_REG_4__2_ <= n3649;
    P2_INSTQUEUE_REG_4__1_ <= n3654;
    P2_INSTQUEUE_REG_4__0_ <= n3659;
    P2_INSTQUEUE_REG_3__7_ <= n3664;
    P2_INSTQUEUE_REG_3__6_ <= n3669;
    P2_INSTQUEUE_REG_3__5_ <= n3674;
    P2_INSTQUEUE_REG_3__4_ <= n3679;
    P2_INSTQUEUE_REG_3__3_ <= n3684;
    P2_INSTQUEUE_REG_3__2_ <= n3689;
    P2_INSTQUEUE_REG_3__1_ <= n3694;
    P2_INSTQUEUE_REG_3__0_ <= n3699;
    P2_INSTQUEUE_REG_2__7_ <= n3704;
    P2_INSTQUEUE_REG_2__6_ <= n3709;
    P2_INSTQUEUE_REG_2__5_ <= n3714;
    P2_INSTQUEUE_REG_2__4_ <= n3719;
    P2_INSTQUEUE_REG_2__3_ <= n3724;
    P2_INSTQUEUE_REG_2__2_ <= n3729;
    P2_INSTQUEUE_REG_2__1_ <= n3734;
    P2_INSTQUEUE_REG_2__0_ <= n3739;
    P2_INSTQUEUE_REG_1__7_ <= n3744;
    P2_INSTQUEUE_REG_1__6_ <= n3749;
    P2_INSTQUEUE_REG_1__5_ <= n3754;
    P2_INSTQUEUE_REG_1__4_ <= n3759;
    P2_INSTQUEUE_REG_1__3_ <= n3764;
    P2_INSTQUEUE_REG_1__2_ <= n3769;
    P2_INSTQUEUE_REG_1__1_ <= n3774;
    P2_INSTQUEUE_REG_1__0_ <= n3779;
    P2_INSTQUEUE_REG_0__7_ <= n3784;
    P2_INSTQUEUE_REG_0__6_ <= n3789;
    P2_INSTQUEUE_REG_0__5_ <= n3794;
    P2_INSTQUEUE_REG_0__4_ <= n3799;
    P2_INSTQUEUE_REG_0__3_ <= n3804;
    P2_INSTQUEUE_REG_0__2_ <= n3809;
    P2_INSTQUEUE_REG_0__1_ <= n3814;
    P2_INSTQUEUE_REG_0__0_ <= n3819;
    P2_INSTQUEUERD_ADDR_REG_4_ <= n3824;
    P2_INSTQUEUERD_ADDR_REG_3_ <= n3829;
    P2_INSTQUEUERD_ADDR_REG_2_ <= n3834;
    P2_INSTQUEUERD_ADDR_REG_1_ <= n3839;
    P2_INSTQUEUERD_ADDR_REG_0_ <= n3844;
    P2_INSTQUEUEWR_ADDR_REG_4_ <= n3849;
    P2_INSTQUEUEWR_ADDR_REG_3_ <= n3854;
    P2_INSTQUEUEWR_ADDR_REG_2_ <= n3859;
    P2_INSTQUEUEWR_ADDR_REG_1_ <= n3864;
    P2_INSTQUEUEWR_ADDR_REG_0_ <= n3869;
    P2_INSTADDRPOINTER_REG_0_ <= n3874;
    P2_INSTADDRPOINTER_REG_1_ <= n3879;
    P2_INSTADDRPOINTER_REG_2_ <= n3884;
    P2_INSTADDRPOINTER_REG_3_ <= n3889;
    P2_INSTADDRPOINTER_REG_4_ <= n3894;
    P2_INSTADDRPOINTER_REG_5_ <= n3899;
    P2_INSTADDRPOINTER_REG_6_ <= n3904;
    P2_INSTADDRPOINTER_REG_7_ <= n3909;
    P2_INSTADDRPOINTER_REG_8_ <= n3914;
    P2_INSTADDRPOINTER_REG_9_ <= n3919;
    P2_INSTADDRPOINTER_REG_10_ <= n3924;
    P2_INSTADDRPOINTER_REG_11_ <= n3929;
    P2_INSTADDRPOINTER_REG_12_ <= n3934;
    P2_INSTADDRPOINTER_REG_13_ <= n3939;
    P2_INSTADDRPOINTER_REG_14_ <= n3944;
    P2_INSTADDRPOINTER_REG_15_ <= n3949;
    P2_INSTADDRPOINTER_REG_16_ <= n3954;
    P2_INSTADDRPOINTER_REG_17_ <= n3959;
    P2_INSTADDRPOINTER_REG_18_ <= n3964;
    P2_INSTADDRPOINTER_REG_19_ <= n3969;
    P2_INSTADDRPOINTER_REG_20_ <= n3974;
    P2_INSTADDRPOINTER_REG_21_ <= n3979;
    P2_INSTADDRPOINTER_REG_22_ <= n3984;
    P2_INSTADDRPOINTER_REG_23_ <= n3989;
    P2_INSTADDRPOINTER_REG_24_ <= n3994;
    P2_INSTADDRPOINTER_REG_25_ <= n3999;
    P2_INSTADDRPOINTER_REG_26_ <= n4004;
    P2_INSTADDRPOINTER_REG_27_ <= n4009;
    P2_INSTADDRPOINTER_REG_28_ <= n4014;
    P2_INSTADDRPOINTER_REG_29_ <= n4019;
    P2_INSTADDRPOINTER_REG_30_ <= n4024;
    P2_INSTADDRPOINTER_REG_31_ <= n4029;
    P2_PHYADDRPOINTER_REG_0_ <= n4034;
    P2_PHYADDRPOINTER_REG_1_ <= n4039;
    P2_PHYADDRPOINTER_REG_2_ <= n4044;
    P2_PHYADDRPOINTER_REG_3_ <= n4049;
    P2_PHYADDRPOINTER_REG_4_ <= n4054;
    P2_PHYADDRPOINTER_REG_5_ <= n4059;
    P2_PHYADDRPOINTER_REG_6_ <= n4064;
    P2_PHYADDRPOINTER_REG_7_ <= n4069;
    P2_PHYADDRPOINTER_REG_8_ <= n4074;
    P2_PHYADDRPOINTER_REG_9_ <= n4079;
    P2_PHYADDRPOINTER_REG_10_ <= n4084;
    P2_PHYADDRPOINTER_REG_11_ <= n4089;
    P2_PHYADDRPOINTER_REG_12_ <= n4094;
    P2_PHYADDRPOINTER_REG_13_ <= n4099;
    P2_PHYADDRPOINTER_REG_14_ <= n4104;
    P2_PHYADDRPOINTER_REG_15_ <= n4109;
    P2_PHYADDRPOINTER_REG_16_ <= n4114;
    P2_PHYADDRPOINTER_REG_17_ <= n4119;
    P2_PHYADDRPOINTER_REG_18_ <= n4124;
    P2_PHYADDRPOINTER_REG_19_ <= n4129;
    P2_PHYADDRPOINTER_REG_20_ <= n4134;
    P2_PHYADDRPOINTER_REG_21_ <= n4139;
    P2_PHYADDRPOINTER_REG_22_ <= n4144;
    P2_PHYADDRPOINTER_REG_23_ <= n4149;
    P2_PHYADDRPOINTER_REG_24_ <= n4154;
    P2_PHYADDRPOINTER_REG_25_ <= n4159;
    P2_PHYADDRPOINTER_REG_26_ <= n4164;
    P2_PHYADDRPOINTER_REG_27_ <= n4169;
    P2_PHYADDRPOINTER_REG_28_ <= n4174;
    P2_PHYADDRPOINTER_REG_29_ <= n4179;
    P2_PHYADDRPOINTER_REG_30_ <= n4184;
    P2_PHYADDRPOINTER_REG_31_ <= n4189;
    P2_LWORD_REG_15_ <= n4194;
    P2_LWORD_REG_14_ <= n4199;
    P2_LWORD_REG_13_ <= n4204;
    P2_LWORD_REG_12_ <= n4209;
    P2_LWORD_REG_11_ <= n4214;
    P2_LWORD_REG_10_ <= n4219;
    P2_LWORD_REG_9_ <= n4224;
    P2_LWORD_REG_8_ <= n4229;
    P2_LWORD_REG_7_ <= n4234;
    P2_LWORD_REG_6_ <= n4239;
    P2_LWORD_REG_5_ <= n4244;
    P2_LWORD_REG_4_ <= n4249;
    P2_LWORD_REG_3_ <= n4254;
    P2_LWORD_REG_2_ <= n4259;
    P2_LWORD_REG_1_ <= n4264;
    P2_LWORD_REG_0_ <= n4269;
    P2_UWORD_REG_14_ <= n4274;
    P2_UWORD_REG_13_ <= n4279;
    P2_UWORD_REG_12_ <= n4284;
    P2_UWORD_REG_11_ <= n4289;
    P2_UWORD_REG_10_ <= n4294;
    P2_UWORD_REG_9_ <= n4299;
    P2_UWORD_REG_8_ <= n4304;
    P2_UWORD_REG_7_ <= n4309;
    P2_UWORD_REG_6_ <= n4314;
    P2_UWORD_REG_5_ <= n4319;
    P2_UWORD_REG_4_ <= n4324;
    P2_UWORD_REG_3_ <= n4329;
    P2_UWORD_REG_2_ <= n4334;
    P2_UWORD_REG_1_ <= n4339;
    P2_UWORD_REG_0_ <= n4344;
    P2_DATAO_REG_0_ <= n4349;
    P2_DATAO_REG_1_ <= n4354;
    P2_DATAO_REG_2_ <= n4359;
    P2_DATAO_REG_3_ <= n4364;
    P2_DATAO_REG_4_ <= n4369;
    P2_DATAO_REG_5_ <= n4374;
    P2_DATAO_REG_6_ <= n4379;
    P2_DATAO_REG_7_ <= n4384;
    P2_DATAO_REG_8_ <= n4389;
    P2_DATAO_REG_9_ <= n4394;
    P2_DATAO_REG_10_ <= n4399;
    P2_DATAO_REG_11_ <= n4404;
    P2_DATAO_REG_12_ <= n4409;
    P2_DATAO_REG_13_ <= n4414;
    P2_DATAO_REG_14_ <= n4419;
    P2_DATAO_REG_15_ <= n4424;
    P2_DATAO_REG_16_ <= n4429;
    P2_DATAO_REG_17_ <= n4434;
    P2_DATAO_REG_18_ <= n4439;
    P2_DATAO_REG_19_ <= n4444;
    P2_DATAO_REG_20_ <= n4449;
    P2_DATAO_REG_21_ <= n4454;
    P2_DATAO_REG_22_ <= n4459;
    P2_DATAO_REG_23_ <= n4464;
    P2_DATAO_REG_24_ <= n4469;
    P2_DATAO_REG_25_ <= n4474;
    P2_DATAO_REG_26_ <= n4479;
    P2_DATAO_REG_27_ <= n4484;
    P2_DATAO_REG_28_ <= n4489;
    P2_DATAO_REG_29_ <= n4494;
    P2_DATAO_REG_30_ <= n4499;
    P2_DATAO_REG_31_ <= n4504;
    P2_EAX_REG_0_ <= n4509;
    P2_EAX_REG_1_ <= n4514;
    P2_EAX_REG_2_ <= n4519;
    P2_EAX_REG_3_ <= n4524;
    P2_EAX_REG_4_ <= n4529;
    P2_EAX_REG_5_ <= n4534;
    P2_EAX_REG_6_ <= n4539;
    P2_EAX_REG_7_ <= n4544;
    P2_EAX_REG_8_ <= n4549;
    P2_EAX_REG_9_ <= n4554;
    P2_EAX_REG_10_ <= n4559;
    P2_EAX_REG_11_ <= n4564;
    P2_EAX_REG_12_ <= n4569;
    P2_EAX_REG_13_ <= n4574;
    P2_EAX_REG_14_ <= n4579;
    P2_EAX_REG_15_ <= n4584;
    P2_EAX_REG_16_ <= n4589;
    P2_EAX_REG_17_ <= n4594;
    P2_EAX_REG_18_ <= n4599;
    P2_EAX_REG_19_ <= n4604;
    P2_EAX_REG_20_ <= n4609;
    P2_EAX_REG_21_ <= n4614;
    P2_EAX_REG_22_ <= n4619;
    P2_EAX_REG_23_ <= n4624;
    P2_EAX_REG_24_ <= n4629;
    P2_EAX_REG_25_ <= n4634;
    P2_EAX_REG_26_ <= n4639;
    P2_EAX_REG_27_ <= n4644;
    P2_EAX_REG_28_ <= n4649;
    P2_EAX_REG_29_ <= n4654;
    P2_EAX_REG_30_ <= n4659;
    P2_EAX_REG_31_ <= n4664;
    P2_EBX_REG_0_ <= n4669;
    P2_EBX_REG_1_ <= n4674;
    P2_EBX_REG_2_ <= n4679;
    P2_EBX_REG_3_ <= n4684;
    P2_EBX_REG_4_ <= n4689;
    P2_EBX_REG_5_ <= n4694;
    P2_EBX_REG_6_ <= n4699;
    P2_EBX_REG_7_ <= n4704;
    P2_EBX_REG_8_ <= n4709;
    P2_EBX_REG_9_ <= n4714;
    P2_EBX_REG_10_ <= n4719;
    P2_EBX_REG_11_ <= n4724;
    P2_EBX_REG_12_ <= n4729;
    P2_EBX_REG_13_ <= n4734;
    P2_EBX_REG_14_ <= n4739;
    P2_EBX_REG_15_ <= n4744;
    P2_EBX_REG_16_ <= n4749;
    P2_EBX_REG_17_ <= n4754;
    P2_EBX_REG_18_ <= n4759;
    P2_EBX_REG_19_ <= n4764;
    P2_EBX_REG_20_ <= n4769;
    P2_EBX_REG_21_ <= n4774;
    P2_EBX_REG_22_ <= n4779;
    P2_EBX_REG_23_ <= n4784;
    P2_EBX_REG_24_ <= n4789;
    P2_EBX_REG_25_ <= n4794;
    P2_EBX_REG_26_ <= n4799;
    P2_EBX_REG_27_ <= n4804;
    P2_EBX_REG_28_ <= n4809;
    P2_EBX_REG_29_ <= n4814;
    P2_EBX_REG_30_ <= n4819;
    P2_EBX_REG_31_ <= n4824;
    P2_REIP_REG_0_ <= n4829;
    P2_REIP_REG_1_ <= n4834;
    P2_REIP_REG_2_ <= n4839;
    P2_REIP_REG_3_ <= n4844;
    P2_REIP_REG_4_ <= n4849;
    P2_REIP_REG_5_ <= n4854;
    P2_REIP_REG_6_ <= n4859;
    P2_REIP_REG_7_ <= n4864;
    P2_REIP_REG_8_ <= n4869;
    P2_REIP_REG_9_ <= n4874;
    P2_REIP_REG_10_ <= n4879;
    P2_REIP_REG_11_ <= n4884;
    P2_REIP_REG_12_ <= n4889;
    P2_REIP_REG_13_ <= n4894;
    P2_REIP_REG_14_ <= n4899;
    P2_REIP_REG_15_ <= n4904;
    P2_REIP_REG_16_ <= n4909;
    P2_REIP_REG_17_ <= n4914;
    P2_REIP_REG_18_ <= n4919;
    P2_REIP_REG_19_ <= n4924;
    P2_REIP_REG_20_ <= n4929;
    P2_REIP_REG_21_ <= n4934;
    P2_REIP_REG_22_ <= n4939;
    P2_REIP_REG_23_ <= n4944;
    P2_REIP_REG_24_ <= n4949;
    P2_REIP_REG_25_ <= n4954;
    P2_REIP_REG_26_ <= n4959;
    P2_REIP_REG_27_ <= n4964;
    P2_REIP_REG_28_ <= n4969;
    P2_REIP_REG_29_ <= n4974;
    P2_REIP_REG_30_ <= n4979;
    P2_REIP_REG_31_ <= n4984;
    P2_BYTEENABLE_REG_3_ <= n4989;
    P2_BYTEENABLE_REG_2_ <= n4994;
    P2_BYTEENABLE_REG_1_ <= n4999;
    P2_BYTEENABLE_REG_0_ <= n5004;
    P2_W_R_N_REG <= n5009;
    P2_FLUSH_REG <= n5014;
    P2_MORE_REG <= n5019;
    P2_STATEBS16_REG <= n5024;
    P2_REQUESTPENDING_REG <= n5029;
    P2_D_C_N_REG <= n5034;
    P2_M_IO_N_REG <= n5039;
    P2_CODEFETCH_REG <= n5044;
    P2_ADS_N_REG <= n5049;
    P2_READREQUEST_REG <= n5054;
    P2_MEMORYFETCH_REG <= n5059;
    P1_BE_N_REG_3_ <= n5064;
    P1_BE_N_REG_2_ <= n5069;
    P1_BE_N_REG_1_ <= n5074;
    P1_BE_N_REG_0_ <= n5079;
    P1_ADDRESS_REG_29_ <= n5084;
    P1_ADDRESS_REG_28_ <= n5088;
    P1_ADDRESS_REG_27_ <= n5092;
    P1_ADDRESS_REG_26_ <= n5096;
    P1_ADDRESS_REG_25_ <= n5100;
    P1_ADDRESS_REG_24_ <= n5104;
    P1_ADDRESS_REG_23_ <= n5108;
    P1_ADDRESS_REG_22_ <= n5112;
    P1_ADDRESS_REG_21_ <= n5116;
    P1_ADDRESS_REG_20_ <= n5120;
    P1_ADDRESS_REG_19_ <= n5124;
    P1_ADDRESS_REG_18_ <= n5128;
    P1_ADDRESS_REG_17_ <= n5132;
    P1_ADDRESS_REG_16_ <= n5136;
    P1_ADDRESS_REG_15_ <= n5140;
    P1_ADDRESS_REG_14_ <= n5144;
    P1_ADDRESS_REG_13_ <= n5148;
    P1_ADDRESS_REG_12_ <= n5152;
    P1_ADDRESS_REG_11_ <= n5156;
    P1_ADDRESS_REG_10_ <= n5160;
    P1_ADDRESS_REG_9_ <= n5164;
    P1_ADDRESS_REG_8_ <= n5168;
    P1_ADDRESS_REG_7_ <= n5172;
    P1_ADDRESS_REG_6_ <= n5176;
    P1_ADDRESS_REG_5_ <= n5180;
    P1_ADDRESS_REG_4_ <= n5184;
    P1_ADDRESS_REG_3_ <= n5188;
    P1_ADDRESS_REG_2_ <= n5192;
    P1_ADDRESS_REG_1_ <= n5196;
    P1_ADDRESS_REG_0_ <= n5200;
    P1_STATE_REG_2_ <= n5204;
    P1_STATE_REG_1_ <= n5209;
    P1_STATE_REG_0_ <= n5214;
    P1_DATAWIDTH_REG_0_ <= n5219;
    P1_DATAWIDTH_REG_1_ <= n5224;
    P1_DATAWIDTH_REG_2_ <= n5229;
    P1_DATAWIDTH_REG_3_ <= n5234;
    P1_DATAWIDTH_REG_4_ <= n5239;
    P1_DATAWIDTH_REG_5_ <= n5244;
    P1_DATAWIDTH_REG_6_ <= n5249;
    P1_DATAWIDTH_REG_7_ <= n5254;
    P1_DATAWIDTH_REG_8_ <= n5259;
    P1_DATAWIDTH_REG_9_ <= n5264;
    P1_DATAWIDTH_REG_10_ <= n5269;
    P1_DATAWIDTH_REG_11_ <= n5274;
    P1_DATAWIDTH_REG_12_ <= n5279;
    P1_DATAWIDTH_REG_13_ <= n5284;
    P1_DATAWIDTH_REG_14_ <= n5289;
    P1_DATAWIDTH_REG_15_ <= n5294;
    P1_DATAWIDTH_REG_16_ <= n5299;
    P1_DATAWIDTH_REG_17_ <= n5304;
    P1_DATAWIDTH_REG_18_ <= n5309;
    P1_DATAWIDTH_REG_19_ <= n5314;
    P1_DATAWIDTH_REG_20_ <= n5319;
    P1_DATAWIDTH_REG_21_ <= n5324;
    P1_DATAWIDTH_REG_22_ <= n5329;
    P1_DATAWIDTH_REG_23_ <= n5334;
    P1_DATAWIDTH_REG_24_ <= n5339;
    P1_DATAWIDTH_REG_25_ <= n5344;
    P1_DATAWIDTH_REG_26_ <= n5349;
    P1_DATAWIDTH_REG_27_ <= n5354;
    P1_DATAWIDTH_REG_28_ <= n5359;
    P1_DATAWIDTH_REG_29_ <= n5364;
    P1_DATAWIDTH_REG_30_ <= n5369;
    P1_DATAWIDTH_REG_31_ <= n5374;
    P1_STATE2_REG_3_ <= n5379;
    P1_STATE2_REG_2_ <= n5384;
    P1_STATE2_REG_1_ <= n5389;
    P1_STATE2_REG_0_ <= n5394;
    P1_INSTQUEUE_REG_15__7_ <= n5399;
    P1_INSTQUEUE_REG_15__6_ <= n5404;
    P1_INSTQUEUE_REG_15__5_ <= n5409;
    P1_INSTQUEUE_REG_15__4_ <= n5414;
    P1_INSTQUEUE_REG_15__3_ <= n5419;
    P1_INSTQUEUE_REG_15__2_ <= n5424;
    P1_INSTQUEUE_REG_15__1_ <= n5429;
    P1_INSTQUEUE_REG_15__0_ <= n5434;
    P1_INSTQUEUE_REG_14__7_ <= n5439;
    P1_INSTQUEUE_REG_14__6_ <= n5444;
    P1_INSTQUEUE_REG_14__5_ <= n5449;
    P1_INSTQUEUE_REG_14__4_ <= n5454;
    P1_INSTQUEUE_REG_14__3_ <= n5459;
    P1_INSTQUEUE_REG_14__2_ <= n5464;
    P1_INSTQUEUE_REG_14__1_ <= n5469;
    P1_INSTQUEUE_REG_14__0_ <= n5474;
    P1_INSTQUEUE_REG_13__7_ <= n5479;
    P1_INSTQUEUE_REG_13__6_ <= n5484;
    P1_INSTQUEUE_REG_13__5_ <= n5489;
    P1_INSTQUEUE_REG_13__4_ <= n5494;
    P1_INSTQUEUE_REG_13__3_ <= n5499;
    P1_INSTQUEUE_REG_13__2_ <= n5504;
    P1_INSTQUEUE_REG_13__1_ <= n5509;
    P1_INSTQUEUE_REG_13__0_ <= n5514;
    P1_INSTQUEUE_REG_12__7_ <= n5519;
    P1_INSTQUEUE_REG_12__6_ <= n5524;
    P1_INSTQUEUE_REG_12__5_ <= n5529;
    P1_INSTQUEUE_REG_12__4_ <= n5534;
    P1_INSTQUEUE_REG_12__3_ <= n5539;
    P1_INSTQUEUE_REG_12__2_ <= n5544;
    P1_INSTQUEUE_REG_12__1_ <= n5549;
    P1_INSTQUEUE_REG_12__0_ <= n5554;
    P1_INSTQUEUE_REG_11__7_ <= n5559;
    P1_INSTQUEUE_REG_11__6_ <= n5564;
    P1_INSTQUEUE_REG_11__5_ <= n5569;
    P1_INSTQUEUE_REG_11__4_ <= n5574;
    P1_INSTQUEUE_REG_11__3_ <= n5579;
    P1_INSTQUEUE_REG_11__2_ <= n5584;
    P1_INSTQUEUE_REG_11__1_ <= n5589;
    P1_INSTQUEUE_REG_11__0_ <= n5594;
    P1_INSTQUEUE_REG_10__7_ <= n5599;
    P1_INSTQUEUE_REG_10__6_ <= n5604;
    P1_INSTQUEUE_REG_10__5_ <= n5609;
    P1_INSTQUEUE_REG_10__4_ <= n5614;
    P1_INSTQUEUE_REG_10__3_ <= n5619;
    P1_INSTQUEUE_REG_10__2_ <= n5624;
    P1_INSTQUEUE_REG_10__1_ <= n5629;
    P1_INSTQUEUE_REG_10__0_ <= n5634;
    P1_INSTQUEUE_REG_9__7_ <= n5639;
    P1_INSTQUEUE_REG_9__6_ <= n5644;
    P1_INSTQUEUE_REG_9__5_ <= n5649;
    P1_INSTQUEUE_REG_9__4_ <= n5654;
    P1_INSTQUEUE_REG_9__3_ <= n5659;
    P1_INSTQUEUE_REG_9__2_ <= n5664;
    P1_INSTQUEUE_REG_9__1_ <= n5669;
    P1_INSTQUEUE_REG_9__0_ <= n5674;
    P1_INSTQUEUE_REG_8__7_ <= n5679;
    P1_INSTQUEUE_REG_8__6_ <= n5684;
    P1_INSTQUEUE_REG_8__5_ <= n5689;
    P1_INSTQUEUE_REG_8__4_ <= n5694;
    P1_INSTQUEUE_REG_8__3_ <= n5699;
    P1_INSTQUEUE_REG_8__2_ <= n5704;
    P1_INSTQUEUE_REG_8__1_ <= n5709;
    P1_INSTQUEUE_REG_8__0_ <= n5714;
    P1_INSTQUEUE_REG_7__7_ <= n5719;
    P1_INSTQUEUE_REG_7__6_ <= n5724;
    P1_INSTQUEUE_REG_7__5_ <= n5729;
    P1_INSTQUEUE_REG_7__4_ <= n5734;
    P1_INSTQUEUE_REG_7__3_ <= n5739;
    P1_INSTQUEUE_REG_7__2_ <= n5744;
    P1_INSTQUEUE_REG_7__1_ <= n5749;
    P1_INSTQUEUE_REG_7__0_ <= n5754;
    P1_INSTQUEUE_REG_6__7_ <= n5759;
    P1_INSTQUEUE_REG_6__6_ <= n5764;
    P1_INSTQUEUE_REG_6__5_ <= n5769;
    P1_INSTQUEUE_REG_6__4_ <= n5774;
    P1_INSTQUEUE_REG_6__3_ <= n5779;
    P1_INSTQUEUE_REG_6__2_ <= n5784;
    P1_INSTQUEUE_REG_6__1_ <= n5789;
    P1_INSTQUEUE_REG_6__0_ <= n5794;
    P1_INSTQUEUE_REG_5__7_ <= n5799;
    P1_INSTQUEUE_REG_5__6_ <= n5804;
    P1_INSTQUEUE_REG_5__5_ <= n5809;
    P1_INSTQUEUE_REG_5__4_ <= n5814;
    P1_INSTQUEUE_REG_5__3_ <= n5819;
    P1_INSTQUEUE_REG_5__2_ <= n5824;
    P1_INSTQUEUE_REG_5__1_ <= n5829;
    P1_INSTQUEUE_REG_5__0_ <= n5834;
    P1_INSTQUEUE_REG_4__7_ <= n5839;
    P1_INSTQUEUE_REG_4__6_ <= n5844;
    P1_INSTQUEUE_REG_4__5_ <= n5849;
    P1_INSTQUEUE_REG_4__4_ <= n5854;
    P1_INSTQUEUE_REG_4__3_ <= n5859;
    P1_INSTQUEUE_REG_4__2_ <= n5864;
    P1_INSTQUEUE_REG_4__1_ <= n5869;
    P1_INSTQUEUE_REG_4__0_ <= n5874;
    P1_INSTQUEUE_REG_3__7_ <= n5879;
    P1_INSTQUEUE_REG_3__6_ <= n5884;
    P1_INSTQUEUE_REG_3__5_ <= n5889;
    P1_INSTQUEUE_REG_3__4_ <= n5894;
    P1_INSTQUEUE_REG_3__3_ <= n5899;
    P1_INSTQUEUE_REG_3__2_ <= n5904;
    P1_INSTQUEUE_REG_3__1_ <= n5909;
    P1_INSTQUEUE_REG_3__0_ <= n5914;
    P1_INSTQUEUE_REG_2__7_ <= n5919;
    P1_INSTQUEUE_REG_2__6_ <= n5924;
    P1_INSTQUEUE_REG_2__5_ <= n5929;
    P1_INSTQUEUE_REG_2__4_ <= n5934;
    P1_INSTQUEUE_REG_2__3_ <= n5939;
    P1_INSTQUEUE_REG_2__2_ <= n5944;
    P1_INSTQUEUE_REG_2__1_ <= n5949;
    P1_INSTQUEUE_REG_2__0_ <= n5954;
    P1_INSTQUEUE_REG_1__7_ <= n5959;
    P1_INSTQUEUE_REG_1__6_ <= n5964;
    P1_INSTQUEUE_REG_1__5_ <= n5969;
    P1_INSTQUEUE_REG_1__4_ <= n5974;
    P1_INSTQUEUE_REG_1__3_ <= n5979;
    P1_INSTQUEUE_REG_1__2_ <= n5984;
    P1_INSTQUEUE_REG_1__1_ <= n5989;
    P1_INSTQUEUE_REG_1__0_ <= n5994;
    P1_INSTQUEUE_REG_0__7_ <= n5999;
    P1_INSTQUEUE_REG_0__6_ <= n6004;
    P1_INSTQUEUE_REG_0__5_ <= n6009;
    P1_INSTQUEUE_REG_0__4_ <= n6014;
    P1_INSTQUEUE_REG_0__3_ <= n6019;
    P1_INSTQUEUE_REG_0__2_ <= n6024;
    P1_INSTQUEUE_REG_0__1_ <= n6029;
    P1_INSTQUEUE_REG_0__0_ <= n6034;
    P1_INSTQUEUERD_ADDR_REG_4_ <= n6039;
    P1_INSTQUEUERD_ADDR_REG_3_ <= n6044;
    P1_INSTQUEUERD_ADDR_REG_2_ <= n6049;
    P1_INSTQUEUERD_ADDR_REG_1_ <= n6054;
    P1_INSTQUEUERD_ADDR_REG_0_ <= n6059;
    P1_INSTQUEUEWR_ADDR_REG_4_ <= n6064;
    P1_INSTQUEUEWR_ADDR_REG_3_ <= n6069;
    P1_INSTQUEUEWR_ADDR_REG_2_ <= n6074;
    P1_INSTQUEUEWR_ADDR_REG_1_ <= n6079;
    P1_INSTQUEUEWR_ADDR_REG_0_ <= n6084;
    P1_INSTADDRPOINTER_REG_0_ <= n6089;
    P1_INSTADDRPOINTER_REG_1_ <= n6094;
    P1_INSTADDRPOINTER_REG_2_ <= n6099;
    P1_INSTADDRPOINTER_REG_3_ <= n6104;
    P1_INSTADDRPOINTER_REG_4_ <= n6109;
    P1_INSTADDRPOINTER_REG_5_ <= n6114;
    P1_INSTADDRPOINTER_REG_6_ <= n6119;
    P1_INSTADDRPOINTER_REG_7_ <= n6124;
    P1_INSTADDRPOINTER_REG_8_ <= n6129;
    P1_INSTADDRPOINTER_REG_9_ <= n6134;
    P1_INSTADDRPOINTER_REG_10_ <= n6139;
    P1_INSTADDRPOINTER_REG_11_ <= n6144;
    P1_INSTADDRPOINTER_REG_12_ <= n6149;
    P1_INSTADDRPOINTER_REG_13_ <= n6154;
    P1_INSTADDRPOINTER_REG_14_ <= n6159;
    P1_INSTADDRPOINTER_REG_15_ <= n6164;
    P1_INSTADDRPOINTER_REG_16_ <= n6169;
    P1_INSTADDRPOINTER_REG_17_ <= n6174;
    P1_INSTADDRPOINTER_REG_18_ <= n6179;
    P1_INSTADDRPOINTER_REG_19_ <= n6184;
    P1_INSTADDRPOINTER_REG_20_ <= n6189;
    P1_INSTADDRPOINTER_REG_21_ <= n6194;
    P1_INSTADDRPOINTER_REG_22_ <= n6199;
    P1_INSTADDRPOINTER_REG_23_ <= n6204;
    P1_INSTADDRPOINTER_REG_24_ <= n6209;
    P1_INSTADDRPOINTER_REG_25_ <= n6214;
    P1_INSTADDRPOINTER_REG_26_ <= n6219;
    P1_INSTADDRPOINTER_REG_27_ <= n6224;
    P1_INSTADDRPOINTER_REG_28_ <= n6229;
    P1_INSTADDRPOINTER_REG_29_ <= n6234;
    P1_INSTADDRPOINTER_REG_30_ <= n6239;
    P1_INSTADDRPOINTER_REG_31_ <= n6244;
    P1_PHYADDRPOINTER_REG_0_ <= n6249;
    P1_PHYADDRPOINTER_REG_1_ <= n6254;
    P1_PHYADDRPOINTER_REG_2_ <= n6259;
    P1_PHYADDRPOINTER_REG_3_ <= n6264;
    P1_PHYADDRPOINTER_REG_4_ <= n6269;
    P1_PHYADDRPOINTER_REG_5_ <= n6274;
    P1_PHYADDRPOINTER_REG_6_ <= n6279;
    P1_PHYADDRPOINTER_REG_7_ <= n6284;
    P1_PHYADDRPOINTER_REG_8_ <= n6289;
    P1_PHYADDRPOINTER_REG_9_ <= n6294;
    P1_PHYADDRPOINTER_REG_10_ <= n6299;
    P1_PHYADDRPOINTER_REG_11_ <= n6304;
    P1_PHYADDRPOINTER_REG_12_ <= n6309;
    P1_PHYADDRPOINTER_REG_13_ <= n6314;
    P1_PHYADDRPOINTER_REG_14_ <= n6319;
    P1_PHYADDRPOINTER_REG_15_ <= n6324;
    P1_PHYADDRPOINTER_REG_16_ <= n6329;
    P1_PHYADDRPOINTER_REG_17_ <= n6334;
    P1_PHYADDRPOINTER_REG_18_ <= n6339;
    P1_PHYADDRPOINTER_REG_19_ <= n6344;
    P1_PHYADDRPOINTER_REG_20_ <= n6349;
    P1_PHYADDRPOINTER_REG_21_ <= n6354;
    P1_PHYADDRPOINTER_REG_22_ <= n6359;
    P1_PHYADDRPOINTER_REG_23_ <= n6364;
    P1_PHYADDRPOINTER_REG_24_ <= n6369;
    P1_PHYADDRPOINTER_REG_25_ <= n6374;
    P1_PHYADDRPOINTER_REG_26_ <= n6379;
    P1_PHYADDRPOINTER_REG_27_ <= n6384;
    P1_PHYADDRPOINTER_REG_28_ <= n6389;
    P1_PHYADDRPOINTER_REG_29_ <= n6394;
    P1_PHYADDRPOINTER_REG_30_ <= n6399;
    P1_PHYADDRPOINTER_REG_31_ <= n6404;
    P1_LWORD_REG_15_ <= n6409;
    P1_LWORD_REG_14_ <= n6414;
    P1_LWORD_REG_13_ <= n6419;
    P1_LWORD_REG_12_ <= n6424;
    P1_LWORD_REG_11_ <= n6429;
    P1_LWORD_REG_10_ <= n6434;
    P1_LWORD_REG_9_ <= n6439;
    P1_LWORD_REG_8_ <= n6444;
    P1_LWORD_REG_7_ <= n6449;
    P1_LWORD_REG_6_ <= n6454;
    P1_LWORD_REG_5_ <= n6459;
    P1_LWORD_REG_4_ <= n6464;
    P1_LWORD_REG_3_ <= n6469;
    P1_LWORD_REG_2_ <= n6474;
    P1_LWORD_REG_1_ <= n6479;
    P1_LWORD_REG_0_ <= n6484;
    P1_UWORD_REG_14_ <= n6489;
    P1_UWORD_REG_13_ <= n6494;
    P1_UWORD_REG_12_ <= n6499;
    P1_UWORD_REG_11_ <= n6504;
    P1_UWORD_REG_10_ <= n6509;
    P1_UWORD_REG_9_ <= n6514;
    P1_UWORD_REG_8_ <= n6519;
    P1_UWORD_REG_7_ <= n6524;
    P1_UWORD_REG_6_ <= n6529;
    P1_UWORD_REG_5_ <= n6534;
    P1_UWORD_REG_4_ <= n6539;
    P1_UWORD_REG_3_ <= n6544;
    P1_UWORD_REG_2_ <= n6549;
    P1_UWORD_REG_1_ <= n6554;
    P1_UWORD_REG_0_ <= n6559;
    P1_DATAO_REG_0_ <= n6564;
    P1_DATAO_REG_1_ <= n6569;
    P1_DATAO_REG_2_ <= n6574;
    P1_DATAO_REG_3_ <= n6579;
    P1_DATAO_REG_4_ <= n6584;
    P1_DATAO_REG_5_ <= n6589;
    P1_DATAO_REG_6_ <= n6594;
    P1_DATAO_REG_7_ <= n6599;
    P1_DATAO_REG_8_ <= n6604;
    P1_DATAO_REG_9_ <= n6609;
    P1_DATAO_REG_10_ <= n6614;
    P1_DATAO_REG_11_ <= n6619;
    P1_DATAO_REG_12_ <= n6624;
    P1_DATAO_REG_13_ <= n6629;
    P1_DATAO_REG_14_ <= n6634;
    P1_DATAO_REG_15_ <= n6639;
    P1_DATAO_REG_16_ <= n6644;
    P1_DATAO_REG_17_ <= n6649;
    P1_DATAO_REG_18_ <= n6654;
    P1_DATAO_REG_19_ <= n6659;
    P1_DATAO_REG_20_ <= n6664;
    P1_DATAO_REG_21_ <= n6669;
    P1_DATAO_REG_22_ <= n6674;
    P1_DATAO_REG_23_ <= n6679;
    P1_DATAO_REG_24_ <= n6684;
    P1_DATAO_REG_25_ <= n6689;
    P1_DATAO_REG_26_ <= n6694;
    P1_DATAO_REG_27_ <= n6699;
    P1_DATAO_REG_28_ <= n6704;
    P1_DATAO_REG_29_ <= n6709;
    P1_DATAO_REG_30_ <= n6714;
    P1_DATAO_REG_31_ <= n6719;
    P1_EAX_REG_0_ <= n6724;
    P1_EAX_REG_1_ <= n6729;
    P1_EAX_REG_2_ <= n6734;
    P1_EAX_REG_3_ <= n6739;
    P1_EAX_REG_4_ <= n6744;
    P1_EAX_REG_5_ <= n6749;
    P1_EAX_REG_6_ <= n6754;
    P1_EAX_REG_7_ <= n6759;
    P1_EAX_REG_8_ <= n6764;
    P1_EAX_REG_9_ <= n6769;
    P1_EAX_REG_10_ <= n6774;
    P1_EAX_REG_11_ <= n6779;
    P1_EAX_REG_12_ <= n6784;
    P1_EAX_REG_13_ <= n6789;
    P1_EAX_REG_14_ <= n6794;
    P1_EAX_REG_15_ <= n6799;
    P1_EAX_REG_16_ <= n6804;
    P1_EAX_REG_17_ <= n6809;
    P1_EAX_REG_18_ <= n6814;
    P1_EAX_REG_19_ <= n6819;
    P1_EAX_REG_20_ <= n6824;
    P1_EAX_REG_21_ <= n6829;
    P1_EAX_REG_22_ <= n6834;
    P1_EAX_REG_23_ <= n6839;
    P1_EAX_REG_24_ <= n6844;
    P1_EAX_REG_25_ <= n6849;
    P1_EAX_REG_26_ <= n6854;
    P1_EAX_REG_27_ <= n6859;
    P1_EAX_REG_28_ <= n6864;
    P1_EAX_REG_29_ <= n6869;
    P1_EAX_REG_30_ <= n6874;
    P1_EAX_REG_31_ <= n6879;
    P1_EBX_REG_0_ <= n6884;
    P1_EBX_REG_1_ <= n6889;
    P1_EBX_REG_2_ <= n6894;
    P1_EBX_REG_3_ <= n6899;
    P1_EBX_REG_4_ <= n6904;
    P1_EBX_REG_5_ <= n6909;
    P1_EBX_REG_6_ <= n6914;
    P1_EBX_REG_7_ <= n6919;
    P1_EBX_REG_8_ <= n6924;
    P1_EBX_REG_9_ <= n6929;
    P1_EBX_REG_10_ <= n6934;
    P1_EBX_REG_11_ <= n6939;
    P1_EBX_REG_12_ <= n6944;
    P1_EBX_REG_13_ <= n6949;
    P1_EBX_REG_14_ <= n6954;
    P1_EBX_REG_15_ <= n6959;
    P1_EBX_REG_16_ <= n6964;
    P1_EBX_REG_17_ <= n6969;
    P1_EBX_REG_18_ <= n6974;
    P1_EBX_REG_19_ <= n6979;
    P1_EBX_REG_20_ <= n6984;
    P1_EBX_REG_21_ <= n6989;
    P1_EBX_REG_22_ <= n6994;
    P1_EBX_REG_23_ <= n6999;
    P1_EBX_REG_24_ <= n7004;
    P1_EBX_REG_25_ <= n7009;
    P1_EBX_REG_26_ <= n7014;
    P1_EBX_REG_27_ <= n7019;
    P1_EBX_REG_28_ <= n7024;
    P1_EBX_REG_29_ <= n7029;
    P1_EBX_REG_30_ <= n7034;
    P1_EBX_REG_31_ <= n7039;
    P1_REIP_REG_0_ <= n7044;
    P1_REIP_REG_1_ <= n7049;
    P1_REIP_REG_2_ <= n7054;
    P1_REIP_REG_3_ <= n7059;
    P1_REIP_REG_4_ <= n7064;
    P1_REIP_REG_5_ <= n7069;
    P1_REIP_REG_6_ <= n7074;
    P1_REIP_REG_7_ <= n7079;
    P1_REIP_REG_8_ <= n7084;
    P1_REIP_REG_9_ <= n7089;
    P1_REIP_REG_10_ <= n7094;
    P1_REIP_REG_11_ <= n7099;
    P1_REIP_REG_12_ <= n7104;
    P1_REIP_REG_13_ <= n7109;
    P1_REIP_REG_14_ <= n7114;
    P1_REIP_REG_15_ <= n7119;
    P1_REIP_REG_16_ <= n7124;
    P1_REIP_REG_17_ <= n7129;
    P1_REIP_REG_18_ <= n7134;
    P1_REIP_REG_19_ <= n7139;
    P1_REIP_REG_20_ <= n7144;
    P1_REIP_REG_21_ <= n7149;
    P1_REIP_REG_22_ <= n7154;
    P1_REIP_REG_23_ <= n7159;
    P1_REIP_REG_24_ <= n7164;
    P1_REIP_REG_25_ <= n7169;
    P1_REIP_REG_26_ <= n7174;
    P1_REIP_REG_27_ <= n7179;
    P1_REIP_REG_28_ <= n7184;
    P1_REIP_REG_29_ <= n7189;
    P1_REIP_REG_30_ <= n7194;
    P1_REIP_REG_31_ <= n7199;
    P1_BYTEENABLE_REG_3_ <= n7204;
    P1_BYTEENABLE_REG_2_ <= n7209;
    P1_BYTEENABLE_REG_1_ <= n7214;
    P1_BYTEENABLE_REG_0_ <= n7219;
    P1_W_R_N_REG <= n7224;
    P1_FLUSH_REG <= n7229;
    P1_MORE_REG <= n7234;
    P1_STATEBS16_REG <= n7239;
    P1_REQUESTPENDING_REG <= n7244;
    P1_D_C_N_REG <= n7249;
    P1_M_IO_N_REG <= n7254;
    P1_CODEFETCH_REG <= n7259;
    P1_ADS_N_REG <= n7264;
    P1_READREQUEST_REG <= n7268;
    P1_MEMORYFETCH_REG <= n7273;
  end
endmodule


