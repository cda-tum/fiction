// Benchmark "top" written by ABC on Mon Feb 19 11:52:41 2024

module top ( 
    txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4, xzfs,
    i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2, p2zzz1,
    qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1, vybb1,
    i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar, psrw,
    xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161, pfin,
    stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4, xz163,
    xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2, txwrd14,
    v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4, v2zzz3, iclr,
    pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11, v1zzz2, v2zzz1,
    axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7, xzfr0, enwin, ofs1,
    pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6, i2zzz5, inybb6, ofs2,
    p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7, p1zzz6, p2zzz5, rpten,
    rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7, i2zzz6, inybb5, p2zzz7,
    inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0, txwrd6, inybb0, txwrd9,
    inybb1, psync, txwrd8, vfin,
    i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p  );
  input  txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4,
    xzfs, i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2,
    p2zzz1, qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1,
    vybb1, i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar,
    psrw, xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161,
    pfin, stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4,
    xz163, xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2,
    txwrd14, v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4,
    v2zzz3, iclr, pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11,
    v1zzz2, v2zzz1, axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7,
    xzfr0, enwin, ofs1, pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6,
    i2zzz5, inybb6, ofs2, p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7,
    p1zzz6, p2zzz5, rpten, rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7,
    i2zzz6, inybb5, p2zzz7, inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0,
    txwrd6, inybb0, txwrd9, inybb1, psync, txwrd8, vfin;
  output i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p;
  wire new_n235, new_n236, new_n237, new_n238, new_n239, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n247, new_n248, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n256, new_n257, new_n258, new_n259,
    new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n274,
    new_n275, new_n277, new_n278, new_n279, new_n280, new_n281, new_n283,
    new_n284, new_n286, new_n287, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n310, new_n311, new_n313, new_n314, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n330, new_n331, new_n332,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n347, new_n348, new_n349,
    new_n350, new_n351, new_n353, new_n354, new_n356, new_n357, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n369, new_n370, new_n372, new_n373, new_n375, new_n376,
    new_n378, new_n379, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n387, new_n388, new_n389, new_n390, new_n391, new_n393,
    new_n394, new_n396, new_n397, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n405, new_n406, new_n407, new_n408, new_n409, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n431, new_n432, new_n434, new_n435,
    new_n437, new_n438, new_n440, new_n441, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n457, new_n458, new_n460, new_n461,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n473, new_n474, new_n475, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n786, new_n787, new_n789, new_n790,
    new_n792, new_n793, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n823, new_n824,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896;
  assign new_n235 = ~inzzze & inybb0;
  assign new_n236 = ~ryz & new_n235;
  assign new_n237 = inybb1 & new_n236;
  assign new_n238 = ~ryz & ~new_n235;
  assign new_n239 = i1zzz0 & new_n238;
  assign i1zzz0_p = new_n237 | new_n239;
  assign new_n241 = vybb0 & ~vzzze;
  assign new_n242 = ~ryz & new_n241;
  assign new_n243 = v1zzz1 & new_n242;
  assign new_n244 = ~ryz & ~new_n241;
  assign new_n245 = v1zzz0 & new_n244;
  assign v1zzz0_p = new_n243 | new_n245;
  assign new_n247 = inybb4 & new_n236;
  assign new_n248 = i1zzz3 & new_n238;
  assign i1zzz3_p = new_n247 | new_n248;
  assign new_n250 = inzzze & inybb0;
  assign new_n251 = ~ryz & new_n250;
  assign new_n252 = inybb3 & new_n251;
  assign new_n253 = ~ryz & ~new_n250;
  assign new_n254 = i2zzz2 & new_n253;
  assign i2zzz2_p = new_n252 | new_n254;
  assign new_n256 = ~infin & ~ryz;
  assign new_n257 = pfin & new_n256;
  assign new_n258 = p2zzz0 & new_n257;
  assign new_n259 = ~pfin & new_n256;
  assign new_n260 = ~b & ~c;
  assign new_n261 = ~txmess_n & ~new_n260;
  assign new_n262 = ~vfin & ~new_n261;
  assign new_n263 = txwrd8 & new_n262;
  assign new_n264 = ~vfin & new_n261;
  assign new_n265 = txwrd9 & new_n264;
  assign new_n266 = v2zzz0 & vfin;
  assign new_n267 = ~new_n263 & ~new_n265;
  assign new_n268 = ~new_n266 & new_n267;
  assign new_n269 = new_n259 & ~new_n268;
  assign new_n270 = infin & ~ryz;
  assign new_n271 = i2zzz0 & new_n270;
  assign new_n272 = ~new_n258 & ~new_n269;
  assign txwrd8_p = new_n271 | ~new_n272;
  assign new_n274 = v1zzz3 & new_n242;
  assign new_n275 = v1zzz2 & new_n244;
  assign v1zzz2_p = new_n274 | new_n275;
  assign new_n277 = vybb0 & vzzze;
  assign new_n278 = ~ryz & new_n277;
  assign new_n279 = v2zzz2 & new_n278;
  assign new_n280 = ~ryz & ~new_n277;
  assign new_n281 = v2zzz1 & new_n280;
  assign v2zzz1_p = new_n279 | new_n281;
  assign new_n283 = inybb5 & new_n236;
  assign new_n284 = i1zzz4 & new_n238;
  assign i1zzz4_p = new_n283 | new_n284;
  assign new_n286 = inybb4 & new_n251;
  assign new_n287 = i2zzz3 & new_n253;
  assign i2zzz3_p = new_n286 | new_n287;
  assign new_n289 = ~infin & ~pfin;
  assign new_n290 = axz1 & axz0;
  assign new_n291 = ~txmess_n & new_n290;
  assign new_n292 = a & new_n291;
  assign new_n293 = ~stw_n & ~new_n292;
  assign new_n294 = new_n289 & ~new_n293;
  assign new_n295 = ~vfin & new_n294;
  assign stw_f = ryz | new_n295;
  assign new_n297 = ~pfin & vfin;
  assign new_n298 = v2zzz1 & new_n297;
  assign new_n299 = ~pfin & new_n262;
  assign new_n300 = txwrd9 & new_n299;
  assign new_n301 = ~pfin & new_n264;
  assign new_n302 = txwrd10 & new_n301;
  assign new_n303 = p2zzz1 & pfin;
  assign new_n304 = ~new_n298 & ~new_n300;
  assign new_n305 = ~new_n302 & ~new_n303;
  assign new_n306 = new_n304 & new_n305;
  assign new_n307 = new_n256 & ~new_n306;
  assign new_n308 = i2zzz1 & new_n270;
  assign txwrd9_p = new_n307 | new_n308;
  assign new_n310 = v1zzz2 & new_n242;
  assign new_n311 = v1zzz1 & new_n244;
  assign v1zzz1_p = new_n310 | new_n311;
  assign new_n313 = v2zzz1 & new_n278;
  assign new_n314 = v2zzz0 & new_n280;
  assign v2zzz0_p = new_n313 | new_n314;
  assign new_n316 = ~iclr & ~psync;
  assign new_n317 = xz321 & xz322;
  assign new_n318 = xz324 & new_n317;
  assign new_n319 = xz323 & new_n318;
  assign new_n320 = ~xz160_n & new_n319;
  assign new_n321 = xz161 & new_n320;
  assign new_n322 = xz320 & new_n321;
  assign new_n323 = xz162 & new_n316;
  assign new_n324 = ~xz163 & new_n323;
  assign new_n325 = new_n322 & new_n324;
  assign new_n326 = xz161 & xz162;
  assign new_n327 = new_n316 & ~new_n326;
  assign new_n328 = new_n316 & ~new_n320;
  assign xz320_p = ~xz320 & new_n316;
  assign new_n330 = ~new_n328 & ~xz320_p;
  assign new_n331 = ~new_n327 & new_n330;
  assign new_n332 = xz163 & ~new_n331;
  assign xz163_p = new_n325 | new_n332;
  assign new_n334 = cbt2 & ~cbt1;
  assign new_n335 = ~cbt0 & new_n334;
  assign new_n336 = ~qpr4 & ~new_n335;
  assign new_n337 = ~qpr1 & qpr2;
  assign new_n338 = qpr0 & new_n337;
  assign new_n339 = ~qpr3 & ~new_n336;
  assign new_n340 = ~txmess_n & new_n338;
  assign new_n341 = new_n339 & new_n340;
  assign new_n342 = ~c & new_n341;
  assign new_n343 = c & ~new_n341;
  assign new_n344 = ~new_n342 & ~new_n343;
  assign c_p = ~ryz & ~new_n344;
  assign ofs1_p = ~iclr & psync;
  assign new_n347 = xzfs & ofs1_p;
  assign new_n348 = ~iclr & enwin;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = ofs1 & ofs2;
  assign new_n351 = ~new_n349 & ~new_n350;
  assign enwin_p = psrw & new_n351;
  assign new_n353 = inybb2 & new_n236;
  assign new_n354 = i1zzz1 & new_n238;
  assign i1zzz1_p = new_n353 | new_n354;
  assign new_n356 = inybb1 & new_n251;
  assign new_n357 = i2zzz0 & new_n253;
  assign i2zzz0_p = new_n356 | new_n357;
  assign new_n359 = p1zzz6 & new_n257;
  assign new_n360 = txwrd6 & new_n262;
  assign new_n361 = txwrd7 & new_n264;
  assign new_n362 = v1zzz6 & vfin;
  assign new_n363 = ~new_n360 & ~new_n361;
  assign new_n364 = ~new_n362 & new_n363;
  assign new_n365 = new_n259 & ~new_n364;
  assign new_n366 = i1zzz6 & new_n270;
  assign new_n367 = ~new_n359 & ~new_n365;
  assign txwrd6_p = new_n366 | ~new_n367;
  assign new_n369 = v1zzz5 & new_n242;
  assign new_n370 = v1zzz4 & new_n244;
  assign v1zzz4_p = new_n369 | new_n370;
  assign new_n372 = v2zzz4 & new_n278;
  assign new_n373 = v2zzz3 & new_n280;
  assign v2zzz3_p = new_n372 | new_n373;
  assign new_n375 = inybb3 & new_n236;
  assign new_n376 = i1zzz2 & new_n238;
  assign i1zzz2_p = new_n375 | new_n376;
  assign new_n378 = inybb2 & new_n251;
  assign new_n379 = i2zzz1 & new_n253;
  assign i2zzz1_p = new_n378 | new_n379;
  assign new_n381 = infin & i1zzz7;
  assign new_n382 = ~infin & pfin;
  assign new_n383 = p1zzz7 & new_n382;
  assign new_n384 = txwrd7 & new_n262;
  assign new_n385 = txwrd8 & new_n264;
  assign new_n386 = v1zzz7 & vfin;
  assign new_n387 = ~new_n384 & ~new_n385;
  assign new_n388 = ~new_n386 & new_n387;
  assign new_n389 = new_n289 & ~new_n388;
  assign new_n390 = ~new_n381 & ~new_n383;
  assign new_n391 = ~new_n389 & new_n390;
  assign txwrd7_p = ~ryz & ~new_n391;
  assign new_n393 = v1zzz4 & new_n242;
  assign new_n394 = v1zzz3 & new_n244;
  assign v1zzz3_p = new_n393 | new_n394;
  assign new_n396 = v2zzz3 & new_n278;
  assign new_n397 = v2zzz2 & new_n280;
  assign v2zzz2_p = new_n396 | new_n397;
  assign new_n399 = ~pzzze & pybb0;
  assign new_n400 = ~ryz & new_n399;
  assign new_n401 = pybb5 & new_n400;
  assign new_n402 = ~ryz & ~new_n399;
  assign new_n403 = p1zzz4 & new_n402;
  assign p1zzz4_p = new_n401 | new_n403;
  assign new_n405 = pzzze & pybb0;
  assign new_n406 = ~ryz & new_n405;
  assign new_n407 = pybb4 & new_n406;
  assign new_n408 = ~ryz & ~new_n405;
  assign new_n409 = p2zzz3 & new_n408;
  assign p2zzz3_p = new_n407 | new_n409;
  assign new_n411 = ~xz162 & new_n316;
  assign new_n412 = new_n322 & new_n411;
  assign new_n413 = ~xz161 & new_n316;
  assign new_n414 = new_n330 & ~new_n413;
  assign new_n415 = xz162 & ~new_n414;
  assign xz162_p = new_n412 | new_n415;
  assign new_n417 = ~cbt1 & ~cbt0;
  assign new_n418 = cbt2 & ~new_n417;
  assign new_n419 = ~qpr4 & ~qpr3;
  assign new_n420 = new_n338 & new_n419;
  assign new_n421 = ~b & new_n420;
  assign new_n422 = new_n418 & new_n421;
  assign new_n423 = ~txmess_n & new_n422;
  assign new_n424 = ~qpr3 & ~new_n418;
  assign new_n425 = new_n338 & ~new_n424;
  assign new_n426 = ~qpr4 & ~txmess_n;
  assign new_n427 = new_n425 & new_n426;
  assign new_n428 = b & ~new_n427;
  assign new_n429 = ~new_n423 & ~new_n428;
  assign b_p = ~ryz & ~new_n429;
  assign new_n431 = pybb4 & new_n400;
  assign new_n432 = p1zzz3 & new_n402;
  assign p1zzz3_p = new_n431 | new_n432;
  assign new_n434 = pybb3 & new_n406;
  assign new_n435 = p2zzz2 & new_n408;
  assign p2zzz2_p = new_n434 | new_n435;
  assign new_n437 = pybb3 & new_n400;
  assign new_n438 = p1zzz2 & new_n402;
  assign p1zzz2_p = new_n437 | new_n438;
  assign new_n440 = pybb2 & new_n406;
  assign new_n441 = p2zzz1 & new_n408;
  assign p2zzz1_p = new_n440 | new_n441;
  assign new_n443 = ~xz163 & new_n319;
  assign new_n444 = ~xz161 & new_n443;
  assign new_n445 = ~xz162 & xz160_n;
  assign new_n446 = new_n444 & new_n445;
  assign new_n447 = xz320 & new_n316;
  assign new_n448 = ~xzfr1 & new_n446;
  assign new_n449 = new_n447 & new_n448;
  assign new_n450 = xzfr0 & new_n449;
  assign new_n451 = ~xzfr0 & new_n316;
  assign new_n452 = new_n316 & ~new_n446;
  assign new_n453 = ~xz320_p & ~new_n452;
  assign new_n454 = ~new_n451 & new_n453;
  assign new_n455 = xzfr1 & ~new_n454;
  assign xzfr1_p = new_n450 | new_n455;
  assign new_n457 = pybb2 & new_n400;
  assign new_n458 = p1zzz1 & new_n402;
  assign p1zzz1_p = new_n457 | new_n458;
  assign new_n460 = pybb1 & new_n406;
  assign new_n461 = p2zzz0 & new_n408;
  assign p2zzz0_p = new_n460 | new_n461;
  assign new_n463 = i2zzz6 & new_n270;
  assign new_n464 = txwrd14 & new_n262;
  assign new_n465 = txwrd15 & new_n264;
  assign new_n466 = v2zzz6 & vfin;
  assign new_n467 = ~new_n464 & ~new_n465;
  assign new_n468 = ~new_n466 & new_n467;
  assign new_n469 = new_n259 & ~new_n468;
  assign new_n470 = p2zzz6 & new_n257;
  assign new_n471 = ~new_n463 & ~new_n469;
  assign txwrd14_p = new_n470 | ~new_n471;
  assign new_n473 = new_n320 & new_n447;
  assign new_n474 = ~xz161 & new_n473;
  assign new_n475 = xz161 & ~new_n330;
  assign xz161_p = new_n474 | new_n475;
  assign new_n477 = ~qpr4 & b;
  assign new_n478 = qpr3 & new_n477;
  assign new_n479 = ~qpr4 & cbt2;
  assign new_n480 = ~qpr3 & ~new_n479;
  assign new_n481 = ~new_n478 & ~new_n480;
  assign new_n482 = new_n338 & ~new_n481;
  assign new_n483 = ~txmess_n & new_n482;
  assign new_n484 = ~a & ~new_n483;
  assign a_p = ~ryz & ~new_n484;
  assign new_n486 = pybb1 & new_n400;
  assign new_n487 = p1zzz0 & new_n402;
  assign p1zzz0_p = new_n486 | new_n487;
  assign new_n489 = ~a & ~new_n482;
  assign new_n490 = ~txmess_n & ~new_n489;
  assign new_n491 = ~axz0 & new_n490;
  assign new_n492 = axz0 & ~new_n490;
  assign new_n493 = ~new_n491 & ~new_n492;
  assign axz0_p = ~ryz & ~new_n493;
  assign new_n495 = txwrd15 & new_n299;
  assign new_n496 = v2zzz7 & new_n297;
  assign new_n497 = pfin & p2zzz7;
  assign new_n498 = ~new_n495 & ~new_n496;
  assign new_n499 = ~new_n497 & new_n498;
  assign new_n500 = new_n256 & ~new_n499;
  assign new_n501 = i2zzz7 & new_n270;
  assign txwrd15_p = new_n500 | new_n501;
  assign new_n503 = ~axz1 & axz0;
  assign new_n504 = new_n490 & new_n503;
  assign new_n505 = axz0 & new_n490;
  assign new_n506 = axz1 & ~new_n505;
  assign new_n507 = ~new_n504 & ~new_n506;
  assign axz1_p = ~ryz & ~new_n507;
  assign new_n509 = rxz0 & ~rxz1;
  assign new_n510 = ~esrsum & new_n509;
  assign new_n511 = ~rxz0 & rxz1;
  assign new_n512 = esrsum & new_n511;
  assign new_n513 = ~new_n510 & ~new_n512;
  assign new_n514 = rpten & ~new_n513;
  assign new_n515 = rptwin & new_n514;
  assign new_n516 = ~axz1 & ~axz0;
  assign new_n517 = a & ~new_n516;
  assign new_n518 = new_n260 & ~new_n517;
  assign new_n519 = ~rptwin & new_n518;
  assign sbuff = rptwin | ~txmess_n;
  assign new_n521 = ~new_n519 & sbuff;
  assign new_n522 = ~qpr0 & slad1;
  assign new_n523 = qpr0 & slad0;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = qpr2 & ~new_n524;
  assign new_n526 = ~qpr1 & new_n525;
  assign new_n527 = ~qpr0 & slad3;
  assign new_n528 = qpr0 & slad2;
  assign new_n529 = ~new_n527 & ~new_n528;
  assign new_n530 = ~qpr2 & ~new_n529;
  assign new_n531 = qpr1 & new_n530;
  assign new_n532 = ~new_n526 & ~new_n531;
  assign new_n533 = ~qpr3 & ~new_n521;
  assign new_n534 = ~qpr4 & new_n533;
  assign new_n535 = ~new_n532 & new_n534;
  assign new_n536 = txwrd0 & ~new_n517;
  assign new_n537 = ~new_n260 & new_n536;
  assign new_n538 = ~mmerr & new_n503;
  assign new_n539 = ~comppar & axz0;
  assign new_n540 = esrsum & ~axz0;
  assign new_n541 = ~new_n539 & ~new_n540;
  assign new_n542 = axz1 & ~new_n541;
  assign new_n543 = ~new_n538 & ~new_n542;
  assign new_n544 = a & ~new_n543;
  assign new_n545 = ~new_n537 & ~new_n544;
  assign new_n546 = ~txmess_n & ~new_n545;
  assign new_n547 = ~rptwin & new_n546;
  assign new_n548 = ~new_n515 & ~new_n535;
  assign new_n549 = ~new_n547 & new_n548;
  assign td_p = ~ryz & ~new_n549;
  assign ofs2_p = ~iclr & ofs1;
  assign new_n552 = ofs2 & ofs2_p;
  assign new_n553 = ~iclr & xzfr1;
  assign fsesr_p = new_n552 | new_n553;
  assign new_n555 = rxz0 & rxz1;
  assign new_n556 = rptwin & ~new_n555;
  assign new_n557 = xzfs & ~slad3;
  assign new_n558 = ~slad2 & psync;
  assign new_n559 = new_n557 & new_n558;
  assign new_n560 = ~slad1 & new_n559;
  assign new_n561 = ~slad0 & new_n560;
  assign new_n562 = ~xz162 & ~slad2;
  assign new_n563 = xz162 & slad2;
  assign new_n564 = ~new_n562 & ~new_n563;
  assign new_n565 = ~xz163 & ~slad3;
  assign new_n566 = xz163 & slad3;
  assign new_n567 = ~new_n565 & ~new_n566;
  assign new_n568 = ~new_n564 & ~new_n567;
  assign new_n569 = ~xz161 & ~slad1;
  assign new_n570 = xz161 & slad1;
  assign new_n571 = ~new_n569 & ~new_n570;
  assign new_n572 = xz323 & new_n317;
  assign new_n573 = xz320 & new_n572;
  assign new_n574 = ~slad0 & xz160_n;
  assign new_n575 = slad0 & ~xz160_n;
  assign new_n576 = ~new_n574 & ~new_n575;
  assign new_n577 = new_n568 & ~new_n571;
  assign new_n578 = enwin & new_n577;
  assign new_n579 = new_n573 & new_n578;
  assign new_n580 = xz324 & new_n579;
  assign new_n581 = ~new_n576 & new_n580;
  assign new_n582 = ~new_n556 & ~new_n561;
  assign new_n583 = ~new_n581 & new_n582;
  assign rptwin_p = ~ryz & ~new_n583;
  assign new_n585 = txwrd12 & new_n262;
  assign new_n586 = txwrd13 & new_n264;
  assign new_n587 = v2zzz4 & vfin;
  assign new_n588 = ~new_n585 & ~new_n586;
  assign new_n589 = ~new_n587 & new_n588;
  assign new_n590 = new_n289 & ~new_n589;
  assign new_n591 = infin & i2zzz4;
  assign new_n592 = p2zzz4 & new_n382;
  assign new_n593 = ~new_n590 & ~new_n591;
  assign new_n594 = ~new_n592 & new_n593;
  assign txwrd12_p = ~ryz & ~new_n594;
  assign new_n596 = txwrd11 & new_n262;
  assign new_n597 = txwrd12 & new_n264;
  assign new_n598 = v2zzz3 & vfin;
  assign new_n599 = ~new_n596 & ~new_n597;
  assign new_n600 = ~new_n598 & new_n599;
  assign new_n601 = new_n289 & ~new_n600;
  assign new_n602 = i2zzz3 & infin;
  assign new_n603 = p2zzz3 & new_n382;
  assign new_n604 = ~new_n601 & ~new_n602;
  assign new_n605 = ~new_n603 & new_n604;
  assign txwrd11_p = ~ryz & ~new_n605;
  assign new_n607 = ~xz322 & new_n447;
  assign new_n608 = xz321 & new_n607;
  assign new_n609 = ~xz321 & new_n316;
  assign new_n610 = ~xz320_p & ~new_n609;
  assign new_n611 = xz322 & ~new_n610;
  assign xz322_p = new_n608 | new_n611;
  assign new_n613 = pybb8 & new_n406;
  assign new_n614 = p2zzz7 & new_n408;
  assign p2zzz7_p = new_n613 | new_n614;
  assign new_n616 = i2zzz5 & new_n270;
  assign new_n617 = txwrd13 & new_n262;
  assign new_n618 = txwrd14 & new_n264;
  assign new_n619 = v2zzz5 & vfin;
  assign new_n620 = ~new_n617 & ~new_n618;
  assign new_n621 = ~new_n619 & new_n620;
  assign new_n622 = new_n259 & ~new_n621;
  assign new_n623 = p2zzz5 & new_n257;
  assign new_n624 = ~new_n616 & ~new_n622;
  assign txwrd13_p = new_n623 | ~new_n624;
  assign new_n626 = new_n316 & new_n573;
  assign new_n627 = ~xz324 & new_n626;
  assign new_n628 = xz323 & xz322;
  assign new_n629 = new_n316 & ~new_n628;
  assign new_n630 = new_n610 & ~new_n629;
  assign new_n631 = xz324 & ~new_n630;
  assign xz324_p = new_n627 | new_n631;
  assign new_n633 = xzfs & ~iclr;
  assign new_n634 = ~ofs1_p & ~new_n633;
  assign new_n635 = ~new_n350 & ~new_n634;
  assign xzfs_p = psrw & new_n635;
  assign new_n637 = pybb8 & new_n400;
  assign new_n638 = p1zzz7 & new_n402;
  assign p1zzz7_p = new_n637 | new_n638;
  assign new_n640 = pybb7 & new_n406;
  assign new_n641 = p2zzz6 & new_n408;
  assign p2zzz6_p = new_n640 | new_n641;
  assign new_n643 = new_n446 & new_n447;
  assign new_n644 = ~xzfr0 & new_n643;
  assign new_n645 = xzfr0 & ~new_n453;
  assign xzfr0_p = new_n644 | new_n645;
  assign new_n647 = pybb7 & new_n400;
  assign new_n648 = p1zzz6 & new_n402;
  assign p1zzz6_p = new_n647 | new_n648;
  assign new_n650 = pybb6 & new_n406;
  assign new_n651 = p2zzz5 & new_n408;
  assign p2zzz5_p = new_n650 | new_n651;
  assign new_n653 = ~slad1 & ~slad2;
  assign new_n654 = xzfs & new_n653;
  assign new_n655 = ~slad0 & new_n654;
  assign new_n656 = ofs1_p & new_n655;
  assign new_n657 = ~slad3 & new_n656;
  assign new_n658 = ~rptwin & ~new_n581;
  assign new_n659 = ~iclr & ~new_n658;
  assign new_n660 = ~new_n657 & ~new_n659;
  assign new_n661 = ~rxz1 & ~new_n660;
  assign new_n662 = rxz0 & new_n661;
  assign new_n663 = ~iclr & ~rxz0;
  assign new_n664 = xz162 & ~slad2;
  assign new_n665 = xz163 & ~slad3;
  assign new_n666 = ~new_n664 & ~new_n665;
  assign new_n667 = ~psync & ~new_n666;
  assign new_n668 = xz161 & ~slad1;
  assign new_n669 = enwin & ~new_n668;
  assign new_n670 = ~slad0 & ~xz160_n;
  assign new_n671 = new_n319 & ~new_n670;
  assign new_n672 = new_n669 & new_n671;
  assign new_n673 = ~new_n559 & ~new_n672;
  assign new_n674 = xz320 & new_n666;
  assign new_n675 = enwin & new_n674;
  assign new_n676 = xz161 & new_n671;
  assign new_n677 = new_n675 & new_n676;
  assign new_n678 = slad1 & ~new_n677;
  assign new_n679 = xz320 & ~new_n664;
  assign new_n680 = xz163 & new_n679;
  assign new_n681 = slad3 & ~new_n680;
  assign new_n682 = xz320 & ~new_n665;
  assign new_n683 = xz162 & new_n682;
  assign new_n684 = slad2 & ~new_n683;
  assign new_n685 = new_n669 & new_n674;
  assign new_n686 = new_n320 & new_n685;
  assign new_n687 = slad0 & ~new_n686;
  assign new_n688 = ~xzfs & ~new_n674;
  assign new_n689 = ~new_n667 & ~new_n673;
  assign new_n690 = ~new_n678 & ~new_n681;
  assign new_n691 = new_n689 & new_n690;
  assign new_n692 = ~new_n684 & ~new_n687;
  assign new_n693 = ~new_n688 & new_n692;
  assign new_n694 = new_n691 & new_n693;
  assign new_n695 = ~iclr & ~new_n694;
  assign new_n696 = ~xz320_p & ~new_n695;
  assign new_n697 = ~rptwin & ~new_n696;
  assign new_n698 = ~new_n663 & ~new_n697;
  assign new_n699 = rxz1 & ~new_n698;
  assign rxz1_p = new_n662 | new_n699;
  assign new_n701 = ~qpr3 & ~new_n532;
  assign new_n702 = ~qpr4 & new_n701;
  assign new_n703 = new_n260 & new_n702;
  assign new_n704 = txwrd0 & ~new_n260;
  assign new_n705 = ~new_n703 & ~new_n704;
  assign new_n706 = ~new_n517 & new_n705;
  assign new_n707 = ~txmess_n & ~new_n706;
  assign new_n708 = comppar & ~new_n707;
  assign new_n709 = ~comppar & ~new_n517;
  assign new_n710 = ~txmess_n & new_n709;
  assign new_n711 = ~new_n705 & new_n710;
  assign new_n712 = ~esrsum & axz1;
  assign new_n713 = mmerr & axz0;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = comppar & ~new_n714;
  assign new_n716 = esrsum & axz1;
  assign new_n717 = ~mmerr & axz0;
  assign new_n718 = ~new_n716 & ~new_n717;
  assign new_n719 = ~comppar & ~txmess_n;
  assign new_n720 = ~new_n718 & new_n719;
  assign new_n721 = ~new_n715 & ~new_n720;
  assign new_n722 = ~new_n291 & new_n721;
  assign new_n723 = a & ~new_n722;
  assign new_n724 = ~new_n708 & ~new_n711;
  assign new_n725 = ~new_n723 & new_n724;
  assign comppar_p = ~ryz & ~new_n725;
  assign new_n727 = pybb6 & new_n400;
  assign new_n728 = p1zzz5 & new_n402;
  assign p1zzz5_p = new_n727 | new_n728;
  assign new_n730 = pybb5 & new_n406;
  assign new_n731 = p2zzz4 & new_n408;
  assign p2zzz4_p = new_n730 | new_n731;
  assign new_n733 = rxz0 & ~new_n696;
  assign new_n734 = ~rptwin & new_n733;
  assign new_n735 = ~rxz0 & ~new_n660;
  assign rxz0_p = new_n734 | new_n735;
  assign new_n737 = new_n317 & new_n447;
  assign new_n738 = ~xz323 & new_n737;
  assign new_n739 = ~xz322 & new_n316;
  assign new_n740 = new_n610 & ~new_n739;
  assign new_n741 = xz323 & ~new_n740;
  assign xz323_p = new_n738 | new_n741;
  assign new_n743 = inybb8 & new_n236;
  assign new_n744 = i1zzz7 & new_n238;
  assign i1zzz7_p = new_n743 | new_n744;
  assign new_n746 = inybb7 & new_n251;
  assign new_n747 = i2zzz6 & new_n253;
  assign i2zzz6_p = new_n746 | new_n747;
  assign ryz_p = iclr | new_n292;
  assign new_n750 = p1zzz4 & new_n257;
  assign new_n751 = txwrd4 & new_n262;
  assign new_n752 = txwrd5 & new_n264;
  assign new_n753 = v1zzz4 & vfin;
  assign new_n754 = ~new_n751 & ~new_n752;
  assign new_n755 = ~new_n753 & new_n754;
  assign new_n756 = new_n259 & ~new_n755;
  assign new_n757 = i1zzz4 & new_n270;
  assign new_n758 = ~new_n750 & ~new_n756;
  assign txwrd4_p = new_n757 | ~new_n758;
  assign new_n760 = v1zzz7 & new_n242;
  assign new_n761 = v1zzz6 & new_n244;
  assign v1zzz6_p = new_n760 | new_n761;
  assign new_n763 = v2zzz6 & new_n278;
  assign new_n764 = v2zzz5 & new_n280;
  assign v2zzz5_p = new_n763 | new_n764;
  assign new_n766 = new_n316 & ~new_n319;
  assign new_n767 = ~xz320_p & ~new_n766;
  assign new_n768 = xz160_n & ~new_n767;
  assign xz160_f = new_n473 | new_n768;
  assign new_n770 = inybb8 & new_n251;
  assign new_n771 = i2zzz7 & new_n253;
  assign i2zzz7_p = new_n770 | new_n771;
  assign new_n773 = p1zzz5 & new_n257;
  assign new_n774 = txwrd5 & new_n262;
  assign new_n775 = txwrd6 & new_n264;
  assign new_n776 = v1zzz5 & vfin;
  assign new_n777 = ~new_n774 & ~new_n775;
  assign new_n778 = ~new_n776 & new_n777;
  assign new_n779 = new_n259 & ~new_n778;
  assign new_n780 = i1zzz5 & new_n270;
  assign new_n781 = ~new_n773 & ~new_n779;
  assign txwrd5_p = new_n780 | ~new_n781;
  assign new_n783 = v1zzz6 & new_n242;
  assign new_n784 = v1zzz5 & new_n244;
  assign v1zzz5_p = new_n783 | new_n784;
  assign new_n786 = v2zzz5 & new_n278;
  assign new_n787 = v2zzz4 & new_n280;
  assign v2zzz4_p = new_n786 | new_n787;
  assign new_n789 = inybb6 & new_n236;
  assign new_n790 = i1zzz5 & new_n238;
  assign i1zzz5_p = new_n789 | new_n790;
  assign new_n792 = inybb5 & new_n251;
  assign new_n793 = i2zzz4 & new_n253;
  assign i2zzz4_p = new_n792 | new_n793;
  assign new_n795 = ~vfin & new_n289;
  assign new_n796 = txmess_n & new_n795;
  assign txmess_f = ryz | new_n796;
  assign new_n798 = qpr0 & ~txmess_f;
  assign new_n799 = qpr1 & new_n798;
  assign new_n800 = qpr3 & new_n799;
  assign new_n801 = ~qpr4 & new_n800;
  assign new_n802 = qpr2 & new_n801;
  assign new_n803 = qpr0 & ~new_n796;
  assign new_n804 = qpr1 & new_n803;
  assign new_n805 = qpr2 & new_n804;
  assign new_n806 = qpr3 & new_n805;
  assign new_n807 = qpr4 & ~ryz;
  assign new_n808 = ~new_n806 & new_n807;
  assign qpr4_p = new_n802 | new_n808;
  assign new_n810 = i1zzz2 & new_n270;
  assign new_n811 = v1zzz2 & new_n297;
  assign new_n812 = txwrd2 & new_n299;
  assign new_n813 = txwrd3 & new_n301;
  assign new_n814 = p1zzz2 & pfin;
  assign new_n815 = ~new_n811 & ~new_n812;
  assign new_n816 = ~new_n813 & ~new_n814;
  assign new_n817 = new_n815 & new_n816;
  assign new_n818 = new_n256 & ~new_n817;
  assign txwrd2_p = new_n810 | new_n818;
  assign new_n820 = vybb1 & new_n278;
  assign new_n821 = v2zzz7 & new_n280;
  assign v2zzz7_p = new_n820 | new_n821;
  assign new_n823 = inybb7 & new_n236;
  assign new_n824 = i1zzz6 & new_n238;
  assign i1zzz6_p = new_n823 | new_n824;
  assign new_n826 = inybb6 & new_n251;
  assign new_n827 = i2zzz5 & new_n253;
  assign i2zzz5_p = new_n826 | new_n827;
  assign new_n829 = p1zzz3 & new_n257;
  assign new_n830 = txwrd3 & new_n262;
  assign new_n831 = txwrd4 & new_n264;
  assign new_n832 = v1zzz3 & vfin;
  assign new_n833 = ~new_n830 & ~new_n831;
  assign new_n834 = ~new_n832 & new_n833;
  assign new_n835 = new_n259 & ~new_n834;
  assign new_n836 = i1zzz3 & new_n270;
  assign new_n837 = ~new_n829 & ~new_n835;
  assign txwrd3_p = new_n836 | ~new_n837;
  assign new_n839 = vybb1 & new_n242;
  assign new_n840 = v1zzz7 & new_n244;
  assign v1zzz7_p = new_n839 | new_n840;
  assign new_n842 = v2zzz7 & new_n278;
  assign new_n843 = v2zzz6 & new_n280;
  assign v2zzz6_p = new_n842 | new_n843;
  assign new_n845 = ~ryz & ~new_n804;
  assign new_n846 = qpr2 & new_n845;
  assign new_n847 = ~qpr2 & new_n799;
  assign qpr2_p = new_n846 | new_n847;
  assign new_n849 = txwrd0 & new_n262;
  assign new_n850 = txwrd1 & new_n264;
  assign new_n851 = v1zzz0 & vfin;
  assign new_n852 = ~new_n849 & ~new_n850;
  assign new_n853 = ~new_n851 & new_n852;
  assign new_n854 = new_n289 & ~new_n853;
  assign new_n855 = p1zzz0 & new_n382;
  assign new_n856 = i1zzz0 & infin;
  assign new_n857 = ~new_n854 & ~new_n855;
  assign new_n858 = ~new_n856 & new_n857;
  assign txwrd0_p = ~ryz & ~new_n858;
  assign new_n860 = ~ryz & ~new_n805;
  assign new_n861 = qpr3 & new_n860;
  assign new_n862 = ~qpr3 & new_n799;
  assign new_n863 = qpr2 & new_n862;
  assign qpr3_p = new_n861 | new_n863;
  assign new_n865 = v1zzz1 & new_n297;
  assign new_n866 = txwrd1 & new_n299;
  assign new_n867 = txwrd2 & new_n301;
  assign new_n868 = p1zzz1 & pfin;
  assign new_n869 = ~new_n865 & ~new_n866;
  assign new_n870 = ~new_n867 & ~new_n868;
  assign new_n871 = new_n869 & new_n870;
  assign new_n872 = new_n256 & ~new_n871;
  assign new_n873 = i1zzz1 & new_n270;
  assign txwrd1_p = new_n872 | new_n873;
  assign new_n875 = xz321 & xz320_p;
  assign new_n876 = ~xz321 & new_n447;
  assign xz321_p = new_n875 | new_n876;
  assign new_n878 = qpr0 & new_n796;
  assign new_n879 = ~ryz & new_n878;
  assign new_n880 = ~qpr0 & ~txmess_f;
  assign qpr0_p = new_n879 | new_n880;
  assign new_n882 = ~ryz & ~new_n803;
  assign new_n883 = qpr1 & new_n882;
  assign new_n884 = ~qpr1 & ~txmess_f;
  assign new_n885 = qpr0 & new_n884;
  assign qpr1_p = new_n883 | new_n885;
  assign new_n887 = txwrd10 & new_n262;
  assign new_n888 = txwrd11 & new_n264;
  assign new_n889 = v2zzz2 & vfin;
  assign new_n890 = ~new_n887 & ~new_n888;
  assign new_n891 = ~new_n889 & new_n890;
  assign new_n892 = new_n289 & ~new_n891;
  assign new_n893 = infin & i2zzz2;
  assign new_n894 = p2zzz2 & new_n382;
  assign new_n895 = ~new_n892 & ~new_n893;
  assign new_n896 = ~new_n894 & new_n895;
  assign txwrd10_p = ~ryz & ~new_n896;
endmodule


