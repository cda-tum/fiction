// Benchmark "top" written by ABC on Mon Feb 19 11:52:44 2024

module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, px,
    py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0, pt0, pu0,
    pv0, pw0, px0  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, px, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po;
  output ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0, pt0, pu0,
    pv0, pw0, px0;
  wire new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57,
    new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n137, new_n138, new_n139, new_n140,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n207, new_n208, new_n209, new_n210,
    new_n211, new_n212, new_n213, new_n214, new_n215, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n287, new_n288,
    new_n289;
  assign new_n51 = ~pp & ~pg0;
  assign new_n52 = ~pf0 & ~pg0;
  assign new_n53 = ~pp & ~pf0;
  assign new_n54 = ~new_n51 & ~new_n52;
  assign new_n55 = ~new_n53 & new_n54;
  assign new_n56 = ~po & ~new_n55;
  assign new_n57 = ~pe0 & ~new_n55;
  assign new_n58 = ~pe0 & ~po;
  assign new_n59 = ~new_n56 & ~new_n57;
  assign new_n60 = ~new_n58 & new_n59;
  assign new_n61 = ~pn & ~new_n60;
  assign new_n62 = ~pd0 & ~new_n60;
  assign new_n63 = ~pd0 & ~pn;
  assign new_n64 = ~new_n61 & ~new_n62;
  assign new_n65 = ~new_n63 & new_n64;
  assign new_n66 = ~pm & ~new_n65;
  assign new_n67 = ~pc0 & ~new_n65;
  assign new_n68 = ~pc0 & ~pm;
  assign new_n69 = ~new_n66 & ~new_n67;
  assign new_n70 = ~new_n68 & new_n69;
  assign new_n71 = ~pl & ~new_n70;
  assign new_n72 = ~pb0 & ~new_n70;
  assign new_n73 = ~pb0 & ~pl;
  assign new_n74 = ~new_n71 & ~new_n72;
  assign new_n75 = ~new_n73 & new_n74;
  assign new_n76 = ~pk & ~new_n75;
  assign new_n77 = ~pa0 & ~new_n75;
  assign new_n78 = ~pa0 & ~pk;
  assign new_n79 = ~new_n76 & ~new_n77;
  assign new_n80 = ~new_n78 & new_n79;
  assign new_n81 = ~pj & ~new_n80;
  assign new_n82 = ~pz & ~new_n80;
  assign new_n83 = ~pz & ~pj;
  assign new_n84 = ~new_n81 & ~new_n82;
  assign new_n85 = ~new_n83 & new_n84;
  assign new_n86 = ~pi & ~new_n85;
  assign new_n87 = ~py & ~new_n85;
  assign new_n88 = ~py & ~pi;
  assign new_n89 = ~new_n86 & ~new_n87;
  assign new_n90 = ~new_n88 & new_n89;
  assign new_n91 = ~ph & ~new_n90;
  assign new_n92 = ~px & ~new_n90;
  assign new_n93 = ~px & ~ph;
  assign new_n94 = ~new_n91 & ~new_n92;
  assign new_n95 = ~new_n93 & new_n94;
  assign new_n96 = ~pg & ~new_n95;
  assign new_n97 = ~pw & ~new_n95;
  assign new_n98 = ~pw & ~pg;
  assign new_n99 = ~new_n96 & ~new_n97;
  assign new_n100 = ~new_n98 & new_n99;
  assign new_n101 = ~pf & ~new_n100;
  assign new_n102 = ~pv & ~new_n100;
  assign new_n103 = ~pv & ~pf;
  assign new_n104 = ~new_n101 & ~new_n102;
  assign new_n105 = ~new_n103 & new_n104;
  assign new_n106 = ~pe & ~new_n105;
  assign new_n107 = ~pu & ~new_n105;
  assign new_n108 = ~pu & ~pe;
  assign new_n109 = ~new_n106 & ~new_n107;
  assign new_n110 = ~new_n108 & new_n109;
  assign new_n111 = ~pd & ~new_n110;
  assign new_n112 = ~pt & ~new_n110;
  assign new_n113 = ~pt & ~pd;
  assign new_n114 = ~new_n111 & ~new_n112;
  assign new_n115 = ~new_n113 & new_n114;
  assign new_n116 = ~pc & ~new_n115;
  assign new_n117 = ~ps & ~new_n115;
  assign new_n118 = ~ps & ~pc;
  assign new_n119 = ~new_n116 & ~new_n117;
  assign new_n120 = ~new_n118 & new_n119;
  assign new_n121 = ~pb & ~new_n120;
  assign new_n122 = ~pr & ~new_n120;
  assign new_n123 = ~pr & ~pb;
  assign new_n124 = ~new_n121 & ~new_n122;
  assign new_n125 = ~new_n123 & new_n124;
  assign new_n126 = ~pq & new_n125;
  assign new_n127 = pa & new_n126;
  assign new_n128 = ~pq & ~new_n125;
  assign new_n129 = ~pa & new_n128;
  assign new_n130 = pq & new_n125;
  assign new_n131 = ~pa & new_n130;
  assign new_n132 = pq & ~new_n125;
  assign new_n133 = pa & new_n132;
  assign new_n134 = ~new_n131 & ~new_n133;
  assign new_n135 = ~new_n127 & ~new_n129;
  assign ph0 = new_n134 & new_n135;
  assign new_n137 = ~pr & new_n120;
  assign new_n138 = pb & new_n137;
  assign new_n139 = ~pb & new_n122;
  assign new_n140 = pr & new_n120;
  assign new_n141 = ~pb & new_n140;
  assign new_n142 = pr & ~new_n120;
  assign new_n143 = pb & new_n142;
  assign new_n144 = ~new_n141 & ~new_n143;
  assign new_n145 = ~new_n138 & ~new_n139;
  assign pi0 = new_n144 & new_n145;
  assign new_n147 = ~ps & new_n115;
  assign new_n148 = pc & new_n147;
  assign new_n149 = ~pc & new_n117;
  assign new_n150 = ps & new_n115;
  assign new_n151 = ~pc & new_n150;
  assign new_n152 = ps & ~new_n115;
  assign new_n153 = pc & new_n152;
  assign new_n154 = ~new_n151 & ~new_n153;
  assign new_n155 = ~new_n148 & ~new_n149;
  assign pj0 = new_n154 & new_n155;
  assign new_n157 = ~pt & new_n110;
  assign new_n158 = pd & new_n157;
  assign new_n159 = ~pd & new_n112;
  assign new_n160 = pt & new_n110;
  assign new_n161 = ~pd & new_n160;
  assign new_n162 = pt & ~new_n110;
  assign new_n163 = pd & new_n162;
  assign new_n164 = ~new_n161 & ~new_n163;
  assign new_n165 = ~new_n158 & ~new_n159;
  assign pk0 = new_n164 & new_n165;
  assign new_n167 = ~pu & new_n105;
  assign new_n168 = pe & new_n167;
  assign new_n169 = ~pe & new_n107;
  assign new_n170 = pu & new_n105;
  assign new_n171 = ~pe & new_n170;
  assign new_n172 = pu & ~new_n105;
  assign new_n173 = pe & new_n172;
  assign new_n174 = ~new_n171 & ~new_n173;
  assign new_n175 = ~new_n168 & ~new_n169;
  assign pl0 = new_n174 & new_n175;
  assign new_n177 = ~pv & new_n100;
  assign new_n178 = pf & new_n177;
  assign new_n179 = ~pf & new_n102;
  assign new_n180 = pv & new_n100;
  assign new_n181 = ~pf & new_n180;
  assign new_n182 = pv & ~new_n100;
  assign new_n183 = pf & new_n182;
  assign new_n184 = ~new_n181 & ~new_n183;
  assign new_n185 = ~new_n178 & ~new_n179;
  assign pm0 = new_n184 & new_n185;
  assign new_n187 = ~pw & new_n95;
  assign new_n188 = pg & new_n187;
  assign new_n189 = ~pg & new_n97;
  assign new_n190 = pw & new_n95;
  assign new_n191 = ~pg & new_n190;
  assign new_n192 = pw & ~new_n95;
  assign new_n193 = pg & new_n192;
  assign new_n194 = ~new_n191 & ~new_n193;
  assign new_n195 = ~new_n188 & ~new_n189;
  assign pn0 = new_n194 & new_n195;
  assign new_n197 = ~px & new_n90;
  assign new_n198 = ph & new_n197;
  assign new_n199 = ~ph & new_n92;
  assign new_n200 = px & new_n90;
  assign new_n201 = ~ph & new_n200;
  assign new_n202 = px & ~new_n90;
  assign new_n203 = ph & new_n202;
  assign new_n204 = ~new_n201 & ~new_n203;
  assign new_n205 = ~new_n198 & ~new_n199;
  assign po0 = new_n204 & new_n205;
  assign new_n207 = ~py & new_n85;
  assign new_n208 = pi & new_n207;
  assign new_n209 = ~pi & new_n87;
  assign new_n210 = py & new_n85;
  assign new_n211 = ~pi & new_n210;
  assign new_n212 = py & ~new_n85;
  assign new_n213 = pi & new_n212;
  assign new_n214 = ~new_n211 & ~new_n213;
  assign new_n215 = ~new_n208 & ~new_n209;
  assign pp0 = new_n214 & new_n215;
  assign new_n217 = ~pz & new_n80;
  assign new_n218 = pj & new_n217;
  assign new_n219 = ~pj & new_n82;
  assign new_n220 = pz & new_n80;
  assign new_n221 = ~pj & new_n220;
  assign new_n222 = pz & ~new_n80;
  assign new_n223 = pj & new_n222;
  assign new_n224 = ~new_n221 & ~new_n223;
  assign new_n225 = ~new_n218 & ~new_n219;
  assign pq0 = new_n224 & new_n225;
  assign new_n227 = ~pa0 & new_n75;
  assign new_n228 = pk & new_n227;
  assign new_n229 = ~pk & new_n77;
  assign new_n230 = pa0 & new_n75;
  assign new_n231 = ~pk & new_n230;
  assign new_n232 = pa0 & ~new_n75;
  assign new_n233 = pk & new_n232;
  assign new_n234 = ~new_n231 & ~new_n233;
  assign new_n235 = ~new_n228 & ~new_n229;
  assign pr0 = new_n234 & new_n235;
  assign new_n237 = ~pb0 & new_n70;
  assign new_n238 = pl & new_n237;
  assign new_n239 = ~pl & new_n72;
  assign new_n240 = pb0 & new_n70;
  assign new_n241 = ~pl & new_n240;
  assign new_n242 = pb0 & ~new_n70;
  assign new_n243 = pl & new_n242;
  assign new_n244 = ~new_n241 & ~new_n243;
  assign new_n245 = ~new_n238 & ~new_n239;
  assign ps0 = new_n244 & new_n245;
  assign new_n247 = ~pc0 & new_n65;
  assign new_n248 = pm & new_n247;
  assign new_n249 = ~pm & new_n67;
  assign new_n250 = pc0 & new_n65;
  assign new_n251 = ~pm & new_n250;
  assign new_n252 = pc0 & ~new_n65;
  assign new_n253 = pm & new_n252;
  assign new_n254 = ~new_n251 & ~new_n253;
  assign new_n255 = ~new_n248 & ~new_n249;
  assign pt0 = new_n254 & new_n255;
  assign new_n257 = ~pd0 & new_n60;
  assign new_n258 = pn & new_n257;
  assign new_n259 = ~pn & new_n62;
  assign new_n260 = pd0 & new_n60;
  assign new_n261 = ~pn & new_n260;
  assign new_n262 = pd0 & ~new_n60;
  assign new_n263 = pn & new_n262;
  assign new_n264 = ~new_n261 & ~new_n263;
  assign new_n265 = ~new_n258 & ~new_n259;
  assign pu0 = new_n264 & new_n265;
  assign new_n267 = ~pe0 & new_n55;
  assign new_n268 = po & new_n267;
  assign new_n269 = ~po & new_n57;
  assign new_n270 = pe0 & new_n55;
  assign new_n271 = ~po & new_n270;
  assign new_n272 = pe0 & ~new_n55;
  assign new_n273 = po & new_n272;
  assign new_n274 = ~new_n271 & ~new_n273;
  assign new_n275 = ~new_n268 & ~new_n269;
  assign pv0 = new_n274 & new_n275;
  assign new_n277 = ~pp & new_n52;
  assign new_n278 = ~pf0 & pg0;
  assign new_n279 = pp & new_n278;
  assign new_n280 = pf0 & ~pg0;
  assign new_n281 = pp & new_n280;
  assign new_n282 = pf0 & pg0;
  assign new_n283 = ~pp & new_n282;
  assign new_n284 = ~new_n281 & ~new_n283;
  assign new_n285 = ~new_n277 & ~new_n279;
  assign pw0 = new_n284 & new_n285;
  assign new_n287 = ~pa & ~new_n125;
  assign new_n288 = ~pq & ~pa;
  assign new_n289 = ~new_n128 & ~new_n287;
  assign px0 = ~new_n288 & new_n289;
endmodule


