// Benchmark "b15" written by ABC on Wed Sep  5 10:17:20 2018

module b15 ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, NA_N, BS16_N, READY_N, HOLD,
    BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, NA_N, BS16_N, READY_N, HOLD;
  output BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_;
  reg BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, STATE_REG_2_, STATE_REG_1_, STATE_REG_0_,
    DATAWIDTH_REG_0_, DATAWIDTH_REG_1_, DATAWIDTH_REG_2_, DATAWIDTH_REG_3_,
    DATAWIDTH_REG_4_, DATAWIDTH_REG_5_, DATAWIDTH_REG_6_, DATAWIDTH_REG_7_,
    DATAWIDTH_REG_8_, DATAWIDTH_REG_9_, DATAWIDTH_REG_10_,
    DATAWIDTH_REG_11_, DATAWIDTH_REG_12_, DATAWIDTH_REG_13_,
    DATAWIDTH_REG_14_, DATAWIDTH_REG_15_, DATAWIDTH_REG_16_,
    DATAWIDTH_REG_17_, DATAWIDTH_REG_18_, DATAWIDTH_REG_19_,
    DATAWIDTH_REG_20_, DATAWIDTH_REG_21_, DATAWIDTH_REG_22_,
    DATAWIDTH_REG_23_, DATAWIDTH_REG_24_, DATAWIDTH_REG_25_,
    DATAWIDTH_REG_26_, DATAWIDTH_REG_27_, DATAWIDTH_REG_28_,
    DATAWIDTH_REG_29_, DATAWIDTH_REG_30_, DATAWIDTH_REG_31_, STATE2_REG_3_,
    STATE2_REG_2_, STATE2_REG_1_, STATE2_REG_0_, INSTQUEUE_REG_15__7_,
    INSTQUEUE_REG_15__6_, INSTQUEUE_REG_15__5_, INSTQUEUE_REG_15__4_,
    INSTQUEUE_REG_15__3_, INSTQUEUE_REG_15__2_, INSTQUEUE_REG_15__1_,
    INSTQUEUE_REG_15__0_, INSTQUEUE_REG_14__7_, INSTQUEUE_REG_14__6_,
    INSTQUEUE_REG_14__5_, INSTQUEUE_REG_14__4_, INSTQUEUE_REG_14__3_,
    INSTQUEUE_REG_14__2_, INSTQUEUE_REG_14__1_, INSTQUEUE_REG_14__0_,
    INSTQUEUE_REG_13__7_, INSTQUEUE_REG_13__6_, INSTQUEUE_REG_13__5_,
    INSTQUEUE_REG_13__4_, INSTQUEUE_REG_13__3_, INSTQUEUE_REG_13__2_,
    INSTQUEUE_REG_13__1_, INSTQUEUE_REG_13__0_, INSTQUEUE_REG_12__7_,
    INSTQUEUE_REG_12__6_, INSTQUEUE_REG_12__5_, INSTQUEUE_REG_12__4_,
    INSTQUEUE_REG_12__3_, INSTQUEUE_REG_12__2_, INSTQUEUE_REG_12__1_,
    INSTQUEUE_REG_12__0_, INSTQUEUE_REG_11__7_, INSTQUEUE_REG_11__6_,
    INSTQUEUE_REG_11__5_, INSTQUEUE_REG_11__4_, INSTQUEUE_REG_11__3_,
    INSTQUEUE_REG_11__2_, INSTQUEUE_REG_11__1_, INSTQUEUE_REG_11__0_,
    INSTQUEUE_REG_10__7_, INSTQUEUE_REG_10__6_, INSTQUEUE_REG_10__5_,
    INSTQUEUE_REG_10__4_, INSTQUEUE_REG_10__3_, INSTQUEUE_REG_10__2_,
    INSTQUEUE_REG_10__1_, INSTQUEUE_REG_10__0_, INSTQUEUE_REG_9__7_,
    INSTQUEUE_REG_9__6_, INSTQUEUE_REG_9__5_, INSTQUEUE_REG_9__4_,
    INSTQUEUE_REG_9__3_, INSTQUEUE_REG_9__2_, INSTQUEUE_REG_9__1_,
    INSTQUEUE_REG_9__0_, INSTQUEUE_REG_8__7_, INSTQUEUE_REG_8__6_,
    INSTQUEUE_REG_8__5_, INSTQUEUE_REG_8__4_, INSTQUEUE_REG_8__3_,
    INSTQUEUE_REG_8__2_, INSTQUEUE_REG_8__1_, INSTQUEUE_REG_8__0_,
    INSTQUEUE_REG_7__7_, INSTQUEUE_REG_7__6_, INSTQUEUE_REG_7__5_,
    INSTQUEUE_REG_7__4_, INSTQUEUE_REG_7__3_, INSTQUEUE_REG_7__2_,
    INSTQUEUE_REG_7__1_, INSTQUEUE_REG_7__0_, INSTQUEUE_REG_6__7_,
    INSTQUEUE_REG_6__6_, INSTQUEUE_REG_6__5_, INSTQUEUE_REG_6__4_,
    INSTQUEUE_REG_6__3_, INSTQUEUE_REG_6__2_, INSTQUEUE_REG_6__1_,
    INSTQUEUE_REG_6__0_, INSTQUEUE_REG_5__7_, INSTQUEUE_REG_5__6_,
    INSTQUEUE_REG_5__5_, INSTQUEUE_REG_5__4_, INSTQUEUE_REG_5__3_,
    INSTQUEUE_REG_5__2_, INSTQUEUE_REG_5__1_, INSTQUEUE_REG_5__0_,
    INSTQUEUE_REG_4__7_, INSTQUEUE_REG_4__6_, INSTQUEUE_REG_4__5_,
    INSTQUEUE_REG_4__4_, INSTQUEUE_REG_4__3_, INSTQUEUE_REG_4__2_,
    INSTQUEUE_REG_4__1_, INSTQUEUE_REG_4__0_, INSTQUEUE_REG_3__7_,
    INSTQUEUE_REG_3__6_, INSTQUEUE_REG_3__5_, INSTQUEUE_REG_3__4_,
    INSTQUEUE_REG_3__3_, INSTQUEUE_REG_3__2_, INSTQUEUE_REG_3__1_,
    INSTQUEUE_REG_3__0_, INSTQUEUE_REG_2__7_, INSTQUEUE_REG_2__6_,
    INSTQUEUE_REG_2__5_, INSTQUEUE_REG_2__4_, INSTQUEUE_REG_2__3_,
    INSTQUEUE_REG_2__2_, INSTQUEUE_REG_2__1_, INSTQUEUE_REG_2__0_,
    INSTQUEUE_REG_1__7_, INSTQUEUE_REG_1__6_, INSTQUEUE_REG_1__5_,
    INSTQUEUE_REG_1__4_, INSTQUEUE_REG_1__3_, INSTQUEUE_REG_1__2_,
    INSTQUEUE_REG_1__1_, INSTQUEUE_REG_1__0_, INSTQUEUE_REG_0__7_,
    INSTQUEUE_REG_0__6_, INSTQUEUE_REG_0__5_, INSTQUEUE_REG_0__4_,
    INSTQUEUE_REG_0__3_, INSTQUEUE_REG_0__2_, INSTQUEUE_REG_0__1_,
    INSTQUEUE_REG_0__0_, INSTQUEUERD_ADDR_REG_4_, INSTQUEUERD_ADDR_REG_3_,
    INSTQUEUERD_ADDR_REG_2_, INSTQUEUERD_ADDR_REG_1_,
    INSTQUEUERD_ADDR_REG_0_, INSTQUEUEWR_ADDR_REG_4_,
    INSTQUEUEWR_ADDR_REG_3_, INSTQUEUEWR_ADDR_REG_2_,
    INSTQUEUEWR_ADDR_REG_1_, INSTQUEUEWR_ADDR_REG_0_,
    INSTADDRPOINTER_REG_0_, INSTADDRPOINTER_REG_1_, INSTADDRPOINTER_REG_2_,
    INSTADDRPOINTER_REG_3_, INSTADDRPOINTER_REG_4_, INSTADDRPOINTER_REG_5_,
    INSTADDRPOINTER_REG_6_, INSTADDRPOINTER_REG_7_, INSTADDRPOINTER_REG_8_,
    INSTADDRPOINTER_REG_9_, INSTADDRPOINTER_REG_10_,
    INSTADDRPOINTER_REG_11_, INSTADDRPOINTER_REG_12_,
    INSTADDRPOINTER_REG_13_, INSTADDRPOINTER_REG_14_,
    INSTADDRPOINTER_REG_15_, INSTADDRPOINTER_REG_16_,
    INSTADDRPOINTER_REG_17_, INSTADDRPOINTER_REG_18_,
    INSTADDRPOINTER_REG_19_, INSTADDRPOINTER_REG_20_,
    INSTADDRPOINTER_REG_21_, INSTADDRPOINTER_REG_22_,
    INSTADDRPOINTER_REG_23_, INSTADDRPOINTER_REG_24_,
    INSTADDRPOINTER_REG_25_, INSTADDRPOINTER_REG_26_,
    INSTADDRPOINTER_REG_27_, INSTADDRPOINTER_REG_28_,
    INSTADDRPOINTER_REG_29_, INSTADDRPOINTER_REG_30_,
    INSTADDRPOINTER_REG_31_, PHYADDRPOINTER_REG_0_, PHYADDRPOINTER_REG_1_,
    PHYADDRPOINTER_REG_2_, PHYADDRPOINTER_REG_3_, PHYADDRPOINTER_REG_4_,
    PHYADDRPOINTER_REG_5_, PHYADDRPOINTER_REG_6_, PHYADDRPOINTER_REG_7_,
    PHYADDRPOINTER_REG_8_, PHYADDRPOINTER_REG_9_, PHYADDRPOINTER_REG_10_,
    PHYADDRPOINTER_REG_11_, PHYADDRPOINTER_REG_12_, PHYADDRPOINTER_REG_13_,
    PHYADDRPOINTER_REG_14_, PHYADDRPOINTER_REG_15_, PHYADDRPOINTER_REG_16_,
    PHYADDRPOINTER_REG_17_, PHYADDRPOINTER_REG_18_, PHYADDRPOINTER_REG_19_,
    PHYADDRPOINTER_REG_20_, PHYADDRPOINTER_REG_21_, PHYADDRPOINTER_REG_22_,
    PHYADDRPOINTER_REG_23_, PHYADDRPOINTER_REG_24_, PHYADDRPOINTER_REG_25_,
    PHYADDRPOINTER_REG_26_, PHYADDRPOINTER_REG_27_, PHYADDRPOINTER_REG_28_,
    PHYADDRPOINTER_REG_29_, PHYADDRPOINTER_REG_30_, PHYADDRPOINTER_REG_31_,
    LWORD_REG_15_, LWORD_REG_14_, LWORD_REG_13_, LWORD_REG_12_,
    LWORD_REG_11_, LWORD_REG_10_, LWORD_REG_9_, LWORD_REG_8_, LWORD_REG_7_,
    LWORD_REG_6_, LWORD_REG_5_, LWORD_REG_4_, LWORD_REG_3_, LWORD_REG_2_,
    LWORD_REG_1_, LWORD_REG_0_, UWORD_REG_14_, UWORD_REG_13_,
    UWORD_REG_12_, UWORD_REG_11_, UWORD_REG_10_, UWORD_REG_9_,
    UWORD_REG_8_, UWORD_REG_7_, UWORD_REG_6_, UWORD_REG_5_, UWORD_REG_4_,
    UWORD_REG_3_, UWORD_REG_2_, UWORD_REG_1_, UWORD_REG_0_, DATAO_REG_0_,
    DATAO_REG_1_, DATAO_REG_2_, DATAO_REG_3_, DATAO_REG_4_, DATAO_REG_5_,
    DATAO_REG_6_, DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_, DATAO_REG_10_,
    DATAO_REG_11_, DATAO_REG_12_, DATAO_REG_13_, DATAO_REG_14_,
    DATAO_REG_15_, DATAO_REG_16_, DATAO_REG_17_, DATAO_REG_18_,
    DATAO_REG_19_, DATAO_REG_20_, DATAO_REG_21_, DATAO_REG_22_,
    DATAO_REG_23_, DATAO_REG_24_, DATAO_REG_25_, DATAO_REG_26_,
    DATAO_REG_27_, DATAO_REG_28_, DATAO_REG_29_, DATAO_REG_30_,
    DATAO_REG_31_, EAX_REG_0_, EAX_REG_1_, EAX_REG_2_, EAX_REG_3_,
    EAX_REG_4_, EAX_REG_5_, EAX_REG_6_, EAX_REG_7_, EAX_REG_8_, EAX_REG_9_,
    EAX_REG_10_, EAX_REG_11_, EAX_REG_12_, EAX_REG_13_, EAX_REG_14_,
    EAX_REG_15_, EAX_REG_16_, EAX_REG_17_, EAX_REG_18_, EAX_REG_19_,
    EAX_REG_20_, EAX_REG_21_, EAX_REG_22_, EAX_REG_23_, EAX_REG_24_,
    EAX_REG_25_, EAX_REG_26_, EAX_REG_27_, EAX_REG_28_, EAX_REG_29_,
    EAX_REG_30_, EAX_REG_31_, EBX_REG_0_, EBX_REG_1_, EBX_REG_2_,
    EBX_REG_3_, EBX_REG_4_, EBX_REG_5_, EBX_REG_6_, EBX_REG_7_, EBX_REG_8_,
    EBX_REG_9_, EBX_REG_10_, EBX_REG_11_, EBX_REG_12_, EBX_REG_13_,
    EBX_REG_14_, EBX_REG_15_, EBX_REG_16_, EBX_REG_17_, EBX_REG_18_,
    EBX_REG_19_, EBX_REG_20_, EBX_REG_21_, EBX_REG_22_, EBX_REG_23_,
    EBX_REG_24_, EBX_REG_25_, EBX_REG_26_, EBX_REG_27_, EBX_REG_28_,
    EBX_REG_29_, EBX_REG_30_, EBX_REG_31_, REIP_REG_0_, REIP_REG_1_,
    REIP_REG_2_, REIP_REG_3_, REIP_REG_4_, REIP_REG_5_, REIP_REG_6_,
    REIP_REG_7_, REIP_REG_8_, REIP_REG_9_, REIP_REG_10_, REIP_REG_11_,
    REIP_REG_12_, REIP_REG_13_, REIP_REG_14_, REIP_REG_15_, REIP_REG_16_,
    REIP_REG_17_, REIP_REG_18_, REIP_REG_19_, REIP_REG_20_, REIP_REG_21_,
    REIP_REG_22_, REIP_REG_23_, REIP_REG_24_, REIP_REG_25_, REIP_REG_26_,
    REIP_REG_27_, REIP_REG_28_, REIP_REG_29_, REIP_REG_30_, REIP_REG_31_,
    BYTEENABLE_REG_3_, BYTEENABLE_REG_2_, BYTEENABLE_REG_1_,
    BYTEENABLE_REG_0_, W_R_N_REG, FLUSH_REG, MORE_REG, STATEBS16_REG,
    REQUESTPENDING_REG, D_C_N_REG, M_IO_N_REG, CODEFETCH_REG, ADS_N_REG,
    READREQUEST_REG, MEMORYFETCH_REG;
  wire n1454, n1455_1, n1456, n1458, n1459, n1461, n1462, n1464, n1465_1,
    n1467, n1468, n1469, n1470_1, n1471, n1472, n1474, n1475_1, n1476,
    n1477, n1479, n1480_1, n1481, n1482, n1484, n1485_1, n1486, n1487,
    n1489, n1490_1, n1491, n1492, n1494, n1495_1, n1496, n1497, n1499,
    n1500_1, n1501, n1502, n1504, n1505_1, n1506, n1507, n1509, n1510_1,
    n1511, n1512, n1514, n1515_1, n1516, n1517, n1519, n1520_1, n1521,
    n1522, n1524, n1525_1, n1526, n1527, n1529, n1530_1, n1531, n1532,
    n1534, n1535_1, n1536, n1537, n1539, n1540_1, n1541, n1542, n1544,
    n1545_1, n1546, n1547, n1549, n1550_1, n1551, n1552, n1554, n1555_1,
    n1556, n1557, n1559, n1560_1, n1561, n1562, n1564, n1565_1, n1566,
    n1567, n1569, n1570_1, n1571, n1572, n1574, n1575_1, n1576, n1577,
    n1579, n1580_1, n1581, n1582, n1584, n1585_1, n1586, n1587, n1589,
    n1590_1, n1591, n1592, n1594, n1595_1, n1596, n1597, n1599, n1600_1,
    n1601, n1602, n1604, n1605_1, n1606, n1607, n1609, n1610_1, n1611,
    n1612, n1614, n1615_1, n1616, n1617, n1619, n1620_1, n1621, n1622,
    n1623, n1624, n1625_1, n1626, n1627, n1628, n1629, n1630_1, n1631,
    n1632, n1633, n1634, n1635_1, n1636, n1637, n1638, n1639, n1640_1,
    n1641, n1643, n1644, n1645_1, n1646, n1647, n1648, n1649, n1650_1,
    n1651, n1652, n1653, n1654, n1655_1, n1657, n1658, n1659, n1660_1,
    n1661, n1662, n1663, n1664, n1665_1, n1667, n1668, n1669, n1670_1,
    n1671, n1672, n1674, n1675_1, n1707, n1708, n1709, n1710_1, n1711,
    n1712, n1713, n1714_1, n1715, n1716, n1717, n1718_1, n1719, n1720,
    n1721, n1722_1, n1723, n1724, n1725, n1726_1, n1727, n1728, n1729,
    n1730_1, n1731, n1732, n1733, n1734_1, n1735, n1736, n1737, n1738_1,
    n1739, n1740, n1741, n1742_1, n1743, n1744, n1745, n1746_1, n1747,
    n1748, n1749, n1750_1, n1751, n1752, n1753, n1754_1, n1755, n1756,
    n1757, n1758_1, n1759, n1760, n1761, n1762_1, n1763, n1764, n1765,
    n1766_1, n1767, n1768, n1769, n1770_1, n1771, n1772, n1773, n1774_1,
    n1775, n1776, n1777, n1778_1, n1779, n1780, n1781, n1782_1, n1783,
    n1784, n1785, n1786_1, n1787, n1788, n1789, n1790_1, n1791, n1792,
    n1793, n1794_1, n1795, n1796, n1797, n1798_1, n1799, n1800, n1801,
    n1802_1, n1803, n1804, n1805, n1806_1, n1807, n1808, n1809, n1810_1,
    n1811, n1812, n1813, n1814_1, n1815, n1816, n1817, n1818_1, n1819,
    n1820, n1821, n1822_1, n1823, n1824, n1825, n1826_1, n1827, n1828,
    n1829, n1830_1, n1831, n1832, n1833, n1834_1, n1835, n1836, n1837,
    n1838_1, n1839, n1840, n1841, n1842, n1843_1, n1844, n1845, n1846,
    n1847, n1848_1, n1849, n1850, n1851, n1852, n1853_1, n1854, n1855,
    n1856, n1857, n1858_1, n1859, n1860, n1861, n1862, n1863_1, n1864,
    n1865, n1866, n1867, n1868_1, n1869, n1870, n1871, n1872, n1873_1,
    n1874, n1875, n1876, n1877, n1878_1, n1879, n1880, n1881, n1882,
    n1883_1, n1884, n1885, n1886, n1887, n1888_1, n1889, n1890, n1891,
    n1892, n1893_1, n1894, n1895, n1896, n1897, n1898_1, n1899, n1900,
    n1901, n1902, n1903_1, n1904, n1905, n1906, n1907, n1908_1, n1909,
    n1910, n1911, n1912, n1913_1, n1914, n1915, n1916, n1917, n1918_1,
    n1919, n1920, n1921, n1922, n1923_1, n1924, n1925, n1926, n1927,
    n1928_1, n1929, n1930, n1931, n1932, n1933_1, n1934, n1935, n1936,
    n1937, n1938_1, n1939, n1940, n1941, n1942, n1943_1, n1944, n1945,
    n1946, n1947, n1948_1, n1949, n1950, n1951, n1952, n1953_1, n1954,
    n1955, n1956, n1957, n1958_1, n1959, n1960, n1961, n1962, n1963_1,
    n1964, n1965, n1966, n1967, n1968_1, n1969, n1970, n1971, n1972,
    n1973_1, n1974, n1975, n1976, n1977, n1978_1, n1979, n1980, n1981,
    n1982, n1983_1, n1984, n1985, n1986, n1987, n1988_1, n1989, n1990,
    n1991, n1992, n1993_1, n1994, n1995, n1996, n1997, n1998_1, n1999,
    n2000, n2001, n2002, n2003_1, n2004, n2005, n2006, n2007, n2008_1,
    n2009, n2010, n2011, n2012, n2013_1, n2014, n2015, n2016, n2017,
    n2018_1, n2019, n2020, n2021, n2022, n2023_1, n2024, n2025, n2026,
    n2027, n2028_1, n2029, n2030, n2031, n2032, n2033_1, n2034, n2035,
    n2036, n2037, n2038_1, n2039, n2040, n2041, n2042, n2043_1, n2044,
    n2045, n2046, n2047, n2048_1, n2049, n2050, n2051, n2052, n2053_1,
    n2054, n2055, n2056, n2057, n2058_1, n2059, n2060, n2061, n2062,
    n2063_1, n2064, n2065, n2066, n2067, n2068_1, n2069, n2070, n2071,
    n2072, n2073_1, n2074, n2075, n2076, n2077, n2078_1, n2079, n2080,
    n2081, n2082, n2083_1, n2084, n2085, n2086, n2087, n2088_1, n2089,
    n2090, n2091, n2092, n2093_1, n2094, n2095, n2096, n2097, n2098_1,
    n2099, n2100, n2101, n2102, n2103_1, n2104, n2105, n2106, n2107,
    n2108_1, n2109, n2110, n2111, n2112, n2113_1, n2114, n2115, n2116,
    n2117, n2118_1, n2119, n2120, n2121, n2122, n2123_1, n2124, n2125,
    n2126, n2127, n2128_1, n2129, n2130, n2131, n2132, n2133_1, n2134,
    n2135, n2136, n2137, n2138_1, n2139, n2140, n2141, n2142, n2143_1,
    n2144, n2145, n2146, n2147, n2148_1, n2149, n2150, n2151, n2152,
    n2153_1, n2154, n2155, n2156, n2157, n2158_1, n2159, n2160, n2161,
    n2162, n2163_1, n2164, n2165, n2166, n2167, n2168_1, n2169, n2170,
    n2171, n2172, n2173_1, n2174, n2175, n2176, n2177, n2178_1, n2179,
    n2180, n2181, n2182, n2183_1, n2184, n2185, n2186, n2187, n2188_1,
    n2189, n2190, n2191, n2192, n2193_1, n2194, n2195, n2196, n2197,
    n2198_1, n2199, n2200, n2201, n2202, n2203_1, n2204, n2205, n2206,
    n2207, n2208_1, n2209, n2210, n2211, n2212, n2213_1, n2214, n2215,
    n2216, n2217, n2218_1, n2219, n2220, n2221, n2222, n2223_1, n2224,
    n2225, n2226, n2227, n2228_1, n2229, n2230, n2231, n2232, n2233_1,
    n2234, n2235, n2236, n2237, n2238_1, n2239, n2240, n2241, n2242,
    n2243_1, n2244, n2245, n2246, n2247, n2248_1, n2249, n2250, n2251,
    n2252, n2253_1, n2254, n2255, n2256, n2257, n2258_1, n2259, n2260,
    n2261, n2262, n2263_1, n2264, n2265, n2266, n2267, n2268_1, n2269,
    n2270, n2271, n2272, n2273_1, n2274, n2275, n2276, n2277, n2278_1,
    n2279, n2280, n2281, n2282, n2283_1, n2284, n2285, n2286, n2287,
    n2288_1, n2289, n2290, n2291, n2292, n2293_1, n2294, n2295, n2296,
    n2297, n2298_1, n2299, n2300, n2301, n2302, n2303_1, n2304, n2305,
    n2306, n2307, n2308_1, n2309, n2310, n2311, n2312, n2313_1, n2314,
    n2315, n2316, n2317, n2318_1, n2319, n2320, n2321, n2322, n2323_1,
    n2324, n2325, n2326, n2327, n2328_1, n2329, n2330, n2331, n2332,
    n2333_1, n2334, n2335, n2336, n2337, n2338_1, n2339, n2340, n2341,
    n2342_1, n2343, n2344, n2345, n2346, n2347_1, n2348, n2349, n2350,
    n2351, n2352_1, n2353, n2354, n2355, n2356, n2357_1, n2358, n2359,
    n2360, n2361, n2362_1, n2363, n2364, n2365, n2366_1, n2367, n2368,
    n2369, n2370_1, n2371, n2372, n2373, n2374, n2375_1, n2376, n2377,
    n2378, n2379_1, n2380, n2381, n2382, n2383, n2384_1, n2385, n2386,
    n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
    n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
    n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
    n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
    n3552, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3701, n3702, n3703, n3704, n3705, n3706,
    n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4063, n4064, n4065, n4066, n4067,
    n4068, n4069, n4070, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4119, n4120, n4121,
    n4122, n4123, n4124, n4125, n4126, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4550, n4551, n4552, n4553, n4554, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4580, n4581, n4582, n4583,
    n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4617,
    n4618, n4619, n4620, n4621, n4622, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
    n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
    n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5233, n5234, n5235, n5236,
    n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
    n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
    n5802, n5803, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
    n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
    n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
    n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
    n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
    n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
    n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6591, n6592, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
    n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
    n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
    n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
    n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
    n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
    n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
    n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
    n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
    n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
    n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
    n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
    n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
    n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
    n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
    n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
    n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
    n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
    n8076, n8077, n8078, n8079, n8080, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
    n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8484, n8485, n8486, n8487, n8488, n8490, n8491, n8492, n8493, n8494,
    n8496, n8497, n8498, n8499, n8500, n8502, n8503, n8504, n8505, n8506,
    n8508, n8509, n8510, n8511, n8512, n8514, n8515, n8516, n8517, n8518,
    n8520, n8521, n8522, n8523, n8524, n8526, n8527, n8528, n8529, n8530,
    n8532, n8533, n8534, n8535, n8536, n8538, n8539, n8540, n8541, n8542,
    n8544, n8545, n8546, n8547, n8548, n8550, n8551, n8552, n8553, n8554,
    n8556, n8557, n8558, n8559, n8560, n8562, n8563, n8564, n8565, n8566,
    n8568, n8569, n8570, n8571, n8572, n8574, n8575, n8576, n8577, n8579,
    n8580, n8581, n8582, n8584, n8585, n8586, n8587, n8589, n8590, n8591,
    n8592, n8594, n8595, n8596, n8597, n8599, n8600, n8601, n8602, n8604,
    n8605, n8606, n8607, n8609, n8610, n8611, n8612, n8614, n8615, n8616,
    n8617, n8619, n8620, n8621, n8622, n8624, n8625, n8626, n8627, n8629,
    n8630, n8631, n8632, n8634, n8635, n8636, n8637, n8639, n8640, n8641,
    n8642, n8644, n8645, n8646, n8647, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8663, n8664,
    n8665, n8666, n8668, n8669, n8670, n8671, n8673, n8674, n8675, n8676,
    n8678, n8679, n8680, n8681, n8683, n8684, n8685, n8686, n8688, n8689,
    n8690, n8691, n8693, n8694, n8695, n8696, n8698, n8699, n8700, n8701,
    n8703, n8704, n8705, n8706, n8708, n8709, n8710, n8711, n8713, n8714,
    n8715, n8716, n8718, n8719, n8720, n8721, n8723, n8724, n8725, n8726,
    n8728, n8729, n8730, n8731, n8733, n8734, n8735, n8736, n8738, n8739,
    n8740, n8741, n8742, n8744, n8745, n8746, n8747, n8749, n8750, n8751,
    n8752, n8754, n8755, n8756, n8757, n8759, n8760, n8761, n8762, n8764,
    n8765, n8766, n8767, n8769, n8770, n8771, n8772, n8774, n8775, n8776,
    n8777, n8779, n8780, n8781, n8782, n8784, n8785, n8786, n8787, n8789,
    n8790, n8791, n8792, n8794, n8795, n8796, n8797, n8799, n8800, n8801,
    n8802, n8804, n8805, n8806, n8807, n8809, n8810, n8811, n8812, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8836,
    n8837, n8838, n8839, n8841, n8842, n8843, n8844, n8846, n8847, n8848,
    n8849, n8851, n8852, n8853, n8854, n8856, n8857, n8858, n8859, n8861,
    n8862, n8863, n8864, n8866, n8867, n8868, n8869, n8871, n8872, n8873,
    n8874, n8876, n8877, n8878, n8879, n8881, n8882, n8883, n8884, n8886,
    n8887, n8888, n8889, n8891, n8892, n8893, n8894, n8896, n8897, n8898,
    n8899, n8901, n8902, n8903, n8904, n8906, n8907, n8908, n8909, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8921, n8922,
    n8923, n8924, n8925, n8926, n8928, n8929, n8930, n8931, n8932, n8933,
    n8935, n8936, n8937, n8938, n8939, n8940, n8942, n8943, n8944, n8945,
    n8946, n8947, n8949, n8950, n8951, n8952, n8953, n8954, n8956, n8957,
    n8958, n8959, n8960, n8961, n8963, n8964, n8965, n8966, n8967, n8968,
    n8970, n8971, n8972, n8973, n8974, n8975, n8977, n8978, n8979, n8980,
    n8981, n8982, n8984, n8985, n8986, n8987, n8988, n8989, n8991, n8992,
    n8993, n8994, n8995, n8996, n8998, n8999, n9000, n9001, n9002, n9003,
    n9005, n9006, n9007, n9008, n9009, n9010, n9012, n9013, n9014, n9015,
    n9016, n9017, n9019, n9020, n9021, n9022, n9023, n9025, n9026, n9027,
    n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
    n9039, n9040, n9041, n9042, n9044, n9045, n9046, n9047, n9049, n9050,
    n9051, n9052, n9054, n9055, n9056, n9057, n9059, n9060, n9061, n9062,
    n9064, n9065, n9066, n9067, n9069, n9070, n9071, n9072, n9074, n9075,
    n9076, n9077, n9079, n9080, n9081, n9082, n9084, n9085, n9086, n9087,
    n9089, n9090, n9091, n9092, n9094, n9095, n9096, n9097, n9099, n9100,
    n9101, n9102, n9104, n9105, n9106, n9107, n9109, n9110, n9111, n9112,
    n9114, n9115, n9116, n9117, n9119, n9120, n9121, n9122, n9124, n9125,
    n9126, n9127, n9129, n9130, n9131, n9132, n9134, n9135, n9136, n9137,
    n9139, n9140, n9141, n9142, n9144, n9145, n9146, n9147, n9149, n9150,
    n9151, n9152, n9154, n9155, n9156, n9157, n9159, n9160, n9161, n9162,
    n9164, n9165, n9166, n9167, n9169, n9170, n9171, n9172, n9174, n9175,
    n9176, n9177, n9179, n9180, n9181, n9182, n9184, n9185, n9186, n9187,
    n9189, n9190, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9479, n9480, n9481, n9482, n9483,
    n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
    n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9621,
    n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
    n9653, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
    n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
    n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9830, n9831, n9832,
    n9833, n9834, n9835, n9836, n9837, n9839, n9840, n9841, n9843, n9844,
    n9845, n9847, n9848, n9850, n9851, n9853, n9854, n9856, n9857, n9858,
    n9859, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
    n9870, n9871, n9872, n9873, n9874, n9875, n9877, n9878, n9879, n9881,
    n9882, n9884, n9885, n9886, n9888, n9890, n9891, n9892, n9893, n9894,
    n9896, n9897, n9898, n9899, n9900, n214, n218, n222, n226, n230, n234,
    n238, n242, n246, n250, n254, n258, n262, n266, n270, n274, n278, n282,
    n286, n290, n294, n298, n302, n306, n310, n314, n318, n322, n326, n330,
    n334, n338, n342, n346, n350, n355, n360, n365, n370, n375, n380, n385,
    n390, n395, n400, n405, n410, n415, n420, n425, n430, n435, n440, n445,
    n450, n455, n460, n465, n470, n475, n480, n485, n490, n495, n500, n505,
    n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560, n565,
    n570, n575, n580, n585, n590, n595, n600, n605, n610, n615, n620, n625,
    n630, n635, n640, n645, n650, n655, n660, n665, n670, n675, n680, n685,
    n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740, n745,
    n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800, n805,
    n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860, n865,
    n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920, n925,
    n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980, n985,
    n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035,
    n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085,
    n1090, n1095, n1100, n1105, n1110, n1115, n1120, n1125, n1130, n1135,
    n1140, n1145, n1150, n1155, n1160, n1165, n1170, n1175, n1180, n1185,
    n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235,
    n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275, n1280, n1285,
    n1290, n1295, n1300, n1305, n1310, n1315, n1320, n1325, n1330, n1335,
    n1340, n1345, n1350, n1355, n1360, n1365, n1370, n1375, n1380, n1385,
    n1390, n1395, n1400, n1405, n1410, n1415, n1420, n1425, n1430, n1435,
    n1440, n1445, n1450, n1455, n1460, n1465, n1470, n1475, n1480, n1485,
    n1490, n1495, n1500, n1505, n1510, n1515, n1520, n1525, n1530, n1535,
    n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575, n1580, n1585,
    n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635,
    n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685,
    n1690, n1695, n1700, n1705, n1710, n1714, n1718, n1722, n1726, n1730,
    n1734, n1738, n1742, n1746, n1750, n1754, n1758, n1762, n1766, n1770,
    n1774, n1778, n1782, n1786, n1790, n1794, n1798, n1802, n1806, n1810,
    n1814, n1818, n1822, n1826, n1830, n1834, n1838, n1843, n1848, n1853,
    n1858, n1863, n1868, n1873, n1878, n1883, n1888, n1893, n1898, n1903,
    n1908, n1913, n1918, n1923, n1928, n1933, n1938, n1943, n1948, n1953,
    n1958, n1963, n1968, n1973, n1978, n1983, n1988, n1993, n1998, n2003,
    n2008, n2013, n2018, n2023, n2028, n2033, n2038, n2043, n2048, n2053,
    n2058, n2063, n2068, n2073, n2078, n2083, n2088, n2093, n2098, n2103,
    n2108, n2113, n2118, n2123, n2128, n2133, n2138, n2143, n2148, n2153,
    n2158, n2163, n2168, n2173, n2178, n2183, n2188, n2193, n2198, n2203,
    n2208, n2213, n2218, n2223, n2228, n2233, n2238, n2243, n2248, n2253,
    n2258, n2263, n2268, n2273, n2278, n2283, n2288, n2293, n2298, n2303,
    n2308, n2313, n2318, n2323, n2328, n2333, n2338, n2342, n2347, n2352,
    n2357, n2362, n2366, n2370, n2375, n2379, n2384;
  assign n1454 = STATE_REG_1_ & ~STATE_REG_0_;
  assign n1455_1 = BYTEENABLE_REG_3_ & n1454;
  assign n1456 = BE_N_REG_3_ & ~n1454;
  assign n214 = n1455_1 | n1456;
  assign n1458 = BYTEENABLE_REG_2_ & n1454;
  assign n1459 = BE_N_REG_2_ & ~n1454;
  assign n218 = n1458 | n1459;
  assign n1461 = BYTEENABLE_REG_1_ & n1454;
  assign n1462 = BE_N_REG_1_ & ~n1454;
  assign n222 = n1461 | n1462;
  assign n1464 = BYTEENABLE_REG_0_ & n1454;
  assign n1465_1 = BE_N_REG_0_ & ~n1454;
  assign n226 = n1464 | n1465_1;
  assign n1467 = STATE_REG_2_ & n1454;
  assign n1468 = REIP_REG_30_ & n1467;
  assign n1469 = ~STATE_REG_2_ & n1454;
  assign n1470_1 = REIP_REG_31_ & n1469;
  assign n1471 = ADDRESS_REG_29_ & ~n1454;
  assign n1472 = ~n1468 & ~n1470_1;
  assign n230 = n1471 | ~n1472;
  assign n1474 = REIP_REG_29_ & n1467;
  assign n1475_1 = REIP_REG_30_ & n1469;
  assign n1476 = ADDRESS_REG_28_ & ~n1454;
  assign n1477 = ~n1474 & ~n1475_1;
  assign n234 = n1476 | ~n1477;
  assign n1479 = REIP_REG_28_ & n1467;
  assign n1480_1 = REIP_REG_29_ & n1469;
  assign n1481 = ADDRESS_REG_27_ & ~n1454;
  assign n1482 = ~n1479 & ~n1480_1;
  assign n238 = n1481 | ~n1482;
  assign n1484 = REIP_REG_27_ & n1467;
  assign n1485_1 = REIP_REG_28_ & n1469;
  assign n1486 = ADDRESS_REG_26_ & ~n1454;
  assign n1487 = ~n1484 & ~n1485_1;
  assign n242 = n1486 | ~n1487;
  assign n1489 = REIP_REG_26_ & n1467;
  assign n1490_1 = REIP_REG_27_ & n1469;
  assign n1491 = ADDRESS_REG_25_ & ~n1454;
  assign n1492 = ~n1489 & ~n1490_1;
  assign n246 = n1491 | ~n1492;
  assign n1494 = REIP_REG_25_ & n1467;
  assign n1495_1 = REIP_REG_26_ & n1469;
  assign n1496 = ADDRESS_REG_24_ & ~n1454;
  assign n1497 = ~n1494 & ~n1495_1;
  assign n250 = n1496 | ~n1497;
  assign n1499 = REIP_REG_24_ & n1467;
  assign n1500_1 = REIP_REG_25_ & n1469;
  assign n1501 = ADDRESS_REG_23_ & ~n1454;
  assign n1502 = ~n1499 & ~n1500_1;
  assign n254 = n1501 | ~n1502;
  assign n1504 = REIP_REG_23_ & n1467;
  assign n1505_1 = REIP_REG_24_ & n1469;
  assign n1506 = ADDRESS_REG_22_ & ~n1454;
  assign n1507 = ~n1504 & ~n1505_1;
  assign n258 = n1506 | ~n1507;
  assign n1509 = REIP_REG_22_ & n1467;
  assign n1510_1 = REIP_REG_23_ & n1469;
  assign n1511 = ADDRESS_REG_21_ & ~n1454;
  assign n1512 = ~n1509 & ~n1510_1;
  assign n262 = n1511 | ~n1512;
  assign n1514 = REIP_REG_21_ & n1467;
  assign n1515_1 = REIP_REG_22_ & n1469;
  assign n1516 = ADDRESS_REG_20_ & ~n1454;
  assign n1517 = ~n1514 & ~n1515_1;
  assign n266 = n1516 | ~n1517;
  assign n1519 = REIP_REG_20_ & n1467;
  assign n1520_1 = REIP_REG_21_ & n1469;
  assign n1521 = ADDRESS_REG_19_ & ~n1454;
  assign n1522 = ~n1519 & ~n1520_1;
  assign n270 = n1521 | ~n1522;
  assign n1524 = REIP_REG_19_ & n1467;
  assign n1525_1 = REIP_REG_20_ & n1469;
  assign n1526 = ADDRESS_REG_18_ & ~n1454;
  assign n1527 = ~n1524 & ~n1525_1;
  assign n274 = n1526 | ~n1527;
  assign n1529 = REIP_REG_18_ & n1467;
  assign n1530_1 = REIP_REG_19_ & n1469;
  assign n1531 = ADDRESS_REG_17_ & ~n1454;
  assign n1532 = ~n1529 & ~n1530_1;
  assign n278 = n1531 | ~n1532;
  assign n1534 = REIP_REG_17_ & n1467;
  assign n1535_1 = REIP_REG_18_ & n1469;
  assign n1536 = ADDRESS_REG_16_ & ~n1454;
  assign n1537 = ~n1534 & ~n1535_1;
  assign n282 = n1536 | ~n1537;
  assign n1539 = REIP_REG_16_ & n1467;
  assign n1540_1 = REIP_REG_17_ & n1469;
  assign n1541 = ADDRESS_REG_15_ & ~n1454;
  assign n1542 = ~n1539 & ~n1540_1;
  assign n286 = n1541 | ~n1542;
  assign n1544 = REIP_REG_15_ & n1467;
  assign n1545_1 = REIP_REG_16_ & n1469;
  assign n1546 = ADDRESS_REG_14_ & ~n1454;
  assign n1547 = ~n1544 & ~n1545_1;
  assign n290 = n1546 | ~n1547;
  assign n1549 = REIP_REG_14_ & n1467;
  assign n1550_1 = REIP_REG_15_ & n1469;
  assign n1551 = ADDRESS_REG_13_ & ~n1454;
  assign n1552 = ~n1549 & ~n1550_1;
  assign n294 = n1551 | ~n1552;
  assign n1554 = REIP_REG_13_ & n1467;
  assign n1555_1 = REIP_REG_14_ & n1469;
  assign n1556 = ADDRESS_REG_12_ & ~n1454;
  assign n1557 = ~n1554 & ~n1555_1;
  assign n298 = n1556 | ~n1557;
  assign n1559 = REIP_REG_12_ & n1467;
  assign n1560_1 = REIP_REG_13_ & n1469;
  assign n1561 = ADDRESS_REG_11_ & ~n1454;
  assign n1562 = ~n1559 & ~n1560_1;
  assign n302 = n1561 | ~n1562;
  assign n1564 = REIP_REG_11_ & n1467;
  assign n1565_1 = REIP_REG_12_ & n1469;
  assign n1566 = ADDRESS_REG_10_ & ~n1454;
  assign n1567 = ~n1564 & ~n1565_1;
  assign n306 = n1566 | ~n1567;
  assign n1569 = REIP_REG_10_ & n1467;
  assign n1570_1 = REIP_REG_11_ & n1469;
  assign n1571 = ADDRESS_REG_9_ & ~n1454;
  assign n1572 = ~n1569 & ~n1570_1;
  assign n310 = n1571 | ~n1572;
  assign n1574 = REIP_REG_9_ & n1467;
  assign n1575_1 = REIP_REG_10_ & n1469;
  assign n1576 = ADDRESS_REG_8_ & ~n1454;
  assign n1577 = ~n1574 & ~n1575_1;
  assign n314 = n1576 | ~n1577;
  assign n1579 = REIP_REG_8_ & n1467;
  assign n1580_1 = REIP_REG_9_ & n1469;
  assign n1581 = ADDRESS_REG_7_ & ~n1454;
  assign n1582 = ~n1579 & ~n1580_1;
  assign n318 = n1581 | ~n1582;
  assign n1584 = REIP_REG_7_ & n1467;
  assign n1585_1 = REIP_REG_8_ & n1469;
  assign n1586 = ADDRESS_REG_6_ & ~n1454;
  assign n1587 = ~n1584 & ~n1585_1;
  assign n322 = n1586 | ~n1587;
  assign n1589 = REIP_REG_6_ & n1467;
  assign n1590_1 = REIP_REG_7_ & n1469;
  assign n1591 = ADDRESS_REG_5_ & ~n1454;
  assign n1592 = ~n1589 & ~n1590_1;
  assign n326 = n1591 | ~n1592;
  assign n1594 = REIP_REG_5_ & n1467;
  assign n1595_1 = REIP_REG_6_ & n1469;
  assign n1596 = ADDRESS_REG_4_ & ~n1454;
  assign n1597 = ~n1594 & ~n1595_1;
  assign n330 = n1596 | ~n1597;
  assign n1599 = REIP_REG_4_ & n1467;
  assign n1600_1 = REIP_REG_5_ & n1469;
  assign n1601 = ADDRESS_REG_3_ & ~n1454;
  assign n1602 = ~n1599 & ~n1600_1;
  assign n334 = n1601 | ~n1602;
  assign n1604 = REIP_REG_3_ & n1467;
  assign n1605_1 = REIP_REG_4_ & n1469;
  assign n1606 = ADDRESS_REG_2_ & ~n1454;
  assign n1607 = ~n1604 & ~n1605_1;
  assign n338 = n1606 | ~n1607;
  assign n1609 = REIP_REG_2_ & n1467;
  assign n1610_1 = REIP_REG_3_ & n1469;
  assign n1611 = ADDRESS_REG_1_ & ~n1454;
  assign n1612 = ~n1609 & ~n1610_1;
  assign n342 = n1611 | ~n1612;
  assign n1614 = REIP_REG_1_ & n1467;
  assign n1615_1 = REIP_REG_2_ & n1469;
  assign n1616 = ADDRESS_REG_0_ & ~n1454;
  assign n1617 = ~n1614 & ~n1615_1;
  assign n346 = n1616 | ~n1617;
  assign n1619 = ~STATE_REG_2_ & STATE_REG_1_;
  assign n1620_1 = NA_N & n1619;
  assign n1621 = READY_N & STATE_REG_1_;
  assign n1622 = ~HOLD & ~REQUESTPENDING_REG;
  assign n1623 = n1621 & ~n1622;
  assign n1624 = ~STATE_REG_2_ & ~STATE_REG_1_;
  assign n1625_1 = HOLD & ~REQUESTPENDING_REG;
  assign n1626 = n1624 & n1625_1;
  assign n1627 = ~n1623 & ~n1626;
  assign n1628 = STATE_REG_0_ & ~n1620_1;
  assign n1629 = ~n1627 & n1628;
  assign n1630_1 = ~n1467 & ~n1629;
  assign n1631 = ~HOLD & REQUESTPENDING_REG;
  assign n1632 = STATE_REG_0_ & ~n1631;
  assign n1633 = ~n1622 & n1632;
  assign n1634 = ~NA_N & ~STATE_REG_0_;
  assign n1635_1 = ~READY_N & n1622;
  assign n1636 = ~READY_N & n1631;
  assign n1637 = STATE_REG_1_ & ~n1635_1;
  assign n1638 = ~n1636 & n1637;
  assign n1639 = ~n1633 & ~n1634;
  assign n1640_1 = ~n1638 & n1639;
  assign n1641 = STATE_REG_2_ & ~n1640_1;
  assign n350 = ~n1630_1 | n1641;
  assign n1643 = STATE_REG_2_ & ~n1632;
  assign n1644 = STATE_REG_0_ & REQUESTPENDING_REG;
  assign n1645_1 = ~STATE_REG_2_ & n1644;
  assign n1646 = ~n1643 & ~n1645_1;
  assign n1647 = ~STATE_REG_1_ & ~n1646;
  assign n1648 = ~READY_N & HOLD;
  assign n1649 = STATE_REG_0_ & ~n1648;
  assign n1650_1 = STATE_REG_2_ & ~n1649;
  assign n1651 = ~n1635_1 & ~n1650_1;
  assign n1652 = STATE_REG_1_ & n1651;
  assign n1653 = READY_N & n1454;
  assign n1654 = ~n1469 & ~n1653;
  assign n1655_1 = ~n1647 & ~n1652;
  assign n355 = ~n1654 | ~n1655_1;
  assign n1657 = STATE_REG_1_ & ~n1636;
  assign n1658 = n1644 & ~n1657;
  assign n1659 = ~STATE_REG_2_ & ~n1658;
  assign n1660_1 = STATE_REG_2_ & n1632;
  assign n1661 = NA_N & ~STATE_REG_0_;
  assign n1662 = STATE_REG_2_ & ~n1631;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~STATE_REG_1_ & ~n1663;
  assign n1665_1 = ~n1659 & ~n1660_1;
  assign n360 = n1664 | ~n1665_1;
  assign n1667 = ~BS16_N & ~n1624;
  assign n1668 = STATE_REG_0_ & n1619;
  assign n1669 = ~STATE_REG_1_ & ~STATE_REG_0_;
  assign n1670_1 = ~n1668 & ~n1669;
  assign n1671 = n1667 & ~n1670_1;
  assign n1672 = DATAWIDTH_REG_0_ & n1670_1;
  assign n365 = n1671 | n1672;
  assign n1674 = DATAWIDTH_REG_1_ & n1670_1;
  assign n1675_1 = ~n1667 & ~n1670_1;
  assign n370 = n1674 | n1675_1;
  assign n375 = DATAWIDTH_REG_2_ & n1670_1;
  assign n380 = DATAWIDTH_REG_3_ & n1670_1;
  assign n385 = DATAWIDTH_REG_4_ & n1670_1;
  assign n390 = DATAWIDTH_REG_5_ & n1670_1;
  assign n395 = DATAWIDTH_REG_6_ & n1670_1;
  assign n400 = DATAWIDTH_REG_7_ & n1670_1;
  assign n405 = DATAWIDTH_REG_8_ & n1670_1;
  assign n410 = DATAWIDTH_REG_9_ & n1670_1;
  assign n415 = DATAWIDTH_REG_10_ & n1670_1;
  assign n420 = DATAWIDTH_REG_11_ & n1670_1;
  assign n425 = DATAWIDTH_REG_12_ & n1670_1;
  assign n430 = DATAWIDTH_REG_13_ & n1670_1;
  assign n435 = DATAWIDTH_REG_14_ & n1670_1;
  assign n440 = DATAWIDTH_REG_15_ & n1670_1;
  assign n445 = DATAWIDTH_REG_16_ & n1670_1;
  assign n450 = DATAWIDTH_REG_17_ & n1670_1;
  assign n455 = DATAWIDTH_REG_18_ & n1670_1;
  assign n460 = DATAWIDTH_REG_19_ & n1670_1;
  assign n465 = DATAWIDTH_REG_20_ & n1670_1;
  assign n470 = DATAWIDTH_REG_21_ & n1670_1;
  assign n475 = DATAWIDTH_REG_22_ & n1670_1;
  assign n480 = DATAWIDTH_REG_23_ & n1670_1;
  assign n485 = DATAWIDTH_REG_24_ & n1670_1;
  assign n490 = DATAWIDTH_REG_25_ & n1670_1;
  assign n495 = DATAWIDTH_REG_26_ & n1670_1;
  assign n500 = DATAWIDTH_REG_27_ & n1670_1;
  assign n505 = DATAWIDTH_REG_28_ & n1670_1;
  assign n510 = DATAWIDTH_REG_29_ & n1670_1;
  assign n515 = DATAWIDTH_REG_30_ & n1670_1;
  assign n520 = DATAWIDTH_REG_31_ & n1670_1;
  assign n1707 = STATE2_REG_2_ & STATE2_REG_1_;
  assign n1708 = READY_N & STATE2_REG_1_;
  assign n1709 = ~STATE2_REG_0_ & ~n1708;
  assign n1710_1 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1711 = INSTQUEUERD_ADDR_REG_1_ & n1710_1;
  assign n1712 = INSTQUEUERD_ADDR_REG_2_ & n1711;
  assign n1713 = INSTQUEUE_REG_15__0_ & n1712;
  assign n1714_1 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_1_;
  assign n1715 = INSTQUEUERD_ADDR_REG_2_ & n1714_1;
  assign n1716 = ~INSTQUEUERD_ADDR_REG_0_ & n1715;
  assign n1717 = INSTQUEUE_REG_14__0_ & n1716;
  assign n1718_1 = INSTQUEUERD_ADDR_REG_2_ & n1710_1;
  assign n1719 = ~INSTQUEUERD_ADDR_REG_1_ & n1718_1;
  assign n1720 = INSTQUEUE_REG_13__0_ & n1719;
  assign n1721 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_2_;
  assign n1722_1 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_0_;
  assign n1723 = n1721 & n1722_1;
  assign n1724 = INSTQUEUE_REG_12__0_ & n1723;
  assign n1725 = ~n1713 & ~n1717;
  assign n1726_1 = ~n1720 & n1725;
  assign n1727 = ~n1724 & n1726_1;
  assign n1728 = ~INSTQUEUERD_ADDR_REG_2_ & n1711;
  assign n1729 = INSTQUEUE_REG_11__0_ & n1728;
  assign n1730_1 = ~INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_0_;
  assign n1731 = n1714_1 & n1730_1;
  assign n1732 = INSTQUEUE_REG_10__0_ & n1731;
  assign n1733 = ~INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_1_;
  assign n1734_1 = n1710_1 & n1733;
  assign n1735 = INSTQUEUE_REG_9__0_ & n1734_1;
  assign n1736 = ~INSTQUEUERD_ADDR_REG_2_ & n1722_1;
  assign n1737 = INSTQUEUERD_ADDR_REG_3_ & n1736;
  assign n1738_1 = INSTQUEUE_REG_8__0_ & n1737;
  assign n1739 = ~n1729 & ~n1732;
  assign n1740 = ~n1735 & n1739;
  assign n1741 = ~n1738_1 & n1740;
  assign n1742_1 = INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_1_;
  assign n1743 = ~INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUERD_ADDR_REG_0_;
  assign n1744 = n1742_1 & n1743;
  assign n1745 = INSTQUEUE_REG_6__0_ & n1744;
  assign n1746_1 = INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1747 = ~INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUERD_ADDR_REG_1_;
  assign n1748 = n1746_1 & n1747;
  assign n1749 = INSTQUEUE_REG_5__0_ & n1748;
  assign n1750_1 = ~INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_2_;
  assign n1751 = n1722_1 & n1750_1;
  assign n1752 = INSTQUEUE_REG_4__0_ & n1751;
  assign n1753 = INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1754_1 = ~INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n1755 = n1753 & n1754_1;
  assign n1756 = INSTQUEUE_REG_3__0_ & n1755;
  assign n1757 = ~n1745 & ~n1749;
  assign n1758_1 = ~n1752 & n1757;
  assign n1759 = ~n1756 & n1758_1;
  assign n1760 = INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_0_;
  assign n1761 = n1754_1 & n1760;
  assign n1762_1 = INSTQUEUE_REG_2__0_ & n1761;
  assign n1763 = ~INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1764 = n1754_1 & n1763;
  assign n1765 = INSTQUEUE_REG_1__0_ & n1764;
  assign n1766_1 = ~INSTQUEUERD_ADDR_REG_3_ & n1736;
  assign n1767 = INSTQUEUE_REG_0__0_ & n1766_1;
  assign n1768 = INSTQUEUERD_ADDR_REG_2_ & n1753;
  assign n1769 = ~INSTQUEUERD_ADDR_REG_3_ & n1768;
  assign n1770_1 = INSTQUEUE_REG_7__0_ & n1769;
  assign n1771 = ~n1762_1 & ~n1765;
  assign n1772 = ~n1767 & n1771;
  assign n1773 = ~n1770_1 & n1772;
  assign n1774_1 = n1727 & n1741;
  assign n1775 = n1759 & n1774_1;
  assign n1776 = n1773 & n1775;
  assign n1777 = INSTQUEUE_REG_15__1_ & n1712;
  assign n1778_1 = INSTQUEUE_REG_14__1_ & n1716;
  assign n1779 = INSTQUEUE_REG_13__1_ & n1719;
  assign n1780 = INSTQUEUE_REG_12__1_ & n1723;
  assign n1781 = ~n1777 & ~n1778_1;
  assign n1782_1 = ~n1779 & n1781;
  assign n1783 = ~n1780 & n1782_1;
  assign n1784 = INSTQUEUE_REG_11__1_ & n1728;
  assign n1785 = INSTQUEUE_REG_10__1_ & n1731;
  assign n1786_1 = INSTQUEUE_REG_9__1_ & n1734_1;
  assign n1787 = INSTQUEUE_REG_8__1_ & n1737;
  assign n1788 = ~n1784 & ~n1785;
  assign n1789 = ~n1786_1 & n1788;
  assign n1790_1 = ~n1787 & n1789;
  assign n1791 = INSTQUEUE_REG_6__1_ & n1744;
  assign n1792 = INSTQUEUE_REG_5__1_ & n1748;
  assign n1793 = INSTQUEUE_REG_4__1_ & n1751;
  assign n1794_1 = INSTQUEUE_REG_3__1_ & n1755;
  assign n1795 = ~n1791 & ~n1792;
  assign n1796 = ~n1793 & n1795;
  assign n1797 = ~n1794_1 & n1796;
  assign n1798_1 = INSTQUEUE_REG_2__1_ & n1761;
  assign n1799 = INSTQUEUE_REG_1__1_ & n1764;
  assign n1800 = INSTQUEUE_REG_0__1_ & n1766_1;
  assign n1801 = INSTQUEUE_REG_7__1_ & n1769;
  assign n1802_1 = ~n1798_1 & ~n1799;
  assign n1803 = ~n1800 & n1802_1;
  assign n1804 = ~n1801 & n1803;
  assign n1805 = n1783 & n1790_1;
  assign n1806_1 = n1797 & n1805;
  assign n1807 = n1804 & n1806_1;
  assign n1808 = n1776 & n1807;
  assign n1809 = INSTQUEUE_REG_15__3_ & n1712;
  assign n1810_1 = INSTQUEUE_REG_14__3_ & n1716;
  assign n1811 = INSTQUEUE_REG_13__3_ & n1719;
  assign n1812 = INSTQUEUE_REG_12__3_ & n1723;
  assign n1813 = ~n1809 & ~n1810_1;
  assign n1814_1 = ~n1811 & n1813;
  assign n1815 = ~n1812 & n1814_1;
  assign n1816 = INSTQUEUE_REG_11__3_ & n1728;
  assign n1817 = INSTQUEUE_REG_10__3_ & n1731;
  assign n1818_1 = INSTQUEUE_REG_9__3_ & n1734_1;
  assign n1819 = INSTQUEUE_REG_8__3_ & n1737;
  assign n1820 = ~n1816 & ~n1817;
  assign n1821 = ~n1818_1 & n1820;
  assign n1822_1 = ~n1819 & n1821;
  assign n1823 = INSTQUEUE_REG_6__3_ & n1744;
  assign n1824 = INSTQUEUE_REG_5__3_ & n1748;
  assign n1825 = INSTQUEUE_REG_4__3_ & n1751;
  assign n1826_1 = INSTQUEUE_REG_3__3_ & n1755;
  assign n1827 = ~n1823 & ~n1824;
  assign n1828 = ~n1825 & n1827;
  assign n1829 = ~n1826_1 & n1828;
  assign n1830_1 = INSTQUEUE_REG_2__3_ & n1761;
  assign n1831 = INSTQUEUE_REG_1__3_ & n1764;
  assign n1832 = INSTQUEUE_REG_0__3_ & n1766_1;
  assign n1833 = INSTQUEUE_REG_7__3_ & n1769;
  assign n1834_1 = ~n1830_1 & ~n1831;
  assign n1835 = ~n1832 & n1834_1;
  assign n1836 = ~n1833 & n1835;
  assign n1837 = n1815 & n1822_1;
  assign n1838_1 = n1829 & n1837;
  assign n1839 = n1836 & n1838_1;
  assign n1840 = n1808 & ~n1839;
  assign n1841 = INSTQUEUE_REG_8__6_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n1842 = ~INSTQUEUERD_ADDR_REG_1_ & n1841;
  assign n1843_1 = ~INSTQUEUERD_ADDR_REG_0_ & n1842;
  assign n1844 = INSTQUEUERD_ADDR_REG_3_ & n1843_1;
  assign n1845 = INSTQUEUE_REG_0__6_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n1846 = ~INSTQUEUERD_ADDR_REG_1_ & n1845;
  assign n1847 = ~INSTQUEUERD_ADDR_REG_0_ & n1846;
  assign n1848_1 = ~INSTQUEUERD_ADDR_REG_3_ & n1847;
  assign n1849 = INSTQUEUE_REG_11__6_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1850 = INSTQUEUERD_ADDR_REG_1_ & n1849;
  assign n1851 = ~INSTQUEUERD_ADDR_REG_2_ & n1850;
  assign n1852 = INSTQUEUERD_ADDR_REG_0_ & n1851;
  assign n1853_1 = INSTQUEUE_REG_10__6_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1854 = INSTQUEUERD_ADDR_REG_1_ & n1853_1;
  assign n1855 = ~INSTQUEUERD_ADDR_REG_2_ & n1854;
  assign n1856 = ~INSTQUEUERD_ADDR_REG_0_ & n1855;
  assign n1857 = ~n1844 & ~n1848_1;
  assign n1858_1 = ~n1852 & n1857;
  assign n1859 = ~n1856 & n1858_1;
  assign n1860 = INSTQUEUE_REG_3__6_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1861 = n1754_1 & n1860;
  assign n1862 = INSTQUEUERD_ADDR_REG_1_ & n1861;
  assign n1863_1 = INSTQUEUE_REG_9__6_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1864 = INSTQUEUERD_ADDR_REG_0_ & n1863_1;
  assign n1865 = ~INSTQUEUERD_ADDR_REG_2_ & n1864;
  assign n1866 = ~INSTQUEUERD_ADDR_REG_1_ & n1865;
  assign n1867 = ~n1862 & ~n1866;
  assign n1868_1 = n1721 & n1760;
  assign n1869 = INSTQUEUE_REG_14__6_ & n1868_1;
  assign n1870 = n1721 & n1763;
  assign n1871 = INSTQUEUE_REG_13__6_ & n1870;
  assign n1872 = n1721 & n1753;
  assign n1873_1 = INSTQUEUE_REG_15__6_ & n1872;
  assign n1874 = ~n1869 & ~n1871;
  assign n1875 = ~n1873_1 & n1874;
  assign n1876 = n1750_1 & n1760;
  assign n1877 = INSTQUEUE_REG_6__6_ & n1876;
  assign n1878_1 = n1750_1 & n1763;
  assign n1879 = INSTQUEUE_REG_5__6_ & n1878_1;
  assign n1880 = INSTQUEUE_REG_12__6_ & n1722_1;
  assign n1881 = n1721 & n1880;
  assign n1882 = ~n1877 & ~n1879;
  assign n1883_1 = ~n1881 & n1882;
  assign n1884 = INSTQUEUE_REG_4__6_ & n1722_1;
  assign n1885 = n1750_1 & n1884;
  assign n1886 = INSTQUEUE_REG_2__6_ & n1754_1;
  assign n1887 = n1760 & n1886;
  assign n1888_1 = INSTQUEUE_REG_1__6_ & n1754_1;
  assign n1889 = n1763 & n1888_1;
  assign n1890 = n1750_1 & n1753;
  assign n1891 = INSTQUEUE_REG_7__6_ & n1890;
  assign n1892 = ~n1885 & ~n1887;
  assign n1893_1 = ~n1889 & n1892;
  assign n1894 = ~n1891 & n1893_1;
  assign n1895 = n1859 & n1867;
  assign n1896 = n1875 & n1895;
  assign n1897 = n1883_1 & n1896;
  assign n1898_1 = n1894 & n1897;
  assign n1899 = INSTQUEUE_REG_15__7_ & n1712;
  assign n1900 = INSTQUEUE_REG_14__7_ & n1716;
  assign n1901 = INSTQUEUE_REG_13__7_ & n1719;
  assign n1902 = INSTQUEUE_REG_12__7_ & n1723;
  assign n1903_1 = ~n1899 & ~n1900;
  assign n1904 = ~n1901 & n1903_1;
  assign n1905 = ~n1902 & n1904;
  assign n1906 = INSTQUEUE_REG_11__7_ & n1728;
  assign n1907 = INSTQUEUE_REG_10__7_ & n1731;
  assign n1908_1 = INSTQUEUE_REG_9__7_ & n1734_1;
  assign n1909 = INSTQUEUE_REG_8__7_ & n1737;
  assign n1910 = ~n1906 & ~n1907;
  assign n1911 = ~n1908_1 & n1910;
  assign n1912 = ~n1909 & n1911;
  assign n1913_1 = INSTQUEUE_REG_6__7_ & n1744;
  assign n1914 = INSTQUEUE_REG_5__7_ & n1748;
  assign n1915 = INSTQUEUE_REG_4__7_ & n1751;
  assign n1916 = INSTQUEUE_REG_3__7_ & n1755;
  assign n1917 = ~n1913_1 & ~n1914;
  assign n1918_1 = ~n1915 & n1917;
  assign n1919 = ~n1916 & n1918_1;
  assign n1920 = INSTQUEUE_REG_2__7_ & n1761;
  assign n1921 = INSTQUEUE_REG_1__7_ & n1764;
  assign n1922 = INSTQUEUE_REG_0__7_ & n1766_1;
  assign n1923_1 = INSTQUEUE_REG_7__7_ & n1769;
  assign n1924 = ~n1920 & ~n1921;
  assign n1925 = ~n1922 & n1924;
  assign n1926 = ~n1923_1 & n1925;
  assign n1927 = n1905 & n1912;
  assign n1928_1 = n1919 & n1927;
  assign n1929 = n1926 & n1928_1;
  assign n1930 = INSTQUEUERD_ADDR_REG_0_ & n1742_1;
  assign n1931 = INSTQUEUE_REG_15__5_ & n1930;
  assign n1932 = INSTQUEUERD_ADDR_REG_3_ & n1931;
  assign n1933_1 = INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_0_;
  assign n1934 = INSTQUEUERD_ADDR_REG_1_ & n1933_1;
  assign n1935 = INSTQUEUE_REG_14__5_ & n1934;
  assign n1936 = INSTQUEUERD_ADDR_REG_3_ & n1935;
  assign n1937 = ~n1932 & ~n1936;
  assign n1938_1 = INSTQUEUE_REG_9__5_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1939 = n1733 & n1938_1;
  assign n1940 = INSTQUEUERD_ADDR_REG_3_ & n1939;
  assign n1941 = INSTQUEUE_REG_3__5_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1942 = INSTQUEUERD_ADDR_REG_1_ & n1941;
  assign n1943_1 = ~INSTQUEUERD_ADDR_REG_2_ & n1942;
  assign n1944 = ~INSTQUEUERD_ADDR_REG_3_ & n1943_1;
  assign n1945 = ~n1940 & ~n1944;
  assign n1946 = INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_1_;
  assign n1947 = INSTQUEUERD_ADDR_REG_0_ & n1946;
  assign n1948_1 = INSTQUEUE_REG_13__5_ & n1947;
  assign n1949 = INSTQUEUERD_ADDR_REG_3_ & n1948_1;
  assign n1950 = INSTQUEUE_REG_12__5_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1951 = INSTQUEUERD_ADDR_REG_2_ & n1722_1;
  assign n1952 = n1950 & n1951;
  assign n1953_1 = ~INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_1_;
  assign n1954 = INSTQUEUERD_ADDR_REG_0_ & n1953_1;
  assign n1955 = INSTQUEUE_REG_11__5_ & n1954;
  assign n1956 = INSTQUEUERD_ADDR_REG_3_ & n1955;
  assign n1957 = INSTQUEUE_REG_10__5_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1958_1 = INSTQUEUERD_ADDR_REG_1_ & n1730_1;
  assign n1959 = n1957 & n1958_1;
  assign n1960 = ~n1949 & ~n1952;
  assign n1961 = ~n1956 & n1960;
  assign n1962 = ~n1959 & n1961;
  assign n1963_1 = INSTQUEUE_REG_8__5_ & INSTQUEUERD_ADDR_REG_3_;
  assign n1964 = n1736 & n1963_1;
  assign n1965 = INSTQUEUE_REG_6__5_ & INSTQUEUERD_ADDR_REG_1_;
  assign n1966 = INSTQUEUERD_ADDR_REG_2_ & n1743;
  assign n1967 = n1965 & n1966;
  assign n1968_1 = INSTQUEUE_REG_5__5_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1969 = INSTQUEUERD_ADDR_REG_2_ & n1747;
  assign n1970 = n1968_1 & n1969;
  assign n1971 = INSTQUEUE_REG_4__5_ & n1722_1;
  assign n1972 = INSTQUEUERD_ADDR_REG_2_ & n1971;
  assign n1973_1 = ~INSTQUEUERD_ADDR_REG_3_ & n1972;
  assign n1974 = ~n1964 & ~n1967;
  assign n1975 = ~n1970 & n1974;
  assign n1976 = ~n1973_1 & n1975;
  assign n1977 = INSTQUEUE_REG_2__5_ & n1754_1;
  assign n1978_1 = INSTQUEUERD_ADDR_REG_1_ & n1977;
  assign n1979 = ~INSTQUEUERD_ADDR_REG_0_ & n1978_1;
  assign n1980 = INSTQUEUE_REG_1__5_ & n1754_1;
  assign n1981 = INSTQUEUERD_ADDR_REG_0_ & n1980;
  assign n1982 = ~INSTQUEUERD_ADDR_REG_1_ & n1981;
  assign n1983_1 = INSTQUEUE_REG_0__5_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign n1984 = n1736 & n1983_1;
  assign n1985 = INSTQUEUERD_ADDR_REG_1_ & n1750_1;
  assign n1986 = INSTQUEUE_REG_7__5_ & n1985;
  assign n1987 = INSTQUEUERD_ADDR_REG_0_ & n1986;
  assign n1988_1 = ~n1979 & ~n1982;
  assign n1989 = ~n1984 & n1988_1;
  assign n1990 = ~n1987 & n1989;
  assign n1991 = n1937 & n1945;
  assign n1992 = n1962 & n1991;
  assign n1993_1 = n1976 & n1992;
  assign n1994 = n1990 & n1993_1;
  assign n1995 = INSTQUEUE_REG_11__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign n1996 = INSTQUEUERD_ADDR_REG_1_ & n1995;
  assign n1997 = ~INSTQUEUERD_ADDR_REG_2_ & n1996;
  assign n1998_1 = INSTQUEUERD_ADDR_REG_3_ & n1997;
  assign n1999 = INSTQUEUE_REG_3__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign n2000 = INSTQUEUERD_ADDR_REG_1_ & n1999;
  assign n2001 = ~INSTQUEUERD_ADDR_REG_2_ & n2000;
  assign n2002 = ~INSTQUEUERD_ADDR_REG_3_ & n2001;
  assign n2003_1 = INSTQUEUE_REG_9__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2004 = n1733 & n2003_1;
  assign n2005 = INSTQUEUERD_ADDR_REG_0_ & n2004;
  assign n2006 = INSTQUEUE_REG_10__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2007 = INSTQUEUERD_ADDR_REG_1_ & n2006;
  assign n2008_1 = ~INSTQUEUERD_ADDR_REG_2_ & n2007;
  assign n2009 = ~INSTQUEUERD_ADDR_REG_0_ & n2008_1;
  assign n2010 = ~n1998_1 & ~n2002;
  assign n2011 = ~n2005 & n2010;
  assign n2012 = ~n2009 & n2011;
  assign n2013_1 = INSTQUEUE_REG_8__4_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n2014 = ~INSTQUEUERD_ADDR_REG_1_ & n2013_1;
  assign n2015 = ~INSTQUEUERD_ADDR_REG_0_ & n2014;
  assign n2016 = INSTQUEUERD_ADDR_REG_3_ & n2015;
  assign n2017 = INSTQUEUE_REG_0__4_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n2018_1 = ~INSTQUEUERD_ADDR_REG_1_ & n2017;
  assign n2019 = ~INSTQUEUERD_ADDR_REG_0_ & n2018_1;
  assign n2020 = ~INSTQUEUERD_ADDR_REG_3_ & n2019;
  assign n2021 = INSTQUEUE_REG_15__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2022 = INSTQUEUERD_ADDR_REG_1_ & n2021;
  assign n2023_1 = INSTQUEUERD_ADDR_REG_2_ & n2022;
  assign n2024 = INSTQUEUERD_ADDR_REG_0_ & n2023_1;
  assign n2025 = INSTQUEUE_REG_14__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2026 = n1742_1 & n2025;
  assign n2027 = ~INSTQUEUERD_ADDR_REG_0_ & n2026;
  assign n2028_1 = ~n2016 & ~n2020;
  assign n2029 = ~n2024 & n2028_1;
  assign n2030 = ~n2027 & n2029;
  assign n2031 = INSTQUEUE_REG_6__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign n2032 = n1743 & n2031;
  assign n2033_1 = INSTQUEUERD_ADDR_REG_1_ & n2032;
  assign n2034 = INSTQUEUE_REG_13__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2035 = n1746_1 & n2034;
  assign n2036 = ~INSTQUEUERD_ADDR_REG_1_ & n2035;
  assign n2037 = INSTQUEUE_REG_12__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign n2038_1 = n1722_1 & n2037;
  assign n2039 = INSTQUEUERD_ADDR_REG_3_ & n2038_1;
  assign n2040 = INSTQUEUE_REG_4__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign n2041 = n1722_1 & n2040;
  assign n2042 = ~INSTQUEUERD_ADDR_REG_3_ & n2041;
  assign n2043_1 = ~n2033_1 & ~n2036;
  assign n2044 = ~n2039 & n2043_1;
  assign n2045 = ~n2042 & n2044;
  assign n2046 = INSTQUEUE_REG_2__4_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign n2047 = ~INSTQUEUERD_ADDR_REG_2_ & n2046;
  assign n2048_1 = ~INSTQUEUERD_ADDR_REG_0_ & n2047;
  assign n2049 = INSTQUEUERD_ADDR_REG_1_ & n2048_1;
  assign n2050 = INSTQUEUE_REG_5__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign n2051 = INSTQUEUERD_ADDR_REG_2_ & n2050;
  assign n2052 = ~INSTQUEUERD_ADDR_REG_3_ & n2051;
  assign n2053_1 = ~INSTQUEUERD_ADDR_REG_1_ & n2052;
  assign n2054 = INSTQUEUE_REG_7__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign n2055 = INSTQUEUERD_ADDR_REG_2_ & n2054;
  assign n2056 = ~INSTQUEUERD_ADDR_REG_3_ & n2055;
  assign n2057 = INSTQUEUERD_ADDR_REG_1_ & n2056;
  assign n2058_1 = INSTQUEUE_REG_1__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign n2059 = n1754_1 & n2058_1;
  assign n2060 = ~INSTQUEUERD_ADDR_REG_1_ & n2059;
  assign n2061 = ~n2049 & ~n2053_1;
  assign n2062 = ~n2057 & n2061;
  assign n2063_1 = ~n2060 & n2062;
  assign n2064 = n2012 & n2030;
  assign n2065 = n2045 & n2064;
  assign n2066 = n2063_1 & n2065;
  assign n2067 = n1898_1 & ~n1929;
  assign n2068_1 = ~n1994 & n2067;
  assign n2069 = ~n2066 & n2068_1;
  assign n2070 = INSTQUEUE_REG_15__2_ & n1712;
  assign n2071 = INSTQUEUE_REG_14__2_ & n1716;
  assign n2072 = INSTQUEUE_REG_13__2_ & n1719;
  assign n2073_1 = INSTQUEUE_REG_12__2_ & n1723;
  assign n2074 = ~n2070 & ~n2071;
  assign n2075 = ~n2072 & n2074;
  assign n2076 = ~n2073_1 & n2075;
  assign n2077 = INSTQUEUE_REG_11__2_ & n1728;
  assign n2078_1 = INSTQUEUE_REG_10__2_ & n1731;
  assign n2079 = INSTQUEUE_REG_9__2_ & n1734_1;
  assign n2080 = INSTQUEUE_REG_8__2_ & n1737;
  assign n2081 = ~n2077 & ~n2078_1;
  assign n2082 = ~n2079 & n2081;
  assign n2083_1 = ~n2080 & n2082;
  assign n2084 = INSTQUEUE_REG_6__2_ & n1744;
  assign n2085 = INSTQUEUE_REG_5__2_ & n1748;
  assign n2086 = INSTQUEUE_REG_4__2_ & n1751;
  assign n2087 = INSTQUEUE_REG_3__2_ & n1755;
  assign n2088_1 = ~n2084 & ~n2085;
  assign n2089 = ~n2086 & n2088_1;
  assign n2090 = ~n2087 & n2089;
  assign n2091 = INSTQUEUE_REG_2__2_ & n1761;
  assign n2092 = INSTQUEUE_REG_1__2_ & n1764;
  assign n2093_1 = INSTQUEUE_REG_0__2_ & n1766_1;
  assign n2094 = INSTQUEUE_REG_7__2_ & n1769;
  assign n2095 = ~n2091 & ~n2092;
  assign n2096 = ~n2093_1 & n2095;
  assign n2097 = ~n2094 & n2096;
  assign n2098_1 = n2076 & n2083_1;
  assign n2099 = n2090 & n2098_1;
  assign n2100 = n2097 & n2099;
  assign n2101 = n2069 & n2100;
  assign n2102 = n1840 & n2101;
  assign n2103_1 = n1776 & ~n1807;
  assign n2104 = n1839 & ~n2100;
  assign n2105 = ~n1898_1 & n2066;
  assign n2106 = ~n1929 & n2105;
  assign n2107 = ~n1994 & n2106;
  assign n2108_1 = n2104 & n2107;
  assign n2109 = n2103_1 & n2108_1;
  assign n2110 = ~n2102 & ~n2109;
  assign n2111 = n1898_1 & n1994;
  assign n2112 = n2100 & n2107;
  assign n2113_1 = ~n1839 & n2112;
  assign n2114 = ~n2111 & ~n2113_1;
  assign n2115 = ~n1776 & ~n1839;
  assign n2116 = n2066 & n2115;
  assign n2117 = n2100 & n2116;
  assign n2118_1 = ~n2114 & n2117;
  assign n2119 = n2110 & ~n2118_1;
  assign n2120 = INSTQUEUERD_ADDR_REG_4_ & ~INSTQUEUEWR_ADDR_REG_4_;
  assign n2121 = ~INSTQUEUERD_ADDR_REG_3_ & INSTQUEUEWR_ADDR_REG_3_;
  assign n2122 = INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUEWR_ADDR_REG_3_;
  assign n2123_1 = ~INSTQUEUERD_ADDR_REG_2_ & INSTQUEUEWR_ADDR_REG_2_;
  assign n2124 = INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUEWR_ADDR_REG_2_;
  assign n2125 = INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUEWR_ADDR_REG_0_;
  assign n2126 = INSTQUEUEWR_ADDR_REG_1_ & ~n2125;
  assign n2127 = ~INSTQUEUEWR_ADDR_REG_1_ & n2125;
  assign n2128_1 = ~INSTQUEUERD_ADDR_REG_1_ & ~n2127;
  assign n2129 = ~n2126 & ~n2128_1;
  assign n2130 = ~n2124 & ~n2129;
  assign n2131 = ~n2123_1 & ~n2130;
  assign n2132 = ~n2122 & ~n2131;
  assign n2133_1 = ~n2121 & ~n2132;
  assign n2134 = ~INSTQUEUERD_ADDR_REG_4_ & INSTQUEUEWR_ADDR_REG_4_;
  assign n2135 = n2133_1 & ~n2134;
  assign n2136 = ~n2120 & ~n2135;
  assign n2137 = STATE2_REG_0_ & ~n2066;
  assign n2138_1 = ~n1776 & n2137;
  assign n2139 = ~n2136 & n2138_1;
  assign n2140 = STATE2_REG_0_ & n1994;
  assign n2141 = n1807 & n2140;
  assign n2142 = ~n2136 & n2141;
  assign n2143_1 = STATE2_REG_0_ & n1776;
  assign n2144 = n1807 & n2143_1;
  assign n2145 = ~n1807 & n2143_1;
  assign n2146 = ~n1807 & n2140;
  assign n2147 = ~n1994 & n2066;
  assign n2148_1 = STATE2_REG_0_ & n2147;
  assign n2149 = ~n1776 & ~n1807;
  assign n2150 = n2148_1 & n2149;
  assign n2151 = STATE2_REG_0_ & ~n1994;
  assign n2152 = ~n1776 & n1807;
  assign n2153_1 = n2151 & n2152;
  assign n2154 = ~n2144 & ~n2145;
  assign n2155 = ~n2146 & n2154;
  assign n2156 = ~n2150 & n2155;
  assign n2157 = ~n2153_1 & n2156;
  assign n2158_1 = ~n2136 & ~n2157;
  assign n2159 = ~n2142 & ~n2158_1;
  assign n2160 = ~STATE2_REG_0_ & INSTQUEUERD_ADDR_REG_4_;
  assign n2161 = ~n2120 & ~n2134;
  assign n2162 = ~n2133_1 & ~n2161;
  assign n2163_1 = n2133_1 & n2161;
  assign n2164 = ~n2162 & ~n2163_1;
  assign n2165 = n2138_1 & ~n2164;
  assign n2166 = ~n2160 & ~n2165;
  assign n2167 = n2141 & ~n2164;
  assign n2168_1 = ~n2157 & ~n2164;
  assign n2169 = ~n2167 & ~n2168_1;
  assign n2170 = ~n2166 & n2169;
  assign n2171 = n2139 & n2159;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173_1 = ~n2121 & ~n2122;
  assign n2174 = ~n2131 & ~n2173_1;
  assign n2175 = n2131 & n2173_1;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n2141 & ~n2176;
  assign n2178_1 = STATE2_REG_0_ & ~n2177;
  assign n2179 = ~n2157 & ~n2176;
  assign n2180 = n2178_1 & ~n2179;
  assign n2181 = ~STATE2_REG_0_ & INSTQUEUERD_ADDR_REG_3_;
  assign n2182 = n2138_1 & ~n2176;
  assign n2183_1 = ~n2181 & ~n2182;
  assign n2184 = ~n2180 & n2183_1;
  assign n2185 = n2166 & ~n2169;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2123_1 & ~n2124;
  assign n2188_1 = ~n2129 & ~n2187;
  assign n2189 = n2129 & n2187;
  assign n2190 = ~n2188_1 & ~n2189;
  assign n2191 = n2138_1 & ~n2190;
  assign n2192 = ~STATE2_REG_0_ & INSTQUEUERD_ADDR_REG_2_;
  assign n2193_1 = ~n2191 & ~n2192;
  assign n2194 = ~n2144 & ~n2151;
  assign n2195 = n1807 & ~n2194;
  assign n2196 = n2193_1 & ~n2195;
  assign n2197 = n2141 & ~n2190;
  assign n2198_1 = ~n1776 & ~n2066;
  assign n2199 = STATE2_REG_0_ & ~n2198_1;
  assign n2200 = ~n2197 & n2199;
  assign n2201 = ~n2157 & ~n2190;
  assign n2202 = n2200 & ~n2201;
  assign n2203_1 = ~n2196 & n2202;
  assign n2204 = n2180 & ~n2183_1;
  assign n2205 = ~n2203_1 & ~n2204;
  assign n2206 = ~INSTQUEUERD_ADDR_REG_1_ & INSTQUEUEWR_ADDR_REG_1_;
  assign n2207 = INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUEWR_ADDR_REG_1_;
  assign n2208_1 = ~n2206 & ~n2207;
  assign n2209 = ~n2125 & ~n2208_1;
  assign n2210 = n2125 & n2208_1;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = n2141 & ~n2211;
  assign n2213_1 = STATE2_REG_0_ & ~n2212;
  assign n2214 = ~n2157 & ~n2211;
  assign n2215 = n2213_1 & ~n2214;
  assign n2216 = ~STATE2_REG_0_ & INSTQUEUERD_ADDR_REG_1_;
  assign n2217 = n2138_1 & ~n2211;
  assign n2218_1 = STATE2_REG_0_ & n2066;
  assign n2219 = ~n1807 & n2218_1;
  assign n2220 = ~n2140 & ~n2219;
  assign n2221 = ~n2216 & ~n2217;
  assign n2222 = n2220 & n2221;
  assign n2223_1 = ~n2145 & n2222;
  assign n2224 = ~n2215 & n2223_1;
  assign n2225 = n2196 & ~n2202;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = n2215 & ~n2223_1;
  assign n2228_1 = ~INSTQUEUERD_ADDR_REG_0_ & INSTQUEUEWR_ADDR_REG_0_;
  assign n2229 = ~n2125 & ~n2228_1;
  assign n2230 = n2141 & ~n2229;
  assign n2231 = n2199 & ~n2230;
  assign n2232 = ~n2157 & ~n2229;
  assign n2233_1 = n2231 & ~n2232;
  assign n2234 = ~n1807 & ~n1994;
  assign n2235 = n2138_1 & n2234;
  assign n2236 = n2233_1 & n2235;
  assign n2237 = ~STATE2_REG_0_ & INSTQUEUERD_ADDR_REG_0_;
  assign n2238_1 = n2138_1 & ~n2229;
  assign n2239 = ~n1776 & n2148_1;
  assign n2240 = ~n2237 & ~n2238_1;
  assign n2241 = ~n2239 & n2240;
  assign n2242 = ~n2195 & n2241;
  assign n2243_1 = n2233_1 & ~n2242;
  assign n2244 = n2235 & ~n2242;
  assign n2245 = ~n2227 & ~n2236;
  assign n2246 = ~n2243_1 & n2245;
  assign n2247 = ~n2244 & n2246;
  assign n2248_1 = n2226 & ~n2247;
  assign n2249 = n2205 & ~n2248_1;
  assign n2250 = n2186 & ~n2249;
  assign n2251 = n2172 & ~n2250;
  assign n2252 = ~n2139 & ~n2159;
  assign n2253_1 = ~n2251 & ~n2252;
  assign n2254 = ~n2159 & ~n2253_1;
  assign n2255 = STATE2_REG_0_ & n2159;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n2139 & ~n2256;
  assign n2258_1 = n2159 & ~n2253_1;
  assign n2259 = ~STATE2_REG_0_ & ~n2159;
  assign n2260 = ~n2258_1 & ~n2259;
  assign n2261 = ~n2139 & ~n2260;
  assign n2262 = ~n2257 & ~n2261;
  assign n2263_1 = ~n2119 & n2262;
  assign n2264 = ~n1807 & ~n1839;
  assign n2265 = ~n1776 & n2264;
  assign n2266 = n2101 & n2265;
  assign n2267 = ~n2262 & n2266;
  assign n2268_1 = n1808 & n2108_1;
  assign n2269 = n2164 & n2176;
  assign n2270 = n2211 & n2269;
  assign n2271 = n2190 & n2270;
  assign n2272 = n2136 & ~n2271;
  assign n2273_1 = n2268_1 & ~n2272;
  assign n2274 = ~n2263_1 & ~n2267;
  assign n2275 = ~n2273_1 & n2274;
  assign n2276 = ~n1929 & ~n2275;
  assign n2277 = ~n1776 & ~n2262;
  assign n2278_1 = n2113_1 & n2277;
  assign n2279 = n2066 & n2111;
  assign n2280 = ~n1839 & ~n1929;
  assign n2281 = n2100 & n2280;
  assign n2282 = n2279 & n2281;
  assign n2283_1 = ~n2262 & n2282;
  assign n2284 = ~n1776 & ~n2283_1;
  assign n2285 = n1807 & ~n2272;
  assign n2286 = n2108_1 & ~n2285;
  assign n2287 = n1776 & ~n2286;
  assign n2288_1 = ~n1807 & n2262;
  assign n2289 = ~n2284 & ~n2287;
  assign n2290 = ~n2288_1 & n2289;
  assign n2291 = STATE_REG_2_ & ~STATE_REG_1_;
  assign n2292 = ~n1619 & ~n2291;
  assign n2293_1 = ~STATE_REG_0_ & ~n2292;
  assign n2294 = ~n2149 & ~n2293_1;
  assign n2295 = ~n1808 & n2294;
  assign n2296 = ~READY_N & ~n2295;
  assign n2297 = n2290 & ~n2296;
  assign n2298_1 = ~FLUSH_REG & ~MORE_REG;
  assign n2299 = n2297 & ~n2298_1;
  assign n2300 = STATE2_REG_1_ & ~FLUSH_REG;
  assign n2301 = INSTQUEUERD_ADDR_REG_2_ & n2300;
  assign n2302 = INSTADDRPOINTER_REG_0_ & INSTADDRPOINTER_REG_31_;
  assign n2303_1 = INSTADDRPOINTER_REG_0_ & ~INSTADDRPOINTER_REG_31_;
  assign n2304 = ~n2302 & ~n2303_1;
  assign n2305 = STATE2_REG_1_ & ~n2304;
  assign n2306 = INSTADDRPOINTER_REG_0_ & ~INSTADDRPOINTER_REG_1_;
  assign n2307 = ~INSTADDRPOINTER_REG_0_ & INSTADDRPOINTER_REG_1_;
  assign n2308_1 = ~n2306 & ~n2307;
  assign n2309 = INSTADDRPOINTER_REG_31_ & ~n2308_1;
  assign n2310 = INSTADDRPOINTER_REG_1_ & ~INSTADDRPOINTER_REG_31_;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = FLUSH_REG & n2305;
  assign n2313_1 = ~n2311 & n2312;
  assign n2314 = ~n2301 & ~n2313_1;
  assign n2315 = n1839 & n2100;
  assign n2316 = n1776 & n2315;
  assign n2317 = n1807 & n2069;
  assign n2318_1 = n2316 & n2317;
  assign n2319 = INSTQUEUERD_ADDR_REG_2_ & ~n1753;
  assign n2320 = ~n1954 & ~n2319;
  assign n2321 = n2318_1 & ~n2320;
  assign n2322 = ~n2102 & ~n2266;
  assign n2323_1 = n2320 & ~n2322;
  assign n2324 = ~n1946 & ~n1953_1;
  assign n2325 = n2109 & ~n2324;
  assign n2326 = ~n2321 & ~n2323_1;
  assign n2327 = ~n2325 & n2326;
  assign n2328_1 = STATE2_REG_0_ & ~n1776;
  assign n2329 = n1807 & ~n2292;
  assign n2330 = n2328_1 & n2329;
  assign n2331 = STATE2_REG_0_ & n2149;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333_1 = n2282 & ~n2332;
  assign n2334 = STATE2_REG_0_ & n1808;
  assign n2335 = n2104 & n2334;
  assign n2336 = n2107 & n2335;
  assign n2337 = ~n2333_1 & ~n2336;
  assign n2338_1 = ~n1898_1 & ~n1929;
  assign n2339 = n2141 & n2338_1;
  assign n2340 = n2316 & n2339;
  assign n2341 = n2337 & ~n2340;
  assign n2342_1 = ~n2100 & n2111;
  assign n2343 = n1929 & n2342_1;
  assign n2344 = n2066 & n2343;
  assign n2345 = STATE2_REG_0_ & n2344;
  assign n2346 = n1994 & n2066;
  assign n2347_1 = n1929 & ~n2346;
  assign n2348 = ~n1898_1 & n1994;
  assign n2349 = n1898_1 & ~n2066;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = n2100 & n2350;
  assign n2352_1 = ~n1839 & ~n2069;
  assign n2353 = ~n2347_1 & ~n2351;
  assign n2354 = ~n2352_1 & n2353;
  assign n2355 = n2144 & ~n2354;
  assign n2356 = ~n2066 & n2067;
  assign n2357_1 = n2315 & n2356;
  assign n2358 = n2144 & n2357_1;
  assign n2359 = ~n2333_1 & ~n2345;
  assign n2360 = ~n2355 & n2359;
  assign n2361 = ~n2358 & n2360;
  assign n2362_1 = n2066 & ~n2348;
  assign n2363 = ~n2067 & n2362_1;
  assign n2364 = ~n2100 & ~n2363;
  assign n2365 = n2144 & n2364;
  assign n2366_1 = n1776 & ~n2264;
  assign n2367 = ~n2100 & ~n2366_1;
  assign n2368 = ~n1967 & ~n1970;
  assign n2369 = ~n1964 & n2368;
  assign n2370_1 = ~n1973_1 & ~n1979;
  assign n2371 = ~n1982 & n2370_1;
  assign n2372 = ~n1987 & n2371;
  assign n2373 = n1992 & n2369;
  assign n2374 = n2372 & n2373;
  assign n2375_1 = n1898_1 & ~n2374;
  assign n2376 = ~n1929 & n2066;
  assign n2377 = ~n2348 & ~n2375_1;
  assign n2378 = n2376 & n2377;
  assign n2379_1 = n2152 & ~n2378;
  assign n2380 = ~n2367 & ~n2379_1;
  assign n2381 = STATE2_REG_0_ & ~n2380;
  assign n2382 = n2107 & n2264;
  assign n2383 = STATE2_REG_0_ & n2382;
  assign n2384_1 = n1807 & n2100;
  assign n2385 = n1994 & n2384_1;
  assign n2386 = n1776 & n2385;
  assign n2387 = n1839 & n2386;
  assign n2388 = ~n2066 & n2338_1;
  assign n2389 = n2387 & n2388;
  assign n2390 = STATE2_REG_0_ & n2389;
  assign n2391 = ~n2365 & ~n2381;
  assign n2392 = ~n2383 & n2391;
  assign n2393 = ~n2390 & n2392;
  assign n2394 = STATE2_REG_0_ & n2265;
  assign n2395 = n1898_1 & ~n1994;
  assign n2396 = ~n2066 & ~n2395;
  assign n2397 = n1898_1 & n2147;
  assign n2398 = ~n1929 & ~n2348;
  assign n2399 = ~n2397 & n2398;
  assign n2400 = ~n2396 & n2399;
  assign n2401 = n2394 & ~n2400;
  assign n2402 = ~n1776 & n1839;
  assign n2403 = STATE2_REG_0_ & n2402;
  assign n2404 = ~n2336 & ~n2403;
  assign n2405 = ~STATE2_REG_3_ & ~STATE2_REG_1_;
  assign n2406 = ~STATE2_REG_0_ & n2405;
  assign n2407 = ~INSTQUEUEWR_ADDR_REG_1_ & INSTQUEUEWR_ADDR_REG_0_;
  assign n2408 = INSTQUEUEWR_ADDR_REG_1_ & ~INSTQUEUEWR_ADDR_REG_0_;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = n2406 & ~n2409;
  assign n2411 = STATE2_REG_2_ & ~STATE2_REG_1_;
  assign n2412 = INSTQUEUEWR_ADDR_REG_1_ & ~n2411;
  assign n2413 = ~n2410 & ~n2412;
  assign n2414 = n1929 & n2066;
  assign n2415 = n2348 & n2414;
  assign n2416 = n2316 & n2415;
  assign n2417 = STATE2_REG_0_ & n2416;
  assign n2418 = n2066 & n2338_1;
  assign n2419 = n2387 & n2418;
  assign n2420 = STATE2_REG_0_ & n2419;
  assign n2421 = n2413 & ~n2417;
  assign n2422 = ~n2420 & n2421;
  assign n2423 = ~n2145 & ~n2401;
  assign n2424 = n2404 & n2423;
  assign n2425 = n2422 & n2424;
  assign n2426 = n2361 & n2393;
  assign n2427 = n2425 & n2426;
  assign n2428 = ~INSTQUEUERD_ADDR_REG_1_ & ~n2412;
  assign n2429 = ~n2410 & n2428;
  assign n2430 = ~n2427 & ~n2429;
  assign n2431 = ~n2341 & n2430;
  assign n2432 = n2354 & ~n2364;
  assign n2433 = n1807 & ~n2432;
  assign n2434 = ~n1807 & ~n2147;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = n1776 & ~n2435;
  assign n2437 = ~n1776 & ~n2100;
  assign n2438 = STATE2_REG_0_ & n2405;
  assign n2439 = n2066 & ~n2395;
  assign n2440 = n2280 & n2439;
  assign n2441 = ~n2348 & n2440;
  assign n2442 = n2152 & ~n2441;
  assign n2443 = n2438 & ~n2442;
  assign n2444 = ~n2356 & ~n2415;
  assign n2445 = n2316 & ~n2444;
  assign n2446 = n1839 & n2344;
  assign n2447 = ~n2382 & ~n2445;
  assign n2448 = ~n2446 & n2447;
  assign n2449 = ~n1776 & ~n2315;
  assign n2450 = n2400 & n2449;
  assign n2451 = ~n1807 & ~n2450;
  assign n2452 = n2448 & ~n2451;
  assign n2453 = ~n2436 & ~n2437;
  assign n2454 = n2443 & n2453;
  assign n2455 = n2452 & n2454;
  assign n2456 = ~n2401 & ~n2403;
  assign n2457 = ~n2357_1 & ~n2364;
  assign n2458 = n2354 & n2457;
  assign n2459 = n2144 & ~n2458;
  assign n2460 = ~n2145 & ~n2417;
  assign n2461 = ~n2420 & n2460;
  assign n2462 = INSTQUEUEWR_ADDR_REG_0_ & ~n2411;
  assign n2463 = ~INSTQUEUEWR_ADDR_REG_0_ & n2406;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = ~n2345 & ~n2383;
  assign n2466 = ~n2390 & n2465;
  assign n2467 = ~n2381 & n2464;
  assign n2468 = n2337 & n2467;
  assign n2469 = n2466 & n2468;
  assign n2470 = n2456 & ~n2459;
  assign n2471 = n2461 & n2470;
  assign n2472 = n2469 & n2471;
  assign n2473 = ~INSTQUEUERD_ADDR_REG_0_ & n2464;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = ~n2455 & n2474;
  assign n2476 = n2341 & ~n2430;
  assign n2477 = n2475 & ~n2476;
  assign n2478 = ~n2431 & ~n2477;
  assign n2479 = INSTQUEUEWR_ADDR_REG_1_ & INSTQUEUEWR_ADDR_REG_0_;
  assign n2480 = ~INSTQUEUEWR_ADDR_REG_2_ & n2479;
  assign n2481 = INSTQUEUEWR_ADDR_REG_2_ & ~n2479;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = n2406 & ~n2482;
  assign n2484 = INSTQUEUEWR_ADDR_REG_2_ & ~n2411;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = n2337 & ~n2381;
  assign n2487 = n2466 & n2486;
  assign n2488 = n2471 & n2487;
  assign n2489 = n2485 & n2488;
  assign n2490 = ~INSTQUEUERD_ADDR_REG_2_ & ~n2484;
  assign n2491 = ~n2483 & n2490;
  assign n2492 = ~n2489 & ~n2491;
  assign n2493 = n2478 & ~n2492;
  assign n2494 = ~n2478 & n2492;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2387 & ~n2446;
  assign n2497 = ~n1807 & n1929;
  assign n2498 = ~n2416 & ~n2497;
  assign n2499 = ~n2268_1 & ~n2382;
  assign n2500 = n2496 & n2499;
  assign n2501 = n2498 & n2500;
  assign n2502 = ~n2282 & n2501;
  assign n2503 = n2264 & ~n2399;
  assign n2504 = ~n2395 & n2398;
  assign n2505 = n2152 & ~n2504;
  assign n2506 = ~n2402 & ~n2505;
  assign n2507 = n1898_1 & ~n2100;
  assign n2508 = ~n2316 & ~n2507;
  assign n2509 = ~n1807 & ~n2508;
  assign n2510 = n2198_1 & ~n2395;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = ~n2367 & ~n2503;
  assign n2513 = n2506 & n2512;
  assign n2514 = n2511 & n2513;
  assign n2515 = ~n2436 & n2514;
  assign n2516 = n2502 & n2515;
  assign n2517 = n2495 & ~n2516;
  assign n2518 = n2327 & ~n2517;
  assign n2519 = ~READY_N & n2149;
  assign n2520 = n2282 & n2519;
  assign n2521 = ~n2102 & ~n2520;
  assign n2522 = ~READY_N & n2293_1;
  assign n2523 = ~n2109 & ~n2282;
  assign n2524 = n2522 & ~n2523;
  assign n2525 = n2521 & ~n2524;
  assign n2526 = ~n2262 & ~n2525;
  assign n2527 = n2262 & n2266;
  assign n2528 = n2100 & n2103_1;
  assign n2529 = ~n2510 & ~n2528;
  assign n2530 = ~READY_N & n2268_1;
  assign n2531 = n2272 & n2530;
  assign n2532 = n2529 & ~n2531;
  assign n2533 = n1776 & n1839;
  assign n2534 = n2107 & n2533;
  assign n2535 = ~n2100 & ~n2534;
  assign n2536 = n1776 & ~n2069;
  assign n2537 = ~n1839 & ~n2536;
  assign n2538 = n2399 & n2537;
  assign n2539 = n2100 & ~n2538;
  assign n2540 = ~n2535 & ~n2539;
  assign n2541 = ~n2505 & n2540;
  assign n2542 = n2532 & n2541;
  assign n2543 = ~n2526 & ~n2527;
  assign n2544 = n2542 & n2543;
  assign n2545 = ~n2518 & ~n2544;
  assign n2546 = INSTQUEUERD_ADDR_REG_2_ & n2544;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = ~STATE2_REG_1_ & ~n2547;
  assign n2549 = n2314 & ~n2548;
  assign n2550 = INSTQUEUERD_ADDR_REG_4_ & n2544;
  assign n2551 = STATE2_REG_0_ & n2103_1;
  assign n2552 = n2108_1 & n2551;
  assign n2553 = ~n2336 & ~n2552;
  assign n2554 = INSTQUEUERD_ADDR_REG_4_ & ~n2553;
  assign n2555 = INSTQUEUEWR_ADDR_REG_3_ & ~INSTQUEUEWR_ADDR_REG_2_;
  assign n2556 = INSTQUEUEWR_ADDR_REG_3_ & ~n2479;
  assign n2557 = ~INSTQUEUEWR_ADDR_REG_3_ & INSTQUEUEWR_ADDR_REG_2_;
  assign n2558 = n2479 & n2557;
  assign n2559 = ~n2555 & ~n2556;
  assign n2560 = ~n2558 & n2559;
  assign n2561 = n2406 & ~n2560;
  assign n2562 = INSTQUEUEWR_ADDR_REG_3_ & ~n2411;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = INSTQUEUERD_ADDR_REG_3_ & ~n2488;
  assign n2565 = n2563 & ~n2564;
  assign n2566 = n2492 & ~n2565;
  assign n2567 = ~n2478 & n2566;
  assign n2568 = n2554 & ~n2567;
  assign n2569 = ~n2554 & n2567;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = n2268_1 & ~n2570;
  assign n2572 = ~n2544 & n2571;
  assign n2573 = ~n2550 & ~n2572;
  assign n2574 = ~STATE2_REG_1_ & ~n2573;
  assign n2575 = INSTQUEUERD_ADDR_REG_4_ & n2300;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = n2549 & n2576;
  assign n2578 = n2494 & n2565;
  assign n2579 = ~n2494 & ~n2565;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = ~n2516 & ~n2580;
  assign n2582 = INSTQUEUERD_ADDR_REG_3_ & ~n1742_1;
  assign n2583 = ~n1985 & ~n2582;
  assign n2584 = n2109 & ~n2583;
  assign n2585 = INSTQUEUERD_ADDR_REG_3_ & ~n1768;
  assign n2586 = ~n1769 & ~n2585;
  assign n2587 = n2318_1 & ~n2586;
  assign n2588 = ~n2584 & ~n2587;
  assign n2589 = ~n1753 & n1754_1;
  assign n2590 = ~INSTQUEUERD_ADDR_REG_2_ & ~n1753;
  assign n2591 = INSTQUEUERD_ADDR_REG_3_ & ~n2590;
  assign n2592 = ~n2589 & ~n2591;
  assign n2593 = ~n2322 & n2592;
  assign n2594 = n2588 & ~n2593;
  assign n2595 = ~n2581 & n2594;
  assign n2596 = ~n2544 & ~n2595;
  assign n2597 = INSTQUEUERD_ADDR_REG_3_ & n2544;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = ~STATE2_REG_1_ & ~n2598;
  assign n2600 = INSTQUEUERD_ADDR_REG_3_ & n2300;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = n2576 & n2601;
  assign n2603 = ~n2577 & ~n2602;
  assign n2604 = ~INSTQUEUEWR_ADDR_REG_4_ & ~n2573;
  assign n2605 = INSTQUEUEWR_ADDR_REG_3_ & n2598;
  assign n2606 = INSTQUEUEWR_ADDR_REG_4_ & n2573;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = ~INSTQUEUEWR_ADDR_REG_2_ & ~n2547;
  assign n2609 = ~INSTQUEUEWR_ADDR_REG_3_ & ~n2598;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = n1808 & n2101;
  assign n2612 = ~n2266 & ~n2611;
  assign n2613 = ~INSTQUEUERD_ADDR_REG_0_ & ~n2612;
  assign n2614 = INSTQUEUERD_ADDR_REG_0_ & n2109;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = n2455 & n2474;
  assign n2617 = ~n2455 & ~n2474;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2516 & ~n2618;
  assign n2620 = n2615 & ~n2619;
  assign n2621 = ~n2544 & ~n2620;
  assign n2622 = INSTQUEUERD_ADDR_REG_0_ & n2544;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = n2479 & n2623;
  assign n2625 = INSTQUEUEWR_ADDR_REG_2_ & n2547;
  assign n2626 = ~INSTQUEUERD_ADDR_REG_1_ & n2109;
  assign n2627 = ~n1722_1 & ~n1753;
  assign n2628 = ~n2612 & n2627;
  assign n2629 = ~n2626 & ~n2628;
  assign n2630 = ~n2431 & ~n2476;
  assign n2631 = ~n2475 & n2630;
  assign n2632 = n2475 & ~n2630;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = ~n2516 & ~n2633;
  assign n2635 = n2629 & ~n2634;
  assign n2636 = ~n2544 & ~n2635;
  assign n2637 = INSTQUEUERD_ADDR_REG_1_ & n2544;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = INSTQUEUEWR_ADDR_REG_1_ & n2638;
  assign n2640 = n2623 & n2638;
  assign n2641 = INSTQUEUEWR_ADDR_REG_0_ & n2640;
  assign n2642 = ~n2624 & ~n2625;
  assign n2643 = ~n2639 & n2642;
  assign n2644 = ~n2641 & n2643;
  assign n2645 = n2610 & ~n2644;
  assign n2646 = n2607 & ~n2645;
  assign n2647 = ~n2604 & ~n2646;
  assign n2648 = ~n2276 & ~n2278_1;
  assign n2649 = ~n2299 & n2648;
  assign n2650 = ~n2603 & n2649;
  assign n2651 = n2647 & n2650;
  assign n2652 = ~STATE2_REG_1_ & n2651;
  assign n2653 = STATE2_REG_0_ & ~n2652;
  assign n2654 = ~READY_N & ~STATEBS16_REG;
  assign n2655 = n2152 & n2654;
  assign n2656 = ~n2262 & n2293_1;
  assign n2657 = n2282 & n2655;
  assign n2658 = n2656 & n2657;
  assign n2659 = STATE2_REG_2_ & ~n2658;
  assign n2660 = ~n1709 & ~n2653;
  assign n2661 = n2659 & n2660;
  assign n2662 = STATE2_REG_0_ & ~n2661;
  assign n2663 = n1707 & n2662;
  assign n2664 = STATE2_REG_3_ & ~n2662;
  assign n525 = n2663 | n2664;
  assign n2666 = ~READY_N & ~STATE2_REG_2_;
  assign n2667 = STATE2_REG_0_ & ~n2666;
  assign n2668 = ~STATE2_REG_0_ & ~STATEBS16_REG;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = STATE2_REG_1_ & n2669;
  assign n2671 = ~n2411 & ~n2670;
  assign n2672 = STATE2_REG_2_ & ~n2662;
  assign n530 = ~n2671 | n2672;
  assign n2674 = STATE2_REG_0_ & n2411;
  assign n2675 = ~n2661 & n2674;
  assign n2676 = READY_N & ~STATE2_REG_2_;
  assign n2677 = STATE2_REG_0_ & n2676;
  assign n2678 = ~n2661 & ~n2677;
  assign n2679 = STATE2_REG_1_ & ~n2678;
  assign n2680 = ~READY_N & n2405;
  assign n2681 = n2662 & n2680;
  assign n2682 = ~STATE2_REG_2_ & ~STATEBS16_REG;
  assign n2683 = STATE2_REG_1_ & ~STATE2_REG_0_;
  assign n2684 = n2682 & n2683;
  assign n2685 = ~n2675 & ~n2679;
  assign n2686 = ~n2681 & n2685;
  assign n535 = n2684 | ~n2686;
  assign n2688 = STATE2_REG_3_ & ~n2262;
  assign n2689 = ~STATE2_REG_2_ & ~STATE2_REG_1_;
  assign n2690 = n2688 & n2689;
  assign n2691 = ~n2661 & ~n2690;
  assign n2692 = ~STATE2_REG_0_ & n2691;
  assign n2693 = FLUSH_REG & n2304;
  assign n2694 = STATE2_REG_1_ & n2693;
  assign n2695 = ~STATE2_REG_1_ & ~n2623;
  assign n2696 = INSTQUEUERD_ADDR_REG_0_ & n2300;
  assign n2697 = ~n2694 & ~n2695;
  assign n2698 = ~n2696 & n2697;
  assign n2699 = INSTQUEUERD_ADDR_REG_1_ & n2300;
  assign n2700 = n2311 & n2312;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = ~STATE2_REG_1_ & ~n2638;
  assign n2703 = n2701 & ~n2702;
  assign n2704 = n2698 & n2703;
  assign n2705 = ~n2549 & ~n2704;
  assign n2706 = ~n2601 & n2705;
  assign n2707 = n2576 & ~n2706;
  assign n2708 = n1707 & n2707;
  assign n2709 = ~n2661 & ~n2708;
  assign n2710 = STATE2_REG_0_ & ~n2709;
  assign n2711 = STATE2_REG_3_ & STATE2_REG_0_;
  assign n2712 = n2689 & n2711;
  assign n2713 = ~n2677 & ~n2712;
  assign n2714 = ~n2651 & n2674;
  assign n2715 = n2713 & ~n2714;
  assign n2716 = ~n2692 & ~n2710;
  assign n540 = ~n2715 | ~n2716;
  assign n2718 = INSTQUEUEWR_ADDR_REG_3_ & INSTQUEUEWR_ADDR_REG_2_;
  assign n2719 = n2479 & n2718;
  assign n2720 = n2495 & ~n2580;
  assign n2721 = ~n2618 & ~n2633;
  assign n2722 = n2720 & n2721;
  assign n2723 = ~n2719 & ~n2722;
  assign n2724 = ~STATE2_REG_3_ & ~STATE2_REG_2_;
  assign n2725 = ~STATEBS16_REG & n2724;
  assign n2726 = n2320 & n2586;
  assign n2727 = INSTQUEUERD_ADDR_REG_0_ & ~n2627;
  assign n2728 = n2726 & n2727;
  assign n2729 = INSTQUEUE_REG_0__7_ & n2728;
  assign n2730 = ~INSTQUEUERD_ADDR_REG_0_ & ~n2627;
  assign n2731 = n2726 & n2730;
  assign n2732 = INSTQUEUE_REG_1__7_ & n2731;
  assign n2733 = INSTQUEUERD_ADDR_REG_0_ & n2627;
  assign n2734 = n2726 & n2733;
  assign n2735 = INSTQUEUE_REG_2__7_ & n2734;
  assign n2736 = ~INSTQUEUERD_ADDR_REG_0_ & n2627;
  assign n2737 = n2726 & n2736;
  assign n2738 = INSTQUEUE_REG_3__7_ & n2737;
  assign n2739 = ~n2729 & ~n2732;
  assign n2740 = ~n2735 & n2739;
  assign n2741 = ~n2738 & n2740;
  assign n2742 = ~n2320 & n2586;
  assign n2743 = n2727 & n2742;
  assign n2744 = INSTQUEUE_REG_4__7_ & n2743;
  assign n2745 = n2730 & n2742;
  assign n2746 = INSTQUEUE_REG_5__7_ & n2745;
  assign n2747 = n2733 & n2742;
  assign n2748 = INSTQUEUE_REG_6__7_ & n2747;
  assign n2749 = n2736 & n2742;
  assign n2750 = INSTQUEUE_REG_7__7_ & n2749;
  assign n2751 = ~n2744 & ~n2746;
  assign n2752 = ~n2748 & n2751;
  assign n2753 = ~n2750 & n2752;
  assign n2754 = n2320 & ~n2586;
  assign n2755 = n2727 & n2754;
  assign n2756 = INSTQUEUE_REG_8__7_ & n2755;
  assign n2757 = n2730 & n2754;
  assign n2758 = INSTQUEUE_REG_9__7_ & n2757;
  assign n2759 = n2733 & n2754;
  assign n2760 = INSTQUEUE_REG_10__7_ & n2759;
  assign n2761 = n2736 & n2754;
  assign n2762 = INSTQUEUE_REG_11__7_ & n2761;
  assign n2763 = ~n2756 & ~n2758;
  assign n2764 = ~n2760 & n2763;
  assign n2765 = ~n2762 & n2764;
  assign n2766 = ~n2320 & ~n2586;
  assign n2767 = n2727 & n2766;
  assign n2768 = INSTQUEUE_REG_12__7_ & n2767;
  assign n2769 = n2730 & n2766;
  assign n2770 = INSTQUEUE_REG_13__7_ & n2769;
  assign n2771 = n2733 & n2766;
  assign n2772 = INSTQUEUE_REG_14__7_ & n2771;
  assign n2773 = n2736 & n2766;
  assign n2774 = INSTQUEUE_REG_15__7_ & n2773;
  assign n2775 = ~n2768 & ~n2770;
  assign n2776 = ~n2772 & n2775;
  assign n2777 = ~n2774 & n2776;
  assign n2778 = n2741 & n2753;
  assign n2779 = n2765 & n2778;
  assign n2780 = n2777 & n2779;
  assign n2781 = n2218_1 & ~n2780;
  assign n2782 = ~STATE2_REG_0_ & ~n2618;
  assign n2783 = n2218_1 & n2780;
  assign n2784 = INSTQUEUE_REG_0__0_ & n2728;
  assign n2785 = INSTQUEUE_REG_1__0_ & n2731;
  assign n2786 = INSTQUEUE_REG_2__0_ & n2734;
  assign n2787 = INSTQUEUE_REG_3__0_ & n2737;
  assign n2788 = ~n2784 & ~n2785;
  assign n2789 = ~n2786 & n2788;
  assign n2790 = ~n2787 & n2789;
  assign n2791 = INSTQUEUE_REG_4__0_ & n2743;
  assign n2792 = INSTQUEUE_REG_5__0_ & n2745;
  assign n2793 = INSTQUEUE_REG_6__0_ & n2747;
  assign n2794 = INSTQUEUE_REG_7__0_ & n2749;
  assign n2795 = ~n2791 & ~n2792;
  assign n2796 = ~n2793 & n2795;
  assign n2797 = ~n2794 & n2796;
  assign n2798 = INSTQUEUE_REG_8__0_ & n2755;
  assign n2799 = INSTQUEUE_REG_9__0_ & n2757;
  assign n2800 = INSTQUEUE_REG_10__0_ & n2759;
  assign n2801 = INSTQUEUE_REG_11__0_ & n2761;
  assign n2802 = ~n2798 & ~n2799;
  assign n2803 = ~n2800 & n2802;
  assign n2804 = ~n2801 & n2803;
  assign n2805 = INSTQUEUE_REG_12__0_ & n2767;
  assign n2806 = INSTQUEUE_REG_13__0_ & n2769;
  assign n2807 = INSTQUEUE_REG_14__0_ & n2771;
  assign n2808 = INSTQUEUE_REG_15__0_ & n2773;
  assign n2809 = ~n2805 & ~n2806;
  assign n2810 = ~n2807 & n2809;
  assign n2811 = ~n2808 & n2810;
  assign n2812 = n2790 & n2797;
  assign n2813 = n2804 & n2812;
  assign n2814 = n2811 & n2813;
  assign n2815 = n2783 & ~n2814;
  assign n2816 = n2781 & n2814;
  assign n2817 = ~n2782 & ~n2815;
  assign n2818 = ~n2816 & n2817;
  assign n2819 = ~n2781 & ~n2818;
  assign n2820 = n2781 & n2818;
  assign n2821 = INSTQUEUE_REG_0__0_ & n2138_1;
  assign n2822 = STATE2_REG_0_ & ~n2821;
  assign n2823 = n2143_1 & ~n2814;
  assign n2824 = n2066 & ~n2780;
  assign n2825 = n2822 & ~n2823;
  assign n2826 = ~n2824 & n2825;
  assign n2827 = ~n2819 & ~n2820;
  assign n2828 = n2826 & n2827;
  assign n2829 = n2781 & ~n2828;
  assign n2830 = ~n2826 & ~n2827;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = ~STATE2_REG_0_ & ~n2633;
  assign n2833 = INSTQUEUE_REG_0__1_ & n2728;
  assign n2834 = INSTQUEUE_REG_1__1_ & n2731;
  assign n2835 = INSTQUEUE_REG_2__1_ & n2734;
  assign n2836 = INSTQUEUE_REG_3__1_ & n2737;
  assign n2837 = ~n2833 & ~n2834;
  assign n2838 = ~n2835 & n2837;
  assign n2839 = ~n2836 & n2838;
  assign n2840 = INSTQUEUE_REG_4__1_ & n2743;
  assign n2841 = INSTQUEUE_REG_5__1_ & n2745;
  assign n2842 = INSTQUEUE_REG_6__1_ & n2747;
  assign n2843 = INSTQUEUE_REG_7__1_ & n2749;
  assign n2844 = ~n2840 & ~n2841;
  assign n2845 = ~n2842 & n2844;
  assign n2846 = ~n2843 & n2845;
  assign n2847 = INSTQUEUE_REG_8__1_ & n2755;
  assign n2848 = INSTQUEUE_REG_9__1_ & n2757;
  assign n2849 = INSTQUEUE_REG_10__1_ & n2759;
  assign n2850 = INSTQUEUE_REG_11__1_ & n2761;
  assign n2851 = ~n2847 & ~n2848;
  assign n2852 = ~n2849 & n2851;
  assign n2853 = ~n2850 & n2852;
  assign n2854 = INSTQUEUE_REG_12__1_ & n2767;
  assign n2855 = INSTQUEUE_REG_13__1_ & n2769;
  assign n2856 = INSTQUEUE_REG_14__1_ & n2771;
  assign n2857 = INSTQUEUE_REG_15__1_ & n2773;
  assign n2858 = ~n2854 & ~n2855;
  assign n2859 = ~n2856 & n2858;
  assign n2860 = ~n2857 & n2859;
  assign n2861 = n2839 & n2846;
  assign n2862 = n2853 & n2861;
  assign n2863 = n2860 & n2862;
  assign n2864 = n2783 & ~n2863;
  assign n2865 = n2781 & n2863;
  assign n2866 = ~n2832 & ~n2864;
  assign n2867 = ~n2865 & n2866;
  assign n2868 = ~n2781 & ~n2867;
  assign n2869 = n2781 & n2867;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = INSTQUEUE_REG_0__1_ & n2138_1;
  assign n2872 = ~n2783 & ~n2871;
  assign n2873 = n2143_1 & ~n2863;
  assign n2874 = n2872 & ~n2873;
  assign n2875 = ~n2870 & n2874;
  assign n2876 = n2870 & ~n2874;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = n2831 & ~n2877;
  assign n2879 = ~n2831 & n2877;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = ~n2828 & ~n2830;
  assign n2882 = ~n2781 & n2881;
  assign n2883 = n2781 & ~n2881;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~n2880 & n2884;
  assign n2886 = n2880 & ~n2884;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = n2884 & ~n2887;
  assign n2889 = ~n2880 & ~n2884;
  assign n2890 = INSTQUEUE_REG_0__2_ & n2138_1;
  assign n2891 = INSTQUEUE_REG_0__2_ & n2728;
  assign n2892 = INSTQUEUE_REG_1__2_ & n2731;
  assign n2893 = INSTQUEUE_REG_2__2_ & n2734;
  assign n2894 = INSTQUEUE_REG_3__2_ & n2737;
  assign n2895 = ~n2891 & ~n2892;
  assign n2896 = ~n2893 & n2895;
  assign n2897 = ~n2894 & n2896;
  assign n2898 = INSTQUEUE_REG_4__2_ & n2743;
  assign n2899 = INSTQUEUE_REG_5__2_ & n2745;
  assign n2900 = INSTQUEUE_REG_6__2_ & n2747;
  assign n2901 = INSTQUEUE_REG_7__2_ & n2749;
  assign n2902 = ~n2898 & ~n2899;
  assign n2903 = ~n2900 & n2902;
  assign n2904 = ~n2901 & n2903;
  assign n2905 = INSTQUEUE_REG_8__2_ & n2755;
  assign n2906 = INSTQUEUE_REG_9__2_ & n2757;
  assign n2907 = INSTQUEUE_REG_10__2_ & n2759;
  assign n2908 = INSTQUEUE_REG_11__2_ & n2761;
  assign n2909 = ~n2905 & ~n2906;
  assign n2910 = ~n2907 & n2909;
  assign n2911 = ~n2908 & n2910;
  assign n2912 = INSTQUEUE_REG_12__2_ & n2767;
  assign n2913 = INSTQUEUE_REG_13__2_ & n2769;
  assign n2914 = INSTQUEUE_REG_14__2_ & n2771;
  assign n2915 = INSTQUEUE_REG_15__2_ & n2773;
  assign n2916 = ~n2912 & ~n2913;
  assign n2917 = ~n2914 & n2916;
  assign n2918 = ~n2915 & n2917;
  assign n2919 = n2897 & n2904;
  assign n2920 = n2911 & n2919;
  assign n2921 = n2918 & n2920;
  assign n2922 = n2143_1 & ~n2921;
  assign n2923 = ~n2890 & ~n2922;
  assign n2924 = n2781 & n2921;
  assign n2925 = n2783 & ~n2921;
  assign n2926 = ~STATE2_REG_0_ & n2495;
  assign n2927 = ~n2924 & ~n2925;
  assign n2928 = ~n2926 & n2927;
  assign n2929 = ~n2781 & ~n2928;
  assign n2930 = n2781 & n2928;
  assign n2931 = ~n2929 & ~n2930;
  assign n2932 = ~n2923 & ~n2931;
  assign n2933 = n2923 & n2931;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~n2870 & ~n2874;
  assign n2936 = n2870 & n2874;
  assign n2937 = ~n2831 & ~n2936;
  assign n2938 = ~n2935 & ~n2937;
  assign n2939 = n2934 & n2938;
  assign n2940 = ~n2934 & ~n2938;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n2889 & n2941;
  assign n2943 = ~n2889 & ~n2941;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2933 & ~n2938;
  assign n2946 = INSTQUEUE_REG_0__3_ & n2138_1;
  assign n2947 = INSTQUEUE_REG_0__3_ & n2728;
  assign n2948 = INSTQUEUE_REG_1__3_ & n2731;
  assign n2949 = INSTQUEUE_REG_2__3_ & n2734;
  assign n2950 = INSTQUEUE_REG_3__3_ & n2737;
  assign n2951 = ~n2947 & ~n2948;
  assign n2952 = ~n2949 & n2951;
  assign n2953 = ~n2950 & n2952;
  assign n2954 = INSTQUEUE_REG_4__3_ & n2743;
  assign n2955 = INSTQUEUE_REG_5__3_ & n2745;
  assign n2956 = INSTQUEUE_REG_6__3_ & n2747;
  assign n2957 = INSTQUEUE_REG_7__3_ & n2749;
  assign n2958 = ~n2954 & ~n2955;
  assign n2959 = ~n2956 & n2958;
  assign n2960 = ~n2957 & n2959;
  assign n2961 = INSTQUEUE_REG_8__3_ & n2755;
  assign n2962 = INSTQUEUE_REG_9__3_ & n2757;
  assign n2963 = INSTQUEUE_REG_10__3_ & n2759;
  assign n2964 = INSTQUEUE_REG_11__3_ & n2761;
  assign n2965 = ~n2961 & ~n2962;
  assign n2966 = ~n2963 & n2965;
  assign n2967 = ~n2964 & n2966;
  assign n2968 = INSTQUEUE_REG_12__3_ & n2767;
  assign n2969 = INSTQUEUE_REG_13__3_ & n2769;
  assign n2970 = INSTQUEUE_REG_14__3_ & n2771;
  assign n2971 = INSTQUEUE_REG_15__3_ & n2773;
  assign n2972 = ~n2968 & ~n2969;
  assign n2973 = ~n2970 & n2972;
  assign n2974 = ~n2971 & n2973;
  assign n2975 = n2953 & n2960;
  assign n2976 = n2967 & n2975;
  assign n2977 = n2974 & n2976;
  assign n2978 = n2143_1 & ~n2977;
  assign n2979 = ~n2946 & ~n2978;
  assign n2980 = n2781 & n2977;
  assign n2981 = n2783 & ~n2977;
  assign n2982 = ~STATE2_REG_0_ & ~n2580;
  assign n2983 = ~n2980 & ~n2981;
  assign n2984 = ~n2982 & n2983;
  assign n2985 = ~n2781 & ~n2984;
  assign n2986 = n2781 & n2984;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2979 & ~n2987;
  assign n2989 = n2979 & n2987;
  assign n2990 = ~n2988 & ~n2989;
  assign n2991 = ~n2932 & ~n2945;
  assign n2992 = ~n2990 & n2991;
  assign n2993 = n2990 & ~n2991;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n2941 & n2994;
  assign n2996 = ~n2889 & n2994;
  assign n2997 = ~n2941 & ~n2994;
  assign n2998 = n2889 & n2997;
  assign n2999 = ~n2995 & ~n2996;
  assign n3000 = ~n2998 & n2999;
  assign n3001 = ~n2944 & ~n3000;
  assign n3002 = n2888 & n3001;
  assign n3003 = ~n2941 & n2994;
  assign n3004 = n2889 & n3003;
  assign n3005 = ~n3002 & ~n3004;
  assign n3006 = STATEBS16_REG & n2724;
  assign n3007 = ~STATE2_REG_2_ & STATE2_REG_1_;
  assign n3008 = ~n2411 & ~n3007;
  assign n3009 = ~n2688 & n3008;
  assign n3010 = ~STATE2_REG_0_ & ~n3009;
  assign n3011 = n3006 & n3010;
  assign n3012 = n3005 & n3011;
  assign n3013 = ~n2725 & ~n3012;
  assign n3014 = n2723 & ~n3013;
  assign n3015 = STATE2_REG_3_ & ~n2719;
  assign n3016 = ~n2482 & ~n2560;
  assign n3017 = ~INSTQUEUEWR_ADDR_REG_0_ & ~n2409;
  assign n3018 = n3016 & n3017;
  assign n3019 = ~n2719 & ~n3018;
  assign n3020 = STATE2_REG_2_ & n3019;
  assign n3021 = ~n3015 & ~n3020;
  assign n3022 = n3010 & n3021;
  assign n3023 = ~n3014 & n3022;
  assign n3024 = INSTQUEUE_REG_15__7_ & ~n3023;
  assign n3025 = DATAI_7_ & n3010;
  assign n3026 = STATE2_REG_2_ & ~n3019;
  assign n3027 = n3005 & n3006;
  assign n3028 = ~n2725 & ~n3027;
  assign n3029 = ~n2723 & ~n3028;
  assign n3030 = ~n3026 & ~n3029;
  assign n3031 = n3025 & ~n3030;
  assign n3032 = DATAI_23_ & n3011;
  assign n3033 = n3004 & n3032;
  assign n3034 = STATE2_REG_3_ & n3010;
  assign n3035 = ~n1929 & n3034;
  assign n3036 = n2719 & n3035;
  assign n3037 = DATAI_31_ & n3011;
  assign n3038 = n3002 & n3037;
  assign n3039 = ~n3033 & ~n3036;
  assign n3040 = ~n3038 & n3039;
  assign n3041 = ~n3024 & ~n3031;
  assign n545 = ~n3040 | ~n3041;
  assign n3043 = INSTQUEUE_REG_15__6_ & ~n3023;
  assign n3044 = DATAI_6_ & n3010;
  assign n3045 = ~n3030 & n3044;
  assign n3046 = DATAI_22_ & n3011;
  assign n3047 = n3004 & n3046;
  assign n3048 = ~n1898_1 & n3034;
  assign n3049 = n2719 & n3048;
  assign n3050 = DATAI_30_ & n3011;
  assign n3051 = n3002 & n3050;
  assign n3052 = ~n3047 & ~n3049;
  assign n3053 = ~n3051 & n3052;
  assign n3054 = ~n3043 & ~n3045;
  assign n550 = ~n3053 | ~n3054;
  assign n3056 = INSTQUEUE_REG_15__5_ & ~n3023;
  assign n3057 = DATAI_5_ & n3010;
  assign n3058 = ~n3030 & n3057;
  assign n3059 = DATAI_21_ & n3011;
  assign n3060 = n3004 & n3059;
  assign n3061 = ~n1994 & n3034;
  assign n3062 = n2719 & n3061;
  assign n3063 = DATAI_29_ & n3011;
  assign n3064 = n3002 & n3063;
  assign n3065 = ~n3060 & ~n3062;
  assign n3066 = ~n3064 & n3065;
  assign n3067 = ~n3056 & ~n3058;
  assign n555 = ~n3066 | ~n3067;
  assign n3069 = INSTQUEUE_REG_15__4_ & ~n3023;
  assign n3070 = DATAI_4_ & n3010;
  assign n3071 = ~n3030 & n3070;
  assign n3072 = DATAI_20_ & n3011;
  assign n3073 = n3004 & n3072;
  assign n3074 = ~n2066 & n3034;
  assign n3075 = n2719 & n3074;
  assign n3076 = DATAI_28_ & n3011;
  assign n3077 = n3002 & n3076;
  assign n3078 = ~n3073 & ~n3075;
  assign n3079 = ~n3077 & n3078;
  assign n3080 = ~n3069 & ~n3071;
  assign n560 = ~n3079 | ~n3080;
  assign n3082 = INSTQUEUE_REG_15__3_ & ~n3023;
  assign n3083 = DATAI_3_ & n3010;
  assign n3084 = ~n3030 & n3083;
  assign n3085 = DATAI_19_ & n3011;
  assign n3086 = n3004 & n3085;
  assign n3087 = ~n1839 & n3034;
  assign n3088 = n2719 & n3087;
  assign n3089 = DATAI_27_ & n3011;
  assign n3090 = n3002 & n3089;
  assign n3091 = ~n3086 & ~n3088;
  assign n3092 = ~n3090 & n3091;
  assign n3093 = ~n3082 & ~n3084;
  assign n565 = ~n3092 | ~n3093;
  assign n3095 = INSTQUEUE_REG_15__2_ & ~n3023;
  assign n3096 = DATAI_2_ & n3010;
  assign n3097 = ~n3030 & n3096;
  assign n3098 = DATAI_18_ & n3011;
  assign n3099 = n3004 & n3098;
  assign n3100 = ~n2100 & n3034;
  assign n3101 = n2719 & n3100;
  assign n3102 = DATAI_26_ & n3011;
  assign n3103 = n3002 & n3102;
  assign n3104 = ~n3099 & ~n3101;
  assign n3105 = ~n3103 & n3104;
  assign n3106 = ~n3095 & ~n3097;
  assign n570 = ~n3105 | ~n3106;
  assign n3108 = INSTQUEUE_REG_15__1_ & ~n3023;
  assign n3109 = DATAI_1_ & n3010;
  assign n3110 = ~n3030 & n3109;
  assign n3111 = DATAI_17_ & n3011;
  assign n3112 = n3004 & n3111;
  assign n3113 = ~n1807 & n3034;
  assign n3114 = n2719 & n3113;
  assign n3115 = DATAI_25_ & n3011;
  assign n3116 = n3002 & n3115;
  assign n3117 = ~n3112 & ~n3114;
  assign n3118 = ~n3116 & n3117;
  assign n3119 = ~n3108 & ~n3110;
  assign n575 = ~n3118 | ~n3119;
  assign n3121 = INSTQUEUE_REG_15__0_ & ~n3023;
  assign n3122 = DATAI_0_ & n3010;
  assign n3123 = ~n3030 & n3122;
  assign n3124 = DATAI_16_ & n3011;
  assign n3125 = n3004 & n3124;
  assign n3126 = ~n1776 & n3034;
  assign n3127 = n2719 & n3126;
  assign n3128 = DATAI_24_ & n3011;
  assign n3129 = n3002 & n3128;
  assign n3130 = ~n3125 & ~n3127;
  assign n3131 = ~n3129 & n3130;
  assign n3132 = ~n3121 & ~n3123;
  assign n580 = ~n3131 | ~n3132;
  assign n3134 = n2408 & n2718;
  assign n3135 = n2618 & ~n2633;
  assign n3136 = n2720 & n3135;
  assign n3137 = ~n3134 & ~n3136;
  assign n3138 = ~n2884 & ~n2887;
  assign n3139 = n3001 & n3138;
  assign n3140 = n2885 & n3003;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = n3011 & n3141;
  assign n3143 = ~n2725 & ~n3142;
  assign n3144 = n3137 & ~n3143;
  assign n3145 = STATE2_REG_3_ & ~n3134;
  assign n3146 = ~n2409 & n3016;
  assign n3147 = STATE2_REG_2_ & ~n3146;
  assign n3148 = ~n3145 & ~n3147;
  assign n3149 = n3010 & n3148;
  assign n3150 = ~n3144 & n3149;
  assign n3151 = INSTQUEUE_REG_14__7_ & ~n3150;
  assign n3152 = STATE2_REG_2_ & n3146;
  assign n3153 = n3006 & n3141;
  assign n3154 = ~n2725 & ~n3153;
  assign n3155 = ~n3137 & ~n3154;
  assign n3156 = ~n3152 & ~n3155;
  assign n3157 = n3025 & ~n3156;
  assign n3158 = n3032 & n3140;
  assign n3159 = n3035 & n3134;
  assign n3160 = n3037 & n3139;
  assign n3161 = ~n3158 & ~n3159;
  assign n3162 = ~n3160 & n3161;
  assign n3163 = ~n3151 & ~n3157;
  assign n585 = ~n3162 | ~n3163;
  assign n3165 = INSTQUEUE_REG_14__6_ & ~n3150;
  assign n3166 = n3044 & ~n3156;
  assign n3167 = n3046 & n3140;
  assign n3168 = n3048 & n3134;
  assign n3169 = n3050 & n3139;
  assign n3170 = ~n3167 & ~n3168;
  assign n3171 = ~n3169 & n3170;
  assign n3172 = ~n3165 & ~n3166;
  assign n590 = ~n3171 | ~n3172;
  assign n3174 = INSTQUEUE_REG_14__5_ & ~n3150;
  assign n3175 = n3057 & ~n3156;
  assign n3176 = n3059 & n3140;
  assign n3177 = n3061 & n3134;
  assign n3178 = n3063 & n3139;
  assign n3179 = ~n3176 & ~n3177;
  assign n3180 = ~n3178 & n3179;
  assign n3181 = ~n3174 & ~n3175;
  assign n595 = ~n3180 | ~n3181;
  assign n3183 = INSTQUEUE_REG_14__4_ & ~n3150;
  assign n3184 = n3070 & ~n3156;
  assign n3185 = n3072 & n3140;
  assign n3186 = n3074 & n3134;
  assign n3187 = n3076 & n3139;
  assign n3188 = ~n3185 & ~n3186;
  assign n3189 = ~n3187 & n3188;
  assign n3190 = ~n3183 & ~n3184;
  assign n600 = ~n3189 | ~n3190;
  assign n3192 = INSTQUEUE_REG_14__3_ & ~n3150;
  assign n3193 = n3083 & ~n3156;
  assign n3194 = n3085 & n3140;
  assign n3195 = n3087 & n3134;
  assign n3196 = n3089 & n3139;
  assign n3197 = ~n3194 & ~n3195;
  assign n3198 = ~n3196 & n3197;
  assign n3199 = ~n3192 & ~n3193;
  assign n605 = ~n3198 | ~n3199;
  assign n3201 = INSTQUEUE_REG_14__2_ & ~n3150;
  assign n3202 = n3096 & ~n3156;
  assign n3203 = n3098 & n3140;
  assign n3204 = n3100 & n3134;
  assign n3205 = n3102 & n3139;
  assign n3206 = ~n3203 & ~n3204;
  assign n3207 = ~n3205 & n3206;
  assign n3208 = ~n3201 & ~n3202;
  assign n610 = ~n3207 | ~n3208;
  assign n3210 = INSTQUEUE_REG_14__1_ & ~n3150;
  assign n3211 = n3109 & ~n3156;
  assign n3212 = n3111 & n3140;
  assign n3213 = n3113 & n3134;
  assign n3214 = n3115 & n3139;
  assign n3215 = ~n3212 & ~n3213;
  assign n3216 = ~n3214 & n3215;
  assign n3217 = ~n3210 & ~n3211;
  assign n615 = ~n3216 | ~n3217;
  assign n3219 = INSTQUEUE_REG_14__0_ & ~n3150;
  assign n3220 = n3122 & ~n3156;
  assign n3221 = n3124 & n3140;
  assign n3222 = n3126 & n3134;
  assign n3223 = n3128 & n3139;
  assign n3224 = ~n3221 & ~n3222;
  assign n3225 = ~n3223 & n3224;
  assign n3226 = ~n3219 & ~n3220;
  assign n620 = ~n3225 | ~n3226;
  assign n3228 = n2407 & n2718;
  assign n3229 = ~n2618 & n2633;
  assign n3230 = n2720 & n3229;
  assign n3231 = ~n3228 & ~n3230;
  assign n3232 = n2884 & n2887;
  assign n3233 = n3001 & n3232;
  assign n3234 = n2886 & n3003;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = n3011 & n3235;
  assign n3237 = ~n2725 & ~n3236;
  assign n3238 = n3231 & ~n3237;
  assign n3239 = STATE2_REG_3_ & ~n3228;
  assign n3240 = ~INSTQUEUEWR_ADDR_REG_0_ & n2409;
  assign n3241 = n3016 & n3240;
  assign n3242 = ~n3228 & ~n3241;
  assign n3243 = STATE2_REG_2_ & n3242;
  assign n3244 = ~n3239 & ~n3243;
  assign n3245 = n3010 & n3244;
  assign n3246 = ~n3238 & n3245;
  assign n3247 = INSTQUEUE_REG_13__7_ & ~n3246;
  assign n3248 = STATE2_REG_2_ & ~n3242;
  assign n3249 = n3006 & n3235;
  assign n3250 = ~n2725 & ~n3249;
  assign n3251 = ~n3231 & ~n3250;
  assign n3252 = ~n3248 & ~n3251;
  assign n3253 = n3025 & ~n3252;
  assign n3254 = n3032 & n3234;
  assign n3255 = n3035 & n3228;
  assign n3256 = n3037 & n3233;
  assign n3257 = ~n3254 & ~n3255;
  assign n3258 = ~n3256 & n3257;
  assign n3259 = ~n3247 & ~n3253;
  assign n625 = ~n3258 | ~n3259;
  assign n3261 = INSTQUEUE_REG_13__6_ & ~n3246;
  assign n3262 = n3044 & ~n3252;
  assign n3263 = n3046 & n3234;
  assign n3264 = n3048 & n3228;
  assign n3265 = n3050 & n3233;
  assign n3266 = ~n3263 & ~n3264;
  assign n3267 = ~n3265 & n3266;
  assign n3268 = ~n3261 & ~n3262;
  assign n630 = ~n3267 | ~n3268;
  assign n3270 = INSTQUEUE_REG_13__5_ & ~n3246;
  assign n3271 = n3057 & ~n3252;
  assign n3272 = n3059 & n3234;
  assign n3273 = n3061 & n3228;
  assign n3274 = n3063 & n3233;
  assign n3275 = ~n3272 & ~n3273;
  assign n3276 = ~n3274 & n3275;
  assign n3277 = ~n3270 & ~n3271;
  assign n635 = ~n3276 | ~n3277;
  assign n3279 = INSTQUEUE_REG_13__4_ & ~n3246;
  assign n3280 = n3070 & ~n3252;
  assign n3281 = n3072 & n3234;
  assign n3282 = n3074 & n3228;
  assign n3283 = n3076 & n3233;
  assign n3284 = ~n3281 & ~n3282;
  assign n3285 = ~n3283 & n3284;
  assign n3286 = ~n3279 & ~n3280;
  assign n640 = ~n3285 | ~n3286;
  assign n3288 = INSTQUEUE_REG_13__3_ & ~n3246;
  assign n3289 = n3083 & ~n3252;
  assign n3290 = n3085 & n3234;
  assign n3291 = n3087 & n3228;
  assign n3292 = n3089 & n3233;
  assign n3293 = ~n3290 & ~n3291;
  assign n3294 = ~n3292 & n3293;
  assign n3295 = ~n3288 & ~n3289;
  assign n645 = ~n3294 | ~n3295;
  assign n3297 = INSTQUEUE_REG_13__2_ & ~n3246;
  assign n3298 = n3096 & ~n3252;
  assign n3299 = n3098 & n3234;
  assign n3300 = n3100 & n3228;
  assign n3301 = n3102 & n3233;
  assign n3302 = ~n3299 & ~n3300;
  assign n3303 = ~n3301 & n3302;
  assign n3304 = ~n3297 & ~n3298;
  assign n650 = ~n3303 | ~n3304;
  assign n3306 = INSTQUEUE_REG_13__1_ & ~n3246;
  assign n3307 = n3109 & ~n3252;
  assign n3308 = n3111 & n3234;
  assign n3309 = n3113 & n3228;
  assign n3310 = n3115 & n3233;
  assign n3311 = ~n3308 & ~n3309;
  assign n3312 = ~n3310 & n3311;
  assign n3313 = ~n3306 & ~n3307;
  assign n655 = ~n3312 | ~n3313;
  assign n3315 = INSTQUEUE_REG_13__0_ & ~n3246;
  assign n3316 = n3122 & ~n3252;
  assign n3317 = n3124 & n3234;
  assign n3318 = n3126 & n3228;
  assign n3319 = n3128 & n3233;
  assign n3320 = ~n3317 & ~n3318;
  assign n3321 = ~n3319 & n3320;
  assign n3322 = ~n3315 & ~n3316;
  assign n660 = ~n3321 | ~n3322;
  assign n3324 = ~INSTQUEUEWR_ADDR_REG_1_ & ~INSTQUEUEWR_ADDR_REG_0_;
  assign n3325 = n2718 & n3324;
  assign n3326 = n2618 & n2633;
  assign n3327 = n2720 & n3326;
  assign n3328 = ~n3325 & ~n3327;
  assign n3329 = ~n2884 & n2887;
  assign n3330 = n3001 & n3329;
  assign n3331 = n2880 & n2884;
  assign n3332 = n3003 & n3331;
  assign n3333 = ~n3330 & ~n3332;
  assign n3334 = n3011 & n3333;
  assign n3335 = ~n2725 & ~n3334;
  assign n3336 = n3328 & ~n3335;
  assign n3337 = STATE2_REG_3_ & ~n3325;
  assign n3338 = n2409 & n3016;
  assign n3339 = STATE2_REG_2_ & ~n3338;
  assign n3340 = ~n3337 & ~n3339;
  assign n3341 = n3010 & n3340;
  assign n3342 = ~n3336 & n3341;
  assign n3343 = INSTQUEUE_REG_12__7_ & ~n3342;
  assign n3344 = STATE2_REG_2_ & n3338;
  assign n3345 = n3006 & n3333;
  assign n3346 = ~n2725 & ~n3345;
  assign n3347 = ~n3328 & ~n3346;
  assign n3348 = ~n3344 & ~n3347;
  assign n3349 = n3025 & ~n3348;
  assign n3350 = n3032 & n3332;
  assign n3351 = n3035 & n3325;
  assign n3352 = n3037 & n3330;
  assign n3353 = ~n3350 & ~n3351;
  assign n3354 = ~n3352 & n3353;
  assign n3355 = ~n3343 & ~n3349;
  assign n665 = ~n3354 | ~n3355;
  assign n3357 = INSTQUEUE_REG_12__6_ & ~n3342;
  assign n3358 = n3044 & ~n3348;
  assign n3359 = n3046 & n3332;
  assign n3360 = n3048 & n3325;
  assign n3361 = n3050 & n3330;
  assign n3362 = ~n3359 & ~n3360;
  assign n3363 = ~n3361 & n3362;
  assign n3364 = ~n3357 & ~n3358;
  assign n670 = ~n3363 | ~n3364;
  assign n3366 = INSTQUEUE_REG_12__5_ & ~n3342;
  assign n3367 = n3057 & ~n3348;
  assign n3368 = n3059 & n3332;
  assign n3369 = n3061 & n3325;
  assign n3370 = n3063 & n3330;
  assign n3371 = ~n3368 & ~n3369;
  assign n3372 = ~n3370 & n3371;
  assign n3373 = ~n3366 & ~n3367;
  assign n675 = ~n3372 | ~n3373;
  assign n3375 = INSTQUEUE_REG_12__4_ & ~n3342;
  assign n3376 = n3070 & ~n3348;
  assign n3377 = n3072 & n3332;
  assign n3378 = n3074 & n3325;
  assign n3379 = n3076 & n3330;
  assign n3380 = ~n3377 & ~n3378;
  assign n3381 = ~n3379 & n3380;
  assign n3382 = ~n3375 & ~n3376;
  assign n680 = ~n3381 | ~n3382;
  assign n3384 = INSTQUEUE_REG_12__3_ & ~n3342;
  assign n3385 = n3083 & ~n3348;
  assign n3386 = n3085 & n3332;
  assign n3387 = n3087 & n3325;
  assign n3388 = n3089 & n3330;
  assign n3389 = ~n3386 & ~n3387;
  assign n3390 = ~n3388 & n3389;
  assign n3391 = ~n3384 & ~n3385;
  assign n685 = ~n3390 | ~n3391;
  assign n3393 = INSTQUEUE_REG_12__2_ & ~n3342;
  assign n3394 = n3096 & ~n3348;
  assign n3395 = n3098 & n3332;
  assign n3396 = n3100 & n3325;
  assign n3397 = n3102 & n3330;
  assign n3398 = ~n3395 & ~n3396;
  assign n3399 = ~n3397 & n3398;
  assign n3400 = ~n3393 & ~n3394;
  assign n690 = ~n3399 | ~n3400;
  assign n3402 = INSTQUEUE_REG_12__1_ & ~n3342;
  assign n3403 = n3109 & ~n3348;
  assign n3404 = n3111 & n3332;
  assign n3405 = n3113 & n3325;
  assign n3406 = n3115 & n3330;
  assign n3407 = ~n3404 & ~n3405;
  assign n3408 = ~n3406 & n3407;
  assign n3409 = ~n3402 & ~n3403;
  assign n695 = ~n3408 | ~n3409;
  assign n3411 = INSTQUEUE_REG_12__0_ & ~n3342;
  assign n3412 = n3122 & ~n3348;
  assign n3413 = n3124 & n3332;
  assign n3414 = n3126 & n3325;
  assign n3415 = n3128 & n3330;
  assign n3416 = ~n3413 & ~n3414;
  assign n3417 = ~n3415 & n3416;
  assign n3418 = ~n3411 & ~n3412;
  assign n700 = ~n3417 | ~n3418;
  assign n3420 = n2479 & n2555;
  assign n3421 = ~n2495 & ~n2580;
  assign n3422 = n2721 & n3421;
  assign n3423 = ~n3420 & ~n3422;
  assign n3424 = n2944 & ~n3000;
  assign n3425 = n2888 & n3424;
  assign n3426 = n2889 & n2995;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n3011 & n3427;
  assign n3429 = ~n2725 & ~n3428;
  assign n3430 = n3423 & ~n3429;
  assign n3431 = STATE2_REG_3_ & ~n3420;
  assign n3432 = n2482 & ~n2560;
  assign n3433 = n3017 & n3432;
  assign n3434 = ~n3420 & ~n3433;
  assign n3435 = STATE2_REG_2_ & n3434;
  assign n3436 = ~n3431 & ~n3435;
  assign n3437 = n3010 & n3436;
  assign n3438 = ~n3430 & n3437;
  assign n3439 = INSTQUEUE_REG_11__7_ & ~n3438;
  assign n3440 = STATE2_REG_2_ & ~n3434;
  assign n3441 = n3006 & n3427;
  assign n3442 = ~n2725 & ~n3441;
  assign n3443 = ~n3423 & ~n3442;
  assign n3444 = ~n3440 & ~n3443;
  assign n3445 = n3025 & ~n3444;
  assign n3446 = n3032 & n3426;
  assign n3447 = n3035 & n3420;
  assign n3448 = n3037 & n3425;
  assign n3449 = ~n3446 & ~n3447;
  assign n3450 = ~n3448 & n3449;
  assign n3451 = ~n3439 & ~n3445;
  assign n705 = ~n3450 | ~n3451;
  assign n3453 = INSTQUEUE_REG_11__6_ & ~n3438;
  assign n3454 = n3044 & ~n3444;
  assign n3455 = n3046 & n3426;
  assign n3456 = n3048 & n3420;
  assign n3457 = n3050 & n3425;
  assign n3458 = ~n3455 & ~n3456;
  assign n3459 = ~n3457 & n3458;
  assign n3460 = ~n3453 & ~n3454;
  assign n710 = ~n3459 | ~n3460;
  assign n3462 = INSTQUEUE_REG_11__5_ & ~n3438;
  assign n3463 = n3057 & ~n3444;
  assign n3464 = n3059 & n3426;
  assign n3465 = n3061 & n3420;
  assign n3466 = n3063 & n3425;
  assign n3467 = ~n3464 & ~n3465;
  assign n3468 = ~n3466 & n3467;
  assign n3469 = ~n3462 & ~n3463;
  assign n715 = ~n3468 | ~n3469;
  assign n3471 = INSTQUEUE_REG_11__4_ & ~n3438;
  assign n3472 = n3070 & ~n3444;
  assign n3473 = n3072 & n3426;
  assign n3474 = n3074 & n3420;
  assign n3475 = n3076 & n3425;
  assign n3476 = ~n3473 & ~n3474;
  assign n3477 = ~n3475 & n3476;
  assign n3478 = ~n3471 & ~n3472;
  assign n720 = ~n3477 | ~n3478;
  assign n3480 = INSTQUEUE_REG_11__3_ & ~n3438;
  assign n3481 = n3083 & ~n3444;
  assign n3482 = n3085 & n3426;
  assign n3483 = n3087 & n3420;
  assign n3484 = n3089 & n3425;
  assign n3485 = ~n3482 & ~n3483;
  assign n3486 = ~n3484 & n3485;
  assign n3487 = ~n3480 & ~n3481;
  assign n725 = ~n3486 | ~n3487;
  assign n3489 = INSTQUEUE_REG_11__2_ & ~n3438;
  assign n3490 = n3096 & ~n3444;
  assign n3491 = n3098 & n3426;
  assign n3492 = n3100 & n3420;
  assign n3493 = n3102 & n3425;
  assign n3494 = ~n3491 & ~n3492;
  assign n3495 = ~n3493 & n3494;
  assign n3496 = ~n3489 & ~n3490;
  assign n730 = ~n3495 | ~n3496;
  assign n3498 = INSTQUEUE_REG_11__1_ & ~n3438;
  assign n3499 = n3109 & ~n3444;
  assign n3500 = n3111 & n3426;
  assign n3501 = n3113 & n3420;
  assign n3502 = n3115 & n3425;
  assign n3503 = ~n3500 & ~n3501;
  assign n3504 = ~n3502 & n3503;
  assign n3505 = ~n3498 & ~n3499;
  assign n735 = ~n3504 | ~n3505;
  assign n3507 = INSTQUEUE_REG_11__0_ & ~n3438;
  assign n3508 = n3122 & ~n3444;
  assign n3509 = n3124 & n3426;
  assign n3510 = n3126 & n3420;
  assign n3511 = n3128 & n3425;
  assign n3512 = ~n3509 & ~n3510;
  assign n3513 = ~n3511 & n3512;
  assign n3514 = ~n3507 & ~n3508;
  assign n740 = ~n3513 | ~n3514;
  assign n3516 = n2408 & n2555;
  assign n3517 = n3135 & n3421;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = n3138 & n3424;
  assign n3520 = n2885 & n2995;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = n3011 & n3521;
  assign n3523 = ~n2725 & ~n3522;
  assign n3524 = n3518 & ~n3523;
  assign n3525 = STATE2_REG_3_ & ~n3516;
  assign n3526 = ~n2409 & n3432;
  assign n3527 = STATE2_REG_2_ & ~n3526;
  assign n3528 = ~n3525 & ~n3527;
  assign n3529 = n3010 & n3528;
  assign n3530 = ~n3524 & n3529;
  assign n3531 = INSTQUEUE_REG_10__7_ & ~n3530;
  assign n3532 = STATE2_REG_2_ & n3526;
  assign n3533 = n3006 & n3521;
  assign n3534 = ~n2725 & ~n3533;
  assign n3535 = ~n3518 & ~n3534;
  assign n3536 = ~n3532 & ~n3535;
  assign n3537 = n3025 & ~n3536;
  assign n3538 = n3032 & n3520;
  assign n3539 = n3035 & n3516;
  assign n3540 = n3037 & n3519;
  assign n3541 = ~n3538 & ~n3539;
  assign n3542 = ~n3540 & n3541;
  assign n3543 = ~n3531 & ~n3537;
  assign n745 = ~n3542 | ~n3543;
  assign n3545 = INSTQUEUE_REG_10__6_ & ~n3530;
  assign n3546 = n3044 & ~n3536;
  assign n3547 = n3046 & n3520;
  assign n3548 = n3048 & n3516;
  assign n3549 = n3050 & n3519;
  assign n3550 = ~n3547 & ~n3548;
  assign n3551 = ~n3549 & n3550;
  assign n3552 = ~n3545 & ~n3546;
  assign n750 = ~n3551 | ~n3552;
  assign n3554 = INSTQUEUE_REG_10__5_ & ~n3530;
  assign n3555 = n3057 & ~n3536;
  assign n3556 = n3059 & n3520;
  assign n3557 = n3061 & n3516;
  assign n3558 = n3063 & n3519;
  assign n3559 = ~n3556 & ~n3557;
  assign n3560 = ~n3558 & n3559;
  assign n3561 = ~n3554 & ~n3555;
  assign n755 = ~n3560 | ~n3561;
  assign n3563 = INSTQUEUE_REG_10__4_ & ~n3530;
  assign n3564 = n3070 & ~n3536;
  assign n3565 = n3072 & n3520;
  assign n3566 = n3074 & n3516;
  assign n3567 = n3076 & n3519;
  assign n3568 = ~n3565 & ~n3566;
  assign n3569 = ~n3567 & n3568;
  assign n3570 = ~n3563 & ~n3564;
  assign n760 = ~n3569 | ~n3570;
  assign n3572 = INSTQUEUE_REG_10__3_ & ~n3530;
  assign n3573 = n3083 & ~n3536;
  assign n3574 = n3085 & n3520;
  assign n3575 = n3087 & n3516;
  assign n3576 = n3089 & n3519;
  assign n3577 = ~n3574 & ~n3575;
  assign n3578 = ~n3576 & n3577;
  assign n3579 = ~n3572 & ~n3573;
  assign n765 = ~n3578 | ~n3579;
  assign n3581 = INSTQUEUE_REG_10__2_ & ~n3530;
  assign n3582 = n3096 & ~n3536;
  assign n3583 = n3098 & n3520;
  assign n3584 = n3100 & n3516;
  assign n3585 = n3102 & n3519;
  assign n3586 = ~n3583 & ~n3584;
  assign n3587 = ~n3585 & n3586;
  assign n3588 = ~n3581 & ~n3582;
  assign n770 = ~n3587 | ~n3588;
  assign n3590 = INSTQUEUE_REG_10__1_ & ~n3530;
  assign n3591 = n3109 & ~n3536;
  assign n3592 = n3111 & n3520;
  assign n3593 = n3113 & n3516;
  assign n3594 = n3115 & n3519;
  assign n3595 = ~n3592 & ~n3593;
  assign n3596 = ~n3594 & n3595;
  assign n3597 = ~n3590 & ~n3591;
  assign n775 = ~n3596 | ~n3597;
  assign n3599 = INSTQUEUE_REG_10__0_ & ~n3530;
  assign n3600 = n3122 & ~n3536;
  assign n3601 = n3124 & n3520;
  assign n3602 = n3126 & n3516;
  assign n3603 = n3128 & n3519;
  assign n3604 = ~n3601 & ~n3602;
  assign n3605 = ~n3603 & n3604;
  assign n3606 = ~n3599 & ~n3600;
  assign n780 = ~n3605 | ~n3606;
  assign n3608 = n2407 & n2555;
  assign n3609 = n3229 & n3421;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = n3232 & n3424;
  assign n3612 = n2886 & n2995;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = n3011 & n3613;
  assign n3615 = ~n2725 & ~n3614;
  assign n3616 = n3610 & ~n3615;
  assign n3617 = STATE2_REG_3_ & ~n3608;
  assign n3618 = n3240 & n3432;
  assign n3619 = ~n3608 & ~n3618;
  assign n3620 = STATE2_REG_2_ & n3619;
  assign n3621 = ~n3617 & ~n3620;
  assign n3622 = n3010 & n3621;
  assign n3623 = ~n3616 & n3622;
  assign n3624 = INSTQUEUE_REG_9__7_ & ~n3623;
  assign n3625 = STATE2_REG_2_ & ~n3619;
  assign n3626 = n3006 & n3613;
  assign n3627 = ~n2725 & ~n3626;
  assign n3628 = ~n3610 & ~n3627;
  assign n3629 = ~n3625 & ~n3628;
  assign n3630 = n3025 & ~n3629;
  assign n3631 = n3032 & n3612;
  assign n3632 = n3035 & n3608;
  assign n3633 = n3037 & n3611;
  assign n3634 = ~n3631 & ~n3632;
  assign n3635 = ~n3633 & n3634;
  assign n3636 = ~n3624 & ~n3630;
  assign n785 = ~n3635 | ~n3636;
  assign n3638 = INSTQUEUE_REG_9__6_ & ~n3623;
  assign n3639 = n3044 & ~n3629;
  assign n3640 = n3046 & n3612;
  assign n3641 = n3048 & n3608;
  assign n3642 = n3050 & n3611;
  assign n3643 = ~n3640 & ~n3641;
  assign n3644 = ~n3642 & n3643;
  assign n3645 = ~n3638 & ~n3639;
  assign n790 = ~n3644 | ~n3645;
  assign n3647 = INSTQUEUE_REG_9__5_ & ~n3623;
  assign n3648 = n3057 & ~n3629;
  assign n3649 = n3059 & n3612;
  assign n3650 = n3061 & n3608;
  assign n3651 = n3063 & n3611;
  assign n3652 = ~n3649 & ~n3650;
  assign n3653 = ~n3651 & n3652;
  assign n3654 = ~n3647 & ~n3648;
  assign n795 = ~n3653 | ~n3654;
  assign n3656 = INSTQUEUE_REG_9__4_ & ~n3623;
  assign n3657 = n3070 & ~n3629;
  assign n3658 = n3072 & n3612;
  assign n3659 = n3074 & n3608;
  assign n3660 = n3076 & n3611;
  assign n3661 = ~n3658 & ~n3659;
  assign n3662 = ~n3660 & n3661;
  assign n3663 = ~n3656 & ~n3657;
  assign n800 = ~n3662 | ~n3663;
  assign n3665 = INSTQUEUE_REG_9__3_ & ~n3623;
  assign n3666 = n3083 & ~n3629;
  assign n3667 = n3085 & n3612;
  assign n3668 = n3087 & n3608;
  assign n3669 = n3089 & n3611;
  assign n3670 = ~n3667 & ~n3668;
  assign n3671 = ~n3669 & n3670;
  assign n3672 = ~n3665 & ~n3666;
  assign n805 = ~n3671 | ~n3672;
  assign n3674 = INSTQUEUE_REG_9__2_ & ~n3623;
  assign n3675 = n3096 & ~n3629;
  assign n3676 = n3098 & n3612;
  assign n3677 = n3100 & n3608;
  assign n3678 = n3102 & n3611;
  assign n3679 = ~n3676 & ~n3677;
  assign n3680 = ~n3678 & n3679;
  assign n3681 = ~n3674 & ~n3675;
  assign n810 = ~n3680 | ~n3681;
  assign n3683 = INSTQUEUE_REG_9__1_ & ~n3623;
  assign n3684 = n3109 & ~n3629;
  assign n3685 = n3111 & n3612;
  assign n3686 = n3113 & n3608;
  assign n3687 = n3115 & n3611;
  assign n3688 = ~n3685 & ~n3686;
  assign n3689 = ~n3687 & n3688;
  assign n3690 = ~n3683 & ~n3684;
  assign n815 = ~n3689 | ~n3690;
  assign n3692 = INSTQUEUE_REG_9__0_ & ~n3623;
  assign n3693 = n3122 & ~n3629;
  assign n3694 = n3124 & n3612;
  assign n3695 = n3126 & n3608;
  assign n3696 = n3128 & n3611;
  assign n3697 = ~n3694 & ~n3695;
  assign n3698 = ~n3696 & n3697;
  assign n3699 = ~n3692 & ~n3693;
  assign n820 = ~n3698 | ~n3699;
  assign n3701 = n2555 & n3324;
  assign n3702 = n3326 & n3421;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = n3329 & n3424;
  assign n3705 = n2995 & n3331;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = n3011 & n3706;
  assign n3708 = ~n2725 & ~n3707;
  assign n3709 = n3703 & ~n3708;
  assign n3710 = STATE2_REG_3_ & ~n3701;
  assign n3711 = n2409 & n3432;
  assign n3712 = STATE2_REG_2_ & ~n3711;
  assign n3713 = ~n3710 & ~n3712;
  assign n3714 = n3010 & n3713;
  assign n3715 = ~n3709 & n3714;
  assign n3716 = INSTQUEUE_REG_8__7_ & ~n3715;
  assign n3717 = STATE2_REG_2_ & n3711;
  assign n3718 = n3006 & n3706;
  assign n3719 = ~n2725 & ~n3718;
  assign n3720 = ~n3703 & ~n3719;
  assign n3721 = ~n3717 & ~n3720;
  assign n3722 = n3025 & ~n3721;
  assign n3723 = n3032 & n3705;
  assign n3724 = n3035 & n3701;
  assign n3725 = n3037 & n3704;
  assign n3726 = ~n3723 & ~n3724;
  assign n3727 = ~n3725 & n3726;
  assign n3728 = ~n3716 & ~n3722;
  assign n825 = ~n3727 | ~n3728;
  assign n3730 = INSTQUEUE_REG_8__6_ & ~n3715;
  assign n3731 = n3044 & ~n3721;
  assign n3732 = n3046 & n3705;
  assign n3733 = n3048 & n3701;
  assign n3734 = n3050 & n3704;
  assign n3735 = ~n3732 & ~n3733;
  assign n3736 = ~n3734 & n3735;
  assign n3737 = ~n3730 & ~n3731;
  assign n830 = ~n3736 | ~n3737;
  assign n3739 = INSTQUEUE_REG_8__5_ & ~n3715;
  assign n3740 = n3057 & ~n3721;
  assign n3741 = n3059 & n3705;
  assign n3742 = n3061 & n3701;
  assign n3743 = n3063 & n3704;
  assign n3744 = ~n3741 & ~n3742;
  assign n3745 = ~n3743 & n3744;
  assign n3746 = ~n3739 & ~n3740;
  assign n835 = ~n3745 | ~n3746;
  assign n3748 = INSTQUEUE_REG_8__4_ & ~n3715;
  assign n3749 = n3070 & ~n3721;
  assign n3750 = n3072 & n3705;
  assign n3751 = n3074 & n3701;
  assign n3752 = n3076 & n3704;
  assign n3753 = ~n3750 & ~n3751;
  assign n3754 = ~n3752 & n3753;
  assign n3755 = ~n3748 & ~n3749;
  assign n840 = ~n3754 | ~n3755;
  assign n3757 = INSTQUEUE_REG_8__3_ & ~n3715;
  assign n3758 = n3083 & ~n3721;
  assign n3759 = n3085 & n3705;
  assign n3760 = n3087 & n3701;
  assign n3761 = n3089 & n3704;
  assign n3762 = ~n3759 & ~n3760;
  assign n3763 = ~n3761 & n3762;
  assign n3764 = ~n3757 & ~n3758;
  assign n845 = ~n3763 | ~n3764;
  assign n3766 = INSTQUEUE_REG_8__2_ & ~n3715;
  assign n3767 = n3096 & ~n3721;
  assign n3768 = n3098 & n3705;
  assign n3769 = n3100 & n3701;
  assign n3770 = n3102 & n3704;
  assign n3771 = ~n3768 & ~n3769;
  assign n3772 = ~n3770 & n3771;
  assign n3773 = ~n3766 & ~n3767;
  assign n850 = ~n3772 | ~n3773;
  assign n3775 = INSTQUEUE_REG_8__1_ & ~n3715;
  assign n3776 = n3109 & ~n3721;
  assign n3777 = n3111 & n3705;
  assign n3778 = n3113 & n3701;
  assign n3779 = n3115 & n3704;
  assign n3780 = ~n3777 & ~n3778;
  assign n3781 = ~n3779 & n3780;
  assign n3782 = ~n3775 & ~n3776;
  assign n855 = ~n3781 | ~n3782;
  assign n3784 = INSTQUEUE_REG_8__0_ & ~n3715;
  assign n3785 = n3122 & ~n3721;
  assign n3786 = n3124 & n3705;
  assign n3787 = n3126 & n3701;
  assign n3788 = n3128 & n3704;
  assign n3789 = ~n3786 & ~n3787;
  assign n3790 = ~n3788 & n3789;
  assign n3791 = ~n3784 & ~n3785;
  assign n860 = ~n3790 | ~n3791;
  assign n3793 = n2495 & n2580;
  assign n3794 = n2721 & n3793;
  assign n3795 = ~n2558 & ~n3794;
  assign n3796 = ~n2944 & n3000;
  assign n3797 = n2888 & n3796;
  assign n3798 = ~n2998 & ~n3797;
  assign n3799 = n3011 & n3798;
  assign n3800 = ~n2725 & ~n3799;
  assign n3801 = n3795 & ~n3800;
  assign n3802 = STATE2_REG_3_ & ~n2558;
  assign n3803 = ~n2482 & n2560;
  assign n3804 = n3017 & n3803;
  assign n3805 = ~n2558 & ~n3804;
  assign n3806 = STATE2_REG_2_ & n3805;
  assign n3807 = ~n3802 & ~n3806;
  assign n3808 = n3010 & n3807;
  assign n3809 = ~n3801 & n3808;
  assign n3810 = INSTQUEUE_REG_7__7_ & ~n3809;
  assign n3811 = STATE2_REG_2_ & ~n3805;
  assign n3812 = n3006 & n3798;
  assign n3813 = ~n2725 & ~n3812;
  assign n3814 = ~n3795 & ~n3813;
  assign n3815 = ~n3811 & ~n3814;
  assign n3816 = n3025 & ~n3815;
  assign n3817 = n2998 & n3032;
  assign n3818 = n2558 & n3035;
  assign n3819 = n3037 & n3797;
  assign n3820 = ~n3817 & ~n3818;
  assign n3821 = ~n3819 & n3820;
  assign n3822 = ~n3810 & ~n3816;
  assign n865 = ~n3821 | ~n3822;
  assign n3824 = INSTQUEUE_REG_7__6_ & ~n3809;
  assign n3825 = n3044 & ~n3815;
  assign n3826 = n2998 & n3046;
  assign n3827 = n2558 & n3048;
  assign n3828 = n3050 & n3797;
  assign n3829 = ~n3826 & ~n3827;
  assign n3830 = ~n3828 & n3829;
  assign n3831 = ~n3824 & ~n3825;
  assign n870 = ~n3830 | ~n3831;
  assign n3833 = INSTQUEUE_REG_7__5_ & ~n3809;
  assign n3834 = n3057 & ~n3815;
  assign n3835 = n2998 & n3059;
  assign n3836 = n2558 & n3061;
  assign n3837 = n3063 & n3797;
  assign n3838 = ~n3835 & ~n3836;
  assign n3839 = ~n3837 & n3838;
  assign n3840 = ~n3833 & ~n3834;
  assign n875 = ~n3839 | ~n3840;
  assign n3842 = INSTQUEUE_REG_7__4_ & ~n3809;
  assign n3843 = n3070 & ~n3815;
  assign n3844 = n2998 & n3072;
  assign n3845 = n2558 & n3074;
  assign n3846 = n3076 & n3797;
  assign n3847 = ~n3844 & ~n3845;
  assign n3848 = ~n3846 & n3847;
  assign n3849 = ~n3842 & ~n3843;
  assign n880 = ~n3848 | ~n3849;
  assign n3851 = INSTQUEUE_REG_7__3_ & ~n3809;
  assign n3852 = n3083 & ~n3815;
  assign n3853 = n2998 & n3085;
  assign n3854 = n2558 & n3087;
  assign n3855 = n3089 & n3797;
  assign n3856 = ~n3853 & ~n3854;
  assign n3857 = ~n3855 & n3856;
  assign n3858 = ~n3851 & ~n3852;
  assign n885 = ~n3857 | ~n3858;
  assign n3860 = INSTQUEUE_REG_7__2_ & ~n3809;
  assign n3861 = n3096 & ~n3815;
  assign n3862 = n2998 & n3098;
  assign n3863 = n2558 & n3100;
  assign n3864 = n3102 & n3797;
  assign n3865 = ~n3862 & ~n3863;
  assign n3866 = ~n3864 & n3865;
  assign n3867 = ~n3860 & ~n3861;
  assign n890 = ~n3866 | ~n3867;
  assign n3869 = INSTQUEUE_REG_7__1_ & ~n3809;
  assign n3870 = n3109 & ~n3815;
  assign n3871 = n2998 & n3111;
  assign n3872 = n2558 & n3113;
  assign n3873 = n3115 & n3797;
  assign n3874 = ~n3871 & ~n3872;
  assign n3875 = ~n3873 & n3874;
  assign n3876 = ~n3869 & ~n3870;
  assign n895 = ~n3875 | ~n3876;
  assign n3878 = INSTQUEUE_REG_7__0_ & ~n3809;
  assign n3879 = n3122 & ~n3815;
  assign n3880 = n2998 & n3124;
  assign n3881 = n2558 & n3126;
  assign n3882 = n3128 & n3797;
  assign n3883 = ~n3880 & ~n3881;
  assign n3884 = ~n3882 & n3883;
  assign n3885 = ~n3878 & ~n3879;
  assign n900 = ~n3884 | ~n3885;
  assign n3887 = n2408 & n2557;
  assign n3888 = n3135 & n3793;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = n3138 & n3796;
  assign n3891 = n2885 & n2997;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = n3011 & n3892;
  assign n3894 = ~n2725 & ~n3893;
  assign n3895 = n3889 & ~n3894;
  assign n3896 = STATE2_REG_3_ & ~n3887;
  assign n3897 = ~n2409 & n3803;
  assign n3898 = STATE2_REG_2_ & ~n3897;
  assign n3899 = ~n3896 & ~n3898;
  assign n3900 = n3010 & n3899;
  assign n3901 = ~n3895 & n3900;
  assign n3902 = INSTQUEUE_REG_6__7_ & ~n3901;
  assign n3903 = STATE2_REG_2_ & n3897;
  assign n3904 = n3006 & n3892;
  assign n3905 = ~n2725 & ~n3904;
  assign n3906 = ~n3889 & ~n3905;
  assign n3907 = ~n3903 & ~n3906;
  assign n3908 = n3025 & ~n3907;
  assign n3909 = n3032 & n3891;
  assign n3910 = n3035 & n3887;
  assign n3911 = n3037 & n3890;
  assign n3912 = ~n3909 & ~n3910;
  assign n3913 = ~n3911 & n3912;
  assign n3914 = ~n3902 & ~n3908;
  assign n905 = ~n3913 | ~n3914;
  assign n3916 = INSTQUEUE_REG_6__6_ & ~n3901;
  assign n3917 = n3044 & ~n3907;
  assign n3918 = n3046 & n3891;
  assign n3919 = n3048 & n3887;
  assign n3920 = n3050 & n3890;
  assign n3921 = ~n3918 & ~n3919;
  assign n3922 = ~n3920 & n3921;
  assign n3923 = ~n3916 & ~n3917;
  assign n910 = ~n3922 | ~n3923;
  assign n3925 = INSTQUEUE_REG_6__5_ & ~n3901;
  assign n3926 = n3057 & ~n3907;
  assign n3927 = n3059 & n3891;
  assign n3928 = n3061 & n3887;
  assign n3929 = n3063 & n3890;
  assign n3930 = ~n3927 & ~n3928;
  assign n3931 = ~n3929 & n3930;
  assign n3932 = ~n3925 & ~n3926;
  assign n915 = ~n3931 | ~n3932;
  assign n3934 = INSTQUEUE_REG_6__4_ & ~n3901;
  assign n3935 = n3070 & ~n3907;
  assign n3936 = n3072 & n3891;
  assign n3937 = n3074 & n3887;
  assign n3938 = n3076 & n3890;
  assign n3939 = ~n3936 & ~n3937;
  assign n3940 = ~n3938 & n3939;
  assign n3941 = ~n3934 & ~n3935;
  assign n920 = ~n3940 | ~n3941;
  assign n3943 = INSTQUEUE_REG_6__3_ & ~n3901;
  assign n3944 = n3083 & ~n3907;
  assign n3945 = n3085 & n3891;
  assign n3946 = n3087 & n3887;
  assign n3947 = n3089 & n3890;
  assign n3948 = ~n3945 & ~n3946;
  assign n3949 = ~n3947 & n3948;
  assign n3950 = ~n3943 & ~n3944;
  assign n925 = ~n3949 | ~n3950;
  assign n3952 = INSTQUEUE_REG_6__2_ & ~n3901;
  assign n3953 = n3096 & ~n3907;
  assign n3954 = n3098 & n3891;
  assign n3955 = n3100 & n3887;
  assign n3956 = n3102 & n3890;
  assign n3957 = ~n3954 & ~n3955;
  assign n3958 = ~n3956 & n3957;
  assign n3959 = ~n3952 & ~n3953;
  assign n930 = ~n3958 | ~n3959;
  assign n3961 = INSTQUEUE_REG_6__1_ & ~n3901;
  assign n3962 = n3109 & ~n3907;
  assign n3963 = n3111 & n3891;
  assign n3964 = n3113 & n3887;
  assign n3965 = n3115 & n3890;
  assign n3966 = ~n3963 & ~n3964;
  assign n3967 = ~n3965 & n3966;
  assign n3968 = ~n3961 & ~n3962;
  assign n935 = ~n3967 | ~n3968;
  assign n3970 = INSTQUEUE_REG_6__0_ & ~n3901;
  assign n3971 = n3122 & ~n3907;
  assign n3972 = n3124 & n3891;
  assign n3973 = n3126 & n3887;
  assign n3974 = n3128 & n3890;
  assign n3975 = ~n3972 & ~n3973;
  assign n3976 = ~n3974 & n3975;
  assign n3977 = ~n3970 & ~n3971;
  assign n940 = ~n3976 | ~n3977;
  assign n3979 = n2407 & n2557;
  assign n3980 = n3229 & n3793;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n3232 & n3796;
  assign n3983 = n2886 & n2997;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = n3011 & n3984;
  assign n3986 = ~n2725 & ~n3985;
  assign n3987 = n3981 & ~n3986;
  assign n3988 = STATE2_REG_3_ & ~n3979;
  assign n3989 = n3240 & n3803;
  assign n3990 = ~n3979 & ~n3989;
  assign n3991 = STATE2_REG_2_ & n3990;
  assign n3992 = ~n3988 & ~n3991;
  assign n3993 = n3010 & n3992;
  assign n3994 = ~n3987 & n3993;
  assign n3995 = INSTQUEUE_REG_5__7_ & ~n3994;
  assign n3996 = STATE2_REG_2_ & ~n3990;
  assign n3997 = n3006 & n3984;
  assign n3998 = ~n2725 & ~n3997;
  assign n3999 = ~n3981 & ~n3998;
  assign n4000 = ~n3996 & ~n3999;
  assign n4001 = n3025 & ~n4000;
  assign n4002 = n3032 & n3983;
  assign n4003 = n3035 & n3979;
  assign n4004 = n3037 & n3982;
  assign n4005 = ~n4002 & ~n4003;
  assign n4006 = ~n4004 & n4005;
  assign n4007 = ~n3995 & ~n4001;
  assign n945 = ~n4006 | ~n4007;
  assign n4009 = INSTQUEUE_REG_5__6_ & ~n3994;
  assign n4010 = n3044 & ~n4000;
  assign n4011 = n3046 & n3983;
  assign n4012 = n3048 & n3979;
  assign n4013 = n3050 & n3982;
  assign n4014 = ~n4011 & ~n4012;
  assign n4015 = ~n4013 & n4014;
  assign n4016 = ~n4009 & ~n4010;
  assign n950 = ~n4015 | ~n4016;
  assign n4018 = INSTQUEUE_REG_5__5_ & ~n3994;
  assign n4019 = n3057 & ~n4000;
  assign n4020 = n3059 & n3983;
  assign n4021 = n3061 & n3979;
  assign n4022 = n3063 & n3982;
  assign n4023 = ~n4020 & ~n4021;
  assign n4024 = ~n4022 & n4023;
  assign n4025 = ~n4018 & ~n4019;
  assign n955 = ~n4024 | ~n4025;
  assign n4027 = INSTQUEUE_REG_5__4_ & ~n3994;
  assign n4028 = n3070 & ~n4000;
  assign n4029 = n3072 & n3983;
  assign n4030 = n3074 & n3979;
  assign n4031 = n3076 & n3982;
  assign n4032 = ~n4029 & ~n4030;
  assign n4033 = ~n4031 & n4032;
  assign n4034 = ~n4027 & ~n4028;
  assign n960 = ~n4033 | ~n4034;
  assign n4036 = INSTQUEUE_REG_5__3_ & ~n3994;
  assign n4037 = n3083 & ~n4000;
  assign n4038 = n3085 & n3983;
  assign n4039 = n3087 & n3979;
  assign n4040 = n3089 & n3982;
  assign n4041 = ~n4038 & ~n4039;
  assign n4042 = ~n4040 & n4041;
  assign n4043 = ~n4036 & ~n4037;
  assign n965 = ~n4042 | ~n4043;
  assign n4045 = INSTQUEUE_REG_5__2_ & ~n3994;
  assign n4046 = n3096 & ~n4000;
  assign n4047 = n3098 & n3983;
  assign n4048 = n3100 & n3979;
  assign n4049 = n3102 & n3982;
  assign n4050 = ~n4047 & ~n4048;
  assign n4051 = ~n4049 & n4050;
  assign n4052 = ~n4045 & ~n4046;
  assign n970 = ~n4051 | ~n4052;
  assign n4054 = INSTQUEUE_REG_5__1_ & ~n3994;
  assign n4055 = n3109 & ~n4000;
  assign n4056 = n3111 & n3983;
  assign n4057 = n3113 & n3979;
  assign n4058 = n3115 & n3982;
  assign n4059 = ~n4056 & ~n4057;
  assign n4060 = ~n4058 & n4059;
  assign n4061 = ~n4054 & ~n4055;
  assign n975 = ~n4060 | ~n4061;
  assign n4063 = INSTQUEUE_REG_5__0_ & ~n3994;
  assign n4064 = n3122 & ~n4000;
  assign n4065 = n3124 & n3983;
  assign n4066 = n3126 & n3979;
  assign n4067 = n3128 & n3982;
  assign n4068 = ~n4065 & ~n4066;
  assign n4069 = ~n4067 & n4068;
  assign n4070 = ~n4063 & ~n4064;
  assign n980 = ~n4069 | ~n4070;
  assign n4072 = n2557 & n3324;
  assign n4073 = n3326 & n3793;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n3329 & n3796;
  assign n4076 = n2997 & n3331;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n3011 & n4077;
  assign n4079 = ~n2725 & ~n4078;
  assign n4080 = n4074 & ~n4079;
  assign n4081 = STATE2_REG_3_ & ~n4072;
  assign n4082 = n2409 & n3803;
  assign n4083 = STATE2_REG_2_ & ~n4082;
  assign n4084 = ~n4081 & ~n4083;
  assign n4085 = n3010 & n4084;
  assign n4086 = ~n4080 & n4085;
  assign n4087 = INSTQUEUE_REG_4__7_ & ~n4086;
  assign n4088 = STATE2_REG_2_ & n4082;
  assign n4089 = n3006 & n4077;
  assign n4090 = ~n2725 & ~n4089;
  assign n4091 = ~n4074 & ~n4090;
  assign n4092 = ~n4088 & ~n4091;
  assign n4093 = n3025 & ~n4092;
  assign n4094 = n3032 & n4076;
  assign n4095 = n3035 & n4072;
  assign n4096 = n3037 & n4075;
  assign n4097 = ~n4094 & ~n4095;
  assign n4098 = ~n4096 & n4097;
  assign n4099 = ~n4087 & ~n4093;
  assign n985 = ~n4098 | ~n4099;
  assign n4101 = INSTQUEUE_REG_4__6_ & ~n4086;
  assign n4102 = n3044 & ~n4092;
  assign n4103 = n3046 & n4076;
  assign n4104 = n3048 & n4072;
  assign n4105 = n3050 & n4075;
  assign n4106 = ~n4103 & ~n4104;
  assign n4107 = ~n4105 & n4106;
  assign n4108 = ~n4101 & ~n4102;
  assign n990 = ~n4107 | ~n4108;
  assign n4110 = INSTQUEUE_REG_4__5_ & ~n4086;
  assign n4111 = n3057 & ~n4092;
  assign n4112 = n3059 & n4076;
  assign n4113 = n3061 & n4072;
  assign n4114 = n3063 & n4075;
  assign n4115 = ~n4112 & ~n4113;
  assign n4116 = ~n4114 & n4115;
  assign n4117 = ~n4110 & ~n4111;
  assign n995 = ~n4116 | ~n4117;
  assign n4119 = INSTQUEUE_REG_4__4_ & ~n4086;
  assign n4120 = n3070 & ~n4092;
  assign n4121 = n3072 & n4076;
  assign n4122 = n3074 & n4072;
  assign n4123 = n3076 & n4075;
  assign n4124 = ~n4121 & ~n4122;
  assign n4125 = ~n4123 & n4124;
  assign n4126 = ~n4119 & ~n4120;
  assign n1000 = ~n4125 | ~n4126;
  assign n4128 = INSTQUEUE_REG_4__3_ & ~n4086;
  assign n4129 = n3083 & ~n4092;
  assign n4130 = n3085 & n4076;
  assign n4131 = n3087 & n4072;
  assign n4132 = n3089 & n4075;
  assign n4133 = ~n4130 & ~n4131;
  assign n4134 = ~n4132 & n4133;
  assign n4135 = ~n4128 & ~n4129;
  assign n1005 = ~n4134 | ~n4135;
  assign n4137 = INSTQUEUE_REG_4__2_ & ~n4086;
  assign n4138 = n3096 & ~n4092;
  assign n4139 = n3098 & n4076;
  assign n4140 = n3100 & n4072;
  assign n4141 = n3102 & n4075;
  assign n4142 = ~n4139 & ~n4140;
  assign n4143 = ~n4141 & n4142;
  assign n4144 = ~n4137 & ~n4138;
  assign n1010 = ~n4143 | ~n4144;
  assign n4146 = INSTQUEUE_REG_4__1_ & ~n4086;
  assign n4147 = n3109 & ~n4092;
  assign n4148 = n3111 & n4076;
  assign n4149 = n3113 & n4072;
  assign n4150 = n3115 & n4075;
  assign n4151 = ~n4148 & ~n4149;
  assign n4152 = ~n4150 & n4151;
  assign n4153 = ~n4146 & ~n4147;
  assign n1015 = ~n4152 | ~n4153;
  assign n4155 = INSTQUEUE_REG_4__0_ & ~n4086;
  assign n4156 = n3122 & ~n4092;
  assign n4157 = n3124 & n4076;
  assign n4158 = n3126 & n4072;
  assign n4159 = n3128 & n4075;
  assign n4160 = ~n4157 & ~n4158;
  assign n4161 = ~n4159 & n4160;
  assign n4162 = ~n4155 & ~n4156;
  assign n1020 = ~n4161 | ~n4162;
  assign n4164 = ~INSTQUEUEWR_ADDR_REG_3_ & ~INSTQUEUEWR_ADDR_REG_2_;
  assign n4165 = n2479 & n4164;
  assign n4166 = ~n2495 & n2580;
  assign n4167 = n2721 & n4166;
  assign n4168 = ~n4165 & ~n4167;
  assign n4169 = n2944 & n3000;
  assign n4170 = n2888 & n4169;
  assign n4171 = n2941 & ~n2994;
  assign n4172 = n2889 & n4171;
  assign n4173 = ~n4170 & ~n4172;
  assign n4174 = n3011 & n4173;
  assign n4175 = ~n2725 & ~n4174;
  assign n4176 = n4168 & ~n4175;
  assign n4177 = STATE2_REG_3_ & ~n4165;
  assign n4178 = n2482 & n2560;
  assign n4179 = n3017 & n4178;
  assign n4180 = ~n4165 & ~n4179;
  assign n4181 = STATE2_REG_2_ & n4180;
  assign n4182 = ~n4177 & ~n4181;
  assign n4183 = n3010 & n4182;
  assign n4184 = ~n4176 & n4183;
  assign n4185 = INSTQUEUE_REG_3__7_ & ~n4184;
  assign n4186 = STATE2_REG_2_ & ~n4180;
  assign n4187 = n3006 & n4173;
  assign n4188 = ~n2725 & ~n4187;
  assign n4189 = ~n4168 & ~n4188;
  assign n4190 = ~n4186 & ~n4189;
  assign n4191 = n3025 & ~n4190;
  assign n4192 = n3032 & n4172;
  assign n4193 = n3035 & n4165;
  assign n4194 = n3037 & n4170;
  assign n4195 = ~n4192 & ~n4193;
  assign n4196 = ~n4194 & n4195;
  assign n4197 = ~n4185 & ~n4191;
  assign n1025 = ~n4196 | ~n4197;
  assign n4199 = INSTQUEUE_REG_3__6_ & ~n4184;
  assign n4200 = n3044 & ~n4190;
  assign n4201 = n3046 & n4172;
  assign n4202 = n3048 & n4165;
  assign n4203 = n3050 & n4170;
  assign n4204 = ~n4201 & ~n4202;
  assign n4205 = ~n4203 & n4204;
  assign n4206 = ~n4199 & ~n4200;
  assign n1030 = ~n4205 | ~n4206;
  assign n4208 = INSTQUEUE_REG_3__5_ & ~n4184;
  assign n4209 = n3057 & ~n4190;
  assign n4210 = n3059 & n4172;
  assign n4211 = n3061 & n4165;
  assign n4212 = n3063 & n4170;
  assign n4213 = ~n4210 & ~n4211;
  assign n4214 = ~n4212 & n4213;
  assign n4215 = ~n4208 & ~n4209;
  assign n1035 = ~n4214 | ~n4215;
  assign n4217 = INSTQUEUE_REG_3__4_ & ~n4184;
  assign n4218 = n3070 & ~n4190;
  assign n4219 = n3072 & n4172;
  assign n4220 = n3074 & n4165;
  assign n4221 = n3076 & n4170;
  assign n4222 = ~n4219 & ~n4220;
  assign n4223 = ~n4221 & n4222;
  assign n4224 = ~n4217 & ~n4218;
  assign n1040 = ~n4223 | ~n4224;
  assign n4226 = INSTQUEUE_REG_3__3_ & ~n4184;
  assign n4227 = n3083 & ~n4190;
  assign n4228 = n3085 & n4172;
  assign n4229 = n3087 & n4165;
  assign n4230 = n3089 & n4170;
  assign n4231 = ~n4228 & ~n4229;
  assign n4232 = ~n4230 & n4231;
  assign n4233 = ~n4226 & ~n4227;
  assign n1045 = ~n4232 | ~n4233;
  assign n4235 = INSTQUEUE_REG_3__2_ & ~n4184;
  assign n4236 = n3096 & ~n4190;
  assign n4237 = n3098 & n4172;
  assign n4238 = n3100 & n4165;
  assign n4239 = n3102 & n4170;
  assign n4240 = ~n4237 & ~n4238;
  assign n4241 = ~n4239 & n4240;
  assign n4242 = ~n4235 & ~n4236;
  assign n1050 = ~n4241 | ~n4242;
  assign n4244 = INSTQUEUE_REG_3__1_ & ~n4184;
  assign n4245 = n3109 & ~n4190;
  assign n4246 = n3111 & n4172;
  assign n4247 = n3113 & n4165;
  assign n4248 = n3115 & n4170;
  assign n4249 = ~n4246 & ~n4247;
  assign n4250 = ~n4248 & n4249;
  assign n4251 = ~n4244 & ~n4245;
  assign n1055 = ~n4250 | ~n4251;
  assign n4253 = INSTQUEUE_REG_3__0_ & ~n4184;
  assign n4254 = n3122 & ~n4190;
  assign n4255 = n3124 & n4172;
  assign n4256 = n3126 & n4165;
  assign n4257 = n3128 & n4170;
  assign n4258 = ~n4255 & ~n4256;
  assign n4259 = ~n4257 & n4258;
  assign n4260 = ~n4253 & ~n4254;
  assign n1060 = ~n4259 | ~n4260;
  assign n4262 = n2408 & n4164;
  assign n4263 = n3135 & n4166;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = n3138 & n4169;
  assign n4266 = n2885 & n4171;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = n3011 & n4267;
  assign n4269 = ~n2725 & ~n4268;
  assign n4270 = n4264 & ~n4269;
  assign n4271 = STATE2_REG_3_ & ~n4262;
  assign n4272 = ~n2409 & n4178;
  assign n4273 = STATE2_REG_2_ & ~n4272;
  assign n4274 = ~n4271 & ~n4273;
  assign n4275 = n3010 & n4274;
  assign n4276 = ~n4270 & n4275;
  assign n4277 = INSTQUEUE_REG_2__7_ & ~n4276;
  assign n4278 = STATE2_REG_2_ & n4272;
  assign n4279 = n3006 & n4267;
  assign n4280 = ~n2725 & ~n4279;
  assign n4281 = ~n4264 & ~n4280;
  assign n4282 = ~n4278 & ~n4281;
  assign n4283 = n3025 & ~n4282;
  assign n4284 = n3032 & n4266;
  assign n4285 = n3035 & n4262;
  assign n4286 = n3037 & n4265;
  assign n4287 = ~n4284 & ~n4285;
  assign n4288 = ~n4286 & n4287;
  assign n4289 = ~n4277 & ~n4283;
  assign n1065 = ~n4288 | ~n4289;
  assign n4291 = INSTQUEUE_REG_2__6_ & ~n4276;
  assign n4292 = n3044 & ~n4282;
  assign n4293 = n3046 & n4266;
  assign n4294 = n3048 & n4262;
  assign n4295 = n3050 & n4265;
  assign n4296 = ~n4293 & ~n4294;
  assign n4297 = ~n4295 & n4296;
  assign n4298 = ~n4291 & ~n4292;
  assign n1070 = ~n4297 | ~n4298;
  assign n4300 = INSTQUEUE_REG_2__5_ & ~n4276;
  assign n4301 = n3057 & ~n4282;
  assign n4302 = n3059 & n4266;
  assign n4303 = n3061 & n4262;
  assign n4304 = n3063 & n4265;
  assign n4305 = ~n4302 & ~n4303;
  assign n4306 = ~n4304 & n4305;
  assign n4307 = ~n4300 & ~n4301;
  assign n1075 = ~n4306 | ~n4307;
  assign n4309 = INSTQUEUE_REG_2__4_ & ~n4276;
  assign n4310 = n3070 & ~n4282;
  assign n4311 = n3072 & n4266;
  assign n4312 = n3074 & n4262;
  assign n4313 = n3076 & n4265;
  assign n4314 = ~n4311 & ~n4312;
  assign n4315 = ~n4313 & n4314;
  assign n4316 = ~n4309 & ~n4310;
  assign n1080 = ~n4315 | ~n4316;
  assign n4318 = INSTQUEUE_REG_2__3_ & ~n4276;
  assign n4319 = n3083 & ~n4282;
  assign n4320 = n3085 & n4266;
  assign n4321 = n3087 & n4262;
  assign n4322 = n3089 & n4265;
  assign n4323 = ~n4320 & ~n4321;
  assign n4324 = ~n4322 & n4323;
  assign n4325 = ~n4318 & ~n4319;
  assign n1085 = ~n4324 | ~n4325;
  assign n4327 = INSTQUEUE_REG_2__2_ & ~n4276;
  assign n4328 = n3096 & ~n4282;
  assign n4329 = n3098 & n4266;
  assign n4330 = n3100 & n4262;
  assign n4331 = n3102 & n4265;
  assign n4332 = ~n4329 & ~n4330;
  assign n4333 = ~n4331 & n4332;
  assign n4334 = ~n4327 & ~n4328;
  assign n1090 = ~n4333 | ~n4334;
  assign n4336 = INSTQUEUE_REG_2__1_ & ~n4276;
  assign n4337 = n3109 & ~n4282;
  assign n4338 = n3111 & n4266;
  assign n4339 = n3113 & n4262;
  assign n4340 = n3115 & n4265;
  assign n4341 = ~n4338 & ~n4339;
  assign n4342 = ~n4340 & n4341;
  assign n4343 = ~n4336 & ~n4337;
  assign n1095 = ~n4342 | ~n4343;
  assign n4345 = INSTQUEUE_REG_2__0_ & ~n4276;
  assign n4346 = n3122 & ~n4282;
  assign n4347 = n3124 & n4266;
  assign n4348 = n3126 & n4262;
  assign n4349 = n3128 & n4265;
  assign n4350 = ~n4347 & ~n4348;
  assign n4351 = ~n4349 & n4350;
  assign n4352 = ~n4345 & ~n4346;
  assign n1100 = ~n4351 | ~n4352;
  assign n4354 = n2407 & n4164;
  assign n4355 = n3229 & n4166;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n3232 & n4169;
  assign n4358 = n2886 & n4171;
  assign n4359 = ~n4357 & ~n4358;
  assign n4360 = n3011 & n4359;
  assign n4361 = ~n2725 & ~n4360;
  assign n4362 = n4356 & ~n4361;
  assign n4363 = STATE2_REG_3_ & ~n4354;
  assign n4364 = n3240 & n4178;
  assign n4365 = ~n4354 & ~n4364;
  assign n4366 = STATE2_REG_2_ & n4365;
  assign n4367 = ~n4363 & ~n4366;
  assign n4368 = n3010 & n4367;
  assign n4369 = ~n4362 & n4368;
  assign n4370 = INSTQUEUE_REG_1__7_ & ~n4369;
  assign n4371 = STATE2_REG_2_ & ~n4365;
  assign n4372 = n3006 & n4359;
  assign n4373 = ~n2725 & ~n4372;
  assign n4374 = ~n4356 & ~n4373;
  assign n4375 = ~n4371 & ~n4374;
  assign n4376 = n3025 & ~n4375;
  assign n4377 = n3032 & n4358;
  assign n4378 = n3035 & n4354;
  assign n4379 = n3037 & n4357;
  assign n4380 = ~n4377 & ~n4378;
  assign n4381 = ~n4379 & n4380;
  assign n4382 = ~n4370 & ~n4376;
  assign n1105 = ~n4381 | ~n4382;
  assign n4384 = INSTQUEUE_REG_1__6_ & ~n4369;
  assign n4385 = n3044 & ~n4375;
  assign n4386 = n3046 & n4358;
  assign n4387 = n3048 & n4354;
  assign n4388 = n3050 & n4357;
  assign n4389 = ~n4386 & ~n4387;
  assign n4390 = ~n4388 & n4389;
  assign n4391 = ~n4384 & ~n4385;
  assign n1110 = ~n4390 | ~n4391;
  assign n4393 = INSTQUEUE_REG_1__5_ & ~n4369;
  assign n4394 = n3057 & ~n4375;
  assign n4395 = n3059 & n4358;
  assign n4396 = n3061 & n4354;
  assign n4397 = n3063 & n4357;
  assign n4398 = ~n4395 & ~n4396;
  assign n4399 = ~n4397 & n4398;
  assign n4400 = ~n4393 & ~n4394;
  assign n1115 = ~n4399 | ~n4400;
  assign n4402 = INSTQUEUE_REG_1__4_ & ~n4369;
  assign n4403 = n3070 & ~n4375;
  assign n4404 = n3072 & n4358;
  assign n4405 = n3074 & n4354;
  assign n4406 = n3076 & n4357;
  assign n4407 = ~n4404 & ~n4405;
  assign n4408 = ~n4406 & n4407;
  assign n4409 = ~n4402 & ~n4403;
  assign n1120 = ~n4408 | ~n4409;
  assign n4411 = INSTQUEUE_REG_1__3_ & ~n4369;
  assign n4412 = n3083 & ~n4375;
  assign n4413 = n3085 & n4358;
  assign n4414 = n3087 & n4354;
  assign n4415 = n3089 & n4357;
  assign n4416 = ~n4413 & ~n4414;
  assign n4417 = ~n4415 & n4416;
  assign n4418 = ~n4411 & ~n4412;
  assign n1125 = ~n4417 | ~n4418;
  assign n4420 = INSTQUEUE_REG_1__2_ & ~n4369;
  assign n4421 = n3096 & ~n4375;
  assign n4422 = n3098 & n4358;
  assign n4423 = n3100 & n4354;
  assign n4424 = n3102 & n4357;
  assign n4425 = ~n4422 & ~n4423;
  assign n4426 = ~n4424 & n4425;
  assign n4427 = ~n4420 & ~n4421;
  assign n1130 = ~n4426 | ~n4427;
  assign n4429 = INSTQUEUE_REG_1__1_ & ~n4369;
  assign n4430 = n3109 & ~n4375;
  assign n4431 = n3111 & n4358;
  assign n4432 = n3113 & n4354;
  assign n4433 = n3115 & n4357;
  assign n4434 = ~n4431 & ~n4432;
  assign n4435 = ~n4433 & n4434;
  assign n4436 = ~n4429 & ~n4430;
  assign n1135 = ~n4435 | ~n4436;
  assign n4438 = INSTQUEUE_REG_1__0_ & ~n4369;
  assign n4439 = n3122 & ~n4375;
  assign n4440 = n3124 & n4358;
  assign n4441 = n3126 & n4354;
  assign n4442 = n3128 & n4357;
  assign n4443 = ~n4440 & ~n4441;
  assign n4444 = ~n4442 & n4443;
  assign n4445 = ~n4438 & ~n4439;
  assign n1140 = ~n4444 | ~n4445;
  assign n4447 = n3324 & n4164;
  assign n4448 = n3326 & n4166;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = n3329 & n4169;
  assign n4451 = n3331 & n4171;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = n3011 & n4452;
  assign n4454 = ~n2725 & ~n4453;
  assign n4455 = n4449 & ~n4454;
  assign n4456 = STATE2_REG_3_ & ~n4447;
  assign n4457 = n2409 & n4178;
  assign n4458 = STATE2_REG_2_ & ~n4457;
  assign n4459 = ~n4456 & ~n4458;
  assign n4460 = n3010 & n4459;
  assign n4461 = ~n4455 & n4460;
  assign n4462 = INSTQUEUE_REG_0__7_ & ~n4461;
  assign n4463 = STATE2_REG_2_ & n4457;
  assign n4464 = n3006 & n4452;
  assign n4465 = ~n2725 & ~n4464;
  assign n4466 = ~n4449 & ~n4465;
  assign n4467 = ~n4463 & ~n4466;
  assign n4468 = n3025 & ~n4467;
  assign n4469 = n3032 & n4451;
  assign n4470 = n3035 & n4447;
  assign n4471 = n3037 & n4450;
  assign n4472 = ~n4469 & ~n4470;
  assign n4473 = ~n4471 & n4472;
  assign n4474 = ~n4462 & ~n4468;
  assign n1145 = ~n4473 | ~n4474;
  assign n4476 = INSTQUEUE_REG_0__6_ & ~n4461;
  assign n4477 = n3044 & ~n4467;
  assign n4478 = n3046 & n4451;
  assign n4479 = n3048 & n4447;
  assign n4480 = n3050 & n4450;
  assign n4481 = ~n4478 & ~n4479;
  assign n4482 = ~n4480 & n4481;
  assign n4483 = ~n4476 & ~n4477;
  assign n1150 = ~n4482 | ~n4483;
  assign n4485 = INSTQUEUE_REG_0__5_ & ~n4461;
  assign n4486 = n3057 & ~n4467;
  assign n4487 = n3059 & n4451;
  assign n4488 = n3061 & n4447;
  assign n4489 = n3063 & n4450;
  assign n4490 = ~n4487 & ~n4488;
  assign n4491 = ~n4489 & n4490;
  assign n4492 = ~n4485 & ~n4486;
  assign n1155 = ~n4491 | ~n4492;
  assign n4494 = INSTQUEUE_REG_0__4_ & ~n4461;
  assign n4495 = n3070 & ~n4467;
  assign n4496 = n3072 & n4451;
  assign n4497 = n3074 & n4447;
  assign n4498 = n3076 & n4450;
  assign n4499 = ~n4496 & ~n4497;
  assign n4500 = ~n4498 & n4499;
  assign n4501 = ~n4494 & ~n4495;
  assign n1160 = ~n4500 | ~n4501;
  assign n4503 = INSTQUEUE_REG_0__3_ & ~n4461;
  assign n4504 = n3083 & ~n4467;
  assign n4505 = n3085 & n4451;
  assign n4506 = n3087 & n4447;
  assign n4507 = n3089 & n4450;
  assign n4508 = ~n4505 & ~n4506;
  assign n4509 = ~n4507 & n4508;
  assign n4510 = ~n4503 & ~n4504;
  assign n1165 = ~n4509 | ~n4510;
  assign n4512 = INSTQUEUE_REG_0__2_ & ~n4461;
  assign n4513 = n3096 & ~n4467;
  assign n4514 = n3098 & n4451;
  assign n4515 = n3100 & n4447;
  assign n4516 = n3102 & n4450;
  assign n4517 = ~n4514 & ~n4515;
  assign n4518 = ~n4516 & n4517;
  assign n4519 = ~n4512 & ~n4513;
  assign n1170 = ~n4518 | ~n4519;
  assign n4521 = INSTQUEUE_REG_0__1_ & ~n4461;
  assign n4522 = n3109 & ~n4467;
  assign n4523 = n3111 & n4451;
  assign n4524 = n3113 & n4447;
  assign n4525 = n3115 & n4450;
  assign n4526 = ~n4523 & ~n4524;
  assign n4527 = ~n4525 & n4526;
  assign n4528 = ~n4521 & ~n4522;
  assign n1175 = ~n4527 | ~n4528;
  assign n4530 = INSTQUEUE_REG_0__0_ & ~n4461;
  assign n4531 = n3122 & ~n4467;
  assign n4532 = n3124 & n4451;
  assign n4533 = n3126 & n4447;
  assign n4534 = n3128 & n4450;
  assign n4535 = ~n4532 & ~n4533;
  assign n4536 = ~n4534 & n4535;
  assign n4537 = ~n4530 & ~n4531;
  assign n1180 = ~n4536 | ~n4537;
  assign n4539 = STATE2_REG_3_ & ~STATE2_REG_0_;
  assign n4540 = STATE2_REG_0_ & FLUSH_REG;
  assign n4541 = n1707 & n4540;
  assign n4542 = ~n4539 & ~n4541;
  assign n4543 = ~n2544 & n2674;
  assign n4544 = n4542 & ~n4543;
  assign n4545 = INSTQUEUERD_ADDR_REG_4_ & n4544;
  assign n4546 = n2268_1 & n2405;
  assign n4547 = ~n2570 & n4546;
  assign n4548 = ~n4544 & n4547;
  assign n1185 = n4545 | n4548;
  assign n4550 = n2405 & ~n2595;
  assign n4551 = ~n2586 & n2688;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4544 & ~n4552;
  assign n4554 = INSTQUEUERD_ADDR_REG_3_ & n4544;
  assign n1190 = n4553 | n4554;
  assign n4556 = n2405 & ~n2518;
  assign n4557 = n2305 & ~n2311;
  assign n4558 = ~n2320 & n2688;
  assign n4559 = ~n4556 & ~n4557;
  assign n4560 = ~n4558 & n4559;
  assign n4561 = ~n4544 & ~n4560;
  assign n4562 = INSTQUEUERD_ADDR_REG_2_ & n4544;
  assign n1195 = n4561 | n4562;
  assign n4564 = n2405 & ~n2635;
  assign n4565 = n2305 & n2311;
  assign n4566 = n2627 & n2688;
  assign n4567 = ~n4564 & ~n4565;
  assign n4568 = ~n4566 & n4567;
  assign n4569 = ~n4544 & ~n4568;
  assign n4570 = INSTQUEUERD_ADDR_REG_1_ & n4544;
  assign n1200 = n4569 | n4570;
  assign n4572 = n2405 & ~n2620;
  assign n4573 = STATE2_REG_1_ & n2304;
  assign n4574 = ~INSTQUEUERD_ADDR_REG_0_ & n2688;
  assign n4575 = ~n4572 & ~n4573;
  assign n4576 = ~n4574 & n4575;
  assign n4577 = ~n4544 & ~n4576;
  assign n4578 = INSTQUEUERD_ADDR_REG_0_ & n4544;
  assign n1205 = n4577 | n4578;
  assign n4580 = STATE2_REG_0_ & n1707;
  assign n4581 = ~n2707 & n4580;
  assign n4582 = ~n3010 & ~n4541;
  assign n4583 = ~n4581 & n4582;
  assign n1210 = INSTQUEUEWR_ADDR_REG_4_ & n4583;
  assign n4585 = ~STATE2_REG_3_ & STATE2_REG_1_;
  assign n4586 = ~n2580 & ~n4585;
  assign n4587 = n2725 & n2994;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = n2888 & ~n2944;
  assign n4590 = ~n3000 & ~n4589;
  assign n4591 = ~n3797 & ~n4590;
  assign n4592 = n3006 & ~n4591;
  assign n4593 = n4588 & ~n4592;
  assign n4594 = ~n4583 & ~n4593;
  assign n4595 = INSTQUEUEWR_ADDR_REG_3_ & n4583;
  assign n1215 = n4594 | n4595;
  assign n4597 = n2495 & ~n4585;
  assign n4598 = n2725 & ~n2941;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = ~n2888 & ~n2944;
  assign n4601 = n2888 & n2944;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = n3006 & ~n4602;
  assign n4604 = n4599 & ~n4603;
  assign n4605 = ~n4583 & ~n4604;
  assign n4606 = INSTQUEUEWR_ADDR_REG_2_ & n4583;
  assign n1220 = n4605 | n4606;
  assign n4608 = ~n2633 & ~n4585;
  assign n4609 = n2725 & ~n2880;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~n3138 & ~n3232;
  assign n4612 = n3006 & ~n4611;
  assign n4613 = n4610 & ~n4612;
  assign n4614 = ~n4583 & ~n4613;
  assign n4615 = INSTQUEUEWR_ADDR_REG_1_ & n4583;
  assign n1225 = n4614 | n4615;
  assign n4617 = ~n2618 & ~n4585;
  assign n4618 = n2724 & ~n2884;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~n2708 & n4619;
  assign n4621 = ~n4583 & ~n4620;
  assign n4622 = INSTQUEUEWR_ADDR_REG_0_ & n4583;
  assign n1230 = n4621 | n4622;
  assign n4624 = ~STATE2_REG_2_ & n2406;
  assign n4625 = ~n2395 & n2411;
  assign n4626 = n2138_1 & n4625;
  assign n4627 = ~n4624 & ~n4626;
  assign n4628 = n2101 & n2288_1;
  assign n4629 = ~n1776 & ~n2338_1;
  assign n4630 = n1807 & ~n2293_1;
  assign n4631 = ~READY_N & ~n4630;
  assign n4632 = n2282 & n4631;
  assign n4633 = n4629 & ~n4632;
  assign n4634 = ~n2262 & ~n4633;
  assign n4635 = n2100 & n4634;
  assign n4636 = ~n1807 & ~n2656;
  assign n4637 = ~n2285 & ~n4636;
  assign n4638 = ~READY_N & n4637;
  assign n4639 = ~n2100 & n4638;
  assign n4640 = n2541 & ~n4628;
  assign n4641 = ~n4635 & n4640;
  assign n4642 = ~n4639 & n4641;
  assign n4643 = n2674 & ~n4642;
  assign n4644 = n4627 & ~n4643;
  assign n4645 = STATE2_REG_2_ & ~n4644;
  assign n4646 = n2266 & n4645;
  assign n4647 = ~INSTADDRPOINTER_REG_0_ & n4646;
  assign n4648 = n2152 & n2814;
  assign n4649 = n1776 & ~n1839;
  assign n4650 = n2234 & ~n2884;
  assign n4651 = ~n4648 & ~n4649;
  assign n4652 = ~n4650 & n4651;
  assign n4653 = ~INSTADDRPOINTER_REG_0_ & n4652;
  assign n4654 = INSTADDRPOINTER_REG_0_ & ~n4652;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = n2112 & n2265;
  assign n4657 = STATE2_REG_2_ & ~n1807;
  assign n4658 = ~n1776 & n4657;
  assign n4659 = n2282 & n4658;
  assign n4660 = ~n4656 & ~n4659;
  assign n4661 = n2113_1 & n2152;
  assign n4662 = ~n2102 & ~n2268_1;
  assign n4663 = ~n2389 & n4662;
  assign n4664 = n4660 & ~n4661;
  assign n4665 = n4663 & n4664;
  assign n4666 = STATE2_REG_2_ & ~n4665;
  assign n4667 = ~n4644 & n4666;
  assign n4668 = n4655 & n4667;
  assign n4669 = ~n4647 & ~n4668;
  assign n4670 = n1776 & n2382;
  assign n4671 = n2356 & n2387;
  assign n4672 = ~n2318_1 & ~n2344;
  assign n4673 = ~n4671 & n4672;
  assign n4674 = n2498 & ~n4670;
  assign n4675 = n4673 & n4674;
  assign n4676 = n2515 & n4675;
  assign n4677 = n4645 & ~n4676;
  assign n4678 = ~INSTADDRPOINTER_REG_0_ & n4677;
  assign n4679 = n2264 & ~n2402;
  assign n4680 = ~n2264 & n2402;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = ~n2264 & ~n2402;
  assign n4683 = EBX_REG_0_ & ~n4682;
  assign n4684 = ~n1776 & ~n2329;
  assign n4685 = INSTADDRPOINTER_REG_0_ & ~n4684;
  assign n4686 = ~n4683 & ~n4685;
  assign n4687 = ~n2264 & ~n4686;
  assign n4688 = n2264 & n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4681 & n4689;
  assign n4691 = n4681 & ~n4689;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = n2152 & n2282;
  assign n4694 = ~n2419 & ~n4693;
  assign n4695 = n4645 & ~n4694;
  assign n4696 = ~n4692 & n4695;
  assign n4697 = ~n4678 & ~n4696;
  assign n4698 = ~STATE2_REG_2_ & ~n4644;
  assign n4699 = REIP_REG_0_ & n4698;
  assign n4700 = INSTADDRPOINTER_REG_0_ & n4644;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = n2109 & n4645;
  assign n4703 = INSTADDRPOINTER_REG_0_ & n4702;
  assign n4704 = n4701 & ~n4703;
  assign n4705 = n4669 & n4697;
  assign n1235 = ~n4704 | ~n4705;
  assign n4707 = ~n2308_1 & n4646;
  assign n4708 = ~n1776 & n1994;
  assign n4709 = n2100 & ~n4708;
  assign n4710 = ~n1839 & n4709;
  assign n4711 = ~n2814 & n2863;
  assign n4712 = n2814 & ~n2863;
  assign n4713 = ~n4711 & ~n4712;
  assign n4714 = n2152 & ~n4713;
  assign n4715 = n2234 & ~n2880;
  assign n4716 = n4710 & ~n4714;
  assign n4717 = ~n4715 & n4716;
  assign n4718 = ~INSTADDRPOINTER_REG_1_ & n4717;
  assign n4719 = INSTADDRPOINTER_REG_1_ & ~n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4654 & n4720;
  assign n4722 = n4654 & ~n4720;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = n4667 & ~n4723;
  assign n4725 = ~n4707 & ~n4724;
  assign n4726 = ~n2308_1 & n4677;
  assign n4727 = n2264 & n2402;
  assign n4728 = ~n4682 & ~n4689;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = EBX_REG_1_ & ~n4682;
  assign n4731 = INSTADDRPOINTER_REG_1_ & ~n4684;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733 = ~n2264 & ~n4732;
  assign n4734 = n2264 & n4732;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = n4684 & ~n4735;
  assign n4737 = ~n4684 & n4735;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = n4729 & ~n4738;
  assign n4740 = ~n4729 & n4738;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = n4695 & ~n4741;
  assign n4743 = ~n4726 & ~n4742;
  assign n4744 = REIP_REG_1_ & n4698;
  assign n4745 = INSTADDRPOINTER_REG_1_ & n4644;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~INSTADDRPOINTER_REG_1_ & n4702;
  assign n4748 = n4746 & ~n4747;
  assign n4749 = n4725 & n4743;
  assign n1240 = ~n4748 | ~n4749;
  assign n4751 = INSTADDRPOINTER_REG_0_ & INSTADDRPOINTER_REG_1_;
  assign n4752 = ~INSTADDRPOINTER_REG_2_ & ~n4751;
  assign n4753 = INSTADDRPOINTER_REG_2_ & n4751;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = n4646 & ~n4754;
  assign n4756 = ~n2814 & ~n2863;
  assign n4757 = n2921 & ~n4756;
  assign n4758 = ~n2921 & n4756;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = n2152 & ~n4759;
  assign n4761 = n2234 & ~n2941;
  assign n4762 = ~n4649 & ~n4760;
  assign n4763 = ~n4761 & n4762;
  assign n4764 = ~INSTADDRPOINTER_REG_2_ & n4763;
  assign n4765 = INSTADDRPOINTER_REG_2_ & ~n4763;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = n4654 & ~n4718;
  assign n4768 = ~n4719 & ~n4767;
  assign n4769 = n4766 & ~n4768;
  assign n4770 = ~n4766 & n4768;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = n4667 & n4771;
  assign n4773 = ~n4755 & ~n4772;
  assign n4774 = ~INSTADDRPOINTER_REG_2_ & n4751;
  assign n4775 = INSTADDRPOINTER_REG_2_ & ~n4751;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n4677 & ~n4776;
  assign n4778 = EBX_REG_2_ & ~n4682;
  assign n4779 = INSTADDRPOINTER_REG_2_ & ~n4684;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n2264 & ~n4780;
  assign n4782 = n2264 & n4780;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = ~n4684 & ~n4735;
  assign n4785 = n4684 & n4735;
  assign n4786 = ~n4729 & ~n4785;
  assign n4787 = ~n4784 & ~n4786;
  assign n4788 = ~n4783 & ~n4787;
  assign n4789 = n4783 & n4787;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = n4695 & n4790;
  assign n4792 = ~n4777 & ~n4791;
  assign n4793 = REIP_REG_2_ & n4698;
  assign n4794 = INSTADDRPOINTER_REG_2_ & n4644;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = INSTADDRPOINTER_REG_1_ & ~INSTADDRPOINTER_REG_2_;
  assign n4797 = ~INSTADDRPOINTER_REG_1_ & INSTADDRPOINTER_REG_2_;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = n4702 & ~n4798;
  assign n4800 = n4795 & ~n4799;
  assign n4801 = n4773 & n4792;
  assign n1245 = ~n4800 | ~n4801;
  assign n4803 = INSTADDRPOINTER_REG_0_ & INSTADDRPOINTER_REG_2_;
  assign n4804 = INSTADDRPOINTER_REG_1_ & n4803;
  assign n4805 = INSTADDRPOINTER_REG_3_ & ~n4804;
  assign n4806 = ~INSTADDRPOINTER_REG_3_ & n4804;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = n4677 & ~n4807;
  assign n4809 = EBX_REG_3_ & ~n4682;
  assign n4810 = INSTADDRPOINTER_REG_3_ & ~n4684;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = ~n2264 & ~n4811;
  assign n4813 = n2264 & n4811;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = ~n4788 & ~n4814;
  assign n4816 = n4788 & n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n4695 & ~n4817;
  assign n4819 = ~INSTADDRPOINTER_REG_3_ & n4752;
  assign n4820 = INSTADDRPOINTER_REG_3_ & ~n4752;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = n4646 & n4821;
  assign n4823 = ~n4808 & ~n4818;
  assign n4824 = ~n4822 & n4823;
  assign n4825 = REIP_REG_3_ & n4698;
  assign n4826 = INSTADDRPOINTER_REG_3_ & n4644;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = INSTADDRPOINTER_REG_1_ & INSTADDRPOINTER_REG_2_;
  assign n4829 = ~INSTADDRPOINTER_REG_3_ & n4828;
  assign n4830 = INSTADDRPOINTER_REG_3_ & ~n4828;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = n4702 & ~n4831;
  assign n4833 = n2977 & n4757;
  assign n4834 = ~n2977 & ~n4757;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = n2152 & n4835;
  assign n4837 = n2234 & n2994;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = ~INSTADDRPOINTER_REG_3_ & n4838;
  assign n4840 = INSTADDRPOINTER_REG_3_ & ~n4838;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = ~n4764 & ~n4768;
  assign n4843 = ~n4765 & ~n4842;
  assign n4844 = n4841 & ~n4843;
  assign n4845 = ~n4841 & n4843;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = n4667 & n4846;
  assign n4848 = n4827 & ~n4832;
  assign n4849 = ~n4847 & n4848;
  assign n1250 = ~n4824 | ~n4849;
  assign n4851 = INSTADDRPOINTER_REG_3_ & n4804;
  assign n4852 = ~INSTADDRPOINTER_REG_4_ & n4851;
  assign n4853 = INSTADDRPOINTER_REG_4_ & ~n4851;
  assign n4854 = ~n4852 & ~n4853;
  assign n4855 = n4677 & ~n4854;
  assign n4856 = EBX_REG_4_ & ~n4682;
  assign n4857 = INSTADDRPOINTER_REG_4_ & ~n4684;
  assign n4858 = ~n4856 & ~n4857;
  assign n4859 = ~n2264 & ~n4858;
  assign n4860 = n2264 & n4858;
  assign n4861 = ~n4859 & ~n4860;
  assign n4862 = ~n4783 & ~n4814;
  assign n4863 = ~n4787 & n4862;
  assign n4864 = ~n4861 & ~n4863;
  assign n4865 = n4861 & n4863;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = n4695 & ~n4866;
  assign n4868 = ~INSTADDRPOINTER_REG_4_ & n4820;
  assign n4869 = INSTADDRPOINTER_REG_4_ & ~n4820;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = n4646 & ~n4870;
  assign n4872 = ~n4855 & ~n4867;
  assign n4873 = ~n4871 & n4872;
  assign n4874 = REIP_REG_4_ & n4698;
  assign n4875 = INSTADDRPOINTER_REG_4_ & n4644;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = INSTADDRPOINTER_REG_3_ & n4828;
  assign n4878 = ~INSTADDRPOINTER_REG_4_ & n4877;
  assign n4879 = INSTADDRPOINTER_REG_4_ & ~n4877;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = n4702 & ~n4880;
  assign n4882 = n4876 & ~n4881;
  assign n4883 = INSTQUEUE_REG_0__4_ & n2728;
  assign n4884 = INSTQUEUE_REG_1__4_ & n2731;
  assign n4885 = INSTQUEUE_REG_2__4_ & n2734;
  assign n4886 = INSTQUEUE_REG_3__4_ & n2737;
  assign n4887 = ~n4883 & ~n4884;
  assign n4888 = ~n4885 & n4887;
  assign n4889 = ~n4886 & n4888;
  assign n4890 = INSTQUEUE_REG_4__4_ & n2743;
  assign n4891 = INSTQUEUE_REG_5__4_ & n2745;
  assign n4892 = INSTQUEUE_REG_6__4_ & n2747;
  assign n4893 = INSTQUEUE_REG_7__4_ & n2749;
  assign n4894 = ~n4890 & ~n4891;
  assign n4895 = ~n4892 & n4894;
  assign n4896 = ~n4893 & n4895;
  assign n4897 = INSTQUEUE_REG_8__4_ & n2755;
  assign n4898 = INSTQUEUE_REG_9__4_ & n2757;
  assign n4899 = INSTQUEUE_REG_10__4_ & n2759;
  assign n4900 = INSTQUEUE_REG_11__4_ & n2761;
  assign n4901 = ~n4897 & ~n4898;
  assign n4902 = ~n4899 & n4901;
  assign n4903 = ~n4900 & n4902;
  assign n4904 = INSTQUEUE_REG_12__4_ & n2767;
  assign n4905 = INSTQUEUE_REG_13__4_ & n2769;
  assign n4906 = INSTQUEUE_REG_14__4_ & n2771;
  assign n4907 = INSTQUEUE_REG_15__4_ & n2773;
  assign n4908 = ~n4904 & ~n4905;
  assign n4909 = ~n4906 & n4908;
  assign n4910 = ~n4907 & n4909;
  assign n4911 = n4889 & n4896;
  assign n4912 = n4903 & n4911;
  assign n4913 = n4910 & n4912;
  assign n4914 = n4834 & n4913;
  assign n4915 = ~n4834 & ~n4913;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = n2152 & ~n4916;
  assign n4918 = INSTQUEUE_REG_0__4_ & n2138_1;
  assign n4919 = n2143_1 & ~n4913;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n2781 & n4913;
  assign n4922 = n2783 & ~n4913;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n2781 & ~n4923;
  assign n4925 = n2781 & n4923;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~n4920 & ~n4926;
  assign n4928 = n4920 & n4926;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n2933 & ~n2989;
  assign n4931 = n2831 & ~n2935;
  assign n4932 = ~n2936 & ~n4931;
  assign n4933 = ~n2932 & ~n4932;
  assign n4934 = n4930 & ~n4933;
  assign n4935 = ~n2988 & ~n4934;
  assign n4936 = n4929 & n4935;
  assign n4937 = ~n4929 & ~n4935;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = n2234 & ~n4938;
  assign n4940 = ~n4917 & ~n4939;
  assign n4941 = ~INSTADDRPOINTER_REG_4_ & n4940;
  assign n4942 = INSTADDRPOINTER_REG_4_ & ~n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4839 & ~n4843;
  assign n4945 = ~n4840 & ~n4944;
  assign n4946 = n4943 & ~n4945;
  assign n4947 = ~n4943 & n4945;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = n4667 & n4948;
  assign n4950 = n4873 & n4882;
  assign n1255 = n4949 | ~n4950;
  assign n4952 = INSTADDRPOINTER_REG_3_ & INSTADDRPOINTER_REG_4_;
  assign n4953 = n4804 & n4952;
  assign n4954 = INSTADDRPOINTER_REG_5_ & ~n4953;
  assign n4955 = ~INSTADDRPOINTER_REG_5_ & n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = n4677 & ~n4956;
  assign n4958 = EBX_REG_5_ & ~n4682;
  assign n4959 = INSTADDRPOINTER_REG_5_ & ~n4684;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = ~n2264 & ~n4960;
  assign n4962 = n2264 & n4960;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = ~n4861 & n4863;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = n4963 & n4964;
  assign n4967 = ~n4965 & ~n4966;
  assign n4968 = n4695 & ~n4967;
  assign n4969 = INSTADDRPOINTER_REG_4_ & n4820;
  assign n4970 = ~INSTADDRPOINTER_REG_5_ & n4969;
  assign n4971 = INSTADDRPOINTER_REG_5_ & ~n4969;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = n4646 & ~n4972;
  assign n4974 = ~n4957 & ~n4968;
  assign n4975 = ~n4973 & n4974;
  assign n4976 = REIP_REG_5_ & n4698;
  assign n4977 = INSTADDRPOINTER_REG_5_ & n4644;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = INSTADDRPOINTER_REG_4_ & n4877;
  assign n4980 = ~INSTADDRPOINTER_REG_5_ & n4979;
  assign n4981 = INSTADDRPOINTER_REG_5_ & ~n4979;
  assign n4982 = ~n4980 & ~n4981;
  assign n4983 = n4702 & ~n4982;
  assign n4984 = n4978 & ~n4983;
  assign n4985 = n4834 & ~n4913;
  assign n4986 = INSTQUEUE_REG_0__5_ & n2728;
  assign n4987 = INSTQUEUE_REG_1__5_ & n2731;
  assign n4988 = INSTQUEUE_REG_2__5_ & n2734;
  assign n4989 = INSTQUEUE_REG_3__5_ & n2737;
  assign n4990 = ~n4986 & ~n4987;
  assign n4991 = ~n4988 & n4990;
  assign n4992 = ~n4989 & n4991;
  assign n4993 = INSTQUEUE_REG_4__5_ & n2743;
  assign n4994 = INSTQUEUE_REG_5__5_ & n2745;
  assign n4995 = INSTQUEUE_REG_6__5_ & n2747;
  assign n4996 = INSTQUEUE_REG_7__5_ & n2749;
  assign n4997 = ~n4993 & ~n4994;
  assign n4998 = ~n4995 & n4997;
  assign n4999 = ~n4996 & n4998;
  assign n5000 = INSTQUEUE_REG_8__5_ & n2755;
  assign n5001 = INSTQUEUE_REG_9__5_ & n2757;
  assign n5002 = INSTQUEUE_REG_10__5_ & n2759;
  assign n5003 = INSTQUEUE_REG_11__5_ & n2761;
  assign n5004 = ~n5000 & ~n5001;
  assign n5005 = ~n5002 & n5004;
  assign n5006 = ~n5003 & n5005;
  assign n5007 = INSTQUEUE_REG_12__5_ & n2767;
  assign n5008 = INSTQUEUE_REG_13__5_ & n2769;
  assign n5009 = INSTQUEUE_REG_14__5_ & n2771;
  assign n5010 = INSTQUEUE_REG_15__5_ & n2773;
  assign n5011 = ~n5007 & ~n5008;
  assign n5012 = ~n5009 & n5011;
  assign n5013 = ~n5010 & n5012;
  assign n5014 = n4992 & n4999;
  assign n5015 = n5006 & n5014;
  assign n5016 = n5013 & n5015;
  assign n5017 = n4985 & n5016;
  assign n5018 = ~n4985 & ~n5016;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = n2152 & ~n5019;
  assign n5021 = INSTQUEUE_REG_0__5_ & n2138_1;
  assign n5022 = n2143_1 & ~n5016;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = n2781 & n5016;
  assign n5025 = n2783 & ~n5016;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = ~n2781 & ~n5026;
  assign n5028 = n2781 & n5026;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = ~n5023 & ~n5029;
  assign n5031 = n5023 & n5029;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = ~n2979 & ~n4928;
  assign n5034 = ~n2987 & n5033;
  assign n5035 = ~n4927 & ~n5034;
  assign n5036 = ~n2933 & ~n4928;
  assign n5037 = ~n2989 & ~n4933;
  assign n5038 = n5036 & n5037;
  assign n5039 = n5035 & ~n5038;
  assign n5040 = n5032 & n5039;
  assign n5041 = ~n5032 & ~n5039;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = n2234 & ~n5042;
  assign n5044 = ~n5020 & ~n5043;
  assign n5045 = ~INSTADDRPOINTER_REG_5_ & n5044;
  assign n5046 = INSTADDRPOINTER_REG_5_ & ~n5044;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = ~n4941 & ~n4945;
  assign n5049 = ~n4942 & ~n5048;
  assign n5050 = n5047 & ~n5049;
  assign n5051 = ~n5047 & n5049;
  assign n5052 = ~n5050 & ~n5051;
  assign n5053 = n4667 & n5052;
  assign n5054 = n4975 & n4984;
  assign n1260 = n5053 | ~n5054;
  assign n5056 = INSTADDRPOINTER_REG_5_ & n4953;
  assign n5057 = ~INSTADDRPOINTER_REG_6_ & n5056;
  assign n5058 = INSTADDRPOINTER_REG_6_ & ~n5056;
  assign n5059 = ~n5057 & ~n5058;
  assign n5060 = n4677 & ~n5059;
  assign n5061 = EBX_REG_6_ & ~n4682;
  assign n5062 = INSTADDRPOINTER_REG_6_ & ~n4684;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = ~n2264 & ~n5063;
  assign n5065 = n2264 & n5063;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = ~n4861 & ~n4963;
  assign n5068 = n4863 & n5067;
  assign n5069 = ~n5066 & ~n5068;
  assign n5070 = n5066 & n5068;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = n4695 & ~n5071;
  assign n5073 = INSTADDRPOINTER_REG_5_ & n4969;
  assign n5074 = ~INSTADDRPOINTER_REG_6_ & n5073;
  assign n5075 = INSTADDRPOINTER_REG_6_ & ~n5073;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = n4646 & ~n5076;
  assign n5078 = ~n5060 & ~n5072;
  assign n5079 = ~n5077 & n5078;
  assign n5080 = REIP_REG_6_ & n4698;
  assign n5081 = INSTADDRPOINTER_REG_6_ & n4644;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = INSTADDRPOINTER_REG_5_ & n4979;
  assign n5084 = ~INSTADDRPOINTER_REG_6_ & n5083;
  assign n5085 = INSTADDRPOINTER_REG_6_ & ~n5083;
  assign n5086 = ~n5084 & ~n5085;
  assign n5087 = n4702 & ~n5086;
  assign n5088 = n5082 & ~n5087;
  assign n5089 = n4985 & ~n5016;
  assign n5090 = INSTQUEUE_REG_0__6_ & n2728;
  assign n5091 = INSTQUEUE_REG_1__6_ & n2731;
  assign n5092 = INSTQUEUE_REG_2__6_ & n2734;
  assign n5093 = INSTQUEUE_REG_3__6_ & n2737;
  assign n5094 = ~n5090 & ~n5091;
  assign n5095 = ~n5092 & n5094;
  assign n5096 = ~n5093 & n5095;
  assign n5097 = INSTQUEUE_REG_4__6_ & n2743;
  assign n5098 = INSTQUEUE_REG_5__6_ & n2745;
  assign n5099 = INSTQUEUE_REG_6__6_ & n2747;
  assign n5100 = INSTQUEUE_REG_7__6_ & n2749;
  assign n5101 = ~n5097 & ~n5098;
  assign n5102 = ~n5099 & n5101;
  assign n5103 = ~n5100 & n5102;
  assign n5104 = INSTQUEUE_REG_8__6_ & n2755;
  assign n5105 = INSTQUEUE_REG_9__6_ & n2757;
  assign n5106 = INSTQUEUE_REG_10__6_ & n2759;
  assign n5107 = INSTQUEUE_REG_11__6_ & n2761;
  assign n5108 = ~n5104 & ~n5105;
  assign n5109 = ~n5106 & n5108;
  assign n5110 = ~n5107 & n5109;
  assign n5111 = INSTQUEUE_REG_12__6_ & n2767;
  assign n5112 = INSTQUEUE_REG_13__6_ & n2769;
  assign n5113 = INSTQUEUE_REG_14__6_ & n2771;
  assign n5114 = INSTQUEUE_REG_15__6_ & n2773;
  assign n5115 = ~n5111 & ~n5112;
  assign n5116 = ~n5113 & n5115;
  assign n5117 = ~n5114 & n5116;
  assign n5118 = n5096 & n5103;
  assign n5119 = n5110 & n5118;
  assign n5120 = n5117 & n5119;
  assign n5121 = n5089 & n5120;
  assign n5122 = ~n5089 & ~n5120;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = n2152 & ~n5123;
  assign n5125 = INSTQUEUE_REG_0__6_ & n2138_1;
  assign n5126 = n2143_1 & ~n5120;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = n2781 & n5120;
  assign n5129 = n2783 & ~n5120;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~n2781 & ~n5130;
  assign n5132 = n2781 & n5130;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = ~n5127 & ~n5133;
  assign n5135 = n5127 & n5133;
  assign n5136 = ~n5134 & ~n5135;
  assign n5137 = ~n5031 & ~n5039;
  assign n5138 = ~n5030 & ~n5137;
  assign n5139 = n5136 & ~n5138;
  assign n5140 = ~n5030 & ~n5136;
  assign n5141 = ~n5137 & n5140;
  assign n5142 = ~n5139 & ~n5141;
  assign n5143 = n2234 & n5142;
  assign n5144 = ~n5124 & ~n5143;
  assign n5145 = INSTADDRPOINTER_REG_6_ & ~n5144;
  assign n5146 = ~INSTADDRPOINTER_REG_6_ & n5144;
  assign n5147 = ~n5145 & ~n5146;
  assign n5148 = ~n5045 & ~n5049;
  assign n5149 = ~n5046 & ~n5148;
  assign n5150 = n5147 & ~n5149;
  assign n5151 = ~n5147 & n5149;
  assign n5152 = ~n5150 & ~n5151;
  assign n5153 = n4667 & n5152;
  assign n5154 = n5079 & n5088;
  assign n1265 = n5153 | ~n5154;
  assign n5156 = INSTADDRPOINTER_REG_5_ & INSTADDRPOINTER_REG_6_;
  assign n5157 = n4953 & n5156;
  assign n5158 = INSTADDRPOINTER_REG_7_ & ~n5157;
  assign n5159 = ~INSTADDRPOINTER_REG_7_ & n5157;
  assign n5160 = ~n5158 & ~n5159;
  assign n5161 = n4677 & ~n5160;
  assign n5162 = EBX_REG_7_ & ~n4682;
  assign n5163 = INSTADDRPOINTER_REG_7_ & ~n4684;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n2264 & ~n5164;
  assign n5166 = n2264 & n5164;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n5066 & n5068;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = n5167 & n5168;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = n4695 & ~n5171;
  assign n5173 = INSTADDRPOINTER_REG_6_ & n5073;
  assign n5174 = ~INSTADDRPOINTER_REG_7_ & n5173;
  assign n5175 = INSTADDRPOINTER_REG_7_ & ~n5173;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = n4646 & ~n5176;
  assign n5178 = ~n5161 & ~n5172;
  assign n5179 = ~n5177 & n5178;
  assign n5180 = REIP_REG_7_ & n4698;
  assign n5181 = INSTADDRPOINTER_REG_7_ & n4644;
  assign n5182 = ~n5180 & ~n5181;
  assign n5183 = INSTADDRPOINTER_REG_6_ & n5083;
  assign n5184 = ~INSTADDRPOINTER_REG_7_ & n5183;
  assign n5185 = INSTADDRPOINTER_REG_7_ & ~n5183;
  assign n5186 = ~n5184 & ~n5185;
  assign n5187 = n4702 & ~n5186;
  assign n5188 = n5182 & ~n5187;
  assign n5189 = n5089 & ~n5120;
  assign n5190 = n2780 & n5189;
  assign n5191 = ~n2780 & ~n5189;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = n2152 & ~n5192;
  assign n5194 = n2780 & n2781;
  assign n5195 = ~n2780 & n2783;
  assign n5196 = ~n5194 & ~n5195;
  assign n5197 = ~n2781 & ~n5196;
  assign n5198 = n2781 & n5196;
  assign n5199 = INSTQUEUE_REG_0__7_ & n2138_1;
  assign n5200 = n2143_1 & ~n2780;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = ~n5197 & ~n5198;
  assign n5203 = n5201 & n5202;
  assign n5204 = ~n5201 & ~n5202;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206 = n5134 & n5205;
  assign n5207 = ~n5030 & ~n5205;
  assign n5208 = ~n5137 & n5207;
  assign n5209 = ~n5134 & n5208;
  assign n5210 = ~n5031 & n5205;
  assign n5211 = ~n4927 & ~n5030;
  assign n5212 = ~n5034 & n5211;
  assign n5213 = ~n5038 & n5212;
  assign n5214 = n5210 & ~n5213;
  assign n5215 = ~n5135 & n5214;
  assign n5216 = n5135 & ~n5205;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5206 & ~n5209;
  assign n5219 = n5217 & n5218;
  assign n5220 = n2234 & n5219;
  assign n5221 = ~n5193 & ~n5220;
  assign n5222 = ~INSTADDRPOINTER_REG_7_ & n5221;
  assign n5223 = INSTADDRPOINTER_REG_7_ & ~n5221;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5146 & ~n5149;
  assign n5226 = ~n5145 & ~n5225;
  assign n5227 = n5224 & ~n5226;
  assign n5228 = ~n5224 & n5226;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = n4667 & n5229;
  assign n5231 = n5179 & n5188;
  assign n1270 = n5230 | ~n5231;
  assign n5233 = INSTADDRPOINTER_REG_7_ & n5157;
  assign n5234 = ~INSTADDRPOINTER_REG_8_ & n5233;
  assign n5235 = INSTADDRPOINTER_REG_8_ & ~n5233;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = n4677 & ~n5236;
  assign n5238 = EBX_REG_8_ & ~n4682;
  assign n5239 = INSTADDRPOINTER_REG_8_ & ~n4684;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = ~n2264 & ~n5240;
  assign n5242 = n2264 & n5240;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = ~n5066 & ~n5167;
  assign n5245 = n5068 & n5244;
  assign n5246 = ~n5243 & ~n5245;
  assign n5247 = n5243 & n5245;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n4695 & ~n5248;
  assign n5250 = INSTADDRPOINTER_REG_7_ & n5173;
  assign n5251 = ~INSTADDRPOINTER_REG_8_ & n5250;
  assign n5252 = INSTADDRPOINTER_REG_8_ & ~n5250;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = n4646 & ~n5253;
  assign n5255 = ~n5237 & ~n5249;
  assign n5256 = ~n5254 & n5255;
  assign n5257 = REIP_REG_8_ & n4698;
  assign n5258 = INSTADDRPOINTER_REG_8_ & n4644;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = INSTADDRPOINTER_REG_7_ & n5183;
  assign n5261 = ~INSTADDRPOINTER_REG_8_ & n5260;
  assign n5262 = INSTADDRPOINTER_REG_8_ & ~n5260;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = n4702 & ~n5263;
  assign n5265 = n5259 & ~n5264;
  assign n5266 = ~n2780 & ~n5120;
  assign n5267 = n5089 & n5266;
  assign n5268 = n2152 & n5267;
  assign n5269 = n2324 & n2583;
  assign n5270 = n1760 & n5269;
  assign n5271 = INSTQUEUE_REG_0__0_ & n5270;
  assign n5272 = n1753 & n5269;
  assign n5273 = INSTQUEUE_REG_1__0_ & n5272;
  assign n5274 = n1722_1 & n5269;
  assign n5275 = INSTQUEUE_REG_2__0_ & n5274;
  assign n5276 = n1763 & n5269;
  assign n5277 = INSTQUEUE_REG_3__0_ & n5276;
  assign n5278 = ~n5271 & ~n5273;
  assign n5279 = ~n5275 & n5278;
  assign n5280 = ~n5277 & n5279;
  assign n5281 = ~n2324 & n2583;
  assign n5282 = n1760 & n5281;
  assign n5283 = INSTQUEUE_REG_4__0_ & n5282;
  assign n5284 = n1753 & n5281;
  assign n5285 = INSTQUEUE_REG_5__0_ & n5284;
  assign n5286 = n1722_1 & n5281;
  assign n5287 = INSTQUEUE_REG_6__0_ & n5286;
  assign n5288 = n1763 & n5281;
  assign n5289 = INSTQUEUE_REG_7__0_ & n5288;
  assign n5290 = ~n5283 & ~n5285;
  assign n5291 = ~n5287 & n5290;
  assign n5292 = ~n5289 & n5291;
  assign n5293 = n2324 & ~n2583;
  assign n5294 = n1760 & n5293;
  assign n5295 = INSTQUEUE_REG_8__0_ & n5294;
  assign n5296 = n1753 & n5293;
  assign n5297 = INSTQUEUE_REG_9__0_ & n5296;
  assign n5298 = n1722_1 & n5293;
  assign n5299 = INSTQUEUE_REG_10__0_ & n5298;
  assign n5300 = n1763 & n5293;
  assign n5301 = INSTQUEUE_REG_11__0_ & n5300;
  assign n5302 = ~n5295 & ~n5297;
  assign n5303 = ~n5299 & n5302;
  assign n5304 = ~n5301 & n5303;
  assign n5305 = ~n2324 & ~n2583;
  assign n5306 = n1760 & n5305;
  assign n5307 = INSTQUEUE_REG_12__0_ & n5306;
  assign n5308 = n1753 & n5305;
  assign n5309 = INSTQUEUE_REG_13__0_ & n5308;
  assign n5310 = n1722_1 & n5305;
  assign n5311 = INSTQUEUE_REG_14__0_ & n5310;
  assign n5312 = n1763 & n5305;
  assign n5313 = INSTQUEUE_REG_15__0_ & n5312;
  assign n5314 = ~n5307 & ~n5309;
  assign n5315 = ~n5311 & n5314;
  assign n5316 = ~n5313 & n5315;
  assign n5317 = n5280 & n5292;
  assign n5318 = n5304 & n5317;
  assign n5319 = n5316 & n5318;
  assign n5320 = ~n2138_1 & ~n2143_1;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = ~n2781 & n5321;
  assign n5323 = n2781 & ~n5321;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5135 & ~n5203;
  assign n5326 = ~n4928 & ~n5031;
  assign n5327 = n5325 & n5326;
  assign n5328 = ~n4935 & n5327;
  assign n5329 = n4927 & ~n5031;
  assign n5330 = n5325 & n5329;
  assign n5331 = n5134 & n5325;
  assign n5332 = n5030 & n5325;
  assign n5333 = ~n5204 & ~n5330;
  assign n5334 = ~n5331 & n5333;
  assign n5335 = ~n5332 & n5334;
  assign n5336 = ~n5328 & n5335;
  assign n5337 = ~n5324 & ~n5336;
  assign n5338 = n5324 & n5336;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = n2234 & n5339;
  assign n5341 = ~n5268 & ~n5340;
  assign n5342 = ~INSTADDRPOINTER_REG_8_ & n5341;
  assign n5343 = INSTADDRPOINTER_REG_8_ & ~n5341;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = n5046 & ~n5222;
  assign n5346 = ~n5146 & n5345;
  assign n5347 = INSTADDRPOINTER_REG_6_ & ~n5222;
  assign n5348 = ~n5144 & n5347;
  assign n5349 = ~n5346 & ~n5348;
  assign n5350 = ~n4941 & ~n5222;
  assign n5351 = ~n5045 & ~n5146;
  assign n5352 = ~n4945 & n5350;
  assign n5353 = n5351 & n5352;
  assign n5354 = n4942 & ~n5045;
  assign n5355 = ~n5146 & n5354;
  assign n5356 = ~n5222 & n5355;
  assign n5357 = ~n5223 & ~n5356;
  assign n5358 = n5349 & ~n5353;
  assign n5359 = n5357 & n5358;
  assign n5360 = n5344 & ~n5359;
  assign n5361 = ~n5344 & n5359;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = n4667 & n5362;
  assign n5364 = n5256 & n5265;
  assign n1275 = n5363 | ~n5364;
  assign n5366 = INSTADDRPOINTER_REG_7_ & INSTADDRPOINTER_REG_8_;
  assign n5367 = n5157 & n5366;
  assign n5368 = INSTADDRPOINTER_REG_9_ & ~n5367;
  assign n5369 = ~INSTADDRPOINTER_REG_9_ & n5367;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371 = n4677 & ~n5370;
  assign n5372 = EBX_REG_9_ & ~n4682;
  assign n5373 = INSTADDRPOINTER_REG_9_ & ~n4684;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n2264 & ~n5374;
  assign n5376 = n2264 & n5374;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5243 & n5245;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = n5377 & n5378;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = n4695 & ~n5381;
  assign n5383 = INSTADDRPOINTER_REG_8_ & n5250;
  assign n5384 = ~INSTADDRPOINTER_REG_9_ & n5383;
  assign n5385 = INSTADDRPOINTER_REG_9_ & ~n5383;
  assign n5386 = ~n5384 & ~n5385;
  assign n5387 = n4646 & ~n5386;
  assign n5388 = ~n5371 & ~n5382;
  assign n5389 = ~n5387 & n5388;
  assign n5390 = REIP_REG_9_ & n4698;
  assign n5391 = INSTADDRPOINTER_REG_9_ & n4644;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = INSTADDRPOINTER_REG_8_ & n5260;
  assign n5394 = ~INSTADDRPOINTER_REG_9_ & n5393;
  assign n5395 = INSTADDRPOINTER_REG_9_ & ~n5393;
  assign n5396 = ~n5394 & ~n5395;
  assign n5397 = n4702 & ~n5396;
  assign n5398 = n5392 & ~n5397;
  assign n5399 = INSTQUEUE_REG_0__1_ & n5270;
  assign n5400 = INSTQUEUE_REG_1__1_ & n5272;
  assign n5401 = INSTQUEUE_REG_2__1_ & n5274;
  assign n5402 = INSTQUEUE_REG_3__1_ & n5276;
  assign n5403 = ~n5399 & ~n5400;
  assign n5404 = ~n5401 & n5403;
  assign n5405 = ~n5402 & n5404;
  assign n5406 = INSTQUEUE_REG_4__1_ & n5282;
  assign n5407 = INSTQUEUE_REG_5__1_ & n5284;
  assign n5408 = INSTQUEUE_REG_6__1_ & n5286;
  assign n5409 = INSTQUEUE_REG_7__1_ & n5288;
  assign n5410 = ~n5406 & ~n5407;
  assign n5411 = ~n5408 & n5410;
  assign n5412 = ~n5409 & n5411;
  assign n5413 = INSTQUEUE_REG_8__1_ & n5294;
  assign n5414 = INSTQUEUE_REG_9__1_ & n5296;
  assign n5415 = INSTQUEUE_REG_10__1_ & n5298;
  assign n5416 = INSTQUEUE_REG_11__1_ & n5300;
  assign n5417 = ~n5413 & ~n5414;
  assign n5418 = ~n5415 & n5417;
  assign n5419 = ~n5416 & n5418;
  assign n5420 = INSTQUEUE_REG_12__1_ & n5306;
  assign n5421 = INSTQUEUE_REG_13__1_ & n5308;
  assign n5422 = INSTQUEUE_REG_14__1_ & n5310;
  assign n5423 = INSTQUEUE_REG_15__1_ & n5312;
  assign n5424 = ~n5420 & ~n5421;
  assign n5425 = ~n5422 & n5424;
  assign n5426 = ~n5423 & n5425;
  assign n5427 = n5405 & n5412;
  assign n5428 = n5419 & n5427;
  assign n5429 = n5426 & n5428;
  assign n5430 = ~n5320 & ~n5429;
  assign n5431 = ~n2781 & n5430;
  assign n5432 = n2781 & ~n5430;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n5337 & ~n5433;
  assign n5435 = n5337 & n5433;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = n2234 & ~n5436;
  assign n5438 = ~INSTADDRPOINTER_REG_9_ & ~n5437;
  assign n5439 = INSTADDRPOINTER_REG_9_ & n5437;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = ~n5342 & ~n5359;
  assign n5442 = ~n5343 & ~n5441;
  assign n5443 = n5440 & ~n5442;
  assign n5444 = ~n5440 & n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n4667 & n5445;
  assign n5447 = n5389 & n5398;
  assign n1280 = n5446 | ~n5447;
  assign n5449 = INSTADDRPOINTER_REG_9_ & n5367;
  assign n5450 = ~INSTADDRPOINTER_REG_10_ & n5449;
  assign n5451 = INSTADDRPOINTER_REG_10_ & ~n5449;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = n4677 & ~n5452;
  assign n5454 = EBX_REG_10_ & ~n4682;
  assign n5455 = INSTADDRPOINTER_REG_10_ & ~n4684;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = ~n2264 & ~n5456;
  assign n5458 = n2264 & n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = ~n5243 & ~n5377;
  assign n5461 = n5245 & n5460;
  assign n5462 = ~n5459 & ~n5461;
  assign n5463 = n5459 & n5461;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = n4695 & ~n5464;
  assign n5466 = INSTADDRPOINTER_REG_9_ & n5383;
  assign n5467 = ~INSTADDRPOINTER_REG_10_ & n5466;
  assign n5468 = INSTADDRPOINTER_REG_10_ & ~n5466;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = n4646 & ~n5469;
  assign n5471 = ~n5453 & ~n5465;
  assign n5472 = ~n5470 & n5471;
  assign n5473 = REIP_REG_10_ & n4698;
  assign n5474 = INSTADDRPOINTER_REG_10_ & n4644;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = INSTADDRPOINTER_REG_9_ & n5393;
  assign n5477 = ~INSTADDRPOINTER_REG_10_ & n5476;
  assign n5478 = INSTADDRPOINTER_REG_10_ & ~n5476;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = n4702 & ~n5479;
  assign n5481 = n5475 & ~n5480;
  assign n5482 = INSTQUEUE_REG_0__2_ & n5270;
  assign n5483 = INSTQUEUE_REG_1__2_ & n5272;
  assign n5484 = INSTQUEUE_REG_2__2_ & n5274;
  assign n5485 = INSTQUEUE_REG_3__2_ & n5276;
  assign n5486 = ~n5482 & ~n5483;
  assign n5487 = ~n5484 & n5486;
  assign n5488 = ~n5485 & n5487;
  assign n5489 = INSTQUEUE_REG_4__2_ & n5282;
  assign n5490 = INSTQUEUE_REG_5__2_ & n5284;
  assign n5491 = INSTQUEUE_REG_6__2_ & n5286;
  assign n5492 = INSTQUEUE_REG_7__2_ & n5288;
  assign n5493 = ~n5489 & ~n5490;
  assign n5494 = ~n5491 & n5493;
  assign n5495 = ~n5492 & n5494;
  assign n5496 = INSTQUEUE_REG_8__2_ & n5294;
  assign n5497 = INSTQUEUE_REG_9__2_ & n5296;
  assign n5498 = INSTQUEUE_REG_10__2_ & n5298;
  assign n5499 = INSTQUEUE_REG_11__2_ & n5300;
  assign n5500 = ~n5496 & ~n5497;
  assign n5501 = ~n5498 & n5500;
  assign n5502 = ~n5499 & n5501;
  assign n5503 = INSTQUEUE_REG_12__2_ & n5306;
  assign n5504 = INSTQUEUE_REG_13__2_ & n5308;
  assign n5505 = INSTQUEUE_REG_14__2_ & n5310;
  assign n5506 = INSTQUEUE_REG_15__2_ & n5312;
  assign n5507 = ~n5503 & ~n5504;
  assign n5508 = ~n5505 & n5507;
  assign n5509 = ~n5506 & n5508;
  assign n5510 = n5488 & n5495;
  assign n5511 = n5502 & n5510;
  assign n5512 = n5509 & n5511;
  assign n5513 = ~n5320 & ~n5512;
  assign n5514 = ~n2781 & n5513;
  assign n5515 = n2781 & ~n5513;
  assign n5516 = ~n5514 & ~n5515;
  assign n5517 = ~n5324 & ~n5433;
  assign n5518 = ~n5336 & n5517;
  assign n5519 = ~n5516 & ~n5518;
  assign n5520 = n5516 & n5518;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = n2234 & ~n5521;
  assign n5523 = INSTADDRPOINTER_REG_10_ & n5522;
  assign n5524 = ~INSTADDRPOINTER_REG_10_ & ~n5522;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = ~n5438 & ~n5442;
  assign n5527 = ~n5439 & ~n5526;
  assign n5528 = n5525 & ~n5527;
  assign n5529 = ~n5525 & n5527;
  assign n5530 = ~n5528 & ~n5529;
  assign n5531 = n4667 & n5530;
  assign n5532 = n5472 & n5481;
  assign n1285 = n5531 | ~n5532;
  assign n5534 = INSTADDRPOINTER_REG_9_ & INSTADDRPOINTER_REG_10_;
  assign n5535 = n5367 & n5534;
  assign n5536 = INSTADDRPOINTER_REG_11_ & ~n5535;
  assign n5537 = ~INSTADDRPOINTER_REG_11_ & n5535;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = n4677 & ~n5538;
  assign n5540 = EBX_REG_11_ & ~n4682;
  assign n5541 = INSTADDRPOINTER_REG_11_ & ~n4684;
  assign n5542 = ~n5540 & ~n5541;
  assign n5543 = ~n2264 & ~n5542;
  assign n5544 = n2264 & n5542;
  assign n5545 = ~n5543 & ~n5544;
  assign n5546 = ~n5459 & n5461;
  assign n5547 = ~n5545 & ~n5546;
  assign n5548 = n5545 & n5546;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = n4695 & ~n5549;
  assign n5551 = INSTADDRPOINTER_REG_10_ & n5466;
  assign n5552 = ~INSTADDRPOINTER_REG_11_ & n5551;
  assign n5553 = INSTADDRPOINTER_REG_11_ & ~n5551;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = n4646 & ~n5554;
  assign n5556 = ~n5539 & ~n5550;
  assign n5557 = ~n5555 & n5556;
  assign n5558 = REIP_REG_11_ & n4698;
  assign n5559 = INSTADDRPOINTER_REG_11_ & n4644;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = INSTADDRPOINTER_REG_10_ & n5476;
  assign n5562 = ~INSTADDRPOINTER_REG_11_ & n5561;
  assign n5563 = INSTADDRPOINTER_REG_11_ & ~n5561;
  assign n5564 = ~n5562 & ~n5563;
  assign n5565 = n4702 & ~n5564;
  assign n5566 = n5560 & ~n5565;
  assign n5567 = INSTQUEUE_REG_0__3_ & n5270;
  assign n5568 = INSTQUEUE_REG_1__3_ & n5272;
  assign n5569 = INSTQUEUE_REG_2__3_ & n5274;
  assign n5570 = INSTQUEUE_REG_3__3_ & n5276;
  assign n5571 = ~n5567 & ~n5568;
  assign n5572 = ~n5569 & n5571;
  assign n5573 = ~n5570 & n5572;
  assign n5574 = INSTQUEUE_REG_4__3_ & n5282;
  assign n5575 = INSTQUEUE_REG_5__3_ & n5284;
  assign n5576 = INSTQUEUE_REG_6__3_ & n5286;
  assign n5577 = INSTQUEUE_REG_7__3_ & n5288;
  assign n5578 = ~n5574 & ~n5575;
  assign n5579 = ~n5576 & n5578;
  assign n5580 = ~n5577 & n5579;
  assign n5581 = INSTQUEUE_REG_8__3_ & n5294;
  assign n5582 = INSTQUEUE_REG_9__3_ & n5296;
  assign n5583 = INSTQUEUE_REG_10__3_ & n5298;
  assign n5584 = INSTQUEUE_REG_11__3_ & n5300;
  assign n5585 = ~n5581 & ~n5582;
  assign n5586 = ~n5583 & n5585;
  assign n5587 = ~n5584 & n5586;
  assign n5588 = INSTQUEUE_REG_12__3_ & n5306;
  assign n5589 = INSTQUEUE_REG_13__3_ & n5308;
  assign n5590 = INSTQUEUE_REG_14__3_ & n5310;
  assign n5591 = INSTQUEUE_REG_15__3_ & n5312;
  assign n5592 = ~n5588 & ~n5589;
  assign n5593 = ~n5590 & n5592;
  assign n5594 = ~n5591 & n5593;
  assign n5595 = n5573 & n5580;
  assign n5596 = n5587 & n5595;
  assign n5597 = n5594 & n5596;
  assign n5598 = ~n5320 & ~n5597;
  assign n5599 = ~n2781 & n5598;
  assign n5600 = n2781 & ~n5598;
  assign n5601 = ~n5599 & ~n5600;
  assign n5602 = ~n5433 & ~n5516;
  assign n5603 = ~n5324 & n5602;
  assign n5604 = ~n5336 & n5603;
  assign n5605 = ~n5601 & ~n5604;
  assign n5606 = n5601 & n5604;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = n2234 & ~n5607;
  assign n5609 = ~INSTADDRPOINTER_REG_11_ & ~n5608;
  assign n5610 = INSTADDRPOINTER_REG_11_ & n5608;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = ~n5524 & ~n5527;
  assign n5613 = ~n5523 & ~n5612;
  assign n5614 = n5611 & ~n5613;
  assign n5615 = ~n5611 & n5613;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = n4667 & n5616;
  assign n5618 = n5557 & n5566;
  assign n1290 = n5617 | ~n5618;
  assign n5620 = INSTADDRPOINTER_REG_11_ & n5535;
  assign n5621 = ~INSTADDRPOINTER_REG_12_ & n5620;
  assign n5622 = INSTADDRPOINTER_REG_12_ & ~n5620;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = n4677 & ~n5623;
  assign n5625 = EBX_REG_12_ & ~n4682;
  assign n5626 = INSTADDRPOINTER_REG_12_ & ~n4684;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = ~n2264 & ~n5627;
  assign n5629 = n2264 & n5627;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = ~n5459 & ~n5545;
  assign n5632 = n5461 & n5631;
  assign n5633 = ~n5630 & ~n5632;
  assign n5634 = n5630 & n5632;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = n4695 & ~n5635;
  assign n5637 = INSTADDRPOINTER_REG_11_ & n5551;
  assign n5638 = ~INSTADDRPOINTER_REG_12_ & n5637;
  assign n5639 = INSTADDRPOINTER_REG_12_ & ~n5637;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = n4646 & ~n5640;
  assign n5642 = ~n5624 & ~n5636;
  assign n5643 = ~n5641 & n5642;
  assign n5644 = REIP_REG_12_ & n4698;
  assign n5645 = INSTADDRPOINTER_REG_12_ & n4644;
  assign n5646 = ~n5644 & ~n5645;
  assign n5647 = INSTADDRPOINTER_REG_11_ & n5561;
  assign n5648 = ~INSTADDRPOINTER_REG_12_ & n5647;
  assign n5649 = INSTADDRPOINTER_REG_12_ & ~n5647;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = n4702 & ~n5650;
  assign n5652 = n5646 & ~n5651;
  assign n5653 = INSTQUEUE_REG_0__4_ & n5270;
  assign n5654 = INSTQUEUE_REG_1__4_ & n5272;
  assign n5655 = INSTQUEUE_REG_2__4_ & n5274;
  assign n5656 = INSTQUEUE_REG_3__4_ & n5276;
  assign n5657 = ~n5653 & ~n5654;
  assign n5658 = ~n5655 & n5657;
  assign n5659 = ~n5656 & n5658;
  assign n5660 = INSTQUEUE_REG_4__4_ & n5282;
  assign n5661 = INSTQUEUE_REG_5__4_ & n5284;
  assign n5662 = INSTQUEUE_REG_6__4_ & n5286;
  assign n5663 = INSTQUEUE_REG_7__4_ & n5288;
  assign n5664 = ~n5660 & ~n5661;
  assign n5665 = ~n5662 & n5664;
  assign n5666 = ~n5663 & n5665;
  assign n5667 = INSTQUEUE_REG_8__4_ & n5294;
  assign n5668 = INSTQUEUE_REG_9__4_ & n5296;
  assign n5669 = INSTQUEUE_REG_10__4_ & n5298;
  assign n5670 = INSTQUEUE_REG_11__4_ & n5300;
  assign n5671 = ~n5667 & ~n5668;
  assign n5672 = ~n5669 & n5671;
  assign n5673 = ~n5670 & n5672;
  assign n5674 = INSTQUEUE_REG_12__4_ & n5306;
  assign n5675 = INSTQUEUE_REG_13__4_ & n5308;
  assign n5676 = INSTQUEUE_REG_14__4_ & n5310;
  assign n5677 = INSTQUEUE_REG_15__4_ & n5312;
  assign n5678 = ~n5674 & ~n5675;
  assign n5679 = ~n5676 & n5678;
  assign n5680 = ~n5677 & n5679;
  assign n5681 = n5659 & n5666;
  assign n5682 = n5673 & n5681;
  assign n5683 = n5680 & n5682;
  assign n5684 = ~n5320 & ~n5683;
  assign n5685 = ~n2781 & n5684;
  assign n5686 = n2781 & ~n5684;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = ~n5516 & ~n5601;
  assign n5689 = ~n5433 & n5688;
  assign n5690 = ~n5324 & n5689;
  assign n5691 = ~n5336 & n5690;
  assign n5692 = ~n5687 & ~n5691;
  assign n5693 = n5687 & n5691;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = n2234 & ~n5694;
  assign n5696 = ~INSTADDRPOINTER_REG_12_ & ~n5695;
  assign n5697 = INSTADDRPOINTER_REG_12_ & n5695;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = ~n5524 & ~n5609;
  assign n5700 = ~n5342 & ~n5438;
  assign n5701 = n5699 & n5700;
  assign n5702 = ~n5223 & ~n5348;
  assign n5703 = ~n5356 & n5702;
  assign n5704 = ~n5346 & ~n5353;
  assign n5705 = n5703 & n5704;
  assign n5706 = n5701 & ~n5705;
  assign n5707 = n5343 & ~n5438;
  assign n5708 = n5699 & n5707;
  assign n5709 = n5523 & n5699;
  assign n5710 = n5439 & n5699;
  assign n5711 = ~n5610 & ~n5708;
  assign n5712 = ~n5709 & n5711;
  assign n5713 = ~n5710 & n5712;
  assign n5714 = ~n5706 & n5713;
  assign n5715 = n5698 & ~n5714;
  assign n5716 = ~n5698 & n5714;
  assign n5717 = ~n5715 & ~n5716;
  assign n5718 = n4667 & n5717;
  assign n5719 = n5643 & n5652;
  assign n1295 = n5718 | ~n5719;
  assign n5721 = REIP_REG_13_ & n4698;
  assign n5722 = INSTADDRPOINTER_REG_13_ & n4644;
  assign n5723 = ~n5721 & ~n5722;
  assign n5724 = INSTADDRPOINTER_REG_12_ & n5647;
  assign n5725 = ~INSTADDRPOINTER_REG_13_ & n5724;
  assign n5726 = INSTADDRPOINTER_REG_13_ & ~n5724;
  assign n5727 = ~n5725 & ~n5726;
  assign n5728 = n4702 & ~n5727;
  assign n5729 = n5723 & ~n5728;
  assign n5730 = INSTADDRPOINTER_REG_11_ & INSTADDRPOINTER_REG_12_;
  assign n5731 = n5535 & n5730;
  assign n5732 = INSTADDRPOINTER_REG_13_ & ~n5731;
  assign n5733 = ~INSTADDRPOINTER_REG_13_ & n5731;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = n4677 & ~n5734;
  assign n5736 = INSTADDRPOINTER_REG_12_ & n5637;
  assign n5737 = ~INSTADDRPOINTER_REG_13_ & n5736;
  assign n5738 = INSTADDRPOINTER_REG_13_ & ~n5736;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = n4646 & ~n5739;
  assign n5741 = ~n5735 & ~n5740;
  assign n5742 = EBX_REG_13_ & ~n4682;
  assign n5743 = INSTADDRPOINTER_REG_13_ & ~n4684;
  assign n5744 = ~n5742 & ~n5743;
  assign n5745 = ~n2264 & ~n5744;
  assign n5746 = n2264 & n5744;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~n5630 & n5632;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = n5747 & n5748;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = n4695 & ~n5751;
  assign n5753 = INSTQUEUE_REG_0__5_ & n5270;
  assign n5754 = INSTQUEUE_REG_1__5_ & n5272;
  assign n5755 = INSTQUEUE_REG_2__5_ & n5274;
  assign n5756 = INSTQUEUE_REG_3__5_ & n5276;
  assign n5757 = ~n5753 & ~n5754;
  assign n5758 = ~n5755 & n5757;
  assign n5759 = ~n5756 & n5758;
  assign n5760 = INSTQUEUE_REG_4__5_ & n5282;
  assign n5761 = INSTQUEUE_REG_5__5_ & n5284;
  assign n5762 = INSTQUEUE_REG_6__5_ & n5286;
  assign n5763 = INSTQUEUE_REG_7__5_ & n5288;
  assign n5764 = ~n5760 & ~n5761;
  assign n5765 = ~n5762 & n5764;
  assign n5766 = ~n5763 & n5765;
  assign n5767 = INSTQUEUE_REG_8__5_ & n5294;
  assign n5768 = INSTQUEUE_REG_9__5_ & n5296;
  assign n5769 = INSTQUEUE_REG_10__5_ & n5298;
  assign n5770 = INSTQUEUE_REG_11__5_ & n5300;
  assign n5771 = ~n5767 & ~n5768;
  assign n5772 = ~n5769 & n5771;
  assign n5773 = ~n5770 & n5772;
  assign n5774 = INSTQUEUE_REG_12__5_ & n5306;
  assign n5775 = INSTQUEUE_REG_13__5_ & n5308;
  assign n5776 = INSTQUEUE_REG_14__5_ & n5310;
  assign n5777 = INSTQUEUE_REG_15__5_ & n5312;
  assign n5778 = ~n5774 & ~n5775;
  assign n5779 = ~n5776 & n5778;
  assign n5780 = ~n5777 & n5779;
  assign n5781 = n5759 & n5766;
  assign n5782 = n5773 & n5781;
  assign n5783 = n5780 & n5782;
  assign n5784 = ~n5320 & ~n5783;
  assign n5785 = ~n2781 & n5784;
  assign n5786 = n2781 & ~n5784;
  assign n5787 = ~n5785 & ~n5786;
  assign n5788 = ~n5687 & n5691;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = n5787 & n5788;
  assign n5791 = ~n5789 & ~n5790;
  assign n5792 = n2234 & ~n5791;
  assign n5793 = ~INSTADDRPOINTER_REG_13_ & ~n5792;
  assign n5794 = INSTADDRPOINTER_REG_13_ & n5792;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = ~n5696 & ~n5714;
  assign n5797 = ~n5697 & ~n5796;
  assign n5798 = n5795 & ~n5797;
  assign n5799 = ~n5795 & n5797;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = n4667 & n5800;
  assign n5802 = n5729 & n5741;
  assign n5803 = ~n5752 & n5802;
  assign n1300 = n5801 | ~n5803;
  assign n5805 = REIP_REG_14_ & n4698;
  assign n5806 = INSTADDRPOINTER_REG_14_ & n4644;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = INSTADDRPOINTER_REG_13_ & n5724;
  assign n5809 = ~INSTADDRPOINTER_REG_14_ & n5808;
  assign n5810 = INSTADDRPOINTER_REG_14_ & ~n5808;
  assign n5811 = ~n5809 & ~n5810;
  assign n5812 = n4702 & ~n5811;
  assign n5813 = n5807 & ~n5812;
  assign n5814 = INSTADDRPOINTER_REG_13_ & n5731;
  assign n5815 = ~INSTADDRPOINTER_REG_14_ & n5814;
  assign n5816 = INSTADDRPOINTER_REG_14_ & ~n5814;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = n4677 & ~n5817;
  assign n5819 = INSTADDRPOINTER_REG_13_ & n5736;
  assign n5820 = ~INSTADDRPOINTER_REG_14_ & n5819;
  assign n5821 = INSTADDRPOINTER_REG_14_ & ~n5819;
  assign n5822 = ~n5820 & ~n5821;
  assign n5823 = n4646 & ~n5822;
  assign n5824 = ~n5818 & ~n5823;
  assign n5825 = EBX_REG_14_ & ~n4682;
  assign n5826 = INSTADDRPOINTER_REG_14_ & ~n4684;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~n2264 & ~n5827;
  assign n5829 = n2264 & n5827;
  assign n5830 = ~n5828 & ~n5829;
  assign n5831 = ~n5630 & ~n5747;
  assign n5832 = n5632 & n5831;
  assign n5833 = ~n5830 & ~n5832;
  assign n5834 = n5830 & n5832;
  assign n5835 = ~n5833 & ~n5834;
  assign n5836 = n4695 & ~n5835;
  assign n5837 = INSTQUEUE_REG_0__6_ & n5270;
  assign n5838 = INSTQUEUE_REG_1__6_ & n5272;
  assign n5839 = INSTQUEUE_REG_2__6_ & n5274;
  assign n5840 = INSTQUEUE_REG_3__6_ & n5276;
  assign n5841 = ~n5837 & ~n5838;
  assign n5842 = ~n5839 & n5841;
  assign n5843 = ~n5840 & n5842;
  assign n5844 = INSTQUEUE_REG_4__6_ & n5282;
  assign n5845 = INSTQUEUE_REG_5__6_ & n5284;
  assign n5846 = INSTQUEUE_REG_6__6_ & n5286;
  assign n5847 = INSTQUEUE_REG_7__6_ & n5288;
  assign n5848 = ~n5844 & ~n5845;
  assign n5849 = ~n5846 & n5848;
  assign n5850 = ~n5847 & n5849;
  assign n5851 = INSTQUEUE_REG_8__6_ & n5294;
  assign n5852 = INSTQUEUE_REG_9__6_ & n5296;
  assign n5853 = INSTQUEUE_REG_10__6_ & n5298;
  assign n5854 = INSTQUEUE_REG_11__6_ & n5300;
  assign n5855 = ~n5851 & ~n5852;
  assign n5856 = ~n5853 & n5855;
  assign n5857 = ~n5854 & n5856;
  assign n5858 = INSTQUEUE_REG_12__6_ & n5306;
  assign n5859 = INSTQUEUE_REG_13__6_ & n5308;
  assign n5860 = INSTQUEUE_REG_14__6_ & n5310;
  assign n5861 = INSTQUEUE_REG_15__6_ & n5312;
  assign n5862 = ~n5858 & ~n5859;
  assign n5863 = ~n5860 & n5862;
  assign n5864 = ~n5861 & n5863;
  assign n5865 = n5843 & n5850;
  assign n5866 = n5857 & n5865;
  assign n5867 = n5864 & n5866;
  assign n5868 = ~n5320 & ~n5867;
  assign n5869 = ~n2781 & n5868;
  assign n5870 = n2781 & ~n5868;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = ~n5687 & ~n5787;
  assign n5873 = n5691 & n5872;
  assign n5874 = ~n5871 & ~n5873;
  assign n5875 = n5871 & n5873;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = n2234 & ~n5876;
  assign n5878 = INSTADDRPOINTER_REG_14_ & n5877;
  assign n5879 = ~INSTADDRPOINTER_REG_14_ & ~n5877;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~n5793 & ~n5797;
  assign n5882 = ~n5794 & ~n5881;
  assign n5883 = n5880 & ~n5882;
  assign n5884 = ~n5880 & n5882;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = n4667 & n5885;
  assign n5887 = n5813 & n5824;
  assign n5888 = ~n5836 & n5887;
  assign n1305 = n5886 | ~n5888;
  assign n5890 = REIP_REG_15_ & n4698;
  assign n5891 = INSTADDRPOINTER_REG_15_ & n4644;
  assign n5892 = ~n5890 & ~n5891;
  assign n5893 = INSTADDRPOINTER_REG_14_ & n5808;
  assign n5894 = ~INSTADDRPOINTER_REG_15_ & n5893;
  assign n5895 = INSTADDRPOINTER_REG_15_ & ~n5893;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = n4702 & ~n5896;
  assign n5898 = n5892 & ~n5897;
  assign n5899 = INSTADDRPOINTER_REG_13_ & INSTADDRPOINTER_REG_14_;
  assign n5900 = n5731 & n5899;
  assign n5901 = INSTADDRPOINTER_REG_15_ & ~n5900;
  assign n5902 = ~INSTADDRPOINTER_REG_15_ & n5900;
  assign n5903 = ~n5901 & ~n5902;
  assign n5904 = n4677 & ~n5903;
  assign n5905 = INSTADDRPOINTER_REG_14_ & n5819;
  assign n5906 = ~INSTADDRPOINTER_REG_15_ & n5905;
  assign n5907 = INSTADDRPOINTER_REG_15_ & ~n5905;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = n4646 & ~n5908;
  assign n5910 = ~n5904 & ~n5909;
  assign n5911 = EBX_REG_15_ & ~n4682;
  assign n5912 = INSTADDRPOINTER_REG_15_ & ~n4684;
  assign n5913 = ~n5911 & ~n5912;
  assign n5914 = ~n2264 & ~n5913;
  assign n5915 = n2264 & n5913;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = ~n5830 & n5832;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = n5916 & n5917;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = n4695 & ~n5920;
  assign n5922 = INSTQUEUE_REG_0__7_ & n5270;
  assign n5923 = INSTQUEUE_REG_1__7_ & n5272;
  assign n5924 = INSTQUEUE_REG_2__7_ & n5274;
  assign n5925 = INSTQUEUE_REG_3__7_ & n5276;
  assign n5926 = ~n5922 & ~n5923;
  assign n5927 = ~n5924 & n5926;
  assign n5928 = ~n5925 & n5927;
  assign n5929 = INSTQUEUE_REG_4__7_ & n5282;
  assign n5930 = INSTQUEUE_REG_5__7_ & n5284;
  assign n5931 = INSTQUEUE_REG_6__7_ & n5286;
  assign n5932 = INSTQUEUE_REG_7__7_ & n5288;
  assign n5933 = ~n5929 & ~n5930;
  assign n5934 = ~n5931 & n5933;
  assign n5935 = ~n5932 & n5934;
  assign n5936 = INSTQUEUE_REG_8__7_ & n5294;
  assign n5937 = INSTQUEUE_REG_9__7_ & n5296;
  assign n5938 = INSTQUEUE_REG_10__7_ & n5298;
  assign n5939 = INSTQUEUE_REG_11__7_ & n5300;
  assign n5940 = ~n5936 & ~n5937;
  assign n5941 = ~n5938 & n5940;
  assign n5942 = ~n5939 & n5941;
  assign n5943 = INSTQUEUE_REG_12__7_ & n5306;
  assign n5944 = INSTQUEUE_REG_13__7_ & n5308;
  assign n5945 = INSTQUEUE_REG_14__7_ & n5310;
  assign n5946 = INSTQUEUE_REG_15__7_ & n5312;
  assign n5947 = ~n5943 & ~n5944;
  assign n5948 = ~n5945 & n5947;
  assign n5949 = ~n5946 & n5948;
  assign n5950 = n5928 & n5935;
  assign n5951 = n5942 & n5950;
  assign n5952 = n5949 & n5951;
  assign n5953 = ~n5320 & ~n5952;
  assign n5954 = ~n2781 & n5953;
  assign n5955 = n2781 & ~n5953;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~n5871 & n5873;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = n5956 & n5957;
  assign n5960 = ~n5958 & ~n5959;
  assign n5961 = n2234 & ~n5960;
  assign n5962 = ~INSTADDRPOINTER_REG_15_ & ~n5961;
  assign n5963 = INSTADDRPOINTER_REG_15_ & n5961;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = ~n5879 & ~n5882;
  assign n5966 = ~n5878 & ~n5965;
  assign n5967 = n5964 & ~n5966;
  assign n5968 = ~n5964 & n5966;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = n4667 & n5969;
  assign n5971 = n5898 & n5910;
  assign n5972 = ~n5921 & n5971;
  assign n1310 = n5970 | ~n5972;
  assign n5974 = REIP_REG_16_ & n4698;
  assign n5975 = INSTADDRPOINTER_REG_16_ & n4644;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = INSTADDRPOINTER_REG_15_ & n5893;
  assign n5978 = ~INSTADDRPOINTER_REG_16_ & n5977;
  assign n5979 = INSTADDRPOINTER_REG_16_ & ~n5977;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = n4702 & ~n5980;
  assign n5982 = n5976 & ~n5981;
  assign n5983 = INSTADDRPOINTER_REG_15_ & n5900;
  assign n5984 = ~INSTADDRPOINTER_REG_16_ & n5983;
  assign n5985 = INSTADDRPOINTER_REG_16_ & ~n5983;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = n4677 & ~n5986;
  assign n5988 = INSTADDRPOINTER_REG_15_ & n5905;
  assign n5989 = ~INSTADDRPOINTER_REG_16_ & n5988;
  assign n5990 = INSTADDRPOINTER_REG_16_ & ~n5988;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = n4646 & ~n5991;
  assign n5993 = ~n5987 & ~n5992;
  assign n5994 = EBX_REG_16_ & ~n4682;
  assign n5995 = INSTADDRPOINTER_REG_16_ & ~n4684;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n2264 & ~n5996;
  assign n5998 = n2264 & n5996;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~n5830 & ~n5916;
  assign n6001 = n5832 & n6000;
  assign n6002 = ~n5999 & ~n6001;
  assign n6003 = n5999 & n6001;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = n4695 & ~n6004;
  assign n6006 = n5872 & ~n5956;
  assign n6007 = ~n5871 & n6006;
  assign n6008 = n5690 & n6007;
  assign n6009 = ~n5336 & n6008;
  assign n6010 = n2781 & ~n6009;
  assign n6011 = ~n2781 & n6009;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = n2234 & ~n6012;
  assign n6014 = ~INSTADDRPOINTER_REG_16_ & ~n6013;
  assign n6015 = INSTADDRPOINTER_REG_16_ & n6013;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = ~n5793 & ~n5879;
  assign n6018 = ~n5696 & n6017;
  assign n6019 = ~n5962 & n6018;
  assign n6020 = ~n5714 & n6019;
  assign n6021 = n5697 & ~n5793;
  assign n6022 = ~n5879 & n6021;
  assign n6023 = ~n5962 & n6022;
  assign n6024 = n5794 & ~n5879;
  assign n6025 = ~n5962 & n6024;
  assign n6026 = n5878 & ~n5962;
  assign n6027 = ~n5963 & ~n6023;
  assign n6028 = ~n6025 & n6027;
  assign n6029 = ~n6026 & n6028;
  assign n6030 = ~n6020 & n6029;
  assign n6031 = n6016 & ~n6030;
  assign n6032 = ~n6016 & n6030;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = n4667 & n6033;
  assign n6035 = n5982 & n5993;
  assign n6036 = ~n6005 & n6035;
  assign n1315 = n6034 | ~n6036;
  assign n6038 = REIP_REG_17_ & n4698;
  assign n6039 = INSTADDRPOINTER_REG_17_ & n4644;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = INSTADDRPOINTER_REG_16_ & n5977;
  assign n6042 = ~INSTADDRPOINTER_REG_17_ & n6041;
  assign n6043 = INSTADDRPOINTER_REG_17_ & ~n6041;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = n4702 & ~n6044;
  assign n6046 = n6040 & ~n6045;
  assign n6047 = INSTADDRPOINTER_REG_15_ & INSTADDRPOINTER_REG_16_;
  assign n6048 = n5900 & n6047;
  assign n6049 = INSTADDRPOINTER_REG_17_ & ~n6048;
  assign n6050 = ~INSTADDRPOINTER_REG_17_ & n6048;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = n4677 & ~n6051;
  assign n6053 = INSTADDRPOINTER_REG_16_ & n5988;
  assign n6054 = ~INSTADDRPOINTER_REG_17_ & n6053;
  assign n6055 = INSTADDRPOINTER_REG_17_ & ~n6053;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = n4646 & ~n6056;
  assign n6058 = ~n6052 & ~n6057;
  assign n6059 = EBX_REG_17_ & ~n4682;
  assign n6060 = INSTADDRPOINTER_REG_17_ & ~n4684;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~n2264 & ~n6061;
  assign n6063 = n2264 & n6061;
  assign n6064 = ~n6062 & ~n6063;
  assign n6065 = ~n5999 & n6001;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = n6064 & n6065;
  assign n6068 = ~n6066 & ~n6067;
  assign n6069 = n4695 & ~n6068;
  assign n6070 = ~n6014 & ~n6030;
  assign n6071 = ~n6015 & ~n6070;
  assign n6072 = n2234 & n6010;
  assign n6073 = ~INSTADDRPOINTER_REG_17_ & ~n6072;
  assign n6074 = INSTADDRPOINTER_REG_17_ & n6072;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = n6071 & ~n6075;
  assign n6077 = ~n6071 & n6075;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = n4667 & n6078;
  assign n6080 = n6046 & n6058;
  assign n6081 = ~n6069 & n6080;
  assign n1320 = n6079 | ~n6081;
  assign n6083 = REIP_REG_18_ & n4698;
  assign n6084 = INSTADDRPOINTER_REG_18_ & n4644;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = INSTADDRPOINTER_REG_17_ & n6041;
  assign n6087 = ~INSTADDRPOINTER_REG_18_ & n6086;
  assign n6088 = INSTADDRPOINTER_REG_18_ & ~n6086;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = n4702 & ~n6089;
  assign n6091 = n6085 & ~n6090;
  assign n6092 = INSTADDRPOINTER_REG_17_ & n6048;
  assign n6093 = ~INSTADDRPOINTER_REG_18_ & n6092;
  assign n6094 = INSTADDRPOINTER_REG_18_ & ~n6092;
  assign n6095 = ~n6093 & ~n6094;
  assign n6096 = n4677 & ~n6095;
  assign n6097 = INSTADDRPOINTER_REG_17_ & n6053;
  assign n6098 = ~INSTADDRPOINTER_REG_18_ & n6097;
  assign n6099 = INSTADDRPOINTER_REG_18_ & ~n6097;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = n4646 & ~n6100;
  assign n6102 = ~n6096 & ~n6101;
  assign n6103 = EBX_REG_18_ & ~n4682;
  assign n6104 = INSTADDRPOINTER_REG_18_ & ~n4684;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = ~n2264 & ~n6105;
  assign n6107 = n2264 & n6105;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n5999 & ~n6064;
  assign n6110 = n6001 & n6109;
  assign n6111 = ~n6108 & ~n6110;
  assign n6112 = n6108 & n6110;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = n4695 & ~n6113;
  assign n6115 = n6015 & ~n6073;
  assign n6116 = ~n6074 & ~n6115;
  assign n6117 = ~n6014 & ~n6073;
  assign n6118 = ~n6030 & n6117;
  assign n6119 = n6116 & ~n6118;
  assign n6120 = ~INSTADDRPOINTER_REG_18_ & ~n6072;
  assign n6121 = INSTADDRPOINTER_REG_18_ & n6072;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = n6119 & ~n6122;
  assign n6124 = ~n6119 & n6122;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = n4667 & n6125;
  assign n6127 = n6091 & n6102;
  assign n6128 = ~n6114 & n6127;
  assign n1325 = n6126 | ~n6128;
  assign n6130 = REIP_REG_19_ & n4698;
  assign n6131 = INSTADDRPOINTER_REG_19_ & n4644;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = INSTADDRPOINTER_REG_18_ & n6086;
  assign n6134 = ~INSTADDRPOINTER_REG_19_ & n6133;
  assign n6135 = INSTADDRPOINTER_REG_19_ & ~n6133;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = n4702 & ~n6136;
  assign n6138 = n6132 & ~n6137;
  assign n6139 = INSTADDRPOINTER_REG_17_ & INSTADDRPOINTER_REG_18_;
  assign n6140 = n6048 & n6139;
  assign n6141 = INSTADDRPOINTER_REG_19_ & ~n6140;
  assign n6142 = ~INSTADDRPOINTER_REG_19_ & n6140;
  assign n6143 = ~n6141 & ~n6142;
  assign n6144 = n4677 & ~n6143;
  assign n6145 = INSTADDRPOINTER_REG_18_ & n6097;
  assign n6146 = ~INSTADDRPOINTER_REG_19_ & n6145;
  assign n6147 = INSTADDRPOINTER_REG_19_ & ~n6145;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = n4646 & ~n6148;
  assign n6150 = ~n6144 & ~n6149;
  assign n6151 = EBX_REG_19_ & ~n4682;
  assign n6152 = INSTADDRPOINTER_REG_19_ & ~n4684;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = ~n2264 & ~n6153;
  assign n6155 = n2264 & n6153;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = ~n6108 & n6110;
  assign n6158 = ~n6156 & ~n6157;
  assign n6159 = n6156 & n6157;
  assign n6160 = ~n6158 & ~n6159;
  assign n6161 = n4695 & ~n6160;
  assign n6162 = ~n6116 & ~n6120;
  assign n6163 = ~n6121 & ~n6162;
  assign n6164 = n6117 & ~n6120;
  assign n6165 = ~n6030 & n6164;
  assign n6166 = n6163 & ~n6165;
  assign n6167 = ~INSTADDRPOINTER_REG_19_ & ~n6072;
  assign n6168 = INSTADDRPOINTER_REG_19_ & n6072;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = n6166 & ~n6169;
  assign n6171 = ~n6166 & n6169;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = n4667 & n6172;
  assign n6174 = n6138 & n6150;
  assign n6175 = ~n6161 & n6174;
  assign n1330 = n6173 | ~n6175;
  assign n6177 = REIP_REG_20_ & n4698;
  assign n6178 = INSTADDRPOINTER_REG_20_ & n4644;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = INSTADDRPOINTER_REG_19_ & n6133;
  assign n6181 = ~INSTADDRPOINTER_REG_20_ & n6180;
  assign n6182 = INSTADDRPOINTER_REG_20_ & ~n6180;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = n4702 & ~n6183;
  assign n6185 = n6179 & ~n6184;
  assign n6186 = INSTADDRPOINTER_REG_19_ & n6140;
  assign n6187 = ~INSTADDRPOINTER_REG_20_ & n6186;
  assign n6188 = INSTADDRPOINTER_REG_20_ & ~n6186;
  assign n6189 = ~n6187 & ~n6188;
  assign n6190 = n4677 & ~n6189;
  assign n6191 = INSTADDRPOINTER_REG_19_ & n6145;
  assign n6192 = ~INSTADDRPOINTER_REG_20_ & n6191;
  assign n6193 = INSTADDRPOINTER_REG_20_ & ~n6191;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = n4646 & ~n6194;
  assign n6196 = ~n6190 & ~n6195;
  assign n6197 = EBX_REG_20_ & ~n4682;
  assign n6198 = INSTADDRPOINTER_REG_20_ & ~n4684;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n2264 & ~n6199;
  assign n6201 = n2264 & n6199;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = ~n6156 & n6157;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = n6202 & n6203;
  assign n6206 = ~n6204 & ~n6205;
  assign n6207 = n4695 & ~n6206;
  assign n6208 = ~n6163 & ~n6167;
  assign n6209 = ~n6168 & ~n6208;
  assign n6210 = n6164 & ~n6167;
  assign n6211 = ~n6030 & n6210;
  assign n6212 = n6209 & ~n6211;
  assign n6213 = ~INSTADDRPOINTER_REG_20_ & ~n6072;
  assign n6214 = INSTADDRPOINTER_REG_20_ & n6072;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = n6212 & ~n6215;
  assign n6217 = ~n6212 & n6215;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = n4667 & n6218;
  assign n6220 = n6185 & n6196;
  assign n6221 = ~n6207 & n6220;
  assign n1335 = n6219 | ~n6221;
  assign n6223 = REIP_REG_21_ & n4698;
  assign n6224 = INSTADDRPOINTER_REG_21_ & n4644;
  assign n6225 = ~n6223 & ~n6224;
  assign n6226 = INSTADDRPOINTER_REG_20_ & n6180;
  assign n6227 = ~INSTADDRPOINTER_REG_21_ & n6226;
  assign n6228 = INSTADDRPOINTER_REG_21_ & ~n6226;
  assign n6229 = ~n6227 & ~n6228;
  assign n6230 = n4702 & ~n6229;
  assign n6231 = n6225 & ~n6230;
  assign n6232 = INSTADDRPOINTER_REG_19_ & INSTADDRPOINTER_REG_20_;
  assign n6233 = n6140 & n6232;
  assign n6234 = INSTADDRPOINTER_REG_21_ & ~n6233;
  assign n6235 = ~INSTADDRPOINTER_REG_21_ & n6233;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = n4677 & ~n6236;
  assign n6238 = INSTADDRPOINTER_REG_20_ & n6191;
  assign n6239 = ~INSTADDRPOINTER_REG_21_ & n6238;
  assign n6240 = INSTADDRPOINTER_REG_21_ & ~n6238;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = n4646 & ~n6241;
  assign n6243 = ~n6237 & ~n6242;
  assign n6244 = EBX_REG_21_ & ~n4682;
  assign n6245 = INSTADDRPOINTER_REG_21_ & ~n4684;
  assign n6246 = ~n6244 & ~n6245;
  assign n6247 = ~n2264 & ~n6246;
  assign n6248 = n2264 & n6246;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = ~n6202 & n6203;
  assign n6251 = ~n6249 & ~n6250;
  assign n6252 = n6249 & n6250;
  assign n6253 = ~n6251 & ~n6252;
  assign n6254 = n4695 & ~n6253;
  assign n6255 = INSTADDRPOINTER_REG_21_ & n6072;
  assign n6256 = ~INSTADDRPOINTER_REG_21_ & ~n6072;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = ~n6212 & ~n6213;
  assign n6259 = ~n6214 & ~n6258;
  assign n6260 = n6257 & ~n6259;
  assign n6261 = ~n6257 & n6259;
  assign n6262 = ~n6260 & ~n6261;
  assign n6263 = n4667 & n6262;
  assign n6264 = n6231 & n6243;
  assign n6265 = ~n6254 & n6264;
  assign n1340 = n6263 | ~n6265;
  assign n6267 = REIP_REG_22_ & n4698;
  assign n6268 = INSTADDRPOINTER_REG_22_ & n4644;
  assign n6269 = ~n6267 & ~n6268;
  assign n6270 = INSTADDRPOINTER_REG_21_ & n6226;
  assign n6271 = ~INSTADDRPOINTER_REG_22_ & n6270;
  assign n6272 = INSTADDRPOINTER_REG_22_ & ~n6270;
  assign n6273 = ~n6271 & ~n6272;
  assign n6274 = n4702 & ~n6273;
  assign n6275 = n6269 & ~n6274;
  assign n6276 = INSTADDRPOINTER_REG_21_ & n6233;
  assign n6277 = ~INSTADDRPOINTER_REG_22_ & n6276;
  assign n6278 = INSTADDRPOINTER_REG_22_ & ~n6276;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = n4677 & ~n6279;
  assign n6281 = INSTADDRPOINTER_REG_21_ & n6238;
  assign n6282 = ~INSTADDRPOINTER_REG_22_ & n6281;
  assign n6283 = INSTADDRPOINTER_REG_22_ & ~n6281;
  assign n6284 = ~n6282 & ~n6283;
  assign n6285 = n4646 & ~n6284;
  assign n6286 = ~n6280 & ~n6285;
  assign n6287 = EBX_REG_22_ & ~n4682;
  assign n6288 = INSTADDRPOINTER_REG_22_ & ~n4684;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~n2264 & ~n6289;
  assign n6291 = n2264 & n6289;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = ~n6249 & n6250;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = n6292 & n6293;
  assign n6296 = ~n6294 & ~n6295;
  assign n6297 = n4695 & ~n6296;
  assign n6298 = INSTADDRPOINTER_REG_22_ & n6072;
  assign n6299 = ~INSTADDRPOINTER_REG_22_ & ~n6072;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 = n6214 & ~n6256;
  assign n6302 = ~n6255 & ~n6301;
  assign n6303 = ~n6213 & ~n6256;
  assign n6304 = ~n6212 & n6303;
  assign n6305 = n6302 & ~n6304;
  assign n6306 = n6300 & ~n6305;
  assign n6307 = ~n6300 & n6305;
  assign n6308 = ~n6306 & ~n6307;
  assign n6309 = n4667 & n6308;
  assign n6310 = n6275 & n6286;
  assign n6311 = ~n6297 & n6310;
  assign n1345 = n6309 | ~n6311;
  assign n6313 = REIP_REG_23_ & n4698;
  assign n6314 = INSTADDRPOINTER_REG_23_ & n4644;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 = INSTADDRPOINTER_REG_22_ & n6270;
  assign n6317 = ~INSTADDRPOINTER_REG_23_ & n6316;
  assign n6318 = INSTADDRPOINTER_REG_23_ & ~n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n4702 & ~n6319;
  assign n6321 = n6315 & ~n6320;
  assign n6322 = INSTADDRPOINTER_REG_21_ & INSTADDRPOINTER_REG_22_;
  assign n6323 = n6233 & n6322;
  assign n6324 = INSTADDRPOINTER_REG_23_ & ~n6323;
  assign n6325 = ~INSTADDRPOINTER_REG_23_ & n6323;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = n4677 & ~n6326;
  assign n6328 = INSTADDRPOINTER_REG_22_ & n6281;
  assign n6329 = ~INSTADDRPOINTER_REG_23_ & n6328;
  assign n6330 = INSTADDRPOINTER_REG_23_ & ~n6328;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = n4646 & ~n6331;
  assign n6333 = ~n6327 & ~n6332;
  assign n6334 = EBX_REG_23_ & ~n4682;
  assign n6335 = INSTADDRPOINTER_REG_23_ & ~n4684;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n2264 & ~n6336;
  assign n6338 = n2264 & n6336;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = ~n6292 & n6293;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = n6339 & n6340;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = n4695 & ~n6343;
  assign n6345 = INSTADDRPOINTER_REG_23_ & n6072;
  assign n6346 = ~INSTADDRPOINTER_REG_23_ & ~n6072;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = ~n6299 & ~n6302;
  assign n6349 = ~n6298 & ~n6348;
  assign n6350 = ~n6299 & n6303;
  assign n6351 = ~n6212 & n6350;
  assign n6352 = n6349 & ~n6351;
  assign n6353 = n6347 & ~n6352;
  assign n6354 = ~n6347 & n6352;
  assign n6355 = ~n6353 & ~n6354;
  assign n6356 = n4667 & n6355;
  assign n6357 = n6321 & n6333;
  assign n6358 = ~n6344 & n6357;
  assign n1350 = n6356 | ~n6358;
  assign n6360 = REIP_REG_24_ & n4698;
  assign n6361 = INSTADDRPOINTER_REG_24_ & n4644;
  assign n6362 = ~n6360 & ~n6361;
  assign n6363 = INSTADDRPOINTER_REG_23_ & n6316;
  assign n6364 = ~INSTADDRPOINTER_REG_24_ & n6363;
  assign n6365 = INSTADDRPOINTER_REG_24_ & ~n6363;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = n4702 & ~n6366;
  assign n6368 = n6362 & ~n6367;
  assign n6369 = INSTADDRPOINTER_REG_23_ & n6323;
  assign n6370 = ~INSTADDRPOINTER_REG_24_ & n6369;
  assign n6371 = INSTADDRPOINTER_REG_24_ & ~n6369;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = n4677 & ~n6372;
  assign n6374 = INSTADDRPOINTER_REG_23_ & n6328;
  assign n6375 = ~INSTADDRPOINTER_REG_24_ & n6374;
  assign n6376 = INSTADDRPOINTER_REG_24_ & ~n6374;
  assign n6377 = ~n6375 & ~n6376;
  assign n6378 = n4646 & ~n6377;
  assign n6379 = ~n6373 & ~n6378;
  assign n6380 = EBX_REG_24_ & ~n4682;
  assign n6381 = INSTADDRPOINTER_REG_24_ & ~n4684;
  assign n6382 = ~n6380 & ~n6381;
  assign n6383 = ~n2264 & ~n6382;
  assign n6384 = n2264 & n6382;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6339 & n6340;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = n6385 & n6386;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = n4695 & ~n6389;
  assign n6391 = INSTADDRPOINTER_REG_24_ & n6072;
  assign n6392 = ~INSTADDRPOINTER_REG_24_ & ~n6072;
  assign n6393 = ~n6391 & ~n6392;
  assign n6394 = ~n6346 & ~n6349;
  assign n6395 = ~n6345 & ~n6394;
  assign n6396 = ~n6346 & n6350;
  assign n6397 = ~n6212 & n6396;
  assign n6398 = n6395 & ~n6397;
  assign n6399 = n6393 & ~n6398;
  assign n6400 = ~n6393 & n6398;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = n4667 & n6401;
  assign n6403 = n6368 & n6379;
  assign n6404 = ~n6390 & n6403;
  assign n1355 = n6402 | ~n6404;
  assign n6406 = REIP_REG_25_ & n4698;
  assign n6407 = INSTADDRPOINTER_REG_25_ & n4644;
  assign n6408 = ~n6406 & ~n6407;
  assign n6409 = INSTADDRPOINTER_REG_24_ & n6363;
  assign n6410 = ~INSTADDRPOINTER_REG_25_ & n6409;
  assign n6411 = INSTADDRPOINTER_REG_25_ & ~n6409;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = n4702 & ~n6412;
  assign n6414 = n6408 & ~n6413;
  assign n6415 = INSTADDRPOINTER_REG_23_ & INSTADDRPOINTER_REG_24_;
  assign n6416 = n6323 & n6415;
  assign n6417 = INSTADDRPOINTER_REG_25_ & ~n6416;
  assign n6418 = ~INSTADDRPOINTER_REG_25_ & n6416;
  assign n6419 = ~n6417 & ~n6418;
  assign n6420 = n4677 & ~n6419;
  assign n6421 = INSTADDRPOINTER_REG_24_ & n6374;
  assign n6422 = ~INSTADDRPOINTER_REG_25_ & n6421;
  assign n6423 = INSTADDRPOINTER_REG_25_ & ~n6421;
  assign n6424 = ~n6422 & ~n6423;
  assign n6425 = n4646 & ~n6424;
  assign n6426 = ~n6420 & ~n6425;
  assign n6427 = EBX_REG_25_ & ~n4682;
  assign n6428 = INSTADDRPOINTER_REG_25_ & ~n4684;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n2264 & ~n6429;
  assign n6431 = n2264 & n6429;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n6385 & n6386;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = n6432 & n6433;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = n4695 & ~n6436;
  assign n6438 = ~INSTADDRPOINTER_REG_25_ & ~n6072;
  assign n6439 = INSTADDRPOINTER_REG_25_ & n6072;
  assign n6440 = ~n6438 & ~n6439;
  assign n6441 = ~n6392 & ~n6395;
  assign n6442 = ~n6391 & ~n6441;
  assign n6443 = ~n6392 & n6396;
  assign n6444 = ~n6212 & n6443;
  assign n6445 = n6442 & ~n6444;
  assign n6446 = n6440 & ~n6445;
  assign n6447 = ~n6440 & n6445;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = n4667 & n6448;
  assign n6450 = n6414 & n6426;
  assign n6451 = ~n6437 & n6450;
  assign n1360 = n6449 | ~n6451;
  assign n6453 = REIP_REG_26_ & n4698;
  assign n6454 = INSTADDRPOINTER_REG_26_ & n4644;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = INSTADDRPOINTER_REG_25_ & n6409;
  assign n6457 = ~INSTADDRPOINTER_REG_26_ & n6456;
  assign n6458 = INSTADDRPOINTER_REG_26_ & ~n6456;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = n4702 & ~n6459;
  assign n6461 = n6455 & ~n6460;
  assign n6462 = INSTADDRPOINTER_REG_25_ & n6416;
  assign n6463 = ~INSTADDRPOINTER_REG_26_ & n6462;
  assign n6464 = INSTADDRPOINTER_REG_26_ & ~n6462;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = n4677 & ~n6465;
  assign n6467 = INSTADDRPOINTER_REG_25_ & n6421;
  assign n6468 = ~INSTADDRPOINTER_REG_26_ & n6467;
  assign n6469 = INSTADDRPOINTER_REG_26_ & ~n6467;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = n4646 & ~n6470;
  assign n6472 = ~n6466 & ~n6471;
  assign n6473 = EBX_REG_26_ & ~n4682;
  assign n6474 = INSTADDRPOINTER_REG_26_ & ~n4684;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~n2264 & ~n6475;
  assign n6477 = n2264 & n6475;
  assign n6478 = ~n6476 & ~n6477;
  assign n6479 = ~n6432 & n6433;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = n6478 & n6479;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = n4695 & ~n6482;
  assign n6484 = ~n6438 & n6443;
  assign n6485 = n6208 & n6484;
  assign n6486 = ~n6438 & ~n6442;
  assign n6487 = n6168 & n6484;
  assign n6488 = ~n6439 & ~n6487;
  assign n6489 = ~n6485 & ~n6486;
  assign n6490 = n6488 & n6489;
  assign n6491 = n6210 & n6484;
  assign n6492 = ~n6030 & n6491;
  assign n6493 = n6490 & ~n6492;
  assign n6494 = ~INSTADDRPOINTER_REG_26_ & ~n6072;
  assign n6495 = INSTADDRPOINTER_REG_26_ & n6072;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = n6493 & ~n6496;
  assign n6498 = ~n6493 & n6496;
  assign n6499 = ~n6497 & ~n6498;
  assign n6500 = n4667 & n6499;
  assign n6501 = n6461 & n6472;
  assign n6502 = ~n6483 & n6501;
  assign n1365 = n6500 | ~n6502;
  assign n6504 = REIP_REG_27_ & n4698;
  assign n6505 = INSTADDRPOINTER_REG_27_ & n4644;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = INSTADDRPOINTER_REG_26_ & n6456;
  assign n6508 = ~INSTADDRPOINTER_REG_27_ & n6507;
  assign n6509 = INSTADDRPOINTER_REG_27_ & ~n6507;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = n4702 & ~n6510;
  assign n6512 = n6506 & ~n6511;
  assign n6513 = INSTADDRPOINTER_REG_25_ & INSTADDRPOINTER_REG_26_;
  assign n6514 = n6416 & n6513;
  assign n6515 = INSTADDRPOINTER_REG_27_ & ~n6514;
  assign n6516 = ~INSTADDRPOINTER_REG_27_ & n6514;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = n4677 & ~n6517;
  assign n6519 = INSTADDRPOINTER_REG_26_ & n6467;
  assign n6520 = ~INSTADDRPOINTER_REG_27_ & n6519;
  assign n6521 = INSTADDRPOINTER_REG_27_ & ~n6519;
  assign n6522 = ~n6520 & ~n6521;
  assign n6523 = n4646 & ~n6522;
  assign n6524 = ~n6518 & ~n6523;
  assign n6525 = EBX_REG_27_ & ~n4682;
  assign n6526 = INSTADDRPOINTER_REG_27_ & ~n4684;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = ~n2264 & ~n6527;
  assign n6529 = n2264 & n6527;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = ~n6478 & n6479;
  assign n6532 = ~n6530 & ~n6531;
  assign n6533 = n6530 & n6531;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = n4695 & ~n6534;
  assign n6536 = ~INSTADDRPOINTER_REG_27_ & ~n6072;
  assign n6537 = INSTADDRPOINTER_REG_27_ & n6072;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = ~n6493 & ~n6494;
  assign n6540 = ~n6495 & ~n6539;
  assign n6541 = n6538 & ~n6540;
  assign n6542 = ~n6538 & n6540;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = n4667 & n6543;
  assign n6545 = n6512 & n6524;
  assign n6546 = ~n6535 & n6545;
  assign n1370 = n6544 | ~n6546;
  assign n6548 = REIP_REG_28_ & n4698;
  assign n6549 = INSTADDRPOINTER_REG_28_ & n4644;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = INSTADDRPOINTER_REG_27_ & n6507;
  assign n6552 = ~INSTADDRPOINTER_REG_28_ & n6551;
  assign n6553 = INSTADDRPOINTER_REG_28_ & ~n6551;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n4702 & ~n6554;
  assign n6556 = n6550 & ~n6555;
  assign n6557 = INSTADDRPOINTER_REG_27_ & n6514;
  assign n6558 = ~INSTADDRPOINTER_REG_28_ & n6557;
  assign n6559 = INSTADDRPOINTER_REG_28_ & ~n6557;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n4677 & ~n6560;
  assign n6562 = INSTADDRPOINTER_REG_27_ & n6519;
  assign n6563 = ~INSTADDRPOINTER_REG_28_ & n6562;
  assign n6564 = INSTADDRPOINTER_REG_28_ & ~n6562;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = n4646 & ~n6565;
  assign n6567 = ~n6561 & ~n6566;
  assign n6568 = EBX_REG_28_ & ~n4682;
  assign n6569 = INSTADDRPOINTER_REG_28_ & ~n4684;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n2264 & ~n6570;
  assign n6572 = n2264 & n6570;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = ~n6530 & n6531;
  assign n6575 = ~n6573 & ~n6574;
  assign n6576 = n6573 & n6574;
  assign n6577 = ~n6575 & ~n6576;
  assign n6578 = n4695 & ~n6577;
  assign n6579 = INSTADDRPOINTER_REG_28_ & ~n6072;
  assign n6580 = ~INSTADDRPOINTER_REG_28_ & n6072;
  assign n6581 = ~n6579 & ~n6580;
  assign n6582 = n6495 & ~n6536;
  assign n6583 = ~n6537 & ~n6582;
  assign n6584 = ~n6494 & ~n6536;
  assign n6585 = ~n6493 & n6584;
  assign n6586 = n6583 & ~n6585;
  assign n6587 = ~n6581 & ~n6586;
  assign n6588 = n6581 & n6586;
  assign n6589 = ~n6587 & ~n6588;
  assign n6590 = n4667 & n6589;
  assign n6591 = n6556 & n6567;
  assign n6592 = ~n6578 & n6591;
  assign n1375 = n6590 | ~n6592;
  assign n6594 = REIP_REG_29_ & n4698;
  assign n6595 = INSTADDRPOINTER_REG_29_ & n4644;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = INSTADDRPOINTER_REG_28_ & n6551;
  assign n6598 = ~INSTADDRPOINTER_REG_29_ & n6597;
  assign n6599 = INSTADDRPOINTER_REG_29_ & ~n6597;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = n4702 & ~n6600;
  assign n6602 = n6596 & ~n6601;
  assign n6603 = INSTADDRPOINTER_REG_27_ & INSTADDRPOINTER_REG_28_;
  assign n6604 = n6514 & n6603;
  assign n6605 = INSTADDRPOINTER_REG_29_ & ~n6604;
  assign n6606 = ~INSTADDRPOINTER_REG_29_ & n6604;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n4677 & ~n6607;
  assign n6609 = INSTADDRPOINTER_REG_28_ & n6562;
  assign n6610 = ~INSTADDRPOINTER_REG_29_ & n6609;
  assign n6611 = INSTADDRPOINTER_REG_29_ & ~n6609;
  assign n6612 = ~n6610 & ~n6611;
  assign n6613 = n4646 & ~n6612;
  assign n6614 = ~n6608 & ~n6613;
  assign n6615 = EBX_REG_29_ & ~n4682;
  assign n6616 = INSTADDRPOINTER_REG_29_ & ~n4684;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n2264 & ~n6617;
  assign n6619 = n2264 & n6617;
  assign n6620 = ~n6618 & ~n6619;
  assign n6621 = ~n6573 & n6574;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = n6620 & n6621;
  assign n6624 = ~n6622 & ~n6623;
  assign n6625 = n4695 & ~n6624;
  assign n6626 = INSTADDRPOINTER_REG_29_ & ~n6072;
  assign n6627 = ~INSTADDRPOINTER_REG_29_ & n6072;
  assign n6628 = ~n6626 & ~n6627;
  assign n6629 = ~INSTADDRPOINTER_REG_28_ & ~n6072;
  assign n6630 = ~n6583 & ~n6629;
  assign n6631 = INSTADDRPOINTER_REG_28_ & n6072;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = n6584 & ~n6629;
  assign n6634 = ~n6493 & n6633;
  assign n6635 = n6632 & ~n6634;
  assign n6636 = ~n6628 & ~n6635;
  assign n6637 = n6628 & n6635;
  assign n6638 = ~n6636 & ~n6637;
  assign n6639 = n4667 & n6638;
  assign n6640 = n6602 & n6614;
  assign n6641 = ~n6625 & n6640;
  assign n1380 = n6639 | ~n6641;
  assign n6643 = REIP_REG_30_ & n4698;
  assign n6644 = INSTADDRPOINTER_REG_30_ & n4644;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = INSTADDRPOINTER_REG_29_ & n6597;
  assign n6647 = ~INSTADDRPOINTER_REG_30_ & n6646;
  assign n6648 = INSTADDRPOINTER_REG_30_ & ~n6646;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = n4702 & ~n6649;
  assign n6651 = n6645 & ~n6650;
  assign n6652 = INSTADDRPOINTER_REG_29_ & n6604;
  assign n6653 = ~INSTADDRPOINTER_REG_30_ & n6652;
  assign n6654 = INSTADDRPOINTER_REG_30_ & ~n6652;
  assign n6655 = ~n6653 & ~n6654;
  assign n6656 = n4677 & ~n6655;
  assign n6657 = INSTADDRPOINTER_REG_29_ & n6609;
  assign n6658 = ~INSTADDRPOINTER_REG_30_ & n6657;
  assign n6659 = INSTADDRPOINTER_REG_30_ & ~n6657;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = n4646 & ~n6660;
  assign n6662 = ~n6656 & ~n6661;
  assign n6663 = EBX_REG_30_ & ~n4682;
  assign n6664 = INSTADDRPOINTER_REG_30_ & ~n4684;
  assign n6665 = ~n6663 & ~n6664;
  assign n6666 = ~n2264 & ~n6665;
  assign n6667 = n2264 & n6665;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = ~n6620 & n6621;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = n6668 & n6669;
  assign n6672 = ~n6670 & ~n6671;
  assign n6673 = n4695 & ~n6672;
  assign n6674 = INSTADDRPOINTER_REG_30_ & ~n6072;
  assign n6675 = ~INSTADDRPOINTER_REG_30_ & n6072;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = ~INSTADDRPOINTER_REG_29_ & ~n6072;
  assign n6678 = ~n6632 & ~n6677;
  assign n6679 = INSTADDRPOINTER_REG_29_ & n6072;
  assign n6680 = ~n6678 & ~n6679;
  assign n6681 = n6633 & ~n6677;
  assign n6682 = ~n6493 & n6681;
  assign n6683 = n6680 & ~n6682;
  assign n6684 = ~n6676 & ~n6683;
  assign n6685 = n6676 & n6683;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = n4667 & n6686;
  assign n6688 = n6651 & n6662;
  assign n6689 = ~n6673 & n6688;
  assign n1385 = n6687 | ~n6689;
  assign n6691 = REIP_REG_31_ & n4698;
  assign n6692 = INSTADDRPOINTER_REG_31_ & n4644;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = INSTADDRPOINTER_REG_30_ & n6646;
  assign n6695 = ~INSTADDRPOINTER_REG_31_ & n6694;
  assign n6696 = INSTADDRPOINTER_REG_31_ & ~n6694;
  assign n6697 = ~n6695 & ~n6696;
  assign n6698 = n4702 & ~n6697;
  assign n6699 = n6693 & ~n6698;
  assign n6700 = INSTADDRPOINTER_REG_30_ & n6652;
  assign n6701 = ~INSTADDRPOINTER_REG_31_ & n6700;
  assign n6702 = INSTADDRPOINTER_REG_31_ & ~n6700;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = n4677 & ~n6703;
  assign n6705 = INSTADDRPOINTER_REG_30_ & n6657;
  assign n6706 = ~INSTADDRPOINTER_REG_31_ & n6705;
  assign n6707 = INSTADDRPOINTER_REG_31_ & ~n6705;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = n4646 & ~n6708;
  assign n6710 = ~n6704 & ~n6709;
  assign n6711 = EBX_REG_31_ & ~n4682;
  assign n6712 = INSTADDRPOINTER_REG_31_ & ~n4684;
  assign n6713 = ~n6711 & ~n6712;
  assign n6714 = ~n2264 & ~n6713;
  assign n6715 = n2264 & n6713;
  assign n6716 = ~n6714 & ~n6715;
  assign n6717 = ~n6620 & ~n6668;
  assign n6718 = n6621 & n6717;
  assign n6719 = ~n6716 & ~n6718;
  assign n6720 = n6716 & n6718;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = n4695 & ~n6721;
  assign n6723 = INSTADDRPOINTER_REG_31_ & ~n6072;
  assign n6724 = ~INSTADDRPOINTER_REG_31_ & n6072;
  assign n6725 = ~n6723 & ~n6724;
  assign n6726 = ~INSTADDRPOINTER_REG_30_ & ~n6072;
  assign n6727 = ~n6680 & ~n6726;
  assign n6728 = INSTADDRPOINTER_REG_30_ & n6072;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = n6681 & ~n6726;
  assign n6731 = ~n6493 & n6730;
  assign n6732 = n6729 & ~n6731;
  assign n6733 = ~n6725 & ~n6732;
  assign n6734 = n6725 & n6732;
  assign n6735 = ~n6733 & ~n6734;
  assign n6736 = n4667 & n6735;
  assign n6737 = n6699 & n6710;
  assign n6738 = ~n6722 & n6737;
  assign n1390 = n6736 | ~n6738;
  assign n6740 = ~STATE2_REG_0_ & n2724;
  assign n6741 = ~n2406 & ~n6740;
  assign n6742 = STATE2_REG_2_ & n2338_1;
  assign n6743 = ~STATE2_REG_1_ & ~n1839;
  assign n6744 = n2100 & n6743;
  assign n6745 = n2148_1 & n6742;
  assign n6746 = n6744 & n6745;
  assign n6747 = n2277 & n6746;
  assign n6748 = n6741 & ~n6747;
  assign n6749 = STATE2_REG_0_ & ~n6748;
  assign n6750 = n4655 & n6749;
  assign n6751 = STATE2_REG_1_ & ~STATEBS16_REG;
  assign n6752 = STATE2_REG_2_ & ~STATE2_REG_0_;
  assign n6753 = ~n6751 & ~n6752;
  assign n6754 = ~n6748 & ~n6753;
  assign n6755 = PHYADDRPOINTER_REG_0_ & n6754;
  assign n6756 = n2689 & ~n6748;
  assign n6757 = REIP_REG_0_ & n6756;
  assign n6758 = PHYADDRPOINTER_REG_0_ & n6748;
  assign n6759 = STATE2_REG_2_ & n1929;
  assign n6760 = n1898_1 & ~n6759;
  assign n6761 = n2884 & n6760;
  assign n6762 = STATE2_REG_2_ & ~n6761;
  assign n6763 = ~STATE2_REG_2_ & STATEBS16_REG;
  assign n6764 = PHYADDRPOINTER_REG_0_ & n6763;
  assign n6765 = STATE2_REG_2_ & n1898_1;
  assign n6766 = ~n4657 & ~n6765;
  assign n6767 = ~n2618 & ~n6766;
  assign n6768 = EAX_REG_0_ & n6759;
  assign n6769 = INSTQUEUERD_ADDR_REG_0_ & n6742;
  assign n6770 = PHYADDRPOINTER_REG_0_ & n2682;
  assign n6771 = ~n6764 & ~n6767;
  assign n6772 = ~n6768 & n6771;
  assign n6773 = ~n6769 & n6772;
  assign n6774 = ~n6770 & n6773;
  assign n6775 = ~n2682 & ~n6774;
  assign n6776 = n2682 & n6774;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = n6762 & ~n6777;
  assign n6779 = ~n6762 & n6777;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = ~n2682 & n6780;
  assign n6782 = n2682 & ~n6780;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = STATE2_REG_1_ & STATEBS16_REG;
  assign n6785 = ~n6748 & n6784;
  assign n6786 = ~n6783 & n6785;
  assign n6787 = ~n6750 & ~n6755;
  assign n6788 = ~n6757 & n6787;
  assign n6789 = ~n6758 & n6788;
  assign n1395 = n6786 | ~n6789;
  assign n6791 = ~n4723 & n6749;
  assign n6792 = ~PHYADDRPOINTER_REG_1_ & n6754;
  assign n6793 = REIP_REG_1_ & n6756;
  assign n6794 = PHYADDRPOINTER_REG_1_ & n6748;
  assign n6795 = ~n2880 & ~n6766;
  assign n6796 = INSTQUEUERD_ADDR_REG_1_ & n6742;
  assign n6797 = ~PHYADDRPOINTER_REG_1_ & n2682;
  assign n6798 = EAX_REG_1_ & n6759;
  assign n6799 = PHYADDRPOINTER_REG_1_ & n6763;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = ~n2633 & ~n6766;
  assign n6802 = ~n6796 & ~n6797;
  assign n6803 = n6800 & n6802;
  assign n6804 = ~n6801 & n6803;
  assign n6805 = ~n2682 & ~n6804;
  assign n6806 = n2682 & n6804;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = n6795 & ~n6807;
  assign n6809 = ~n6795 & n6807;
  assign n6810 = ~n6808 & ~n6809;
  assign n6811 = n2682 & ~n6779;
  assign n6812 = ~n6778 & ~n6811;
  assign n6813 = n6810 & n6812;
  assign n6814 = ~n6810 & ~n6812;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = n6785 & ~n6815;
  assign n6817 = ~n6791 & ~n6792;
  assign n6818 = ~n6793 & n6817;
  assign n6819 = ~n6794 & n6818;
  assign n1400 = n6816 | ~n6819;
  assign n6821 = REIP_REG_2_ & n6756;
  assign n6822 = ~PHYADDRPOINTER_REG_1_ & PHYADDRPOINTER_REG_2_;
  assign n6823 = PHYADDRPOINTER_REG_1_ & ~PHYADDRPOINTER_REG_2_;
  assign n6824 = ~n6822 & ~n6823;
  assign n6825 = n6754 & ~n6824;
  assign n6826 = n4771 & n6749;
  assign n6827 = PHYADDRPOINTER_REG_2_ & n6748;
  assign n6828 = ~n6809 & ~n6812;
  assign n6829 = ~n6808 & ~n6828;
  assign n6830 = INSTQUEUERD_ADDR_REG_2_ & n6742;
  assign n6831 = n2682 & ~n6824;
  assign n6832 = EAX_REG_2_ & n6759;
  assign n6833 = PHYADDRPOINTER_REG_2_ & n6763;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = n2495 & ~n6766;
  assign n6836 = ~n6830 & ~n6831;
  assign n6837 = n6834 & n6836;
  assign n6838 = ~n6835 & n6837;
  assign n6839 = ~n2682 & ~n6838;
  assign n6840 = n2682 & n6838;
  assign n6841 = ~n2941 & ~n6766;
  assign n6842 = ~n6763 & ~n6841;
  assign n6843 = ~n6839 & ~n6840;
  assign n6844 = n6842 & n6843;
  assign n6845 = ~n6829 & ~n6844;
  assign n6846 = ~n6842 & ~n6843;
  assign n6847 = n6845 & ~n6846;
  assign n6848 = ~n6844 & ~n6846;
  assign n6849 = n6829 & ~n6848;
  assign n6850 = ~n6847 & ~n6849;
  assign n6851 = n6785 & n6850;
  assign n6852 = ~n6821 & ~n6825;
  assign n6853 = ~n6826 & n6852;
  assign n6854 = ~n6827 & n6853;
  assign n1405 = n6851 | ~n6854;
  assign n6856 = REIP_REG_3_ & n6756;
  assign n6857 = PHYADDRPOINTER_REG_1_ & PHYADDRPOINTER_REG_2_;
  assign n6858 = ~PHYADDRPOINTER_REG_3_ & n6857;
  assign n6859 = PHYADDRPOINTER_REG_3_ & ~n6857;
  assign n6860 = ~n6858 & ~n6859;
  assign n6861 = n6754 & ~n6860;
  assign n6862 = n4846 & n6749;
  assign n6863 = PHYADDRPOINTER_REG_3_ & n6748;
  assign n6864 = INSTQUEUERD_ADDR_REG_3_ & n6742;
  assign n6865 = n2682 & ~n6860;
  assign n6866 = EAX_REG_3_ & n6759;
  assign n6867 = PHYADDRPOINTER_REG_3_ & n6763;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = ~n2580 & ~n6766;
  assign n6870 = ~n6864 & ~n6865;
  assign n6871 = n6868 & n6870;
  assign n6872 = ~n6869 & n6871;
  assign n6873 = ~n2682 & ~n6872;
  assign n6874 = n2682 & n6872;
  assign n6875 = n2994 & ~n6766;
  assign n6876 = ~n6873 & ~n6874;
  assign n6877 = ~n6875 & n6876;
  assign n6878 = n6875 & ~n6876;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = ~n6845 & ~n6846;
  assign n6881 = ~n6879 & n6880;
  assign n6882 = n6879 & ~n6880;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = n6785 & n6883;
  assign n6885 = ~n6856 & ~n6861;
  assign n6886 = ~n6862 & n6885;
  assign n6887 = ~n6863 & n6886;
  assign n1410 = n6884 | ~n6887;
  assign n6889 = REIP_REG_4_ & n6756;
  assign n6890 = PHYADDRPOINTER_REG_1_ & PHYADDRPOINTER_REG_3_;
  assign n6891 = PHYADDRPOINTER_REG_2_ & n6890;
  assign n6892 = ~PHYADDRPOINTER_REG_4_ & n6891;
  assign n6893 = PHYADDRPOINTER_REG_4_ & ~n6891;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = n6754 & ~n6894;
  assign n6896 = n4948 & n6749;
  assign n6897 = PHYADDRPOINTER_REG_4_ & n6748;
  assign n6898 = ~n4938 & ~n6766;
  assign n6899 = INSTQUEUERD_ADDR_REG_4_ & n6742;
  assign n6900 = n2682 & ~n6894;
  assign n6901 = EAX_REG_4_ & n6759;
  assign n6902 = PHYADDRPOINTER_REG_4_ & n6763;
  assign n6903 = ~n6901 & ~n6902;
  assign n6904 = ~n2570 & ~n6766;
  assign n6905 = ~n6899 & ~n6900;
  assign n6906 = n6903 & n6905;
  assign n6907 = ~n6904 & n6906;
  assign n6908 = ~n2682 & ~n6907;
  assign n6909 = n2682 & n6907;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = n6898 & ~n6910;
  assign n6912 = ~n6898 & n6910;
  assign n6913 = ~n6911 & ~n6912;
  assign n6914 = ~n6844 & ~n6877;
  assign n6915 = ~n6779 & ~n6809;
  assign n6916 = ~n2682 & ~n6778;
  assign n6917 = n6915 & ~n6916;
  assign n6918 = ~n6808 & ~n6917;
  assign n6919 = ~n6846 & n6918;
  assign n6920 = n6914 & ~n6919;
  assign n6921 = ~n6878 & ~n6920;
  assign n6922 = n6913 & n6921;
  assign n6923 = ~n6913 & ~n6921;
  assign n6924 = ~n6922 & ~n6923;
  assign n6925 = n6785 & ~n6924;
  assign n6926 = ~n6889 & ~n6895;
  assign n6927 = ~n6896 & n6926;
  assign n6928 = ~n6897 & n6927;
  assign n1415 = n6925 | ~n6928;
  assign n6930 = REIP_REG_5_ & n6756;
  assign n6931 = PHYADDRPOINTER_REG_4_ & n6891;
  assign n6932 = ~PHYADDRPOINTER_REG_5_ & n6931;
  assign n6933 = PHYADDRPOINTER_REG_5_ & ~n6931;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = n6754 & ~n6934;
  assign n6936 = n5052 & n6749;
  assign n6937 = PHYADDRPOINTER_REG_5_ & n6748;
  assign n6938 = ~n5042 & ~n6766;
  assign n6939 = n2554 & n2567;
  assign n6940 = ~n6766 & n6939;
  assign n6941 = EAX_REG_5_ & n6759;
  assign n6942 = n2682 & ~n6934;
  assign n6943 = PHYADDRPOINTER_REG_5_ & n6763;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = ~n6941 & n6944;
  assign n6946 = ~n6940 & n6945;
  assign n6947 = ~n2682 & ~n6946;
  assign n6948 = n2682 & n6946;
  assign n6949 = ~n6947 & ~n6948;
  assign n6950 = n6938 & ~n6949;
  assign n6951 = ~n6938 & n6949;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = ~n6912 & ~n6921;
  assign n6954 = ~n6911 & ~n6953;
  assign n6955 = n6952 & n6954;
  assign n6956 = ~n6952 & ~n6954;
  assign n6957 = ~n6955 & ~n6956;
  assign n6958 = n6785 & ~n6957;
  assign n6959 = ~n6930 & ~n6935;
  assign n6960 = ~n6936 & n6959;
  assign n6961 = ~n6937 & n6960;
  assign n1420 = n6958 | ~n6961;
  assign n6963 = REIP_REG_6_ & n6756;
  assign n6964 = PHYADDRPOINTER_REG_1_ & PHYADDRPOINTER_REG_5_;
  assign n6965 = PHYADDRPOINTER_REG_4_ & n6964;
  assign n6966 = PHYADDRPOINTER_REG_2_ & n6965;
  assign n6967 = PHYADDRPOINTER_REG_3_ & n6966;
  assign n6968 = ~PHYADDRPOINTER_REG_6_ & n6967;
  assign n6969 = PHYADDRPOINTER_REG_6_ & ~n6967;
  assign n6970 = ~n6968 & ~n6969;
  assign n6971 = n6754 & ~n6970;
  assign n6972 = n5152 & n6749;
  assign n6973 = PHYADDRPOINTER_REG_6_ & n6748;
  assign n6974 = EAX_REG_6_ & n6759;
  assign n6975 = n2682 & ~n6970;
  assign n6976 = PHYADDRPOINTER_REG_6_ & n6763;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = ~n6974 & n6977;
  assign n6979 = ~n2682 & ~n6978;
  assign n6980 = n2682 & n6978;
  assign n6981 = ~n6979 & ~n6980;
  assign n6982 = n5142 & ~n6766;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = n6981 & n6982;
  assign n6985 = ~n6983 & ~n6984;
  assign n6986 = ~n6951 & ~n6954;
  assign n6987 = ~n6950 & ~n6986;
  assign n6988 = ~n6985 & n6987;
  assign n6989 = n6981 & ~n6982;
  assign n6990 = ~n6981 & n6982;
  assign n6991 = ~n6989 & ~n6990;
  assign n6992 = ~n6987 & ~n6991;
  assign n6993 = ~n6988 & ~n6992;
  assign n6994 = n6785 & ~n6993;
  assign n6995 = ~n6963 & ~n6971;
  assign n6996 = ~n6972 & n6995;
  assign n6997 = ~n6973 & n6996;
  assign n1425 = n6994 | ~n6997;
  assign n6999 = REIP_REG_7_ & n6756;
  assign n7000 = PHYADDRPOINTER_REG_6_ & n6967;
  assign n7001 = ~PHYADDRPOINTER_REG_7_ & n7000;
  assign n7002 = PHYADDRPOINTER_REG_7_ & ~n7000;
  assign n7003 = ~n7001 & ~n7002;
  assign n7004 = n6754 & ~n7003;
  assign n7005 = n5229 & n6749;
  assign n7006 = PHYADDRPOINTER_REG_7_ & n6748;
  assign n7007 = n5219 & ~n6766;
  assign n7008 = EAX_REG_7_ & n6759;
  assign n7009 = n2682 & ~n7003;
  assign n7010 = PHYADDRPOINTER_REG_7_ & n6763;
  assign n7011 = ~n7009 & ~n7010;
  assign n7012 = ~n7008 & n7011;
  assign n7013 = ~n2682 & ~n7012;
  assign n7014 = n2682 & n7012;
  assign n7015 = ~n7013 & ~n7014;
  assign n7016 = n7007 & ~n7015;
  assign n7017 = ~n7007 & n7015;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = ~n6990 & ~n7018;
  assign n7020 = ~n6987 & ~n6989;
  assign n7021 = n7019 & ~n7020;
  assign n7022 = n6982 & ~n7017;
  assign n7023 = ~n6981 & ~n7017;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = ~n7016 & ~n7024;
  assign n7026 = n6987 & ~n6990;
  assign n7027 = n7025 & ~n7026;
  assign n7028 = ~n7021 & ~n7027;
  assign n7029 = n6785 & n7028;
  assign n7030 = ~n6999 & ~n7004;
  assign n7031 = ~n7005 & n7030;
  assign n7032 = ~n7006 & n7031;
  assign n1430 = n7029 | ~n7032;
  assign n7034 = REIP_REG_8_ & n6756;
  assign n7035 = PHYADDRPOINTER_REG_6_ & PHYADDRPOINTER_REG_7_;
  assign n7036 = n6967 & n7035;
  assign n7037 = ~PHYADDRPOINTER_REG_8_ & n7036;
  assign n7038 = PHYADDRPOINTER_REG_8_ & ~n7036;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = n6754 & ~n7039;
  assign n7041 = PHYADDRPOINTER_REG_8_ & n6748;
  assign n7042 = n5362 & n6749;
  assign n7043 = n5339 & ~n6766;
  assign n7044 = EAX_REG_8_ & n6759;
  assign n7045 = n2682 & ~n7039;
  assign n7046 = PHYADDRPOINTER_REG_8_ & n6763;
  assign n7047 = ~n7045 & ~n7046;
  assign n7048 = ~n7044 & n7047;
  assign n7049 = ~n2682 & ~n7048;
  assign n7050 = n2682 & n7048;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = n7043 & ~n7051;
  assign n7053 = ~n7043 & n7051;
  assign n7054 = ~n7052 & ~n7053;
  assign n7055 = n6990 & ~n7017;
  assign n7056 = ~n6912 & ~n6951;
  assign n7057 = ~n6921 & n7056;
  assign n7058 = ~n7024 & n7057;
  assign n7059 = ~n6911 & ~n6950;
  assign n7060 = ~n6951 & ~n7059;
  assign n7061 = ~n7024 & n7060;
  assign n7062 = ~n7016 & ~n7061;
  assign n7063 = ~n7055 & ~n7058;
  assign n7064 = n7062 & n7063;
  assign n7065 = n7054 & n7064;
  assign n7066 = ~n7054 & ~n7064;
  assign n7067 = ~n7065 & ~n7066;
  assign n7068 = n6785 & ~n7067;
  assign n7069 = ~n7034 & ~n7040;
  assign n7070 = ~n7041 & n7069;
  assign n7071 = ~n7042 & n7070;
  assign n1435 = n7068 | ~n7071;
  assign n7073 = REIP_REG_9_ & n6756;
  assign n7074 = PHYADDRPOINTER_REG_8_ & n7036;
  assign n7075 = ~PHYADDRPOINTER_REG_9_ & n7074;
  assign n7076 = PHYADDRPOINTER_REG_9_ & ~n7074;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = n6754 & ~n7077;
  assign n7079 = PHYADDRPOINTER_REG_9_ & n6748;
  assign n7080 = n5445 & n6749;
  assign n7081 = ~n7053 & ~n7064;
  assign n7082 = ~n7052 & ~n7081;
  assign n7083 = EAX_REG_9_ & n6759;
  assign n7084 = n2682 & ~n7077;
  assign n7085 = PHYADDRPOINTER_REG_9_ & n6763;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = ~n7083 & n7086;
  assign n7088 = ~n2682 & ~n7087;
  assign n7089 = n2682 & n7087;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = ~n5436 & ~n6766;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = n7090 & n7091;
  assign n7094 = ~n7092 & ~n7093;
  assign n7095 = n7082 & ~n7094;
  assign n7096 = ~n7082 & n7094;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = n6785 & ~n7097;
  assign n7099 = ~n7073 & ~n7078;
  assign n7100 = ~n7079 & n7099;
  assign n7101 = ~n7080 & n7100;
  assign n1440 = n7098 | ~n7101;
  assign n7103 = REIP_REG_10_ & n6756;
  assign n7104 = PHYADDRPOINTER_REG_8_ & PHYADDRPOINTER_REG_9_;
  assign n7105 = n7036 & n7104;
  assign n7106 = ~PHYADDRPOINTER_REG_10_ & n7105;
  assign n7107 = PHYADDRPOINTER_REG_10_ & ~n7105;
  assign n7108 = ~n7106 & ~n7107;
  assign n7109 = n6754 & ~n7108;
  assign n7110 = PHYADDRPOINTER_REG_10_ & n6748;
  assign n7111 = n5530 & n6749;
  assign n7112 = n7090 & ~n7091;
  assign n7113 = n7052 & ~n7112;
  assign n7114 = ~n7090 & n7091;
  assign n7115 = ~n7113 & ~n7114;
  assign n7116 = ~n7053 & ~n7112;
  assign n7117 = ~n7064 & n7116;
  assign n7118 = n7115 & ~n7117;
  assign n7119 = EAX_REG_10_ & n6759;
  assign n7120 = n2682 & ~n7108;
  assign n7121 = PHYADDRPOINTER_REG_10_ & n6763;
  assign n7122 = ~n7120 & ~n7121;
  assign n7123 = ~n7119 & n7122;
  assign n7124 = ~n2682 & ~n7123;
  assign n7125 = n2682 & n7123;
  assign n7126 = ~n5521 & ~n6766;
  assign n7127 = ~n7124 & ~n7125;
  assign n7128 = ~n7126 & n7127;
  assign n7129 = ~n7118 & ~n7128;
  assign n7130 = n7126 & ~n7127;
  assign n7131 = n7129 & ~n7130;
  assign n7132 = ~n7128 & ~n7130;
  assign n7133 = n7118 & ~n7132;
  assign n7134 = ~n7131 & ~n7133;
  assign n7135 = n6785 & n7134;
  assign n7136 = ~n7103 & ~n7109;
  assign n7137 = ~n7110 & n7136;
  assign n7138 = ~n7111 & n7137;
  assign n1445 = n7135 | ~n7138;
  assign n7140 = REIP_REG_11_ & n6756;
  assign n7141 = PHYADDRPOINTER_REG_10_ & n7105;
  assign n7142 = ~PHYADDRPOINTER_REG_11_ & n7141;
  assign n7143 = PHYADDRPOINTER_REG_11_ & ~n7141;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = n6754 & ~n7144;
  assign n7146 = PHYADDRPOINTER_REG_11_ & n6748;
  assign n7147 = n5616 & n6749;
  assign n7148 = EAX_REG_11_ & n6759;
  assign n7149 = PHYADDRPOINTER_REG_11_ & n6763;
  assign n7150 = n2682 & ~n7144;
  assign n7151 = ~n7148 & ~n7149;
  assign n7152 = ~n7150 & n7151;
  assign n7153 = ~n2682 & ~n7152;
  assign n7154 = n2682 & n7152;
  assign n7155 = ~n5607 & ~n6766;
  assign n7156 = ~n7153 & ~n7154;
  assign n7157 = ~n7155 & n7156;
  assign n7158 = n7155 & ~n7156;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~n7130 & ~n7159;
  assign n7161 = ~n7129 & n7160;
  assign n7162 = ~n7129 & ~n7130;
  assign n7163 = n7159 & ~n7162;
  assign n7164 = ~n7161 & ~n7163;
  assign n7165 = n6785 & n7164;
  assign n7166 = ~n7140 & ~n7145;
  assign n7167 = ~n7146 & n7166;
  assign n7168 = ~n7147 & n7167;
  assign n1450 = n7165 | ~n7168;
  assign n7170 = REIP_REG_12_ & n6756;
  assign n7171 = PHYADDRPOINTER_REG_10_ & PHYADDRPOINTER_REG_11_;
  assign n7172 = n7105 & n7171;
  assign n7173 = ~PHYADDRPOINTER_REG_12_ & n7172;
  assign n7174 = PHYADDRPOINTER_REG_12_ & ~n7172;
  assign n7175 = ~n7173 & ~n7174;
  assign n7176 = n6754 & ~n7175;
  assign n7177 = PHYADDRPOINTER_REG_12_ & n6748;
  assign n7178 = n5717 & n6749;
  assign n7179 = EAX_REG_12_ & n6759;
  assign n7180 = PHYADDRPOINTER_REG_12_ & n6763;
  assign n7181 = n2682 & ~n7175;
  assign n7182 = ~n7179 & ~n7180;
  assign n7183 = ~n7181 & n7182;
  assign n7184 = ~n2682 & ~n7183;
  assign n7185 = n2682 & n7183;
  assign n7186 = ~n5694 & ~n6766;
  assign n7187 = ~n7184 & ~n7185;
  assign n7188 = ~n7186 & n7187;
  assign n7189 = n7186 & ~n7187;
  assign n7190 = ~n7188 & ~n7189;
  assign n7191 = ~n7128 & ~n7157;
  assign n7192 = ~n7115 & n7191;
  assign n7193 = ~n7130 & ~n7158;
  assign n7194 = ~n7157 & ~n7193;
  assign n7195 = ~n7192 & ~n7194;
  assign n7196 = n7116 & n7191;
  assign n7197 = ~n7064 & n7196;
  assign n7198 = n7195 & ~n7197;
  assign n7199 = n7190 & n7198;
  assign n7200 = ~n7190 & ~n7198;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = n6785 & ~n7201;
  assign n7203 = ~n7170 & ~n7176;
  assign n7204 = ~n7177 & n7203;
  assign n7205 = ~n7178 & n7204;
  assign n1455 = n7202 | ~n7205;
  assign n7207 = REIP_REG_13_ & n6756;
  assign n7208 = PHYADDRPOINTER_REG_12_ & n7172;
  assign n7209 = ~PHYADDRPOINTER_REG_13_ & n7208;
  assign n7210 = PHYADDRPOINTER_REG_13_ & ~n7208;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = n6754 & ~n7211;
  assign n7213 = PHYADDRPOINTER_REG_13_ & n6748;
  assign n7214 = n5800 & n6749;
  assign n7215 = ~n7188 & ~n7198;
  assign n7216 = ~n7189 & ~n7215;
  assign n7217 = EAX_REG_13_ & n6759;
  assign n7218 = PHYADDRPOINTER_REG_13_ & n6763;
  assign n7219 = n2682 & ~n7211;
  assign n7220 = ~n7217 & ~n7218;
  assign n7221 = ~n7219 & n7220;
  assign n7222 = ~n2682 & ~n7221;
  assign n7223 = n2682 & n7221;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = ~n5791 & ~n6766;
  assign n7226 = ~n7224 & ~n7225;
  assign n7227 = n7224 & n7225;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = n7216 & ~n7228;
  assign n7230 = n7224 & ~n7225;
  assign n7231 = ~n7224 & n7225;
  assign n7232 = ~n7230 & ~n7231;
  assign n7233 = ~n7216 & ~n7232;
  assign n7234 = ~n7229 & ~n7233;
  assign n7235 = n6785 & ~n7234;
  assign n7236 = ~n7207 & ~n7212;
  assign n7237 = ~n7213 & n7236;
  assign n7238 = ~n7214 & n7237;
  assign n1460 = n7235 | ~n7238;
  assign n7240 = REIP_REG_14_ & n6756;
  assign n7241 = PHYADDRPOINTER_REG_12_ & PHYADDRPOINTER_REG_13_;
  assign n7242 = n7172 & n7241;
  assign n7243 = ~PHYADDRPOINTER_REG_14_ & n7242;
  assign n7244 = PHYADDRPOINTER_REG_14_ & ~n7242;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = n6754 & ~n7245;
  assign n7247 = PHYADDRPOINTER_REG_14_ & n6748;
  assign n7248 = n5885 & n6749;
  assign n7249 = EAX_REG_14_ & n6759;
  assign n7250 = PHYADDRPOINTER_REG_14_ & n6763;
  assign n7251 = n2682 & ~n7245;
  assign n7252 = ~n7249 & ~n7250;
  assign n7253 = ~n7251 & n7252;
  assign n7254 = ~n2682 & ~n7253;
  assign n7255 = n2682 & n7253;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = ~n5876 & ~n6766;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = n7256 & n7257;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = ~n7216 & ~n7230;
  assign n7262 = ~n7231 & ~n7261;
  assign n7263 = ~n7260 & n7262;
  assign n7264 = ~n7256 & n7257;
  assign n7265 = n7256 & ~n7257;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = ~n7262 & ~n7266;
  assign n7268 = ~n7263 & ~n7267;
  assign n7269 = n6785 & ~n7268;
  assign n7270 = ~n7240 & ~n7246;
  assign n7271 = ~n7247 & n7270;
  assign n7272 = ~n7248 & n7271;
  assign n1465 = n7269 | ~n7272;
  assign n7274 = REIP_REG_15_ & n6756;
  assign n7275 = PHYADDRPOINTER_REG_14_ & n7242;
  assign n7276 = ~PHYADDRPOINTER_REG_15_ & n7275;
  assign n7277 = PHYADDRPOINTER_REG_15_ & ~n7275;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = n6754 & ~n7278;
  assign n7280 = PHYADDRPOINTER_REG_15_ & n6748;
  assign n7281 = n5969 & n6749;
  assign n7282 = ~n5960 & ~n6766;
  assign n7283 = EAX_REG_15_ & n6759;
  assign n7284 = PHYADDRPOINTER_REG_15_ & n6763;
  assign n7285 = n2682 & ~n7278;
  assign n7286 = ~n7283 & ~n7284;
  assign n7287 = ~n7285 & n7286;
  assign n7288 = ~n2682 & ~n7287;
  assign n7289 = n2682 & n7287;
  assign n7290 = ~n7288 & ~n7289;
  assign n7291 = n7282 & ~n7290;
  assign n7292 = ~n7282 & n7290;
  assign n7293 = ~n7291 & ~n7292;
  assign n7294 = ~n7264 & ~n7293;
  assign n7295 = ~n7262 & ~n7265;
  assign n7296 = n7294 & ~n7295;
  assign n7297 = ~n7265 & ~n7292;
  assign n7298 = ~n7291 & n7297;
  assign n7299 = n7262 & ~n7264;
  assign n7300 = n7298 & ~n7299;
  assign n7301 = ~n7296 & ~n7300;
  assign n7302 = n6785 & n7301;
  assign n7303 = ~n7274 & ~n7279;
  assign n7304 = ~n7280 & n7303;
  assign n7305 = ~n7281 & n7304;
  assign n1470 = n7302 | ~n7305;
  assign n7307 = REIP_REG_16_ & n6756;
  assign n7308 = PHYADDRPOINTER_REG_14_ & PHYADDRPOINTER_REG_15_;
  assign n7309 = n7242 & n7308;
  assign n7310 = ~PHYADDRPOINTER_REG_16_ & n7309;
  assign n7311 = PHYADDRPOINTER_REG_16_ & ~n7309;
  assign n7312 = ~n7310 & ~n7311;
  assign n7313 = n6754 & ~n7312;
  assign n7314 = PHYADDRPOINTER_REG_16_ & n6748;
  assign n7315 = n6033 & n6749;
  assign n7316 = INSTQUEUERD_ADDR_REG_2_ & ~n1722_1;
  assign n7317 = ~INSTQUEUERD_ADDR_REG_3_ & n7316;
  assign n7318 = INSTQUEUERD_ADDR_REG_3_ & ~n7316;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = ~n1736 & ~n7316;
  assign n7321 = n7319 & n7320;
  assign n7322 = n2730 & n7321;
  assign n7323 = INSTQUEUE_REG_7__0_ & n7322;
  assign n7324 = n2727 & n7321;
  assign n7325 = INSTQUEUE_REG_6__0_ & n7324;
  assign n7326 = n2736 & n7321;
  assign n7327 = INSTQUEUE_REG_5__0_ & n7326;
  assign n7328 = n2733 & n7321;
  assign n7329 = INSTQUEUE_REG_4__0_ & n7328;
  assign n7330 = ~n7323 & ~n7325;
  assign n7331 = ~n7327 & n7330;
  assign n7332 = ~n7329 & n7331;
  assign n7333 = n7319 & ~n7320;
  assign n7334 = n2730 & n7333;
  assign n7335 = INSTQUEUE_REG_3__0_ & n7334;
  assign n7336 = n2727 & n7333;
  assign n7337 = INSTQUEUE_REG_2__0_ & n7336;
  assign n7338 = n2736 & n7333;
  assign n7339 = INSTQUEUE_REG_1__0_ & n7338;
  assign n7340 = n2733 & n7333;
  assign n7341 = INSTQUEUE_REG_0__0_ & n7340;
  assign n7342 = ~n7335 & ~n7337;
  assign n7343 = ~n7339 & n7342;
  assign n7344 = ~n7341 & n7343;
  assign n7345 = ~n7319 & n7320;
  assign n7346 = n2730 & n7345;
  assign n7347 = INSTQUEUE_REG_15__0_ & n7346;
  assign n7348 = n2727 & n7345;
  assign n7349 = INSTQUEUE_REG_14__0_ & n7348;
  assign n7350 = n2736 & n7345;
  assign n7351 = INSTQUEUE_REG_13__0_ & n7350;
  assign n7352 = n2733 & n7345;
  assign n7353 = INSTQUEUE_REG_12__0_ & n7352;
  assign n7354 = ~n7347 & ~n7349;
  assign n7355 = ~n7351 & n7354;
  assign n7356 = ~n7353 & n7355;
  assign n7357 = ~n7319 & ~n7320;
  assign n7358 = n2730 & n7357;
  assign n7359 = INSTQUEUE_REG_11__0_ & n7358;
  assign n7360 = n2727 & n7357;
  assign n7361 = INSTQUEUE_REG_10__0_ & n7360;
  assign n7362 = n2736 & n7357;
  assign n7363 = INSTQUEUE_REG_9__0_ & n7362;
  assign n7364 = n2733 & n7357;
  assign n7365 = INSTQUEUE_REG_8__0_ & n7364;
  assign n7366 = ~n7359 & ~n7361;
  assign n7367 = ~n7363 & n7366;
  assign n7368 = ~n7365 & n7367;
  assign n7369 = n7332 & n7344;
  assign n7370 = n7356 & n7369;
  assign n7371 = n7368 & n7370;
  assign n7372 = STATE2_REG_0_ & n2266;
  assign n7373 = n2101 & n2144;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = ~n7371 & ~n7374;
  assign n7376 = ~n6766 & n7375;
  assign n7377 = EAX_REG_16_ & n6759;
  assign n7378 = PHYADDRPOINTER_REG_16_ & n6763;
  assign n7379 = n2682 & ~n7312;
  assign n7380 = ~n7377 & ~n7378;
  assign n7381 = ~n7379 & n7380;
  assign n7382 = ~n7376 & n7381;
  assign n7383 = ~n2682 & ~n7382;
  assign n7384 = n2682 & n7382;
  assign n7385 = ~n6012 & ~n6766;
  assign n7386 = ~n7383 & ~n7384;
  assign n7387 = ~n7385 & n7386;
  assign n7388 = n7231 & ~n7265;
  assign n7389 = ~n7292 & n7388;
  assign n7390 = ~n7188 & ~n7265;
  assign n7391 = ~n7230 & ~n7292;
  assign n7392 = ~n7198 & n7390;
  assign n7393 = n7391 & n7392;
  assign n7394 = ~n7264 & ~n7282;
  assign n7395 = ~n7264 & n7290;
  assign n7396 = ~n7292 & ~n7394;
  assign n7397 = ~n7395 & n7396;
  assign n7398 = n7189 & ~n7230;
  assign n7399 = ~n7265 & n7398;
  assign n7400 = ~n7292 & n7399;
  assign n7401 = ~n7397 & ~n7400;
  assign n7402 = ~n7389 & ~n7393;
  assign n7403 = n7401 & n7402;
  assign n7404 = ~n7387 & ~n7403;
  assign n7405 = n7385 & ~n7386;
  assign n7406 = n7404 & ~n7405;
  assign n7407 = ~n7387 & ~n7405;
  assign n7408 = n7403 & ~n7407;
  assign n7409 = ~n7406 & ~n7408;
  assign n7410 = n6785 & n7409;
  assign n7411 = ~n7307 & ~n7313;
  assign n7412 = ~n7314 & n7411;
  assign n7413 = ~n7315 & n7412;
  assign n1475 = n7410 | ~n7413;
  assign n7415 = REIP_REG_17_ & n6756;
  assign n7416 = PHYADDRPOINTER_REG_16_ & n7309;
  assign n7417 = ~PHYADDRPOINTER_REG_17_ & n7416;
  assign n7418 = PHYADDRPOINTER_REG_17_ & ~n7416;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = n6754 & ~n7419;
  assign n7421 = PHYADDRPOINTER_REG_17_ & n6748;
  assign n7422 = n6078 & n6749;
  assign n7423 = n6010 & ~n6766;
  assign n7424 = INSTQUEUE_REG_7__1_ & n7322;
  assign n7425 = INSTQUEUE_REG_6__1_ & n7324;
  assign n7426 = INSTQUEUE_REG_5__1_ & n7326;
  assign n7427 = INSTQUEUE_REG_4__1_ & n7328;
  assign n7428 = ~n7424 & ~n7425;
  assign n7429 = ~n7426 & n7428;
  assign n7430 = ~n7427 & n7429;
  assign n7431 = INSTQUEUE_REG_3__1_ & n7334;
  assign n7432 = INSTQUEUE_REG_2__1_ & n7336;
  assign n7433 = INSTQUEUE_REG_1__1_ & n7338;
  assign n7434 = INSTQUEUE_REG_0__1_ & n7340;
  assign n7435 = ~n7431 & ~n7432;
  assign n7436 = ~n7433 & n7435;
  assign n7437 = ~n7434 & n7436;
  assign n7438 = INSTQUEUE_REG_15__1_ & n7346;
  assign n7439 = INSTQUEUE_REG_14__1_ & n7348;
  assign n7440 = INSTQUEUE_REG_13__1_ & n7350;
  assign n7441 = INSTQUEUE_REG_12__1_ & n7352;
  assign n7442 = ~n7438 & ~n7439;
  assign n7443 = ~n7440 & n7442;
  assign n7444 = ~n7441 & n7443;
  assign n7445 = INSTQUEUE_REG_11__1_ & n7358;
  assign n7446 = INSTQUEUE_REG_10__1_ & n7360;
  assign n7447 = INSTQUEUE_REG_9__1_ & n7362;
  assign n7448 = INSTQUEUE_REG_8__1_ & n7364;
  assign n7449 = ~n7445 & ~n7446;
  assign n7450 = ~n7447 & n7449;
  assign n7451 = ~n7448 & n7450;
  assign n7452 = n7430 & n7437;
  assign n7453 = n7444 & n7452;
  assign n7454 = n7451 & n7453;
  assign n7455 = ~n7374 & ~n7454;
  assign n7456 = ~n6766 & n7455;
  assign n7457 = EAX_REG_17_ & n6759;
  assign n7458 = PHYADDRPOINTER_REG_17_ & n6763;
  assign n7459 = n2682 & ~n7419;
  assign n7460 = ~n7457 & ~n7458;
  assign n7461 = ~n7459 & n7460;
  assign n7462 = ~n7456 & n7461;
  assign n7463 = ~n2682 & ~n7462;
  assign n7464 = n2682 & n7462;
  assign n7465 = ~n7463 & ~n7464;
  assign n7466 = n7423 & ~n7465;
  assign n7467 = ~n7423 & n7465;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = ~n7404 & ~n7405;
  assign n7470 = n7468 & n7469;
  assign n7471 = ~n7468 & ~n7469;
  assign n7472 = ~n7470 & ~n7471;
  assign n7473 = n6785 & ~n7472;
  assign n7474 = ~n7415 & ~n7420;
  assign n7475 = ~n7421 & n7474;
  assign n7476 = ~n7422 & n7475;
  assign n1480 = n7473 | ~n7476;
  assign n7478 = REIP_REG_18_ & n6756;
  assign n7479 = PHYADDRPOINTER_REG_16_ & PHYADDRPOINTER_REG_17_;
  assign n7480 = n7309 & n7479;
  assign n7481 = ~PHYADDRPOINTER_REG_18_ & n7480;
  assign n7482 = PHYADDRPOINTER_REG_18_ & ~n7480;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = n6754 & ~n7483;
  assign n7485 = PHYADDRPOINTER_REG_18_ & n6748;
  assign n7486 = n6125 & n6749;
  assign n7487 = INSTQUEUE_REG_7__2_ & n7322;
  assign n7488 = INSTQUEUE_REG_6__2_ & n7324;
  assign n7489 = INSTQUEUE_REG_5__2_ & n7326;
  assign n7490 = INSTQUEUE_REG_4__2_ & n7328;
  assign n7491 = ~n7487 & ~n7488;
  assign n7492 = ~n7489 & n7491;
  assign n7493 = ~n7490 & n7492;
  assign n7494 = INSTQUEUE_REG_3__2_ & n7334;
  assign n7495 = INSTQUEUE_REG_2__2_ & n7336;
  assign n7496 = INSTQUEUE_REG_1__2_ & n7338;
  assign n7497 = INSTQUEUE_REG_0__2_ & n7340;
  assign n7498 = ~n7494 & ~n7495;
  assign n7499 = ~n7496 & n7498;
  assign n7500 = ~n7497 & n7499;
  assign n7501 = INSTQUEUE_REG_15__2_ & n7346;
  assign n7502 = INSTQUEUE_REG_14__2_ & n7348;
  assign n7503 = INSTQUEUE_REG_13__2_ & n7350;
  assign n7504 = INSTQUEUE_REG_12__2_ & n7352;
  assign n7505 = ~n7501 & ~n7502;
  assign n7506 = ~n7503 & n7505;
  assign n7507 = ~n7504 & n7506;
  assign n7508 = INSTQUEUE_REG_11__2_ & n7358;
  assign n7509 = INSTQUEUE_REG_10__2_ & n7360;
  assign n7510 = INSTQUEUE_REG_9__2_ & n7362;
  assign n7511 = INSTQUEUE_REG_8__2_ & n7364;
  assign n7512 = ~n7508 & ~n7509;
  assign n7513 = ~n7510 & n7512;
  assign n7514 = ~n7511 & n7513;
  assign n7515 = n7493 & n7500;
  assign n7516 = n7507 & n7515;
  assign n7517 = n7514 & n7516;
  assign n7518 = ~n7374 & ~n7517;
  assign n7519 = ~n6766 & n7518;
  assign n7520 = EAX_REG_18_ & n6759;
  assign n7521 = PHYADDRPOINTER_REG_18_ & n6763;
  assign n7522 = n2682 & ~n7483;
  assign n7523 = ~n7520 & ~n7521;
  assign n7524 = ~n7522 & n7523;
  assign n7525 = ~n7519 & n7524;
  assign n7526 = ~n2682 & ~n7525;
  assign n7527 = n2682 & n7525;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = n7423 & ~n7528;
  assign n7530 = ~n7423 & n7528;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = ~n7467 & ~n7469;
  assign n7533 = ~n7466 & ~n7532;
  assign n7534 = n7531 & n7533;
  assign n7535 = ~n7531 & ~n7533;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = n6785 & ~n7536;
  assign n7538 = ~n7478 & ~n7484;
  assign n7539 = ~n7485 & n7538;
  assign n7540 = ~n7486 & n7539;
  assign n1485 = n7537 | ~n7540;
  assign n7542 = REIP_REG_19_ & n6756;
  assign n7543 = PHYADDRPOINTER_REG_18_ & n7480;
  assign n7544 = ~PHYADDRPOINTER_REG_19_ & n7543;
  assign n7545 = PHYADDRPOINTER_REG_19_ & ~n7543;
  assign n7546 = ~n7544 & ~n7545;
  assign n7547 = n6754 & ~n7546;
  assign n7548 = PHYADDRPOINTER_REG_19_ & n6748;
  assign n7549 = n6172 & n6749;
  assign n7550 = INSTQUEUE_REG_7__3_ & n7322;
  assign n7551 = INSTQUEUE_REG_6__3_ & n7324;
  assign n7552 = INSTQUEUE_REG_5__3_ & n7326;
  assign n7553 = INSTQUEUE_REG_4__3_ & n7328;
  assign n7554 = ~n7550 & ~n7551;
  assign n7555 = ~n7552 & n7554;
  assign n7556 = ~n7553 & n7555;
  assign n7557 = INSTQUEUE_REG_3__3_ & n7334;
  assign n7558 = INSTQUEUE_REG_2__3_ & n7336;
  assign n7559 = INSTQUEUE_REG_1__3_ & n7338;
  assign n7560 = INSTQUEUE_REG_0__3_ & n7340;
  assign n7561 = ~n7557 & ~n7558;
  assign n7562 = ~n7559 & n7561;
  assign n7563 = ~n7560 & n7562;
  assign n7564 = INSTQUEUE_REG_15__3_ & n7346;
  assign n7565 = INSTQUEUE_REG_14__3_ & n7348;
  assign n7566 = INSTQUEUE_REG_13__3_ & n7350;
  assign n7567 = INSTQUEUE_REG_12__3_ & n7352;
  assign n7568 = ~n7564 & ~n7565;
  assign n7569 = ~n7566 & n7568;
  assign n7570 = ~n7567 & n7569;
  assign n7571 = INSTQUEUE_REG_11__3_ & n7358;
  assign n7572 = INSTQUEUE_REG_10__3_ & n7360;
  assign n7573 = INSTQUEUE_REG_9__3_ & n7362;
  assign n7574 = INSTQUEUE_REG_8__3_ & n7364;
  assign n7575 = ~n7571 & ~n7572;
  assign n7576 = ~n7573 & n7575;
  assign n7577 = ~n7574 & n7576;
  assign n7578 = n7556 & n7563;
  assign n7579 = n7570 & n7578;
  assign n7580 = n7577 & n7579;
  assign n7581 = ~n7374 & ~n7580;
  assign n7582 = ~n6766 & n7581;
  assign n7583 = EAX_REG_19_ & n6759;
  assign n7584 = PHYADDRPOINTER_REG_19_ & n6763;
  assign n7585 = n2682 & ~n7546;
  assign n7586 = ~n7583 & ~n7584;
  assign n7587 = ~n7585 & n7586;
  assign n7588 = ~n7582 & n7587;
  assign n7589 = ~n2682 & ~n7588;
  assign n7590 = n2682 & n7588;
  assign n7591 = ~n7589 & ~n7590;
  assign n7592 = ~n7423 & n7591;
  assign n7593 = n7423 & ~n7591;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = ~n7467 & ~n7530;
  assign n7596 = n7466 & n7595;
  assign n7597 = n7405 & n7595;
  assign n7598 = ~n7529 & ~n7596;
  assign n7599 = ~n7597 & n7598;
  assign n7600 = ~n7387 & n7595;
  assign n7601 = ~n7403 & n7600;
  assign n7602 = n7599 & ~n7601;
  assign n7603 = n7594 & n7602;
  assign n7604 = ~n7594 & ~n7602;
  assign n7605 = ~n7603 & ~n7604;
  assign n7606 = n6785 & ~n7605;
  assign n7607 = ~n7542 & ~n7547;
  assign n7608 = ~n7548 & n7607;
  assign n7609 = ~n7549 & n7608;
  assign n1490 = n7606 | ~n7609;
  assign n7611 = REIP_REG_20_ & n6756;
  assign n7612 = PHYADDRPOINTER_REG_18_ & PHYADDRPOINTER_REG_19_;
  assign n7613 = n7480 & n7612;
  assign n7614 = ~PHYADDRPOINTER_REG_20_ & n7613;
  assign n7615 = PHYADDRPOINTER_REG_20_ & ~n7613;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = n6754 & ~n7616;
  assign n7618 = PHYADDRPOINTER_REG_20_ & n6748;
  assign n7619 = n6218 & n6749;
  assign n7620 = INSTQUEUE_REG_0__4_ & n7340;
  assign n7621 = INSTQUEUE_REG_7__4_ & n7322;
  assign n7622 = INSTQUEUE_REG_6__4_ & n7324;
  assign n7623 = INSTQUEUE_REG_5__4_ & n7326;
  assign n7624 = ~n7620 & ~n7621;
  assign n7625 = ~n7622 & n7624;
  assign n7626 = ~n7623 & n7625;
  assign n7627 = INSTQUEUE_REG_4__4_ & n7328;
  assign n7628 = INSTQUEUE_REG_3__4_ & n7334;
  assign n7629 = INSTQUEUE_REG_2__4_ & n7336;
  assign n7630 = INSTQUEUE_REG_1__4_ & n7338;
  assign n7631 = ~n7627 & ~n7628;
  assign n7632 = ~n7629 & n7631;
  assign n7633 = ~n7630 & n7632;
  assign n7634 = INSTQUEUE_REG_15__4_ & n7346;
  assign n7635 = INSTQUEUE_REG_14__4_ & n7348;
  assign n7636 = INSTQUEUE_REG_13__4_ & n7350;
  assign n7637 = INSTQUEUE_REG_12__4_ & n7352;
  assign n7638 = ~n7634 & ~n7635;
  assign n7639 = ~n7636 & n7638;
  assign n7640 = ~n7637 & n7639;
  assign n7641 = INSTQUEUE_REG_11__4_ & n7358;
  assign n7642 = INSTQUEUE_REG_10__4_ & n7360;
  assign n7643 = INSTQUEUE_REG_9__4_ & n7362;
  assign n7644 = INSTQUEUE_REG_8__4_ & n7364;
  assign n7645 = ~n7641 & ~n7642;
  assign n7646 = ~n7643 & n7645;
  assign n7647 = ~n7644 & n7646;
  assign n7648 = n7626 & n7633;
  assign n7649 = n7640 & n7648;
  assign n7650 = n7647 & n7649;
  assign n7651 = ~n7374 & ~n7650;
  assign n7652 = ~n6766 & n7651;
  assign n7653 = EAX_REG_20_ & n6759;
  assign n7654 = PHYADDRPOINTER_REG_20_ & n6763;
  assign n7655 = n2682 & ~n7616;
  assign n7656 = ~n7653 & ~n7654;
  assign n7657 = ~n7655 & n7656;
  assign n7658 = ~n7652 & n7657;
  assign n7659 = ~n2682 & ~n7658;
  assign n7660 = n2682 & n7658;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7423 & ~n7661;
  assign n7663 = n7423 & n7661;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = ~n7592 & ~n7599;
  assign n7666 = ~n7593 & ~n7665;
  assign n7667 = ~n7387 & ~n7592;
  assign n7668 = n7595 & n7667;
  assign n7669 = ~n7403 & n7668;
  assign n7670 = n7666 & ~n7669;
  assign n7671 = ~n7664 & n7670;
  assign n7672 = ~n7423 & n7661;
  assign n7673 = n7423 & ~n7661;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = ~n7670 & ~n7674;
  assign n7676 = ~n7671 & ~n7675;
  assign n7677 = n6785 & ~n7676;
  assign n7678 = ~n7611 & ~n7617;
  assign n7679 = ~n7618 & n7678;
  assign n7680 = ~n7619 & n7679;
  assign n1495 = n7677 | ~n7680;
  assign n7682 = REIP_REG_21_ & n6756;
  assign n7683 = PHYADDRPOINTER_REG_20_ & n7613;
  assign n7684 = ~PHYADDRPOINTER_REG_21_ & n7683;
  assign n7685 = PHYADDRPOINTER_REG_21_ & ~n7683;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = n6754 & ~n7686;
  assign n7688 = PHYADDRPOINTER_REG_21_ & n6748;
  assign n7689 = n6262 & n6749;
  assign n7690 = n7666 & ~n7673;
  assign n7691 = ~n7669 & n7690;
  assign n7692 = ~n7672 & ~n7691;
  assign n7693 = INSTQUEUE_REG_7__5_ & n7322;
  assign n7694 = INSTQUEUE_REG_6__5_ & n7324;
  assign n7695 = INSTQUEUE_REG_5__5_ & n7326;
  assign n7696 = INSTQUEUE_REG_4__5_ & n7328;
  assign n7697 = ~n7693 & ~n7694;
  assign n7698 = ~n7695 & n7697;
  assign n7699 = ~n7696 & n7698;
  assign n7700 = INSTQUEUE_REG_3__5_ & n7334;
  assign n7701 = INSTQUEUE_REG_2__5_ & n7336;
  assign n7702 = INSTQUEUE_REG_1__5_ & n7338;
  assign n7703 = INSTQUEUE_REG_0__5_ & n7340;
  assign n7704 = ~n7700 & ~n7701;
  assign n7705 = ~n7702 & n7704;
  assign n7706 = ~n7703 & n7705;
  assign n7707 = INSTQUEUE_REG_15__5_ & n7346;
  assign n7708 = INSTQUEUE_REG_14__5_ & n7348;
  assign n7709 = INSTQUEUE_REG_13__5_ & n7350;
  assign n7710 = INSTQUEUE_REG_12__5_ & n7352;
  assign n7711 = ~n7707 & ~n7708;
  assign n7712 = ~n7709 & n7711;
  assign n7713 = ~n7710 & n7712;
  assign n7714 = INSTQUEUE_REG_11__5_ & n7358;
  assign n7715 = INSTQUEUE_REG_10__5_ & n7360;
  assign n7716 = INSTQUEUE_REG_9__5_ & n7362;
  assign n7717 = INSTQUEUE_REG_8__5_ & n7364;
  assign n7718 = ~n7714 & ~n7715;
  assign n7719 = ~n7716 & n7718;
  assign n7720 = ~n7717 & n7719;
  assign n7721 = n7699 & n7706;
  assign n7722 = n7713 & n7721;
  assign n7723 = n7720 & n7722;
  assign n7724 = ~n7374 & ~n7723;
  assign n7725 = ~n6766 & n7724;
  assign n7726 = EAX_REG_21_ & n6759;
  assign n7727 = PHYADDRPOINTER_REG_21_ & n6763;
  assign n7728 = n2682 & ~n7686;
  assign n7729 = ~n7726 & ~n7727;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = ~n7725 & n7730;
  assign n7732 = ~n2682 & ~n7731;
  assign n7733 = n2682 & n7731;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = n7423 & ~n7734;
  assign n7736 = ~n7423 & n7734;
  assign n7737 = ~n7735 & ~n7736;
  assign n7738 = ~n7692 & ~n7737;
  assign n7739 = ~n7672 & ~n7736;
  assign n7740 = ~n7735 & n7739;
  assign n7741 = n7670 & ~n7673;
  assign n7742 = n7740 & ~n7741;
  assign n7743 = ~n7738 & ~n7742;
  assign n7744 = n6785 & n7743;
  assign n7745 = ~n7682 & ~n7687;
  assign n7746 = ~n7688 & n7745;
  assign n7747 = ~n7689 & n7746;
  assign n1500 = n7744 | ~n7747;
  assign n7749 = REIP_REG_22_ & n6756;
  assign n7750 = PHYADDRPOINTER_REG_20_ & PHYADDRPOINTER_REG_21_;
  assign n7751 = n7613 & n7750;
  assign n7752 = ~PHYADDRPOINTER_REG_22_ & n7751;
  assign n7753 = PHYADDRPOINTER_REG_22_ & ~n7751;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = n6754 & ~n7754;
  assign n7756 = PHYADDRPOINTER_REG_22_ & n6748;
  assign n7757 = n6308 & n6749;
  assign n7758 = INSTQUEUE_REG_7__6_ & n7322;
  assign n7759 = INSTQUEUE_REG_6__6_ & n7324;
  assign n7760 = INSTQUEUE_REG_5__6_ & n7326;
  assign n7761 = INSTQUEUE_REG_4__6_ & n7328;
  assign n7762 = ~n7758 & ~n7759;
  assign n7763 = ~n7760 & n7762;
  assign n7764 = ~n7761 & n7763;
  assign n7765 = INSTQUEUE_REG_3__6_ & n7334;
  assign n7766 = INSTQUEUE_REG_2__6_ & n7336;
  assign n7767 = INSTQUEUE_REG_1__6_ & n7338;
  assign n7768 = INSTQUEUE_REG_0__6_ & n7340;
  assign n7769 = ~n7765 & ~n7766;
  assign n7770 = ~n7767 & n7769;
  assign n7771 = ~n7768 & n7770;
  assign n7772 = INSTQUEUE_REG_15__6_ & n7346;
  assign n7773 = INSTQUEUE_REG_14__6_ & n7348;
  assign n7774 = INSTQUEUE_REG_13__6_ & n7350;
  assign n7775 = INSTQUEUE_REG_12__6_ & n7352;
  assign n7776 = ~n7772 & ~n7773;
  assign n7777 = ~n7774 & n7776;
  assign n7778 = ~n7775 & n7777;
  assign n7779 = INSTQUEUE_REG_11__6_ & n7358;
  assign n7780 = INSTQUEUE_REG_10__6_ & n7360;
  assign n7781 = INSTQUEUE_REG_9__6_ & n7362;
  assign n7782 = INSTQUEUE_REG_8__6_ & n7364;
  assign n7783 = ~n7779 & ~n7780;
  assign n7784 = ~n7781 & n7783;
  assign n7785 = ~n7782 & n7784;
  assign n7786 = n7764 & n7771;
  assign n7787 = n7778 & n7786;
  assign n7788 = n7785 & n7787;
  assign n7789 = ~n7374 & ~n7788;
  assign n7790 = ~n6766 & n7789;
  assign n7791 = EAX_REG_22_ & n6759;
  assign n7792 = PHYADDRPOINTER_REG_22_ & n6763;
  assign n7793 = n2682 & ~n7754;
  assign n7794 = ~n7791 & ~n7792;
  assign n7795 = ~n7793 & n7794;
  assign n7796 = ~n7790 & n7795;
  assign n7797 = ~n2682 & ~n7796;
  assign n7798 = n2682 & n7796;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = ~n7423 & n7799;
  assign n7801 = n7423 & ~n7799;
  assign n7802 = ~n7800 & ~n7801;
  assign n7803 = ~n7692 & ~n7735;
  assign n7804 = ~n7736 & ~n7803;
  assign n7805 = n7802 & ~n7804;
  assign n7806 = ~n7802 & n7804;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = n6785 & ~n7807;
  assign n7809 = ~n7749 & ~n7755;
  assign n7810 = ~n7756 & n7809;
  assign n7811 = ~n7757 & n7810;
  assign n1505 = n7808 | ~n7811;
  assign n7813 = REIP_REG_23_ & n6756;
  assign n7814 = PHYADDRPOINTER_REG_22_ & n7751;
  assign n7815 = ~PHYADDRPOINTER_REG_23_ & n7814;
  assign n7816 = PHYADDRPOINTER_REG_23_ & ~n7814;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = n6754 & ~n7817;
  assign n7819 = PHYADDRPOINTER_REG_23_ & n6748;
  assign n7820 = n6355 & n6749;
  assign n7821 = INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign n7822 = ~n1750_1 & ~n7821;
  assign n7823 = n1954 & n7822;
  assign n7824 = INSTQUEUE_REG_7__0_ & n7823;
  assign n7825 = n1958_1 & n7822;
  assign n7826 = INSTQUEUE_REG_6__0_ & n7825;
  assign n7827 = INSTQUEUERD_ADDR_REG_0_ & n1733;
  assign n7828 = n7822 & n7827;
  assign n7829 = INSTQUEUE_REG_5__0_ & n7828;
  assign n7830 = n1736 & n7822;
  assign n7831 = INSTQUEUE_REG_4__0_ & n7830;
  assign n7832 = ~n7824 & ~n7826;
  assign n7833 = ~n7829 & n7832;
  assign n7834 = ~n7831 & n7833;
  assign n7835 = INSTQUEUERD_ADDR_REG_2_ & n7822;
  assign n7836 = n1753 & n7835;
  assign n7837 = INSTQUEUE_REG_3__0_ & n7836;
  assign n7838 = n1760 & n7835;
  assign n7839 = INSTQUEUE_REG_2__0_ & n7838;
  assign n7840 = n1763 & n7835;
  assign n7841 = INSTQUEUE_REG_1__0_ & n7840;
  assign n7842 = n1722_1 & n7835;
  assign n7843 = INSTQUEUE_REG_0__0_ & n7842;
  assign n7844 = ~n7837 & ~n7839;
  assign n7845 = ~n7841 & n7844;
  assign n7846 = ~n7843 & n7845;
  assign n7847 = n1954 & ~n7822;
  assign n7848 = INSTQUEUE_REG_15__0_ & n7847;
  assign n7849 = n1958_1 & ~n7822;
  assign n7850 = INSTQUEUE_REG_14__0_ & n7849;
  assign n7851 = ~n7822 & n7827;
  assign n7852 = INSTQUEUE_REG_13__0_ & n7851;
  assign n7853 = n1736 & ~n7822;
  assign n7854 = INSTQUEUE_REG_12__0_ & n7853;
  assign n7855 = ~n7848 & ~n7850;
  assign n7856 = ~n7852 & n7855;
  assign n7857 = ~n7854 & n7856;
  assign n7858 = INSTQUEUERD_ADDR_REG_2_ & ~n7822;
  assign n7859 = n1753 & n7858;
  assign n7860 = INSTQUEUE_REG_11__0_ & n7859;
  assign n7861 = n1760 & n7858;
  assign n7862 = INSTQUEUE_REG_10__0_ & n7861;
  assign n7863 = n1763 & n7858;
  assign n7864 = INSTQUEUE_REG_9__0_ & n7863;
  assign n7865 = n1722_1 & n7858;
  assign n7866 = INSTQUEUE_REG_8__0_ & n7865;
  assign n7867 = ~n7860 & ~n7862;
  assign n7868 = ~n7864 & n7867;
  assign n7869 = ~n7866 & n7868;
  assign n7870 = n7834 & n7846;
  assign n7871 = n7857 & n7870;
  assign n7872 = n7869 & n7871;
  assign n7873 = ~n7374 & ~n7872;
  assign n7874 = INSTQUEUE_REG_7__7_ & n7322;
  assign n7875 = INSTQUEUE_REG_6__7_ & n7324;
  assign n7876 = INSTQUEUE_REG_5__7_ & n7326;
  assign n7877 = INSTQUEUE_REG_4__7_ & n7328;
  assign n7878 = ~n7874 & ~n7875;
  assign n7879 = ~n7876 & n7878;
  assign n7880 = ~n7877 & n7879;
  assign n7881 = INSTQUEUE_REG_3__7_ & n7334;
  assign n7882 = INSTQUEUE_REG_2__7_ & n7336;
  assign n7883 = INSTQUEUE_REG_1__7_ & n7338;
  assign n7884 = INSTQUEUE_REG_0__7_ & n7340;
  assign n7885 = ~n7881 & ~n7882;
  assign n7886 = ~n7883 & n7885;
  assign n7887 = ~n7884 & n7886;
  assign n7888 = INSTQUEUE_REG_15__7_ & n7346;
  assign n7889 = INSTQUEUE_REG_14__7_ & n7348;
  assign n7890 = INSTQUEUE_REG_13__7_ & n7350;
  assign n7891 = INSTQUEUE_REG_12__7_ & n7352;
  assign n7892 = ~n7888 & ~n7889;
  assign n7893 = ~n7890 & n7892;
  assign n7894 = ~n7891 & n7893;
  assign n7895 = INSTQUEUE_REG_11__7_ & n7358;
  assign n7896 = INSTQUEUE_REG_10__7_ & n7360;
  assign n7897 = INSTQUEUE_REG_9__7_ & n7362;
  assign n7898 = INSTQUEUE_REG_8__7_ & n7364;
  assign n7899 = ~n7895 & ~n7896;
  assign n7900 = ~n7897 & n7899;
  assign n7901 = ~n7898 & n7900;
  assign n7902 = n7880 & n7887;
  assign n7903 = n7894 & n7902;
  assign n7904 = n7901 & n7903;
  assign n7905 = ~n7374 & ~n7904;
  assign n7906 = ~n7873 & ~n7905;
  assign n7907 = n7873 & n7905;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = ~n6766 & n7908;
  assign n7910 = EAX_REG_23_ & n6759;
  assign n7911 = PHYADDRPOINTER_REG_23_ & n6763;
  assign n7912 = n2682 & ~n7817;
  assign n7913 = ~n7910 & ~n7911;
  assign n7914 = ~n7912 & n7913;
  assign n7915 = ~n7909 & n7914;
  assign n7916 = ~n2682 & ~n7915;
  assign n7917 = n2682 & n7915;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = ~n7423 & n7918;
  assign n7920 = n7423 & ~n7918;
  assign n7921 = ~n7919 & ~n7920;
  assign n7922 = n7403 & n7666;
  assign n7923 = n7739 & ~n7800;
  assign n7924 = n7666 & ~n7668;
  assign n7925 = n7923 & ~n7924;
  assign n7926 = ~n7922 & n7925;
  assign n7927 = ~n7735 & ~n7801;
  assign n7928 = n7673 & ~n7736;
  assign n7929 = n7927 & ~n7928;
  assign n7930 = ~n7800 & ~n7929;
  assign n7931 = ~n7926 & ~n7930;
  assign n7932 = n7921 & n7931;
  assign n7933 = ~n7921 & ~n7931;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = n6785 & ~n7934;
  assign n7936 = ~n7813 & ~n7818;
  assign n7937 = ~n7819 & n7936;
  assign n7938 = ~n7820 & n7937;
  assign n1510 = n7935 | ~n7938;
  assign n7940 = REIP_REG_24_ & n6756;
  assign n7941 = PHYADDRPOINTER_REG_22_ & PHYADDRPOINTER_REG_23_;
  assign n7942 = n7751 & n7941;
  assign n7943 = ~PHYADDRPOINTER_REG_24_ & n7942;
  assign n7944 = PHYADDRPOINTER_REG_24_ & ~n7942;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n6754 & ~n7945;
  assign n7947 = PHYADDRPOINTER_REG_24_ & n6748;
  assign n7948 = n6401 & n6749;
  assign n7949 = INSTQUEUE_REG_7__1_ & n7823;
  assign n7950 = INSTQUEUE_REG_6__1_ & n7825;
  assign n7951 = INSTQUEUE_REG_5__1_ & n7828;
  assign n7952 = INSTQUEUE_REG_4__1_ & n7830;
  assign n7953 = ~n7949 & ~n7950;
  assign n7954 = ~n7951 & n7953;
  assign n7955 = ~n7952 & n7954;
  assign n7956 = INSTQUEUE_REG_3__1_ & n7836;
  assign n7957 = INSTQUEUE_REG_2__1_ & n7838;
  assign n7958 = INSTQUEUE_REG_1__1_ & n7840;
  assign n7959 = INSTQUEUE_REG_0__1_ & n7842;
  assign n7960 = ~n7956 & ~n7957;
  assign n7961 = ~n7958 & n7960;
  assign n7962 = ~n7959 & n7961;
  assign n7963 = INSTQUEUE_REG_15__1_ & n7847;
  assign n7964 = INSTQUEUE_REG_14__1_ & n7849;
  assign n7965 = INSTQUEUE_REG_13__1_ & n7851;
  assign n7966 = INSTQUEUE_REG_12__1_ & n7853;
  assign n7967 = ~n7963 & ~n7964;
  assign n7968 = ~n7965 & n7967;
  assign n7969 = ~n7966 & n7968;
  assign n7970 = INSTQUEUE_REG_11__1_ & n7859;
  assign n7971 = INSTQUEUE_REG_10__1_ & n7861;
  assign n7972 = INSTQUEUE_REG_9__1_ & n7863;
  assign n7973 = INSTQUEUE_REG_8__1_ & n7865;
  assign n7974 = ~n7970 & ~n7971;
  assign n7975 = ~n7972 & n7974;
  assign n7976 = ~n7973 & n7975;
  assign n7977 = n7955 & n7962;
  assign n7978 = n7969 & n7977;
  assign n7979 = n7976 & n7978;
  assign n7980 = ~n7374 & ~n7979;
  assign n7981 = ~n7907 & n7980;
  assign n7982 = n7907 & ~n7980;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = ~n6766 & ~n7983;
  assign n7985 = EAX_REG_24_ & n6759;
  assign n7986 = PHYADDRPOINTER_REG_24_ & n6763;
  assign n7987 = n2682 & ~n7945;
  assign n7988 = ~n7985 & ~n7986;
  assign n7989 = ~n7987 & n7988;
  assign n7990 = ~n7984 & n7989;
  assign n7991 = ~n2682 & ~n7990;
  assign n7992 = n2682 & n7990;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = n7423 & ~n7993;
  assign n7995 = ~n7423 & n7993;
  assign n7996 = ~n7994 & ~n7995;
  assign n7997 = ~n7919 & ~n7931;
  assign n7998 = ~n7920 & ~n7997;
  assign n7999 = n7996 & n7998;
  assign n8000 = ~n7996 & ~n7998;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = n6785 & ~n8001;
  assign n8003 = ~n7940 & ~n7946;
  assign n8004 = ~n7947 & n8003;
  assign n8005 = ~n7948 & n8004;
  assign n1515 = n8002 | ~n8005;
  assign n8007 = REIP_REG_25_ & n6756;
  assign n8008 = PHYADDRPOINTER_REG_24_ & n7942;
  assign n8009 = ~PHYADDRPOINTER_REG_25_ & n8008;
  assign n8010 = PHYADDRPOINTER_REG_25_ & ~n8008;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = n6754 & ~n8011;
  assign n8013 = PHYADDRPOINTER_REG_25_ & n6748;
  assign n8014 = n6448 & n6749;
  assign n8015 = n7907 & n7980;
  assign n8016 = INSTQUEUE_REG_7__2_ & n7823;
  assign n8017 = INSTQUEUE_REG_6__2_ & n7825;
  assign n8018 = INSTQUEUE_REG_5__2_ & n7828;
  assign n8019 = INSTQUEUE_REG_4__2_ & n7830;
  assign n8020 = ~n8016 & ~n8017;
  assign n8021 = ~n8018 & n8020;
  assign n8022 = ~n8019 & n8021;
  assign n8023 = INSTQUEUE_REG_3__2_ & n7836;
  assign n8024 = INSTQUEUE_REG_2__2_ & n7838;
  assign n8025 = INSTQUEUE_REG_1__2_ & n7840;
  assign n8026 = INSTQUEUE_REG_0__2_ & n7842;
  assign n8027 = ~n8023 & ~n8024;
  assign n8028 = ~n8025 & n8027;
  assign n8029 = ~n8026 & n8028;
  assign n8030 = INSTQUEUE_REG_15__2_ & n7847;
  assign n8031 = INSTQUEUE_REG_14__2_ & n7849;
  assign n8032 = INSTQUEUE_REG_13__2_ & n7851;
  assign n8033 = INSTQUEUE_REG_12__2_ & n7853;
  assign n8034 = ~n8030 & ~n8031;
  assign n8035 = ~n8032 & n8034;
  assign n8036 = ~n8033 & n8035;
  assign n8037 = INSTQUEUE_REG_11__2_ & n7859;
  assign n8038 = INSTQUEUE_REG_10__2_ & n7861;
  assign n8039 = INSTQUEUE_REG_9__2_ & n7863;
  assign n8040 = INSTQUEUE_REG_8__2_ & n7865;
  assign n8041 = ~n8037 & ~n8038;
  assign n8042 = ~n8039 & n8041;
  assign n8043 = ~n8040 & n8042;
  assign n8044 = n8022 & n8029;
  assign n8045 = n8036 & n8044;
  assign n8046 = n8043 & n8045;
  assign n8047 = ~n7374 & ~n8046;
  assign n8048 = n8015 & ~n8047;
  assign n8049 = ~n8015 & n8047;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = ~n6766 & ~n8050;
  assign n8052 = EAX_REG_25_ & n6759;
  assign n8053 = PHYADDRPOINTER_REG_25_ & n6763;
  assign n8054 = n2682 & ~n8011;
  assign n8055 = ~n8052 & ~n8053;
  assign n8056 = ~n8054 & n8055;
  assign n8057 = ~n8051 & n8056;
  assign n8058 = ~n2682 & ~n8057;
  assign n8059 = n2682 & n8057;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = ~n7423 & n8060;
  assign n8062 = n7423 & ~n8060;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n7919 & ~n7995;
  assign n8065 = n7923 & n8064;
  assign n8066 = ~n7666 & n8065;
  assign n8067 = ~n7920 & ~n7930;
  assign n8068 = n8064 & ~n8067;
  assign n8069 = ~n7994 & ~n8068;
  assign n8070 = ~n8066 & n8069;
  assign n8071 = n7668 & n8065;
  assign n8072 = ~n7403 & n8071;
  assign n8073 = n8070 & ~n8072;
  assign n8074 = n8063 & n8073;
  assign n8075 = ~n8063 & ~n8073;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = n6785 & ~n8076;
  assign n8078 = ~n8007 & ~n8012;
  assign n8079 = ~n8013 & n8078;
  assign n8080 = ~n8014 & n8079;
  assign n1520 = n8077 | ~n8080;
  assign n8082 = REIP_REG_26_ & n6756;
  assign n8083 = PHYADDRPOINTER_REG_24_ & PHYADDRPOINTER_REG_25_;
  assign n8084 = n7942 & n8083;
  assign n8085 = ~PHYADDRPOINTER_REG_26_ & n8084;
  assign n8086 = PHYADDRPOINTER_REG_26_ & ~n8084;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = n6754 & ~n8087;
  assign n8089 = PHYADDRPOINTER_REG_26_ & n6748;
  assign n8090 = n6499 & n6749;
  assign n8091 = INSTQUEUE_REG_7__3_ & n7823;
  assign n8092 = INSTQUEUE_REG_6__3_ & n7825;
  assign n8093 = INSTQUEUE_REG_5__3_ & n7828;
  assign n8094 = INSTQUEUE_REG_4__3_ & n7830;
  assign n8095 = ~n8091 & ~n8092;
  assign n8096 = ~n8093 & n8095;
  assign n8097 = ~n8094 & n8096;
  assign n8098 = INSTQUEUE_REG_3__3_ & n7836;
  assign n8099 = INSTQUEUE_REG_2__3_ & n7838;
  assign n8100 = INSTQUEUE_REG_1__3_ & n7840;
  assign n8101 = INSTQUEUE_REG_0__3_ & n7842;
  assign n8102 = ~n8098 & ~n8099;
  assign n8103 = ~n8100 & n8102;
  assign n8104 = ~n8101 & n8103;
  assign n8105 = INSTQUEUE_REG_15__3_ & n7847;
  assign n8106 = INSTQUEUE_REG_14__3_ & n7849;
  assign n8107 = INSTQUEUE_REG_13__3_ & n7851;
  assign n8108 = INSTQUEUE_REG_12__3_ & n7853;
  assign n8109 = ~n8105 & ~n8106;
  assign n8110 = ~n8107 & n8109;
  assign n8111 = ~n8108 & n8110;
  assign n8112 = INSTQUEUE_REG_11__3_ & n7859;
  assign n8113 = INSTQUEUE_REG_10__3_ & n7861;
  assign n8114 = INSTQUEUE_REG_9__3_ & n7863;
  assign n8115 = INSTQUEUE_REG_8__3_ & n7865;
  assign n8116 = ~n8112 & ~n8113;
  assign n8117 = ~n8114 & n8116;
  assign n8118 = ~n8115 & n8117;
  assign n8119 = n8097 & n8104;
  assign n8120 = n8111 & n8119;
  assign n8121 = n8118 & n8120;
  assign n8122 = ~n7374 & ~n8121;
  assign n8123 = n7980 & n8047;
  assign n8124 = n7907 & n8123;
  assign n8125 = n8122 & ~n8124;
  assign n8126 = ~n8122 & n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~n6766 & ~n8127;
  assign n8129 = EAX_REG_26_ & n6759;
  assign n8130 = PHYADDRPOINTER_REG_26_ & n6763;
  assign n8131 = n2682 & ~n8087;
  assign n8132 = ~n8129 & ~n8130;
  assign n8133 = ~n8131 & n8132;
  assign n8134 = ~n8128 & n8133;
  assign n8135 = ~n2682 & ~n8134;
  assign n8136 = n2682 & n8134;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~n7423 & n8137;
  assign n8139 = n7423 & ~n8137;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n8061 & ~n8073;
  assign n8142 = ~n8062 & ~n8141;
  assign n8143 = n8140 & n8142;
  assign n8144 = ~n8140 & ~n8142;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = n6785 & ~n8145;
  assign n8147 = ~n8082 & ~n8088;
  assign n8148 = ~n8089 & n8147;
  assign n8149 = ~n8090 & n8148;
  assign n1525 = n8146 | ~n8149;
  assign n8151 = REIP_REG_27_ & n6756;
  assign n8152 = PHYADDRPOINTER_REG_26_ & n8084;
  assign n8153 = ~PHYADDRPOINTER_REG_27_ & n8152;
  assign n8154 = PHYADDRPOINTER_REG_27_ & ~n8152;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = n6754 & ~n8155;
  assign n8157 = PHYADDRPOINTER_REG_27_ & n6748;
  assign n8158 = n6543 & n6749;
  assign n8159 = n8122 & n8124;
  assign n8160 = INSTQUEUE_REG_0__4_ & n7842;
  assign n8161 = INSTQUEUE_REG_7__4_ & n7823;
  assign n8162 = INSTQUEUE_REG_6__4_ & n7825;
  assign n8163 = INSTQUEUE_REG_5__4_ & n7828;
  assign n8164 = ~n8162 & ~n8163;
  assign n8165 = ~n8160 & ~n8161;
  assign n8166 = n8164 & n8165;
  assign n8167 = INSTQUEUE_REG_4__4_ & n7830;
  assign n8168 = INSTQUEUE_REG_3__4_ & n7836;
  assign n8169 = INSTQUEUE_REG_2__4_ & n7838;
  assign n8170 = INSTQUEUE_REG_1__4_ & n7840;
  assign n8171 = ~n8167 & ~n8168;
  assign n8172 = ~n8169 & n8171;
  assign n8173 = ~n8170 & n8172;
  assign n8174 = INSTQUEUE_REG_15__4_ & n7847;
  assign n8175 = INSTQUEUE_REG_14__4_ & n7849;
  assign n8176 = INSTQUEUE_REG_13__4_ & n7851;
  assign n8177 = INSTQUEUE_REG_12__4_ & n7853;
  assign n8178 = ~n8174 & ~n8175;
  assign n8179 = ~n8176 & n8178;
  assign n8180 = ~n8177 & n8179;
  assign n8181 = INSTQUEUE_REG_11__4_ & n7859;
  assign n8182 = INSTQUEUE_REG_10__4_ & n7861;
  assign n8183 = INSTQUEUE_REG_9__4_ & n7863;
  assign n8184 = INSTQUEUE_REG_8__4_ & n7865;
  assign n8185 = ~n8181 & ~n8182;
  assign n8186 = ~n8183 & n8185;
  assign n8187 = ~n8184 & n8186;
  assign n8188 = n8166 & n8173;
  assign n8189 = n8180 & n8188;
  assign n8190 = n8187 & n8189;
  assign n8191 = ~n7374 & ~n8190;
  assign n8192 = n8159 & ~n8191;
  assign n8193 = ~n8159 & n8191;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = ~n6766 & ~n8194;
  assign n8196 = EAX_REG_27_ & n6759;
  assign n8197 = PHYADDRPOINTER_REG_27_ & n6763;
  assign n8198 = n2682 & ~n8155;
  assign n8199 = ~n8196 & ~n8197;
  assign n8200 = ~n8198 & n8199;
  assign n8201 = ~n8195 & n8200;
  assign n8202 = ~n2682 & ~n8201;
  assign n8203 = n2682 & n8201;
  assign n8204 = ~n8202 & ~n8203;
  assign n8205 = n7423 & ~n8204;
  assign n8206 = ~n7423 & n8204;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n8062 & ~n8139;
  assign n8209 = ~n8141 & n8208;
  assign n8210 = ~n8138 & ~n8209;
  assign n8211 = n8207 & ~n8210;
  assign n8212 = ~n8207 & n8210;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = n6785 & ~n8213;
  assign n8215 = ~n8151 & ~n8156;
  assign n8216 = ~n8157 & n8215;
  assign n8217 = ~n8158 & n8216;
  assign n1530 = n8214 | ~n8217;
  assign n8219 = REIP_REG_28_ & n6756;
  assign n8220 = PHYADDRPOINTER_REG_27_ & n8152;
  assign n8221 = ~PHYADDRPOINTER_REG_28_ & n8220;
  assign n8222 = PHYADDRPOINTER_REG_28_ & ~n8220;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = n6754 & ~n8223;
  assign n8225 = PHYADDRPOINTER_REG_28_ & n6748;
  assign n8226 = n6589 & n6749;
  assign n8227 = INSTQUEUE_REG_7__5_ & n7823;
  assign n8228 = INSTQUEUE_REG_6__5_ & n7825;
  assign n8229 = INSTQUEUE_REG_5__5_ & n7828;
  assign n8230 = INSTQUEUE_REG_4__5_ & n7830;
  assign n8231 = ~n8227 & ~n8228;
  assign n8232 = ~n8229 & n8231;
  assign n8233 = ~n8230 & n8232;
  assign n8234 = INSTQUEUE_REG_3__5_ & n7836;
  assign n8235 = INSTQUEUE_REG_2__5_ & n7838;
  assign n8236 = INSTQUEUE_REG_1__5_ & n7840;
  assign n8237 = INSTQUEUE_REG_0__5_ & n7842;
  assign n8238 = ~n8234 & ~n8235;
  assign n8239 = ~n8236 & n8238;
  assign n8240 = ~n8237 & n8239;
  assign n8241 = INSTQUEUE_REG_15__5_ & n7847;
  assign n8242 = INSTQUEUE_REG_14__5_ & n7849;
  assign n8243 = INSTQUEUE_REG_13__5_ & n7851;
  assign n8244 = INSTQUEUE_REG_12__5_ & n7853;
  assign n8245 = ~n8241 & ~n8242;
  assign n8246 = ~n8243 & n8245;
  assign n8247 = ~n8244 & n8246;
  assign n8248 = INSTQUEUE_REG_11__5_ & n7859;
  assign n8249 = INSTQUEUE_REG_10__5_ & n7861;
  assign n8250 = INSTQUEUE_REG_9__5_ & n7863;
  assign n8251 = INSTQUEUE_REG_8__5_ & n7865;
  assign n8252 = ~n8248 & ~n8249;
  assign n8253 = ~n8250 & n8252;
  assign n8254 = ~n8251 & n8253;
  assign n8255 = n8233 & n8240;
  assign n8256 = n8247 & n8255;
  assign n8257 = n8254 & n8256;
  assign n8258 = ~n7374 & ~n8257;
  assign n8259 = n8122 & n8191;
  assign n8260 = n8124 & n8259;
  assign n8261 = n8258 & ~n8260;
  assign n8262 = ~n8258 & n8260;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = ~n6766 & ~n8263;
  assign n8265 = EAX_REG_28_ & n6759;
  assign n8266 = PHYADDRPOINTER_REG_28_ & n6763;
  assign n8267 = n2682 & ~n8223;
  assign n8268 = ~n8265 & ~n8266;
  assign n8269 = ~n8267 & n8268;
  assign n8270 = ~n8264 & n8269;
  assign n8271 = ~n2682 & ~n8270;
  assign n8272 = n2682 & n8270;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = n7423 & ~n8273;
  assign n8275 = ~n7423 & n8273;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n8138 & ~n8206;
  assign n8278 = ~n8208 & n8277;
  assign n8279 = ~n8205 & ~n8278;
  assign n8280 = ~n8061 & n8277;
  assign n8281 = ~n8073 & n8280;
  assign n8282 = n8279 & ~n8281;
  assign n8283 = n8276 & n8282;
  assign n8284 = ~n8276 & ~n8282;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = n6785 & ~n8285;
  assign n8287 = ~n8219 & ~n8224;
  assign n8288 = ~n8225 & n8287;
  assign n8289 = ~n8226 & n8288;
  assign n1535 = n8286 | ~n8289;
  assign n8291 = REIP_REG_29_ & n6756;
  assign n8292 = PHYADDRPOINTER_REG_28_ & n8220;
  assign n8293 = ~PHYADDRPOINTER_REG_29_ & n8292;
  assign n8294 = PHYADDRPOINTER_REG_29_ & ~n8292;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = n6754 & ~n8295;
  assign n8297 = PHYADDRPOINTER_REG_29_ & n6748;
  assign n8298 = n6638 & n6749;
  assign n8299 = n8258 & n8260;
  assign n8300 = INSTQUEUE_REG_7__6_ & n7823;
  assign n8301 = INSTQUEUE_REG_6__6_ & n7825;
  assign n8302 = INSTQUEUE_REG_5__6_ & n7828;
  assign n8303 = INSTQUEUE_REG_4__6_ & n7830;
  assign n8304 = ~n8300 & ~n8301;
  assign n8305 = ~n8302 & n8304;
  assign n8306 = ~n8303 & n8305;
  assign n8307 = INSTQUEUE_REG_3__6_ & n7836;
  assign n8308 = INSTQUEUE_REG_2__6_ & n7838;
  assign n8309 = INSTQUEUE_REG_1__6_ & n7840;
  assign n8310 = INSTQUEUE_REG_0__6_ & n7842;
  assign n8311 = ~n8307 & ~n8308;
  assign n8312 = ~n8309 & n8311;
  assign n8313 = ~n8310 & n8312;
  assign n8314 = INSTQUEUE_REG_15__6_ & n7847;
  assign n8315 = INSTQUEUE_REG_14__6_ & n7849;
  assign n8316 = INSTQUEUE_REG_13__6_ & n7851;
  assign n8317 = INSTQUEUE_REG_12__6_ & n7853;
  assign n8318 = ~n8314 & ~n8315;
  assign n8319 = ~n8316 & n8318;
  assign n8320 = ~n8317 & n8319;
  assign n8321 = INSTQUEUE_REG_11__6_ & n7859;
  assign n8322 = INSTQUEUE_REG_10__6_ & n7861;
  assign n8323 = INSTQUEUE_REG_9__6_ & n7863;
  assign n8324 = INSTQUEUE_REG_8__6_ & n7865;
  assign n8325 = ~n8321 & ~n8322;
  assign n8326 = ~n8323 & n8325;
  assign n8327 = ~n8324 & n8326;
  assign n8328 = n8306 & n8313;
  assign n8329 = n8320 & n8328;
  assign n8330 = n8327 & n8329;
  assign n8331 = ~n7374 & ~n8330;
  assign n8332 = n8299 & ~n8331;
  assign n8333 = ~n8299 & n8331;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~n6766 & ~n8334;
  assign n8336 = EAX_REG_29_ & n6759;
  assign n8337 = PHYADDRPOINTER_REG_29_ & n6763;
  assign n8338 = n2682 & ~n8295;
  assign n8339 = ~n8336 & ~n8337;
  assign n8340 = ~n8338 & n8339;
  assign n8341 = ~n8335 & n8340;
  assign n8342 = ~n2682 & ~n8341;
  assign n8343 = n2682 & n8341;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = n7423 & ~n8344;
  assign n8346 = ~n7423 & n8344;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = ~n8061 & ~n8138;
  assign n8349 = ~n8206 & n8348;
  assign n8350 = ~n8275 & n8349;
  assign n8351 = ~n8073 & n8350;
  assign n8352 = ~n8205 & ~n8274;
  assign n8353 = ~n8278 & n8352;
  assign n8354 = ~n8275 & ~n8353;
  assign n8355 = ~n8351 & ~n8354;
  assign n8356 = n8347 & n8355;
  assign n8357 = ~n8347 & ~n8355;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = n6785 & ~n8358;
  assign n8360 = ~n8291 & ~n8296;
  assign n8361 = ~n8297 & n8360;
  assign n8362 = ~n8298 & n8361;
  assign n1540 = n8359 | ~n8362;
  assign n8364 = REIP_REG_30_ & n6756;
  assign n8365 = PHYADDRPOINTER_REG_29_ & n8292;
  assign n8366 = ~PHYADDRPOINTER_REG_30_ & n8365;
  assign n8367 = PHYADDRPOINTER_REG_30_ & ~n8365;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = n6754 & ~n8368;
  assign n8370 = PHYADDRPOINTER_REG_30_ & n6748;
  assign n8371 = n6686 & n6749;
  assign n8372 = n8299 & n8331;
  assign n8373 = INSTQUEUE_REG_7__7_ & n7823;
  assign n8374 = INSTQUEUE_REG_6__7_ & n7825;
  assign n8375 = INSTQUEUE_REG_5__7_ & n7828;
  assign n8376 = INSTQUEUE_REG_4__7_ & n7830;
  assign n8377 = ~n8373 & ~n8374;
  assign n8378 = ~n8375 & n8377;
  assign n8379 = ~n8376 & n8378;
  assign n8380 = INSTQUEUE_REG_3__7_ & n7836;
  assign n8381 = INSTQUEUE_REG_2__7_ & n7838;
  assign n8382 = INSTQUEUE_REG_1__7_ & n7840;
  assign n8383 = INSTQUEUE_REG_0__7_ & n7842;
  assign n8384 = ~n8380 & ~n8381;
  assign n8385 = ~n8382 & n8384;
  assign n8386 = ~n8383 & n8385;
  assign n8387 = INSTQUEUE_REG_15__7_ & n7847;
  assign n8388 = INSTQUEUE_REG_14__7_ & n7849;
  assign n8389 = INSTQUEUE_REG_13__7_ & n7851;
  assign n8390 = INSTQUEUE_REG_12__7_ & n7853;
  assign n8391 = ~n8387 & ~n8388;
  assign n8392 = ~n8389 & n8391;
  assign n8393 = ~n8390 & n8392;
  assign n8394 = INSTQUEUE_REG_11__7_ & n7859;
  assign n8395 = INSTQUEUE_REG_10__7_ & n7861;
  assign n8396 = INSTQUEUE_REG_9__7_ & n7863;
  assign n8397 = INSTQUEUE_REG_8__7_ & n7865;
  assign n8398 = ~n8394 & ~n8395;
  assign n8399 = ~n8396 & n8398;
  assign n8400 = ~n8397 & n8399;
  assign n8401 = n8379 & n8386;
  assign n8402 = n8393 & n8401;
  assign n8403 = n8400 & n8402;
  assign n8404 = ~n7374 & ~n8403;
  assign n8405 = n8372 & ~n8404;
  assign n8406 = ~n8372 & n8404;
  assign n8407 = ~n8405 & ~n8406;
  assign n8408 = ~n6766 & ~n8407;
  assign n8409 = EAX_REG_30_ & n6759;
  assign n8410 = PHYADDRPOINTER_REG_30_ & n6763;
  assign n8411 = n2682 & ~n8368;
  assign n8412 = ~n8409 & ~n8410;
  assign n8413 = ~n8411 & n8412;
  assign n8414 = ~n8408 & n8413;
  assign n8415 = ~n2682 & ~n8414;
  assign n8416 = n2682 & n8414;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n7423 & ~n8417;
  assign n8419 = ~n7423 & n8417;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~n8275 & ~n8346;
  assign n8422 = ~n8353 & n8421;
  assign n8423 = ~n8345 & ~n8422;
  assign n8424 = ~n8346 & n8350;
  assign n8425 = ~n8073 & n8424;
  assign n8426 = n8423 & ~n8425;
  assign n8427 = n8420 & n8426;
  assign n8428 = ~n8420 & ~n8426;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = n6785 & ~n8429;
  assign n8431 = ~n8364 & ~n8369;
  assign n8432 = ~n8370 & n8431;
  assign n8433 = ~n8371 & n8432;
  assign n1545 = n8430 | ~n8433;
  assign n8435 = REIP_REG_31_ & n6756;
  assign n8436 = PHYADDRPOINTER_REG_30_ & n8365;
  assign n8437 = ~PHYADDRPOINTER_REG_31_ & n8436;
  assign n8438 = PHYADDRPOINTER_REG_31_ & ~n8436;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = n6754 & ~n8439;
  assign n8441 = PHYADDRPOINTER_REG_31_ & n6748;
  assign n8442 = n6735 & n6749;
  assign n8443 = ~n8419 & ~n8423;
  assign n8444 = ~n8418 & ~n8443;
  assign n8445 = ~n8346 & ~n8419;
  assign n8446 = n8350 & n8445;
  assign n8447 = ~n8069 & n8446;
  assign n8448 = n8065 & n8446;
  assign n8449 = ~n7666 & n8448;
  assign n8450 = n8444 & ~n8447;
  assign n8451 = ~n8449 & n8450;
  assign n8452 = n7668 & n8448;
  assign n8453 = ~n7403 & n8452;
  assign n8454 = n8451 & ~n8453;
  assign n8455 = PHYADDRPOINTER_REG_31_ & n6763;
  assign n8456 = EAX_REG_31_ & n6759;
  assign n8457 = n2682 & ~n8439;
  assign n8458 = ~n8455 & ~n8456;
  assign n8459 = ~n8457 & n8458;
  assign n8460 = ~n2682 & ~n8459;
  assign n8461 = n2682 & n8459;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = n8454 & ~n8462;
  assign n8464 = ~n8454 & n8462;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = n6785 & ~n8465;
  assign n8467 = ~n8435 & ~n8440;
  assign n8468 = ~n8441 & n8467;
  assign n8469 = ~n8442 & n8468;
  assign n1550 = n8466 | ~n8469;
  assign n8471 = READY_N & ~n2152;
  assign n8472 = ~n1776 & n2674;
  assign n8473 = ~n8471 & n8472;
  assign n8474 = ~n2262 & n8473;
  assign n8475 = ~n1807 & n8474;
  assign n8476 = DATAI_15_ & n8475;
  assign n8477 = n1807 & n8474;
  assign n8478 = EAX_REG_15_ & n8477;
  assign n8479 = ~n8476 & ~n8478;
  assign n8480 = n2282 & ~n8479;
  assign n8481 = n2282 & n8474;
  assign n8482 = LWORD_REG_15_ & ~n8481;
  assign n1555 = n8480 | n8482;
  assign n8484 = DATAI_14_ & n8475;
  assign n8485 = EAX_REG_14_ & n8477;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = n2282 & ~n8486;
  assign n8488 = LWORD_REG_14_ & ~n8481;
  assign n1560 = n8487 | n8488;
  assign n8490 = DATAI_13_ & n8475;
  assign n8491 = EAX_REG_13_ & n8477;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = n2282 & ~n8492;
  assign n8494 = LWORD_REG_13_ & ~n8481;
  assign n1565 = n8493 | n8494;
  assign n8496 = DATAI_12_ & n8475;
  assign n8497 = EAX_REG_12_ & n8477;
  assign n8498 = ~n8496 & ~n8497;
  assign n8499 = n2282 & ~n8498;
  assign n8500 = LWORD_REG_12_ & ~n8481;
  assign n1570 = n8499 | n8500;
  assign n8502 = DATAI_11_ & n8475;
  assign n8503 = EAX_REG_11_ & n8477;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = n2282 & ~n8504;
  assign n8506 = LWORD_REG_11_ & ~n8481;
  assign n1575 = n8505 | n8506;
  assign n8508 = DATAI_10_ & n8475;
  assign n8509 = EAX_REG_10_ & n8477;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = n2282 & ~n8510;
  assign n8512 = LWORD_REG_10_ & ~n8481;
  assign n1580 = n8511 | n8512;
  assign n8514 = DATAI_9_ & n8475;
  assign n8515 = EAX_REG_9_ & n8477;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = n2282 & ~n8516;
  assign n8518 = LWORD_REG_9_ & ~n8481;
  assign n1585 = n8517 | n8518;
  assign n8520 = DATAI_8_ & n8475;
  assign n8521 = EAX_REG_8_ & n8477;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = n2282 & ~n8522;
  assign n8524 = LWORD_REG_8_ & ~n8481;
  assign n1590 = n8523 | n8524;
  assign n8526 = DATAI_7_ & n8475;
  assign n8527 = EAX_REG_7_ & n8477;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = n2282 & ~n8528;
  assign n8530 = LWORD_REG_7_ & ~n8481;
  assign n1595 = n8529 | n8530;
  assign n8532 = DATAI_6_ & n8475;
  assign n8533 = EAX_REG_6_ & n8477;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = n2282 & ~n8534;
  assign n8536 = LWORD_REG_6_ & ~n8481;
  assign n1600 = n8535 | n8536;
  assign n8538 = DATAI_5_ & n8475;
  assign n8539 = EAX_REG_5_ & n8477;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = n2282 & ~n8540;
  assign n8542 = LWORD_REG_5_ & ~n8481;
  assign n1605 = n8541 | n8542;
  assign n8544 = DATAI_4_ & n8475;
  assign n8545 = EAX_REG_4_ & n8477;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = n2282 & ~n8546;
  assign n8548 = LWORD_REG_4_ & ~n8481;
  assign n1610 = n8547 | n8548;
  assign n8550 = DATAI_3_ & n8475;
  assign n8551 = EAX_REG_3_ & n8477;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = n2282 & ~n8552;
  assign n8554 = LWORD_REG_3_ & ~n8481;
  assign n1615 = n8553 | n8554;
  assign n8556 = DATAI_2_ & n8475;
  assign n8557 = EAX_REG_2_ & n8477;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = n2282 & ~n8558;
  assign n8560 = LWORD_REG_2_ & ~n8481;
  assign n1620 = n8559 | n8560;
  assign n8562 = DATAI_1_ & n8475;
  assign n8563 = EAX_REG_1_ & n8477;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = n2282 & ~n8564;
  assign n8566 = LWORD_REG_1_ & ~n8481;
  assign n1625 = n8565 | n8566;
  assign n8568 = DATAI_0_ & n8475;
  assign n8569 = EAX_REG_0_ & n8477;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = n2282 & ~n8570;
  assign n8572 = LWORD_REG_0_ & ~n8481;
  assign n1630 = n8571 | n8572;
  assign n8574 = EAX_REG_30_ & n8477;
  assign n8575 = ~n8484 & ~n8574;
  assign n8576 = n2282 & ~n8575;
  assign n8577 = UWORD_REG_14_ & ~n8481;
  assign n1635 = n8576 | n8577;
  assign n8579 = EAX_REG_29_ & n8477;
  assign n8580 = ~n8490 & ~n8579;
  assign n8581 = n2282 & ~n8580;
  assign n8582 = UWORD_REG_13_ & ~n8481;
  assign n1640 = n8581 | n8582;
  assign n8584 = EAX_REG_28_ & n8477;
  assign n8585 = ~n8496 & ~n8584;
  assign n8586 = n2282 & ~n8585;
  assign n8587 = UWORD_REG_12_ & ~n8481;
  assign n1645 = n8586 | n8587;
  assign n8589 = EAX_REG_27_ & n8477;
  assign n8590 = ~n8502 & ~n8589;
  assign n8591 = n2282 & ~n8590;
  assign n8592 = UWORD_REG_11_ & ~n8481;
  assign n1650 = n8591 | n8592;
  assign n8594 = EAX_REG_26_ & n8477;
  assign n8595 = ~n8508 & ~n8594;
  assign n8596 = n2282 & ~n8595;
  assign n8597 = UWORD_REG_10_ & ~n8481;
  assign n1655 = n8596 | n8597;
  assign n8599 = EAX_REG_25_ & n8477;
  assign n8600 = ~n8514 & ~n8599;
  assign n8601 = n2282 & ~n8600;
  assign n8602 = UWORD_REG_9_ & ~n8481;
  assign n1660 = n8601 | n8602;
  assign n8604 = EAX_REG_24_ & n8477;
  assign n8605 = ~n8520 & ~n8604;
  assign n8606 = n2282 & ~n8605;
  assign n8607 = UWORD_REG_8_ & ~n8481;
  assign n1665 = n8606 | n8607;
  assign n8609 = EAX_REG_23_ & n8477;
  assign n8610 = ~n8526 & ~n8609;
  assign n8611 = n2282 & ~n8610;
  assign n8612 = UWORD_REG_7_ & ~n8481;
  assign n1670 = n8611 | n8612;
  assign n8614 = EAX_REG_22_ & n8477;
  assign n8615 = ~n8532 & ~n8614;
  assign n8616 = n2282 & ~n8615;
  assign n8617 = UWORD_REG_6_ & ~n8481;
  assign n1675 = n8616 | n8617;
  assign n8619 = EAX_REG_21_ & n8477;
  assign n8620 = ~n8538 & ~n8619;
  assign n8621 = n2282 & ~n8620;
  assign n8622 = UWORD_REG_5_ & ~n8481;
  assign n1680 = n8621 | n8622;
  assign n8624 = EAX_REG_20_ & n8477;
  assign n8625 = ~n8544 & ~n8624;
  assign n8626 = n2282 & ~n8625;
  assign n8627 = UWORD_REG_4_ & ~n8481;
  assign n1685 = n8626 | n8627;
  assign n8629 = EAX_REG_19_ & n8477;
  assign n8630 = ~n8550 & ~n8629;
  assign n8631 = n2282 & ~n8630;
  assign n8632 = UWORD_REG_3_ & ~n8481;
  assign n1690 = n8631 | n8632;
  assign n8634 = EAX_REG_18_ & n8477;
  assign n8635 = ~n8556 & ~n8634;
  assign n8636 = n2282 & ~n8635;
  assign n8637 = UWORD_REG_2_ & ~n8481;
  assign n1695 = n8636 | n8637;
  assign n8639 = EAX_REG_17_ & n8477;
  assign n8640 = ~n8562 & ~n8639;
  assign n8641 = n2282 & ~n8640;
  assign n8642 = UWORD_REG_1_ & ~n8481;
  assign n1700 = n8641 | n8642;
  assign n8644 = EAX_REG_16_ & n8477;
  assign n8645 = ~n8568 & ~n8644;
  assign n8646 = n2282 & ~n8645;
  assign n8647 = UWORD_REG_0_ & ~n8481;
  assign n1705 = n8646 | n8647;
  assign n8649 = ~STATE2_REG_0_ & n1707;
  assign n8650 = n2152 & n2674;
  assign n8651 = n2282 & n8650;
  assign n8652 = ~n2552 & ~n8651;
  assign n8653 = n2411 & ~n8652;
  assign n8654 = n2656 & n8653;
  assign n8655 = ~n8649 & ~n8654;
  assign n8656 = STATE2_REG_0_ & ~n8655;
  assign n8657 = EAX_REG_0_ & n8656;
  assign n8658 = ~STATE2_REG_0_ & ~n8655;
  assign n8659 = LWORD_REG_0_ & n8658;
  assign n8660 = DATAO_REG_0_ & n8655;
  assign n8661 = ~n8657 & ~n8659;
  assign n1710 = n8660 | ~n8661;
  assign n8663 = EAX_REG_1_ & n8656;
  assign n8664 = LWORD_REG_1_ & n8658;
  assign n8665 = DATAO_REG_1_ & n8655;
  assign n8666 = ~n8663 & ~n8664;
  assign n1714 = n8665 | ~n8666;
  assign n8668 = EAX_REG_2_ & n8656;
  assign n8669 = LWORD_REG_2_ & n8658;
  assign n8670 = DATAO_REG_2_ & n8655;
  assign n8671 = ~n8668 & ~n8669;
  assign n1718 = n8670 | ~n8671;
  assign n8673 = EAX_REG_3_ & n8656;
  assign n8674 = LWORD_REG_3_ & n8658;
  assign n8675 = DATAO_REG_3_ & n8655;
  assign n8676 = ~n8673 & ~n8674;
  assign n1722 = n8675 | ~n8676;
  assign n8678 = EAX_REG_4_ & n8656;
  assign n8679 = LWORD_REG_4_ & n8658;
  assign n8680 = DATAO_REG_4_ & n8655;
  assign n8681 = ~n8678 & ~n8679;
  assign n1726 = n8680 | ~n8681;
  assign n8683 = EAX_REG_5_ & n8656;
  assign n8684 = LWORD_REG_5_ & n8658;
  assign n8685 = DATAO_REG_5_ & n8655;
  assign n8686 = ~n8683 & ~n8684;
  assign n1730 = n8685 | ~n8686;
  assign n8688 = EAX_REG_6_ & n8656;
  assign n8689 = LWORD_REG_6_ & n8658;
  assign n8690 = DATAO_REG_6_ & n8655;
  assign n8691 = ~n8688 & ~n8689;
  assign n1734 = n8690 | ~n8691;
  assign n8693 = EAX_REG_7_ & n8656;
  assign n8694 = LWORD_REG_7_ & n8658;
  assign n8695 = DATAO_REG_7_ & n8655;
  assign n8696 = ~n8693 & ~n8694;
  assign n1738 = n8695 | ~n8696;
  assign n8698 = EAX_REG_8_ & n8656;
  assign n8699 = LWORD_REG_8_ & n8658;
  assign n8700 = DATAO_REG_8_ & n8655;
  assign n8701 = ~n8698 & ~n8699;
  assign n1742 = n8700 | ~n8701;
  assign n8703 = EAX_REG_9_ & n8656;
  assign n8704 = LWORD_REG_9_ & n8658;
  assign n8705 = DATAO_REG_9_ & n8655;
  assign n8706 = ~n8703 & ~n8704;
  assign n1746 = n8705 | ~n8706;
  assign n8708 = EAX_REG_10_ & n8656;
  assign n8709 = LWORD_REG_10_ & n8658;
  assign n8710 = DATAO_REG_10_ & n8655;
  assign n8711 = ~n8708 & ~n8709;
  assign n1750 = n8710 | ~n8711;
  assign n8713 = EAX_REG_11_ & n8656;
  assign n8714 = LWORD_REG_11_ & n8658;
  assign n8715 = DATAO_REG_11_ & n8655;
  assign n8716 = ~n8713 & ~n8714;
  assign n1754 = n8715 | ~n8716;
  assign n8718 = EAX_REG_12_ & n8656;
  assign n8719 = LWORD_REG_12_ & n8658;
  assign n8720 = DATAO_REG_12_ & n8655;
  assign n8721 = ~n8718 & ~n8719;
  assign n1758 = n8720 | ~n8721;
  assign n8723 = EAX_REG_13_ & n8656;
  assign n8724 = LWORD_REG_13_ & n8658;
  assign n8725 = DATAO_REG_13_ & n8655;
  assign n8726 = ~n8723 & ~n8724;
  assign n1762 = n8725 | ~n8726;
  assign n8728 = EAX_REG_14_ & n8656;
  assign n8729 = LWORD_REG_14_ & n8658;
  assign n8730 = DATAO_REG_14_ & n8655;
  assign n8731 = ~n8728 & ~n8729;
  assign n1766 = n8730 | ~n8731;
  assign n8733 = EAX_REG_15_ & n8656;
  assign n8734 = LWORD_REG_15_ & n8658;
  assign n8735 = DATAO_REG_15_ & n8655;
  assign n8736 = ~n8733 & ~n8734;
  assign n1770 = n8735 | ~n8736;
  assign n8738 = UWORD_REG_0_ & n8658;
  assign n8739 = DATAO_REG_16_ & n8655;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~n1776 & n8656;
  assign n8742 = EAX_REG_16_ & n8741;
  assign n1774 = ~n8740 | n8742;
  assign n8744 = UWORD_REG_1_ & n8658;
  assign n8745 = DATAO_REG_17_ & n8655;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = EAX_REG_17_ & n8741;
  assign n1778 = ~n8746 | n8747;
  assign n8749 = UWORD_REG_2_ & n8658;
  assign n8750 = DATAO_REG_18_ & n8655;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = EAX_REG_18_ & n8741;
  assign n1782 = ~n8751 | n8752;
  assign n8754 = UWORD_REG_3_ & n8658;
  assign n8755 = DATAO_REG_19_ & n8655;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = EAX_REG_19_ & n8741;
  assign n1786 = ~n8756 | n8757;
  assign n8759 = UWORD_REG_4_ & n8658;
  assign n8760 = DATAO_REG_20_ & n8655;
  assign n8761 = ~n8759 & ~n8760;
  assign n8762 = EAX_REG_20_ & n8741;
  assign n1790 = ~n8761 | n8762;
  assign n8764 = UWORD_REG_5_ & n8658;
  assign n8765 = DATAO_REG_21_ & n8655;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = EAX_REG_21_ & n8741;
  assign n1794 = ~n8766 | n8767;
  assign n8769 = UWORD_REG_6_ & n8658;
  assign n8770 = DATAO_REG_22_ & n8655;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = EAX_REG_22_ & n8741;
  assign n1798 = ~n8771 | n8772;
  assign n8774 = UWORD_REG_7_ & n8658;
  assign n8775 = DATAO_REG_23_ & n8655;
  assign n8776 = ~n8774 & ~n8775;
  assign n8777 = EAX_REG_23_ & n8741;
  assign n1802 = ~n8776 | n8777;
  assign n8779 = UWORD_REG_8_ & n8658;
  assign n8780 = DATAO_REG_24_ & n8655;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = EAX_REG_24_ & n8741;
  assign n1806 = ~n8781 | n8782;
  assign n8784 = UWORD_REG_9_ & n8658;
  assign n8785 = DATAO_REG_25_ & n8655;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = EAX_REG_25_ & n8741;
  assign n1810 = ~n8786 | n8787;
  assign n8789 = UWORD_REG_10_ & n8658;
  assign n8790 = DATAO_REG_26_ & n8655;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = EAX_REG_26_ & n8741;
  assign n1814 = ~n8791 | n8792;
  assign n8794 = UWORD_REG_11_ & n8658;
  assign n8795 = DATAO_REG_27_ & n8655;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = EAX_REG_27_ & n8741;
  assign n1818 = ~n8796 | n8797;
  assign n8799 = UWORD_REG_12_ & n8658;
  assign n8800 = DATAO_REG_28_ & n8655;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = EAX_REG_28_ & n8741;
  assign n1822 = ~n8801 | n8802;
  assign n8804 = UWORD_REG_13_ & n8658;
  assign n8805 = DATAO_REG_29_ & n8655;
  assign n8806 = ~n8804 & ~n8805;
  assign n8807 = EAX_REG_29_ & n8741;
  assign n1826 = ~n8806 | n8807;
  assign n8809 = UWORD_REG_14_ & n8658;
  assign n8810 = DATAO_REG_30_ & n8655;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = EAX_REG_30_ & n8741;
  assign n1830 = ~n8811 | n8812;
  assign n1834 = DATAO_REG_31_ & n8655;
  assign n8815 = ~n1839 & n7373;
  assign n8816 = ~n2262 & n8815;
  assign n8817 = n2315 & n2415;
  assign n8818 = n2144 & n8817;
  assign n8819 = ~n8816 & ~n8818;
  assign n8820 = n2282 & n2331;
  assign n8821 = ~n2262 & n8820;
  assign n8822 = n2108_1 & n2144;
  assign n8823 = n2272 & n8822;
  assign n8824 = ~n8821 & ~n8823;
  assign n8825 = ~READY_N & ~n8824;
  assign n8826 = n8819 & ~n8825;
  assign n8827 = n2411 & ~n8826;
  assign n8828 = ~n1929 & ~n2395;
  assign n8829 = n8827 & ~n8828;
  assign n8830 = ~n6783 & n8829;
  assign n8831 = n8827 & n8828;
  assign n8832 = DATAI_0_ & n8831;
  assign n8833 = EAX_REG_0_ & ~n8827;
  assign n8834 = ~n8830 & ~n8832;
  assign n1838 = n8833 | ~n8834;
  assign n8836 = ~n6815 & n8829;
  assign n8837 = DATAI_1_ & n8831;
  assign n8838 = EAX_REG_1_ & ~n8827;
  assign n8839 = ~n8836 & ~n8837;
  assign n1843 = n8838 | ~n8839;
  assign n8841 = EAX_REG_2_ & ~n8827;
  assign n8842 = DATAI_2_ & n8831;
  assign n8843 = n6850 & n8829;
  assign n8844 = ~n8841 & ~n8842;
  assign n1848 = n8843 | ~n8844;
  assign n8846 = EAX_REG_3_ & ~n8827;
  assign n8847 = DATAI_3_ & n8831;
  assign n8848 = n6883 & n8829;
  assign n8849 = ~n8846 & ~n8847;
  assign n1853 = n8848 | ~n8849;
  assign n8851 = EAX_REG_4_ & ~n8827;
  assign n8852 = DATAI_4_ & n8831;
  assign n8853 = ~n6924 & n8829;
  assign n8854 = ~n8851 & ~n8852;
  assign n1858 = n8853 | ~n8854;
  assign n8856 = EAX_REG_5_ & ~n8827;
  assign n8857 = DATAI_5_ & n8831;
  assign n8858 = ~n6957 & n8829;
  assign n8859 = ~n8856 & ~n8857;
  assign n1863 = n8858 | ~n8859;
  assign n8861 = EAX_REG_6_ & ~n8827;
  assign n8862 = DATAI_6_ & n8831;
  assign n8863 = ~n6993 & n8829;
  assign n8864 = ~n8861 & ~n8862;
  assign n1868 = n8863 | ~n8864;
  assign n8866 = EAX_REG_7_ & ~n8827;
  assign n8867 = DATAI_7_ & n8831;
  assign n8868 = n7028 & n8829;
  assign n8869 = ~n8866 & ~n8867;
  assign n1873 = n8868 | ~n8869;
  assign n8871 = EAX_REG_8_ & ~n8827;
  assign n8872 = DATAI_8_ & n8831;
  assign n8873 = ~n7067 & n8829;
  assign n8874 = ~n8871 & ~n8872;
  assign n1878 = n8873 | ~n8874;
  assign n8876 = EAX_REG_9_ & ~n8827;
  assign n8877 = DATAI_9_ & n8831;
  assign n8878 = ~n7097 & n8829;
  assign n8879 = ~n8876 & ~n8877;
  assign n1883 = n8878 | ~n8879;
  assign n8881 = EAX_REG_10_ & ~n8827;
  assign n8882 = DATAI_10_ & n8831;
  assign n8883 = n7134 & n8829;
  assign n8884 = ~n8881 & ~n8882;
  assign n1888 = n8883 | ~n8884;
  assign n8886 = EAX_REG_11_ & ~n8827;
  assign n8887 = DATAI_11_ & n8831;
  assign n8888 = n7164 & n8829;
  assign n8889 = ~n8886 & ~n8887;
  assign n1893 = n8888 | ~n8889;
  assign n8891 = EAX_REG_12_ & ~n8827;
  assign n8892 = DATAI_12_ & n8831;
  assign n8893 = ~n7201 & n8829;
  assign n8894 = ~n8891 & ~n8892;
  assign n1898 = n8893 | ~n8894;
  assign n8896 = EAX_REG_13_ & ~n8827;
  assign n8897 = DATAI_13_ & n8831;
  assign n8898 = ~n7234 & n8829;
  assign n8899 = ~n8896 & ~n8897;
  assign n1903 = n8898 | ~n8899;
  assign n8901 = EAX_REG_14_ & ~n8827;
  assign n8902 = DATAI_14_ & n8831;
  assign n8903 = ~n7268 & n8829;
  assign n8904 = ~n8901 & ~n8902;
  assign n1908 = n8903 | ~n8904;
  assign n8906 = EAX_REG_15_ & ~n8827;
  assign n8907 = DATAI_15_ & n8831;
  assign n8908 = n7301 & n8829;
  assign n8909 = ~n8906 & ~n8907;
  assign n1913 = n8908 | ~n8909;
  assign n8911 = ~n1929 & n1994;
  assign n8912 = n8827 & n8911;
  assign n8913 = DATAI_0_ & n8912;
  assign n8914 = n2338_1 & n8827;
  assign n8915 = DATAI_16_ & n8914;
  assign n8916 = EAX_REG_16_ & ~n8827;
  assign n8917 = n7409 & n8829;
  assign n8918 = ~n8913 & ~n8915;
  assign n8919 = ~n8916 & n8918;
  assign n1918 = n8917 | ~n8919;
  assign n8921 = DATAI_1_ & n8912;
  assign n8922 = DATAI_17_ & n8914;
  assign n8923 = EAX_REG_17_ & ~n8827;
  assign n8924 = ~n7472 & n8829;
  assign n8925 = ~n8921 & ~n8922;
  assign n8926 = ~n8923 & n8925;
  assign n1923 = n8924 | ~n8926;
  assign n8928 = DATAI_2_ & n8912;
  assign n8929 = DATAI_18_ & n8914;
  assign n8930 = EAX_REG_18_ & ~n8827;
  assign n8931 = ~n7536 & n8829;
  assign n8932 = ~n8928 & ~n8929;
  assign n8933 = ~n8930 & n8932;
  assign n1928 = n8931 | ~n8933;
  assign n8935 = DATAI_3_ & n8912;
  assign n8936 = DATAI_19_ & n8914;
  assign n8937 = EAX_REG_19_ & ~n8827;
  assign n8938 = ~n7605 & n8829;
  assign n8939 = ~n8935 & ~n8936;
  assign n8940 = ~n8937 & n8939;
  assign n1933 = n8938 | ~n8940;
  assign n8942 = DATAI_4_ & n8912;
  assign n8943 = DATAI_20_ & n8914;
  assign n8944 = EAX_REG_20_ & ~n8827;
  assign n8945 = ~n7676 & n8829;
  assign n8946 = ~n8942 & ~n8943;
  assign n8947 = ~n8944 & n8946;
  assign n1938 = n8945 | ~n8947;
  assign n8949 = DATAI_5_ & n8912;
  assign n8950 = DATAI_21_ & n8914;
  assign n8951 = EAX_REG_21_ & ~n8827;
  assign n8952 = n7743 & n8829;
  assign n8953 = ~n8949 & ~n8950;
  assign n8954 = ~n8951 & n8953;
  assign n1943 = n8952 | ~n8954;
  assign n8956 = DATAI_6_ & n8912;
  assign n8957 = DATAI_22_ & n8914;
  assign n8958 = EAX_REG_22_ & ~n8827;
  assign n8959 = ~n7807 & n8829;
  assign n8960 = ~n8956 & ~n8957;
  assign n8961 = ~n8958 & n8960;
  assign n1948 = n8959 | ~n8961;
  assign n8963 = DATAI_7_ & n8912;
  assign n8964 = DATAI_23_ & n8914;
  assign n8965 = EAX_REG_23_ & ~n8827;
  assign n8966 = ~n7934 & n8829;
  assign n8967 = ~n8963 & ~n8964;
  assign n8968 = ~n8965 & n8967;
  assign n1953 = n8966 | ~n8968;
  assign n8970 = DATAI_8_ & n8912;
  assign n8971 = DATAI_24_ & n8914;
  assign n8972 = EAX_REG_24_ & ~n8827;
  assign n8973 = ~n8001 & n8829;
  assign n8974 = ~n8970 & ~n8971;
  assign n8975 = ~n8972 & n8974;
  assign n1958 = n8973 | ~n8975;
  assign n8977 = DATAI_9_ & n8912;
  assign n8978 = DATAI_25_ & n8914;
  assign n8979 = EAX_REG_25_ & ~n8827;
  assign n8980 = ~n8076 & n8829;
  assign n8981 = ~n8977 & ~n8978;
  assign n8982 = ~n8979 & n8981;
  assign n1963 = n8980 | ~n8982;
  assign n8984 = DATAI_10_ & n8912;
  assign n8985 = DATAI_26_ & n8914;
  assign n8986 = EAX_REG_26_ & ~n8827;
  assign n8987 = ~n8145 & n8829;
  assign n8988 = ~n8984 & ~n8985;
  assign n8989 = ~n8986 & n8988;
  assign n1968 = n8987 | ~n8989;
  assign n8991 = DATAI_11_ & n8912;
  assign n8992 = DATAI_27_ & n8914;
  assign n8993 = EAX_REG_27_ & ~n8827;
  assign n8994 = ~n8213 & n8829;
  assign n8995 = ~n8991 & ~n8992;
  assign n8996 = ~n8993 & n8995;
  assign n1973 = n8994 | ~n8996;
  assign n8998 = DATAI_12_ & n8912;
  assign n8999 = DATAI_28_ & n8914;
  assign n9000 = EAX_REG_28_ & ~n8827;
  assign n9001 = ~n8285 & n8829;
  assign n9002 = ~n8998 & ~n8999;
  assign n9003 = ~n9000 & n9002;
  assign n1978 = n9001 | ~n9003;
  assign n9005 = DATAI_13_ & n8912;
  assign n9006 = DATAI_29_ & n8914;
  assign n9007 = EAX_REG_29_ & ~n8827;
  assign n9008 = ~n8358 & n8829;
  assign n9009 = ~n9005 & ~n9006;
  assign n9010 = ~n9007 & n9009;
  assign n1983 = n9008 | ~n9010;
  assign n9012 = DATAI_14_ & n8912;
  assign n9013 = DATAI_30_ & n8914;
  assign n9014 = EAX_REG_30_ & ~n8827;
  assign n9015 = ~n8429 & n8829;
  assign n9016 = ~n9012 & ~n9013;
  assign n9017 = ~n9014 & n9016;
  assign n1988 = n9015 | ~n9017;
  assign n9019 = n1929 & ~n8465;
  assign n9020 = n8827 & n9019;
  assign n9021 = EAX_REG_31_ & ~n8827;
  assign n9022 = ~n9020 & ~n9021;
  assign n9023 = DATAI_31_ & n8914;
  assign n1993 = ~n9022 | n9023;
  assign n9025 = STATE2_REG_0_ & ~n1807;
  assign n9026 = n2100 & n9025;
  assign n9027 = n2402 & n9026;
  assign n9028 = n2415 & n9027;
  assign n9029 = n2262 & n7372;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = n2411 & ~n9030;
  assign n9032 = n1929 & n9031;
  assign n9033 = ~n4692 & n9032;
  assign n9034 = ~n1929 & n9031;
  assign n9035 = ~n6783 & n9034;
  assign n9036 = EBX_REG_0_ & ~n9031;
  assign n9037 = ~n9033 & ~n9035;
  assign n1998 = n9036 | ~n9037;
  assign n9039 = ~n4741 & n9032;
  assign n9040 = EBX_REG_1_ & ~n9031;
  assign n9041 = ~n6815 & n9034;
  assign n9042 = ~n9039 & ~n9040;
  assign n2003 = n9041 | ~n9042;
  assign n9044 = n4790 & n9032;
  assign n9045 = EBX_REG_2_ & ~n9031;
  assign n9046 = n6850 & n9034;
  assign n9047 = ~n9044 & ~n9045;
  assign n2008 = n9046 | ~n9047;
  assign n9049 = ~n4817 & n9032;
  assign n9050 = EBX_REG_3_ & ~n9031;
  assign n9051 = n6883 & n9034;
  assign n9052 = ~n9049 & ~n9050;
  assign n2013 = n9051 | ~n9052;
  assign n9054 = ~n4866 & n9032;
  assign n9055 = EBX_REG_4_ & ~n9031;
  assign n9056 = ~n6924 & n9034;
  assign n9057 = ~n9054 & ~n9055;
  assign n2018 = n9056 | ~n9057;
  assign n9059 = ~n4967 & n9032;
  assign n9060 = EBX_REG_5_ & ~n9031;
  assign n9061 = ~n6957 & n9034;
  assign n9062 = ~n9059 & ~n9060;
  assign n2023 = n9061 | ~n9062;
  assign n9064 = ~n5071 & n9032;
  assign n9065 = EBX_REG_6_ & ~n9031;
  assign n9066 = ~n6993 & n9034;
  assign n9067 = ~n9064 & ~n9065;
  assign n2028 = n9066 | ~n9067;
  assign n9069 = ~n5171 & n9032;
  assign n9070 = EBX_REG_7_ & ~n9031;
  assign n9071 = n7028 & n9034;
  assign n9072 = ~n9069 & ~n9070;
  assign n2033 = n9071 | ~n9072;
  assign n9074 = ~n5248 & n9032;
  assign n9075 = EBX_REG_8_ & ~n9031;
  assign n9076 = ~n7067 & n9034;
  assign n9077 = ~n9074 & ~n9075;
  assign n2038 = n9076 | ~n9077;
  assign n9079 = ~n5381 & n9032;
  assign n9080 = EBX_REG_9_ & ~n9031;
  assign n9081 = ~n7097 & n9034;
  assign n9082 = ~n9079 & ~n9080;
  assign n2043 = n9081 | ~n9082;
  assign n9084 = ~n5464 & n9032;
  assign n9085 = EBX_REG_10_ & ~n9031;
  assign n9086 = n7134 & n9034;
  assign n9087 = ~n9084 & ~n9085;
  assign n2048 = n9086 | ~n9087;
  assign n9089 = ~n5549 & n9032;
  assign n9090 = EBX_REG_11_ & ~n9031;
  assign n9091 = n7164 & n9034;
  assign n9092 = ~n9089 & ~n9090;
  assign n2053 = n9091 | ~n9092;
  assign n9094 = ~n5635 & n9032;
  assign n9095 = EBX_REG_12_ & ~n9031;
  assign n9096 = ~n7201 & n9034;
  assign n9097 = ~n9094 & ~n9095;
  assign n2058 = n9096 | ~n9097;
  assign n9099 = ~n5751 & n9032;
  assign n9100 = EBX_REG_13_ & ~n9031;
  assign n9101 = ~n7234 & n9034;
  assign n9102 = ~n9099 & ~n9100;
  assign n2063 = n9101 | ~n9102;
  assign n9104 = ~n5835 & n9032;
  assign n9105 = EBX_REG_14_ & ~n9031;
  assign n9106 = ~n7268 & n9034;
  assign n9107 = ~n9104 & ~n9105;
  assign n2068 = n9106 | ~n9107;
  assign n9109 = ~n5920 & n9032;
  assign n9110 = EBX_REG_15_ & ~n9031;
  assign n9111 = n7301 & n9034;
  assign n9112 = ~n9109 & ~n9110;
  assign n2073 = n9111 | ~n9112;
  assign n9114 = ~n6004 & n9032;
  assign n9115 = EBX_REG_16_ & ~n9031;
  assign n9116 = n7409 & n9034;
  assign n9117 = ~n9114 & ~n9115;
  assign n2078 = n9116 | ~n9117;
  assign n9119 = ~n6068 & n9032;
  assign n9120 = EBX_REG_17_ & ~n9031;
  assign n9121 = ~n7472 & n9034;
  assign n9122 = ~n9119 & ~n9120;
  assign n2083 = n9121 | ~n9122;
  assign n9124 = ~n6113 & n9032;
  assign n9125 = EBX_REG_18_ & ~n9031;
  assign n9126 = ~n7536 & n9034;
  assign n9127 = ~n9124 & ~n9125;
  assign n2088 = n9126 | ~n9127;
  assign n9129 = ~n6160 & n9032;
  assign n9130 = EBX_REG_19_ & ~n9031;
  assign n9131 = ~n7605 & n9034;
  assign n9132 = ~n9129 & ~n9130;
  assign n2093 = n9131 | ~n9132;
  assign n9134 = ~n6206 & n9032;
  assign n9135 = EBX_REG_20_ & ~n9031;
  assign n9136 = ~n7676 & n9034;
  assign n9137 = ~n9134 & ~n9135;
  assign n2098 = n9136 | ~n9137;
  assign n9139 = ~n6253 & n9032;
  assign n9140 = EBX_REG_21_ & ~n9031;
  assign n9141 = n7743 & n9034;
  assign n9142 = ~n9139 & ~n9140;
  assign n2103 = n9141 | ~n9142;
  assign n9144 = ~n6296 & n9032;
  assign n9145 = EBX_REG_22_ & ~n9031;
  assign n9146 = ~n7807 & n9034;
  assign n9147 = ~n9144 & ~n9145;
  assign n2108 = n9146 | ~n9147;
  assign n9149 = ~n6343 & n9032;
  assign n9150 = EBX_REG_23_ & ~n9031;
  assign n9151 = ~n7934 & n9034;
  assign n9152 = ~n9149 & ~n9150;
  assign n2113 = n9151 | ~n9152;
  assign n9154 = ~n6389 & n9032;
  assign n9155 = EBX_REG_24_ & ~n9031;
  assign n9156 = ~n8001 & n9034;
  assign n9157 = ~n9154 & ~n9155;
  assign n2118 = n9156 | ~n9157;
  assign n9159 = ~n6436 & n9032;
  assign n9160 = EBX_REG_25_ & ~n9031;
  assign n9161 = ~n8076 & n9034;
  assign n9162 = ~n9159 & ~n9160;
  assign n2123 = n9161 | ~n9162;
  assign n9164 = ~n6482 & n9032;
  assign n9165 = EBX_REG_26_ & ~n9031;
  assign n9166 = ~n8145 & n9034;
  assign n9167 = ~n9164 & ~n9165;
  assign n2128 = n9166 | ~n9167;
  assign n9169 = ~n6534 & n9032;
  assign n9170 = EBX_REG_27_ & ~n9031;
  assign n9171 = ~n8213 & n9034;
  assign n9172 = ~n9169 & ~n9170;
  assign n2133 = n9171 | ~n9172;
  assign n9174 = ~n6577 & n9032;
  assign n9175 = EBX_REG_28_ & ~n9031;
  assign n9176 = ~n8285 & n9034;
  assign n9177 = ~n9174 & ~n9175;
  assign n2138 = n9176 | ~n9177;
  assign n9179 = ~n6624 & n9032;
  assign n9180 = EBX_REG_29_ & ~n9031;
  assign n9181 = ~n8358 & n9034;
  assign n9182 = ~n9179 & ~n9180;
  assign n2143 = n9181 | ~n9182;
  assign n9184 = ~n6672 & n9032;
  assign n9185 = EBX_REG_30_ & ~n9031;
  assign n9186 = ~n8429 & n9034;
  assign n9187 = ~n9184 & ~n9185;
  assign n2148 = n9186 | ~n9187;
  assign n9189 = EBX_REG_31_ & ~n9031;
  assign n9190 = ~n6721 & n9032;
  assign n2153 = n9189 | n9190;
  assign n9192 = ~n2262 & n2552;
  assign n9193 = n2272 & n2336;
  assign n9194 = n2277 & n2674;
  assign n9195 = n2282 & n9194;
  assign n9196 = ~n9192 & ~n9193;
  assign n9197 = ~n9195 & n9196;
  assign n9198 = n2411 & ~n9197;
  assign n9199 = ~n2684 & ~n2712;
  assign n9200 = ~n4624 & n9199;
  assign n9201 = ~n9198 & n9200;
  assign n9202 = STATE2_REG_2_ & ~n9201;
  assign n9203 = n2152 & n9202;
  assign n9204 = n2293_1 & n9203;
  assign n9205 = n2654 & n9204;
  assign n9206 = n2149 & n9202;
  assign n9207 = n2654 & n9206;
  assign n9208 = ~n9205 & ~n9207;
  assign n9209 = REIP_REG_0_ & ~n9208;
  assign n9210 = ~n2654 & n9206;
  assign n9211 = EBX_REG_31_ & n9210;
  assign n9212 = ~n4692 & n9211;
  assign n9213 = ~EBX_REG_31_ & n9210;
  assign n9214 = ~n2293_1 & n9203;
  assign n9215 = ~n2654 & n9204;
  assign n9216 = ~n9213 & ~n9214;
  assign n9217 = ~n9215 & n9216;
  assign n9218 = EBX_REG_0_ & ~n9217;
  assign n9219 = STATE2_REG_3_ & ~n9201;
  assign n9220 = PHYADDRPOINTER_REG_0_ & n9219;
  assign n9221 = n1776 & n4657;
  assign n9222 = ~n9201 & n9221;
  assign n9223 = ~n2618 & n9222;
  assign n9224 = REIP_REG_0_ & n9201;
  assign n9225 = STATE2_REG_1_ & ~n9201;
  assign n9226 = n8439 & n9225;
  assign n9227 = PHYADDRPOINTER_REG_0_ & n9226;
  assign n9228 = STATE2_REG_1_ & ~n8439;
  assign n9229 = STATE2_REG_2_ & n1808;
  assign n9230 = ~n9228 & ~n9229;
  assign n9231 = ~n9201 & ~n9230;
  assign n9232 = ~n6783 & n9231;
  assign n9233 = ~n9220 & ~n9223;
  assign n9234 = ~n9224 & n9233;
  assign n9235 = ~n9227 & n9234;
  assign n9236 = ~n9232 & n9235;
  assign n9237 = ~n9209 & ~n9212;
  assign n9238 = ~n9218 & n9237;
  assign n2158 = ~n9236 | ~n9238;
  assign n9240 = ~REIP_REG_1_ & ~n9208;
  assign n9241 = ~n4741 & n9211;
  assign n9242 = EBX_REG_1_ & ~n9217;
  assign n9243 = PHYADDRPOINTER_REG_1_ & n9219;
  assign n9244 = ~n2633 & n9222;
  assign n9245 = REIP_REG_1_ & n9201;
  assign n9246 = ~PHYADDRPOINTER_REG_1_ & n9226;
  assign n9247 = ~n6815 & n9231;
  assign n9248 = ~n9243 & ~n9244;
  assign n9249 = ~n9245 & n9248;
  assign n9250 = ~n9246 & n9249;
  assign n9251 = ~n9247 & n9250;
  assign n9252 = ~n9240 & ~n9241;
  assign n9253 = ~n9242 & n9252;
  assign n2163 = ~n9251 | ~n9253;
  assign n9255 = REIP_REG_1_ & ~REIP_REG_2_;
  assign n9256 = ~REIP_REG_1_ & REIP_REG_2_;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = ~n9208 & ~n9257;
  assign n9259 = n4790 & n9211;
  assign n9260 = EBX_REG_2_ & ~n9217;
  assign n9261 = PHYADDRPOINTER_REG_2_ & n9219;
  assign n9262 = n2495 & n9222;
  assign n9263 = REIP_REG_2_ & n9201;
  assign n9264 = ~n6824 & n9226;
  assign n9265 = n6850 & n9231;
  assign n9266 = ~n9261 & ~n9262;
  assign n9267 = ~n9263 & n9266;
  assign n9268 = ~n9264 & n9267;
  assign n9269 = ~n9265 & n9268;
  assign n9270 = ~n9258 & ~n9259;
  assign n9271 = ~n9260 & n9270;
  assign n2168 = ~n9269 | ~n9271;
  assign n9273 = REIP_REG_1_ & REIP_REG_2_;
  assign n9274 = ~REIP_REG_3_ & n9273;
  assign n9275 = REIP_REG_3_ & ~n9273;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = ~n9208 & ~n9276;
  assign n9278 = ~n4817 & n9211;
  assign n9279 = EBX_REG_3_ & ~n9217;
  assign n9280 = PHYADDRPOINTER_REG_3_ & n9219;
  assign n9281 = ~n2580 & n9222;
  assign n9282 = REIP_REG_3_ & n9201;
  assign n9283 = ~n6860 & n9226;
  assign n9284 = n6883 & n9231;
  assign n9285 = ~n9280 & ~n9281;
  assign n9286 = ~n9282 & n9285;
  assign n9287 = ~n9283 & n9286;
  assign n9288 = ~n9284 & n9287;
  assign n9289 = ~n9277 & ~n9278;
  assign n9290 = ~n9279 & n9289;
  assign n2173 = ~n9288 | ~n9290;
  assign n9292 = ~n4866 & n9211;
  assign n9293 = ~STATE2_REG_1_ & n2724;
  assign n9294 = ~n9201 & n9293;
  assign n9295 = ~n9292 & ~n9294;
  assign n9296 = REIP_REG_3_ & n9273;
  assign n9297 = ~REIP_REG_4_ & n9296;
  assign n9298 = REIP_REG_4_ & ~n9296;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = ~n9208 & ~n9299;
  assign n9301 = PHYADDRPOINTER_REG_4_ & n9219;
  assign n9302 = ~n2570 & n9222;
  assign n9303 = REIP_REG_4_ & n9201;
  assign n9304 = ~n6894 & n9226;
  assign n9305 = ~n9301 & ~n9302;
  assign n9306 = ~n9303 & n9305;
  assign n9307 = ~n9304 & n9306;
  assign n9308 = ~n6924 & n9231;
  assign n9309 = EBX_REG_4_ & ~n9217;
  assign n9310 = n9295 & ~n9300;
  assign n9311 = n9307 & n9310;
  assign n9312 = ~n9308 & n9311;
  assign n2178 = n9309 | ~n9312;
  assign n9314 = ~n4967 & n9211;
  assign n9315 = ~n9294 & ~n9314;
  assign n9316 = REIP_REG_4_ & n9296;
  assign n9317 = ~REIP_REG_5_ & n9316;
  assign n9318 = REIP_REG_5_ & ~n9316;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = ~n9208 & ~n9319;
  assign n9321 = EBX_REG_5_ & ~n9217;
  assign n9322 = PHYADDRPOINTER_REG_5_ & n9219;
  assign n9323 = n6939 & n9222;
  assign n9324 = REIP_REG_5_ & n9201;
  assign n9325 = ~n6934 & n9226;
  assign n9326 = ~n6957 & n9231;
  assign n9327 = ~n9322 & ~n9323;
  assign n9328 = ~n9324 & n9327;
  assign n9329 = ~n9325 & n9328;
  assign n9330 = ~n9326 & n9329;
  assign n9331 = n9315 & ~n9320;
  assign n9332 = ~n9321 & n9331;
  assign n2183 = ~n9330 | ~n9332;
  assign n9334 = REIP_REG_6_ & n9201;
  assign n9335 = PHYADDRPOINTER_REG_6_ & n9219;
  assign n9336 = ~n6970 & n9226;
  assign n9337 = ~n9334 & ~n9335;
  assign n9338 = ~n9336 & n9337;
  assign n9339 = EBX_REG_6_ & ~n9217;
  assign n9340 = ~n5071 & n9211;
  assign n9341 = ~n9294 & ~n9340;
  assign n9342 = REIP_REG_5_ & n9316;
  assign n9343 = ~REIP_REG_6_ & n9342;
  assign n9344 = REIP_REG_6_ & ~n9342;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = ~n9208 & ~n9345;
  assign n9347 = ~n8439 & n9225;
  assign n9348 = ~n6993 & n9347;
  assign n9349 = n9338 & ~n9339;
  assign n9350 = n9341 & n9349;
  assign n9351 = ~n9346 & n9350;
  assign n2188 = n9348 | ~n9351;
  assign n9353 = REIP_REG_7_ & n9201;
  assign n9354 = PHYADDRPOINTER_REG_7_ & n9219;
  assign n9355 = ~n7003 & n9226;
  assign n9356 = ~n9353 & ~n9354;
  assign n9357 = ~n9355 & n9356;
  assign n9358 = EBX_REG_7_ & ~n9217;
  assign n9359 = ~n5171 & n9211;
  assign n9360 = ~n9294 & ~n9359;
  assign n9361 = REIP_REG_6_ & n9342;
  assign n9362 = ~REIP_REG_7_ & n9361;
  assign n9363 = REIP_REG_7_ & ~n9361;
  assign n9364 = ~n9362 & ~n9363;
  assign n9365 = ~n9208 & ~n9364;
  assign n9366 = n7028 & n9347;
  assign n9367 = n9357 & ~n9358;
  assign n9368 = n9360 & n9367;
  assign n9369 = ~n9365 & n9368;
  assign n2193 = n9366 | ~n9369;
  assign n9371 = REIP_REG_8_ & n9201;
  assign n9372 = PHYADDRPOINTER_REG_8_ & n9219;
  assign n9373 = ~n7039 & n9226;
  assign n9374 = ~n9371 & ~n9372;
  assign n9375 = ~n9373 & n9374;
  assign n9376 = EBX_REG_8_ & ~n9217;
  assign n9377 = ~n5248 & n9211;
  assign n9378 = ~n9294 & ~n9377;
  assign n9379 = REIP_REG_7_ & n9361;
  assign n9380 = ~REIP_REG_8_ & n9379;
  assign n9381 = REIP_REG_8_ & ~n9379;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = ~n9208 & ~n9382;
  assign n9384 = ~n7067 & n9347;
  assign n9385 = n9375 & ~n9376;
  assign n9386 = n9378 & n9385;
  assign n9387 = ~n9383 & n9386;
  assign n2198 = n9384 | ~n9387;
  assign n9389 = REIP_REG_9_ & n9201;
  assign n9390 = PHYADDRPOINTER_REG_9_ & n9219;
  assign n9391 = ~n7077 & n9226;
  assign n9392 = ~n9389 & ~n9390;
  assign n9393 = ~n9391 & n9392;
  assign n9394 = EBX_REG_9_ & ~n9217;
  assign n9395 = ~n5381 & n9211;
  assign n9396 = ~n9294 & ~n9395;
  assign n9397 = REIP_REG_8_ & n9379;
  assign n9398 = ~REIP_REG_9_ & n9397;
  assign n9399 = REIP_REG_9_ & ~n9397;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = ~n9208 & ~n9400;
  assign n9402 = ~n7097 & n9347;
  assign n9403 = n9393 & ~n9394;
  assign n9404 = n9396 & n9403;
  assign n9405 = ~n9401 & n9404;
  assign n2203 = n9402 | ~n9405;
  assign n9407 = REIP_REG_10_ & n9201;
  assign n9408 = PHYADDRPOINTER_REG_10_ & n9219;
  assign n9409 = ~n7108 & n9226;
  assign n9410 = ~n9407 & ~n9408;
  assign n9411 = ~n9409 & n9410;
  assign n9412 = EBX_REG_10_ & ~n9217;
  assign n9413 = ~n5464 & n9211;
  assign n9414 = ~n9294 & ~n9413;
  assign n9415 = REIP_REG_9_ & n9397;
  assign n9416 = ~REIP_REG_10_ & n9415;
  assign n9417 = REIP_REG_10_ & ~n9415;
  assign n9418 = ~n9416 & ~n9417;
  assign n9419 = ~n9208 & ~n9418;
  assign n9420 = n7134 & n9347;
  assign n9421 = n9411 & ~n9412;
  assign n9422 = n9414 & n9421;
  assign n9423 = ~n9419 & n9422;
  assign n2208 = n9420 | ~n9423;
  assign n9425 = REIP_REG_11_ & n9201;
  assign n9426 = PHYADDRPOINTER_REG_11_ & n9219;
  assign n9427 = ~n7144 & n9226;
  assign n9428 = ~n9425 & ~n9426;
  assign n9429 = ~n9427 & n9428;
  assign n9430 = EBX_REG_11_ & ~n9217;
  assign n9431 = ~n5549 & n9211;
  assign n9432 = ~n9294 & ~n9431;
  assign n9433 = REIP_REG_10_ & n9415;
  assign n9434 = ~REIP_REG_11_ & n9433;
  assign n9435 = REIP_REG_11_ & ~n9433;
  assign n9436 = ~n9434 & ~n9435;
  assign n9437 = ~n9208 & ~n9436;
  assign n9438 = n7164 & n9347;
  assign n9439 = n9429 & ~n9430;
  assign n9440 = n9432 & n9439;
  assign n9441 = ~n9437 & n9440;
  assign n2213 = n9438 | ~n9441;
  assign n9443 = REIP_REG_12_ & n9201;
  assign n9444 = PHYADDRPOINTER_REG_12_ & n9219;
  assign n9445 = ~n7175 & n9226;
  assign n9446 = ~n9443 & ~n9444;
  assign n9447 = ~n9445 & n9446;
  assign n9448 = EBX_REG_12_ & ~n9217;
  assign n9449 = ~n5635 & n9211;
  assign n9450 = ~n9294 & ~n9449;
  assign n9451 = REIP_REG_11_ & n9433;
  assign n9452 = ~REIP_REG_12_ & n9451;
  assign n9453 = REIP_REG_12_ & ~n9451;
  assign n9454 = ~n9452 & ~n9453;
  assign n9455 = ~n9208 & ~n9454;
  assign n9456 = ~n7201 & n9347;
  assign n9457 = n9447 & ~n9448;
  assign n9458 = n9450 & n9457;
  assign n9459 = ~n9455 & n9458;
  assign n2218 = n9456 | ~n9459;
  assign n9461 = REIP_REG_13_ & n9201;
  assign n9462 = PHYADDRPOINTER_REG_13_ & n9219;
  assign n9463 = ~n7211 & n9226;
  assign n9464 = ~n9461 & ~n9462;
  assign n9465 = ~n9463 & n9464;
  assign n9466 = EBX_REG_13_ & ~n9217;
  assign n9467 = ~n5751 & n9211;
  assign n9468 = ~n9294 & ~n9467;
  assign n9469 = REIP_REG_12_ & n9451;
  assign n9470 = ~REIP_REG_13_ & n9469;
  assign n9471 = REIP_REG_13_ & ~n9469;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = ~n9208 & ~n9472;
  assign n9474 = ~n7234 & n9347;
  assign n9475 = n9465 & ~n9466;
  assign n9476 = n9468 & n9475;
  assign n9477 = ~n9473 & n9476;
  assign n2223 = n9474 | ~n9477;
  assign n9479 = REIP_REG_14_ & n9201;
  assign n9480 = PHYADDRPOINTER_REG_14_ & n9219;
  assign n9481 = ~n7245 & n9226;
  assign n9482 = ~n9479 & ~n9480;
  assign n9483 = ~n9481 & n9482;
  assign n9484 = EBX_REG_14_ & ~n9217;
  assign n9485 = ~n5835 & n9211;
  assign n9486 = ~n9294 & ~n9485;
  assign n9487 = REIP_REG_13_ & n9469;
  assign n9488 = ~REIP_REG_14_ & n9487;
  assign n9489 = REIP_REG_14_ & ~n9487;
  assign n9490 = ~n9488 & ~n9489;
  assign n9491 = ~n9208 & ~n9490;
  assign n9492 = ~n7268 & n9347;
  assign n9493 = n9483 & ~n9484;
  assign n9494 = n9486 & n9493;
  assign n9495 = ~n9491 & n9494;
  assign n2228 = n9492 | ~n9495;
  assign n9497 = EBX_REG_15_ & ~n9217;
  assign n9498 = REIP_REG_14_ & n9487;
  assign n9499 = ~REIP_REG_15_ & n9498;
  assign n9500 = REIP_REG_15_ & ~n9498;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = ~n9208 & ~n9501;
  assign n9503 = REIP_REG_15_ & n9201;
  assign n9504 = PHYADDRPOINTER_REG_15_ & n9219;
  assign n9505 = ~n7278 & n9226;
  assign n9506 = ~n9503 & ~n9504;
  assign n9507 = ~n9505 & n9506;
  assign n9508 = ~n5920 & n9211;
  assign n9509 = ~n9294 & ~n9508;
  assign n9510 = n7301 & n9347;
  assign n9511 = ~n9497 & ~n9502;
  assign n9512 = n9507 & n9511;
  assign n9513 = n9509 & n9512;
  assign n2233 = n9510 | ~n9513;
  assign n9515 = EBX_REG_16_ & ~n9217;
  assign n9516 = REIP_REG_15_ & n9498;
  assign n9517 = ~REIP_REG_16_ & n9516;
  assign n9518 = REIP_REG_16_ & ~n9516;
  assign n9519 = ~n9517 & ~n9518;
  assign n9520 = ~n9208 & ~n9519;
  assign n9521 = REIP_REG_16_ & n9201;
  assign n9522 = PHYADDRPOINTER_REG_16_ & n9219;
  assign n9523 = ~n7312 & n9226;
  assign n9524 = ~n9521 & ~n9522;
  assign n9525 = ~n9523 & n9524;
  assign n9526 = ~n6004 & n9211;
  assign n9527 = ~n9294 & ~n9526;
  assign n9528 = n7409 & n9347;
  assign n9529 = ~n9515 & ~n9520;
  assign n9530 = n9525 & n9529;
  assign n9531 = n9527 & n9530;
  assign n2238 = n9528 | ~n9531;
  assign n9533 = REIP_REG_16_ & n9516;
  assign n9534 = ~REIP_REG_17_ & n9533;
  assign n9535 = REIP_REG_17_ & ~n9533;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = ~n9208 & ~n9536;
  assign n9538 = ~n9294 & ~n9537;
  assign n9539 = EBX_REG_17_ & ~n9217;
  assign n9540 = REIP_REG_17_ & n9201;
  assign n9541 = PHYADDRPOINTER_REG_17_ & n9219;
  assign n9542 = ~n7419 & n9226;
  assign n9543 = ~n9540 & ~n9541;
  assign n9544 = ~n9542 & n9543;
  assign n9545 = ~n6068 & n9211;
  assign n9546 = ~n7472 & n9347;
  assign n9547 = n9538 & ~n9539;
  assign n9548 = n9544 & n9547;
  assign n9549 = ~n9545 & n9548;
  assign n2243 = n9546 | ~n9549;
  assign n9551 = REIP_REG_17_ & n9533;
  assign n9552 = ~REIP_REG_18_ & n9551;
  assign n9553 = REIP_REG_18_ & ~n9551;
  assign n9554 = ~n9552 & ~n9553;
  assign n9555 = ~n9208 & ~n9554;
  assign n9556 = ~n9294 & ~n9555;
  assign n9557 = EBX_REG_18_ & ~n9217;
  assign n9558 = REIP_REG_18_ & n9201;
  assign n9559 = PHYADDRPOINTER_REG_18_ & n9219;
  assign n9560 = ~n7483 & n9226;
  assign n9561 = ~n9558 & ~n9559;
  assign n9562 = ~n9560 & n9561;
  assign n9563 = ~n6113 & n9211;
  assign n9564 = ~n7536 & n9347;
  assign n9565 = n9556 & ~n9557;
  assign n9566 = n9562 & n9565;
  assign n9567 = ~n9563 & n9566;
  assign n2248 = n9564 | ~n9567;
  assign n9569 = REIP_REG_18_ & n9551;
  assign n9570 = ~REIP_REG_19_ & n9569;
  assign n9571 = REIP_REG_19_ & ~n9569;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = ~n9208 & ~n9572;
  assign n9574 = ~n9294 & ~n9573;
  assign n9575 = EBX_REG_19_ & ~n9217;
  assign n9576 = REIP_REG_19_ & n9201;
  assign n9577 = PHYADDRPOINTER_REG_19_ & n9219;
  assign n9578 = ~n7546 & n9226;
  assign n9579 = ~n9576 & ~n9577;
  assign n9580 = ~n9578 & n9579;
  assign n9581 = ~n6160 & n9211;
  assign n9582 = ~n7605 & n9347;
  assign n9583 = n9574 & ~n9575;
  assign n9584 = n9580 & n9583;
  assign n9585 = ~n9581 & n9584;
  assign n2253 = n9582 | ~n9585;
  assign n9587 = EBX_REG_20_ & ~n9217;
  assign n9588 = PHYADDRPOINTER_REG_20_ & n9219;
  assign n9589 = REIP_REG_19_ & n9569;
  assign n9590 = ~REIP_REG_20_ & n9589;
  assign n9591 = REIP_REG_20_ & ~n9589;
  assign n9592 = ~n9590 & ~n9591;
  assign n9593 = ~n9208 & ~n9592;
  assign n9594 = ~n9588 & ~n9593;
  assign n9595 = ~n7616 & n9226;
  assign n9596 = REIP_REG_20_ & n9201;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = ~n6206 & n9211;
  assign n9599 = ~n7676 & n9347;
  assign n9600 = ~n9587 & n9594;
  assign n9601 = n9597 & n9600;
  assign n9602 = ~n9598 & n9601;
  assign n2258 = n9599 | ~n9602;
  assign n9604 = EBX_REG_21_ & ~n9217;
  assign n9605 = PHYADDRPOINTER_REG_21_ & n9219;
  assign n9606 = REIP_REG_20_ & n9589;
  assign n9607 = ~REIP_REG_21_ & n9606;
  assign n9608 = REIP_REG_21_ & ~n9606;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = ~n9208 & ~n9609;
  assign n9611 = ~n9605 & ~n9610;
  assign n9612 = ~n7686 & n9226;
  assign n9613 = REIP_REG_21_ & n9201;
  assign n9614 = ~n9612 & ~n9613;
  assign n9615 = ~n6253 & n9211;
  assign n9616 = n7743 & n9347;
  assign n9617 = ~n9604 & n9611;
  assign n9618 = n9614 & n9617;
  assign n9619 = ~n9615 & n9618;
  assign n2263 = n9616 | ~n9619;
  assign n9621 = EBX_REG_22_ & ~n9217;
  assign n9622 = PHYADDRPOINTER_REG_22_ & n9219;
  assign n9623 = REIP_REG_21_ & n9606;
  assign n9624 = ~REIP_REG_22_ & n9623;
  assign n9625 = REIP_REG_22_ & ~n9623;
  assign n9626 = ~n9624 & ~n9625;
  assign n9627 = ~n9208 & ~n9626;
  assign n9628 = ~n9622 & ~n9627;
  assign n9629 = ~n7754 & n9226;
  assign n9630 = REIP_REG_22_ & n9201;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = ~n6296 & n9211;
  assign n9633 = ~n7807 & n9347;
  assign n9634 = ~n9621 & n9628;
  assign n9635 = n9631 & n9634;
  assign n9636 = ~n9632 & n9635;
  assign n2268 = n9633 | ~n9636;
  assign n9638 = EBX_REG_23_ & ~n9217;
  assign n9639 = PHYADDRPOINTER_REG_23_ & n9219;
  assign n9640 = REIP_REG_22_ & n9623;
  assign n9641 = ~REIP_REG_23_ & n9640;
  assign n9642 = REIP_REG_23_ & ~n9640;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = ~n9208 & ~n9643;
  assign n9645 = ~n9639 & ~n9644;
  assign n9646 = ~n7817 & n9226;
  assign n9647 = REIP_REG_23_ & n9201;
  assign n9648 = ~n9646 & ~n9647;
  assign n9649 = ~n6343 & n9211;
  assign n9650 = ~n7934 & n9347;
  assign n9651 = ~n9638 & n9645;
  assign n9652 = n9648 & n9651;
  assign n9653 = ~n9649 & n9652;
  assign n2273 = n9650 | ~n9653;
  assign n9655 = EBX_REG_24_ & ~n9217;
  assign n9656 = PHYADDRPOINTER_REG_24_ & n9219;
  assign n9657 = REIP_REG_23_ & n9640;
  assign n9658 = ~REIP_REG_24_ & n9657;
  assign n9659 = REIP_REG_24_ & ~n9657;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = ~n9208 & ~n9660;
  assign n9662 = ~n9656 & ~n9661;
  assign n9663 = ~n7945 & n9226;
  assign n9664 = REIP_REG_24_ & n9201;
  assign n9665 = ~n9663 & ~n9664;
  assign n9666 = ~n6389 & n9211;
  assign n9667 = ~n8001 & n9347;
  assign n9668 = ~n9655 & n9662;
  assign n9669 = n9665 & n9668;
  assign n9670 = ~n9666 & n9669;
  assign n2278 = n9667 | ~n9670;
  assign n9672 = EBX_REG_25_ & ~n9217;
  assign n9673 = PHYADDRPOINTER_REG_25_ & n9219;
  assign n9674 = REIP_REG_24_ & n9657;
  assign n9675 = ~REIP_REG_25_ & n9674;
  assign n9676 = REIP_REG_25_ & ~n9674;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = ~n9208 & ~n9677;
  assign n9679 = ~n9673 & ~n9678;
  assign n9680 = ~n8011 & n9226;
  assign n9681 = REIP_REG_25_ & n9201;
  assign n9682 = ~n9680 & ~n9681;
  assign n9683 = ~n6436 & n9211;
  assign n9684 = ~n8076 & n9347;
  assign n9685 = ~n9672 & n9679;
  assign n9686 = n9682 & n9685;
  assign n9687 = ~n9683 & n9686;
  assign n2283 = n9684 | ~n9687;
  assign n9689 = EBX_REG_26_ & ~n9217;
  assign n9690 = PHYADDRPOINTER_REG_26_ & n9219;
  assign n9691 = REIP_REG_25_ & n9674;
  assign n9692 = ~REIP_REG_26_ & n9691;
  assign n9693 = REIP_REG_26_ & ~n9691;
  assign n9694 = ~n9692 & ~n9693;
  assign n9695 = ~n9208 & ~n9694;
  assign n9696 = ~n9690 & ~n9695;
  assign n9697 = ~n8087 & n9226;
  assign n9698 = REIP_REG_26_ & n9201;
  assign n9699 = ~n9697 & ~n9698;
  assign n9700 = ~n6482 & n9211;
  assign n9701 = ~n8145 & n9347;
  assign n9702 = ~n9689 & n9696;
  assign n9703 = n9699 & n9702;
  assign n9704 = ~n9700 & n9703;
  assign n2288 = n9701 | ~n9704;
  assign n9706 = EBX_REG_27_ & ~n9217;
  assign n9707 = PHYADDRPOINTER_REG_27_ & n9219;
  assign n9708 = REIP_REG_26_ & n9691;
  assign n9709 = ~REIP_REG_27_ & n9708;
  assign n9710 = REIP_REG_27_ & ~n9708;
  assign n9711 = ~n9709 & ~n9710;
  assign n9712 = ~n9208 & ~n9711;
  assign n9713 = ~n9707 & ~n9712;
  assign n9714 = ~n8155 & n9226;
  assign n9715 = REIP_REG_27_ & n9201;
  assign n9716 = ~n9714 & ~n9715;
  assign n9717 = ~n6534 & n9211;
  assign n9718 = ~n8213 & n9347;
  assign n9719 = ~n9706 & n9713;
  assign n9720 = n9716 & n9719;
  assign n9721 = ~n9717 & n9720;
  assign n2293 = n9718 | ~n9721;
  assign n9723 = EBX_REG_28_ & ~n9217;
  assign n9724 = PHYADDRPOINTER_REG_28_ & n9219;
  assign n9725 = REIP_REG_27_ & n9708;
  assign n9726 = ~REIP_REG_28_ & n9725;
  assign n9727 = REIP_REG_28_ & ~n9725;
  assign n9728 = ~n9726 & ~n9727;
  assign n9729 = ~n9208 & ~n9728;
  assign n9730 = ~n9724 & ~n9729;
  assign n9731 = ~n8223 & n9226;
  assign n9732 = REIP_REG_28_ & n9201;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = ~n6577 & n9211;
  assign n9735 = ~n8285 & n9347;
  assign n9736 = ~n9723 & n9730;
  assign n9737 = n9733 & n9736;
  assign n9738 = ~n9734 & n9737;
  assign n2298 = n9735 | ~n9738;
  assign n9740 = EBX_REG_29_ & ~n9217;
  assign n9741 = PHYADDRPOINTER_REG_29_ & n9219;
  assign n9742 = REIP_REG_28_ & n9725;
  assign n9743 = ~REIP_REG_29_ & n9742;
  assign n9744 = REIP_REG_29_ & ~n9742;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = ~n9208 & ~n9745;
  assign n9747 = ~n9741 & ~n9746;
  assign n9748 = ~n8295 & n9226;
  assign n9749 = REIP_REG_29_ & n9201;
  assign n9750 = ~n9748 & ~n9749;
  assign n9751 = ~n6624 & n9211;
  assign n9752 = ~n8358 & n9347;
  assign n9753 = ~n9740 & n9747;
  assign n9754 = n9750 & n9753;
  assign n9755 = ~n9751 & n9754;
  assign n2303 = n9752 | ~n9755;
  assign n9757 = EBX_REG_30_ & ~n9217;
  assign n9758 = PHYADDRPOINTER_REG_30_ & n9219;
  assign n9759 = REIP_REG_29_ & n9742;
  assign n9760 = ~REIP_REG_30_ & n9759;
  assign n9761 = REIP_REG_30_ & ~n9759;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = ~n9208 & ~n9762;
  assign n9764 = ~n9758 & ~n9763;
  assign n9765 = ~n8368 & n9226;
  assign n9766 = REIP_REG_30_ & n9201;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = ~n6672 & n9211;
  assign n9769 = ~n8429 & n9347;
  assign n9770 = ~n9757 & n9764;
  assign n9771 = n9767 & n9770;
  assign n9772 = ~n9768 & n9771;
  assign n2308 = n9769 | ~n9772;
  assign n9774 = EBX_REG_31_ & ~n9217;
  assign n9775 = PHYADDRPOINTER_REG_31_ & n9219;
  assign n9776 = REIP_REG_30_ & n9759;
  assign n9777 = ~REIP_REG_31_ & n9776;
  assign n9778 = REIP_REG_31_ & ~n9776;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = ~n9208 & ~n9779;
  assign n9781 = ~n9775 & ~n9780;
  assign n9782 = ~n8439 & n9226;
  assign n9783 = REIP_REG_31_ & n9201;
  assign n9784 = ~n9782 & ~n9783;
  assign n9785 = ~n6721 & n9211;
  assign n9786 = ~n8465 & n9347;
  assign n9787 = ~n9774 & n9781;
  assign n9788 = n9784 & n9787;
  assign n9789 = ~n9785 & n9788;
  assign n2313 = n9786 | ~n9789;
  assign n9791 = ~DATAWIDTH_REG_1_ & ~REIP_REG_1_;
  assign n9792 = ~DATAWIDTH_REG_30_ & ~DATAWIDTH_REG_31_;
  assign n9793 = DATAWIDTH_REG_0_ & DATAWIDTH_REG_1_;
  assign n9794 = ~DATAWIDTH_REG_28_ & ~DATAWIDTH_REG_29_;
  assign n9795 = ~DATAWIDTH_REG_26_ & ~DATAWIDTH_REG_27_;
  assign n9796 = n9792 & ~n9793;
  assign n9797 = n9794 & n9796;
  assign n9798 = n9795 & n9797;
  assign n9799 = ~DATAWIDTH_REG_22_ & ~DATAWIDTH_REG_23_;
  assign n9800 = ~DATAWIDTH_REG_24_ & n9799;
  assign n9801 = ~DATAWIDTH_REG_25_ & n9800;
  assign n9802 = ~DATAWIDTH_REG_18_ & ~DATAWIDTH_REG_19_;
  assign n9803 = ~DATAWIDTH_REG_20_ & n9802;
  assign n9804 = ~DATAWIDTH_REG_21_ & n9803;
  assign n9805 = n9801 & n9804;
  assign n9806 = ~DATAWIDTH_REG_14_ & ~DATAWIDTH_REG_15_;
  assign n9807 = ~DATAWIDTH_REG_16_ & n9806;
  assign n9808 = ~DATAWIDTH_REG_17_ & n9807;
  assign n9809 = ~DATAWIDTH_REG_10_ & ~DATAWIDTH_REG_11_;
  assign n9810 = ~DATAWIDTH_REG_12_ & n9809;
  assign n9811 = ~DATAWIDTH_REG_13_ & n9810;
  assign n9812 = n9808 & n9811;
  assign n9813 = ~DATAWIDTH_REG_6_ & ~DATAWIDTH_REG_7_;
  assign n9814 = ~DATAWIDTH_REG_8_ & n9813;
  assign n9815 = ~DATAWIDTH_REG_9_ & n9814;
  assign n9816 = ~DATAWIDTH_REG_2_ & ~DATAWIDTH_REG_3_;
  assign n9817 = ~DATAWIDTH_REG_4_ & n9816;
  assign n9818 = ~DATAWIDTH_REG_5_ & n9817;
  assign n9819 = n9815 & n9818;
  assign n9820 = n9798 & n9805;
  assign n9821 = n9812 & n9820;
  assign n9822 = n9819 & n9821;
  assign n9823 = n9791 & n9822;
  assign n9824 = BYTEENABLE_REG_3_ & ~n9822;
  assign n9825 = ~DATAWIDTH_REG_0_ & ~REIP_REG_0_;
  assign n9826 = ~DATAWIDTH_REG_1_ & n9825;
  assign n9827 = n9822 & n9826;
  assign n9828 = ~n9823 & ~n9824;
  assign n2318 = n9827 | ~n9828;
  assign n9830 = REIP_REG_0_ & REIP_REG_1_;
  assign n9831 = DATAWIDTH_REG_0_ & ~REIP_REG_0_;
  assign n9832 = ~DATAWIDTH_REG_0_ & ~DATAWIDTH_REG_1_;
  assign n9833 = ~n9831 & ~n9832;
  assign n9834 = ~REIP_REG_1_ & ~n9833;
  assign n9835 = ~n9830 & ~n9834;
  assign n9836 = n9822 & ~n9835;
  assign n9837 = BYTEENABLE_REG_2_ & ~n9822;
  assign n2323 = n9836 | n9837;
  assign n9839 = REIP_REG_1_ & n9822;
  assign n9840 = BYTEENABLE_REG_1_ & ~n9822;
  assign n9841 = ~n9839 & ~n9840;
  assign n2328 = n9827 | ~n9841;
  assign n9843 = ~REIP_REG_0_ & ~REIP_REG_1_;
  assign n9844 = n9822 & ~n9843;
  assign n9845 = BYTEENABLE_REG_0_ & ~n9822;
  assign n2333 = n9844 | n9845;
  assign n9847 = W_R_N_REG & ~n1454;
  assign n9848 = ~READREQUEST_REG & n1454;
  assign n2338 = n9847 | n9848;
  assign n9850 = ~n2297 & n2674;
  assign n9851 = FLUSH_REG & ~n9850;
  assign n2342 = n6747 | n9851;
  assign n9853 = n2276 & n9850;
  assign n9854 = MORE_REG & ~n9850;
  assign n2347 = n9853 | n9854;
  assign n9856 = BS16_N & ~n1670_1;
  assign n9857 = STATEBS16_REG & n1670_1;
  assign n9858 = ~STATE_REG_0_ & n1624;
  assign n9859 = ~n9856 & ~n9857;
  assign n2352 = n9858 | ~n9859;
  assign n9861 = n2145 & ~n2293_1;
  assign n9862 = ~n2689 & ~n9861;
  assign n9863 = ~READY_N & STATE2_REG_2_;
  assign n9864 = STATEBS16_REG & n2293_1;
  assign n9865 = n2152 & ~n9864;
  assign n9866 = n9863 & ~n9865;
  assign n9867 = STATE2_REG_0_ & ~n9866;
  assign n9868 = n9862 & ~n9867;
  assign n9869 = ~READY_N & ~STATE2_REG_0_;
  assign n9870 = n1707 & n9869;
  assign n9871 = ~n2406 & ~n2724;
  assign n9872 = ~n9870 & n9871;
  assign n9873 = ~n9198 & n9872;
  assign n9874 = ~n9868 & ~n9873;
  assign n9875 = REQUESTPENDING_REG & n9873;
  assign n2357 = n9874 | n9875;
  assign n9877 = D_C_N_REG & ~n1454;
  assign n9878 = ~CODEFETCH_REG & n1454;
  assign n9879 = ~n9877 & ~n9878;
  assign n2362 = n9858 | ~n9879;
  assign n9881 = MEMORYFETCH_REG & n1454;
  assign n9882 = M_IO_N_REG & ~n1454;
  assign n2366 = n9881 | n9882;
  assign n9884 = STATE2_REG_0_ & n9293;
  assign n9885 = n2290 & n2674;
  assign n9886 = CODEFETCH_REG & ~n9885;
  assign n2370 = n9884 | n9886;
  assign n9888 = STATE_REG_0_ & ADS_N_REG;
  assign n2375 = ~n1670_1 | n9888;
  assign n9890 = STATE2_REG_2_ & ~n1808;
  assign n9891 = ~n2265 & n9890;
  assign n9892 = ~n9198 & ~n9293;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = READREQUEST_REG & n9892;
  assign n2379 = n9893 | n9894;
  assign n9896 = n2143_1 & n2411;
  assign n9897 = n2286 & n9896;
  assign n9898 = ~n2288_1 & n9897;
  assign n9899 = MEMORYFETCH_REG & ~n9898;
  assign n9900 = ~n9293 & ~n9899;
  assign n2384 = n9195 | ~n9900;
  always @ (posedge clock) begin
    BE_N_REG_3_ <= n214;
    BE_N_REG_2_ <= n218;
    BE_N_REG_1_ <= n222;
    BE_N_REG_0_ <= n226;
    ADDRESS_REG_29_ <= n230;
    ADDRESS_REG_28_ <= n234;
    ADDRESS_REG_27_ <= n238;
    ADDRESS_REG_26_ <= n242;
    ADDRESS_REG_25_ <= n246;
    ADDRESS_REG_24_ <= n250;
    ADDRESS_REG_23_ <= n254;
    ADDRESS_REG_22_ <= n258;
    ADDRESS_REG_21_ <= n262;
    ADDRESS_REG_20_ <= n266;
    ADDRESS_REG_19_ <= n270;
    ADDRESS_REG_18_ <= n274;
    ADDRESS_REG_17_ <= n278;
    ADDRESS_REG_16_ <= n282;
    ADDRESS_REG_15_ <= n286;
    ADDRESS_REG_14_ <= n290;
    ADDRESS_REG_13_ <= n294;
    ADDRESS_REG_12_ <= n298;
    ADDRESS_REG_11_ <= n302;
    ADDRESS_REG_10_ <= n306;
    ADDRESS_REG_9_ <= n310;
    ADDRESS_REG_8_ <= n314;
    ADDRESS_REG_7_ <= n318;
    ADDRESS_REG_6_ <= n322;
    ADDRESS_REG_5_ <= n326;
    ADDRESS_REG_4_ <= n330;
    ADDRESS_REG_3_ <= n334;
    ADDRESS_REG_2_ <= n338;
    ADDRESS_REG_1_ <= n342;
    ADDRESS_REG_0_ <= n346;
    STATE_REG_2_ <= n350;
    STATE_REG_1_ <= n355;
    STATE_REG_0_ <= n360;
    DATAWIDTH_REG_0_ <= n365;
    DATAWIDTH_REG_1_ <= n370;
    DATAWIDTH_REG_2_ <= n375;
    DATAWIDTH_REG_3_ <= n380;
    DATAWIDTH_REG_4_ <= n385;
    DATAWIDTH_REG_5_ <= n390;
    DATAWIDTH_REG_6_ <= n395;
    DATAWIDTH_REG_7_ <= n400;
    DATAWIDTH_REG_8_ <= n405;
    DATAWIDTH_REG_9_ <= n410;
    DATAWIDTH_REG_10_ <= n415;
    DATAWIDTH_REG_11_ <= n420;
    DATAWIDTH_REG_12_ <= n425;
    DATAWIDTH_REG_13_ <= n430;
    DATAWIDTH_REG_14_ <= n435;
    DATAWIDTH_REG_15_ <= n440;
    DATAWIDTH_REG_16_ <= n445;
    DATAWIDTH_REG_17_ <= n450;
    DATAWIDTH_REG_18_ <= n455;
    DATAWIDTH_REG_19_ <= n460;
    DATAWIDTH_REG_20_ <= n465;
    DATAWIDTH_REG_21_ <= n470;
    DATAWIDTH_REG_22_ <= n475;
    DATAWIDTH_REG_23_ <= n480;
    DATAWIDTH_REG_24_ <= n485;
    DATAWIDTH_REG_25_ <= n490;
    DATAWIDTH_REG_26_ <= n495;
    DATAWIDTH_REG_27_ <= n500;
    DATAWIDTH_REG_28_ <= n505;
    DATAWIDTH_REG_29_ <= n510;
    DATAWIDTH_REG_30_ <= n515;
    DATAWIDTH_REG_31_ <= n520;
    STATE2_REG_3_ <= n525;
    STATE2_REG_2_ <= n530;
    STATE2_REG_1_ <= n535;
    STATE2_REG_0_ <= n540;
    INSTQUEUE_REG_15__7_ <= n545;
    INSTQUEUE_REG_15__6_ <= n550;
    INSTQUEUE_REG_15__5_ <= n555;
    INSTQUEUE_REG_15__4_ <= n560;
    INSTQUEUE_REG_15__3_ <= n565;
    INSTQUEUE_REG_15__2_ <= n570;
    INSTQUEUE_REG_15__1_ <= n575;
    INSTQUEUE_REG_15__0_ <= n580;
    INSTQUEUE_REG_14__7_ <= n585;
    INSTQUEUE_REG_14__6_ <= n590;
    INSTQUEUE_REG_14__5_ <= n595;
    INSTQUEUE_REG_14__4_ <= n600;
    INSTQUEUE_REG_14__3_ <= n605;
    INSTQUEUE_REG_14__2_ <= n610;
    INSTQUEUE_REG_14__1_ <= n615;
    INSTQUEUE_REG_14__0_ <= n620;
    INSTQUEUE_REG_13__7_ <= n625;
    INSTQUEUE_REG_13__6_ <= n630;
    INSTQUEUE_REG_13__5_ <= n635;
    INSTQUEUE_REG_13__4_ <= n640;
    INSTQUEUE_REG_13__3_ <= n645;
    INSTQUEUE_REG_13__2_ <= n650;
    INSTQUEUE_REG_13__1_ <= n655;
    INSTQUEUE_REG_13__0_ <= n660;
    INSTQUEUE_REG_12__7_ <= n665;
    INSTQUEUE_REG_12__6_ <= n670;
    INSTQUEUE_REG_12__5_ <= n675;
    INSTQUEUE_REG_12__4_ <= n680;
    INSTQUEUE_REG_12__3_ <= n685;
    INSTQUEUE_REG_12__2_ <= n690;
    INSTQUEUE_REG_12__1_ <= n695;
    INSTQUEUE_REG_12__0_ <= n700;
    INSTQUEUE_REG_11__7_ <= n705;
    INSTQUEUE_REG_11__6_ <= n710;
    INSTQUEUE_REG_11__5_ <= n715;
    INSTQUEUE_REG_11__4_ <= n720;
    INSTQUEUE_REG_11__3_ <= n725;
    INSTQUEUE_REG_11__2_ <= n730;
    INSTQUEUE_REG_11__1_ <= n735;
    INSTQUEUE_REG_11__0_ <= n740;
    INSTQUEUE_REG_10__7_ <= n745;
    INSTQUEUE_REG_10__6_ <= n750;
    INSTQUEUE_REG_10__5_ <= n755;
    INSTQUEUE_REG_10__4_ <= n760;
    INSTQUEUE_REG_10__3_ <= n765;
    INSTQUEUE_REG_10__2_ <= n770;
    INSTQUEUE_REG_10__1_ <= n775;
    INSTQUEUE_REG_10__0_ <= n780;
    INSTQUEUE_REG_9__7_ <= n785;
    INSTQUEUE_REG_9__6_ <= n790;
    INSTQUEUE_REG_9__5_ <= n795;
    INSTQUEUE_REG_9__4_ <= n800;
    INSTQUEUE_REG_9__3_ <= n805;
    INSTQUEUE_REG_9__2_ <= n810;
    INSTQUEUE_REG_9__1_ <= n815;
    INSTQUEUE_REG_9__0_ <= n820;
    INSTQUEUE_REG_8__7_ <= n825;
    INSTQUEUE_REG_8__6_ <= n830;
    INSTQUEUE_REG_8__5_ <= n835;
    INSTQUEUE_REG_8__4_ <= n840;
    INSTQUEUE_REG_8__3_ <= n845;
    INSTQUEUE_REG_8__2_ <= n850;
    INSTQUEUE_REG_8__1_ <= n855;
    INSTQUEUE_REG_8__0_ <= n860;
    INSTQUEUE_REG_7__7_ <= n865;
    INSTQUEUE_REG_7__6_ <= n870;
    INSTQUEUE_REG_7__5_ <= n875;
    INSTQUEUE_REG_7__4_ <= n880;
    INSTQUEUE_REG_7__3_ <= n885;
    INSTQUEUE_REG_7__2_ <= n890;
    INSTQUEUE_REG_7__1_ <= n895;
    INSTQUEUE_REG_7__0_ <= n900;
    INSTQUEUE_REG_6__7_ <= n905;
    INSTQUEUE_REG_6__6_ <= n910;
    INSTQUEUE_REG_6__5_ <= n915;
    INSTQUEUE_REG_6__4_ <= n920;
    INSTQUEUE_REG_6__3_ <= n925;
    INSTQUEUE_REG_6__2_ <= n930;
    INSTQUEUE_REG_6__1_ <= n935;
    INSTQUEUE_REG_6__0_ <= n940;
    INSTQUEUE_REG_5__7_ <= n945;
    INSTQUEUE_REG_5__6_ <= n950;
    INSTQUEUE_REG_5__5_ <= n955;
    INSTQUEUE_REG_5__4_ <= n960;
    INSTQUEUE_REG_5__3_ <= n965;
    INSTQUEUE_REG_5__2_ <= n970;
    INSTQUEUE_REG_5__1_ <= n975;
    INSTQUEUE_REG_5__0_ <= n980;
    INSTQUEUE_REG_4__7_ <= n985;
    INSTQUEUE_REG_4__6_ <= n990;
    INSTQUEUE_REG_4__5_ <= n995;
    INSTQUEUE_REG_4__4_ <= n1000;
    INSTQUEUE_REG_4__3_ <= n1005;
    INSTQUEUE_REG_4__2_ <= n1010;
    INSTQUEUE_REG_4__1_ <= n1015;
    INSTQUEUE_REG_4__0_ <= n1020;
    INSTQUEUE_REG_3__7_ <= n1025;
    INSTQUEUE_REG_3__6_ <= n1030;
    INSTQUEUE_REG_3__5_ <= n1035;
    INSTQUEUE_REG_3__4_ <= n1040;
    INSTQUEUE_REG_3__3_ <= n1045;
    INSTQUEUE_REG_3__2_ <= n1050;
    INSTQUEUE_REG_3__1_ <= n1055;
    INSTQUEUE_REG_3__0_ <= n1060;
    INSTQUEUE_REG_2__7_ <= n1065;
    INSTQUEUE_REG_2__6_ <= n1070;
    INSTQUEUE_REG_2__5_ <= n1075;
    INSTQUEUE_REG_2__4_ <= n1080;
    INSTQUEUE_REG_2__3_ <= n1085;
    INSTQUEUE_REG_2__2_ <= n1090;
    INSTQUEUE_REG_2__1_ <= n1095;
    INSTQUEUE_REG_2__0_ <= n1100;
    INSTQUEUE_REG_1__7_ <= n1105;
    INSTQUEUE_REG_1__6_ <= n1110;
    INSTQUEUE_REG_1__5_ <= n1115;
    INSTQUEUE_REG_1__4_ <= n1120;
    INSTQUEUE_REG_1__3_ <= n1125;
    INSTQUEUE_REG_1__2_ <= n1130;
    INSTQUEUE_REG_1__1_ <= n1135;
    INSTQUEUE_REG_1__0_ <= n1140;
    INSTQUEUE_REG_0__7_ <= n1145;
    INSTQUEUE_REG_0__6_ <= n1150;
    INSTQUEUE_REG_0__5_ <= n1155;
    INSTQUEUE_REG_0__4_ <= n1160;
    INSTQUEUE_REG_0__3_ <= n1165;
    INSTQUEUE_REG_0__2_ <= n1170;
    INSTQUEUE_REG_0__1_ <= n1175;
    INSTQUEUE_REG_0__0_ <= n1180;
    INSTQUEUERD_ADDR_REG_4_ <= n1185;
    INSTQUEUERD_ADDR_REG_3_ <= n1190;
    INSTQUEUERD_ADDR_REG_2_ <= n1195;
    INSTQUEUERD_ADDR_REG_1_ <= n1200;
    INSTQUEUERD_ADDR_REG_0_ <= n1205;
    INSTQUEUEWR_ADDR_REG_4_ <= n1210;
    INSTQUEUEWR_ADDR_REG_3_ <= n1215;
    INSTQUEUEWR_ADDR_REG_2_ <= n1220;
    INSTQUEUEWR_ADDR_REG_1_ <= n1225;
    INSTQUEUEWR_ADDR_REG_0_ <= n1230;
    INSTADDRPOINTER_REG_0_ <= n1235;
    INSTADDRPOINTER_REG_1_ <= n1240;
    INSTADDRPOINTER_REG_2_ <= n1245;
    INSTADDRPOINTER_REG_3_ <= n1250;
    INSTADDRPOINTER_REG_4_ <= n1255;
    INSTADDRPOINTER_REG_5_ <= n1260;
    INSTADDRPOINTER_REG_6_ <= n1265;
    INSTADDRPOINTER_REG_7_ <= n1270;
    INSTADDRPOINTER_REG_8_ <= n1275;
    INSTADDRPOINTER_REG_9_ <= n1280;
    INSTADDRPOINTER_REG_10_ <= n1285;
    INSTADDRPOINTER_REG_11_ <= n1290;
    INSTADDRPOINTER_REG_12_ <= n1295;
    INSTADDRPOINTER_REG_13_ <= n1300;
    INSTADDRPOINTER_REG_14_ <= n1305;
    INSTADDRPOINTER_REG_15_ <= n1310;
    INSTADDRPOINTER_REG_16_ <= n1315;
    INSTADDRPOINTER_REG_17_ <= n1320;
    INSTADDRPOINTER_REG_18_ <= n1325;
    INSTADDRPOINTER_REG_19_ <= n1330;
    INSTADDRPOINTER_REG_20_ <= n1335;
    INSTADDRPOINTER_REG_21_ <= n1340;
    INSTADDRPOINTER_REG_22_ <= n1345;
    INSTADDRPOINTER_REG_23_ <= n1350;
    INSTADDRPOINTER_REG_24_ <= n1355;
    INSTADDRPOINTER_REG_25_ <= n1360;
    INSTADDRPOINTER_REG_26_ <= n1365;
    INSTADDRPOINTER_REG_27_ <= n1370;
    INSTADDRPOINTER_REG_28_ <= n1375;
    INSTADDRPOINTER_REG_29_ <= n1380;
    INSTADDRPOINTER_REG_30_ <= n1385;
    INSTADDRPOINTER_REG_31_ <= n1390;
    PHYADDRPOINTER_REG_0_ <= n1395;
    PHYADDRPOINTER_REG_1_ <= n1400;
    PHYADDRPOINTER_REG_2_ <= n1405;
    PHYADDRPOINTER_REG_3_ <= n1410;
    PHYADDRPOINTER_REG_4_ <= n1415;
    PHYADDRPOINTER_REG_5_ <= n1420;
    PHYADDRPOINTER_REG_6_ <= n1425;
    PHYADDRPOINTER_REG_7_ <= n1430;
    PHYADDRPOINTER_REG_8_ <= n1435;
    PHYADDRPOINTER_REG_9_ <= n1440;
    PHYADDRPOINTER_REG_10_ <= n1445;
    PHYADDRPOINTER_REG_11_ <= n1450;
    PHYADDRPOINTER_REG_12_ <= n1455;
    PHYADDRPOINTER_REG_13_ <= n1460;
    PHYADDRPOINTER_REG_14_ <= n1465;
    PHYADDRPOINTER_REG_15_ <= n1470;
    PHYADDRPOINTER_REG_16_ <= n1475;
    PHYADDRPOINTER_REG_17_ <= n1480;
    PHYADDRPOINTER_REG_18_ <= n1485;
    PHYADDRPOINTER_REG_19_ <= n1490;
    PHYADDRPOINTER_REG_20_ <= n1495;
    PHYADDRPOINTER_REG_21_ <= n1500;
    PHYADDRPOINTER_REG_22_ <= n1505;
    PHYADDRPOINTER_REG_23_ <= n1510;
    PHYADDRPOINTER_REG_24_ <= n1515;
    PHYADDRPOINTER_REG_25_ <= n1520;
    PHYADDRPOINTER_REG_26_ <= n1525;
    PHYADDRPOINTER_REG_27_ <= n1530;
    PHYADDRPOINTER_REG_28_ <= n1535;
    PHYADDRPOINTER_REG_29_ <= n1540;
    PHYADDRPOINTER_REG_30_ <= n1545;
    PHYADDRPOINTER_REG_31_ <= n1550;
    LWORD_REG_15_ <= n1555;
    LWORD_REG_14_ <= n1560;
    LWORD_REG_13_ <= n1565;
    LWORD_REG_12_ <= n1570;
    LWORD_REG_11_ <= n1575;
    LWORD_REG_10_ <= n1580;
    LWORD_REG_9_ <= n1585;
    LWORD_REG_8_ <= n1590;
    LWORD_REG_7_ <= n1595;
    LWORD_REG_6_ <= n1600;
    LWORD_REG_5_ <= n1605;
    LWORD_REG_4_ <= n1610;
    LWORD_REG_3_ <= n1615;
    LWORD_REG_2_ <= n1620;
    LWORD_REG_1_ <= n1625;
    LWORD_REG_0_ <= n1630;
    UWORD_REG_14_ <= n1635;
    UWORD_REG_13_ <= n1640;
    UWORD_REG_12_ <= n1645;
    UWORD_REG_11_ <= n1650;
    UWORD_REG_10_ <= n1655;
    UWORD_REG_9_ <= n1660;
    UWORD_REG_8_ <= n1665;
    UWORD_REG_7_ <= n1670;
    UWORD_REG_6_ <= n1675;
    UWORD_REG_5_ <= n1680;
    UWORD_REG_4_ <= n1685;
    UWORD_REG_3_ <= n1690;
    UWORD_REG_2_ <= n1695;
    UWORD_REG_1_ <= n1700;
    UWORD_REG_0_ <= n1705;
    DATAO_REG_0_ <= n1710;
    DATAO_REG_1_ <= n1714;
    DATAO_REG_2_ <= n1718;
    DATAO_REG_3_ <= n1722;
    DATAO_REG_4_ <= n1726;
    DATAO_REG_5_ <= n1730;
    DATAO_REG_6_ <= n1734;
    DATAO_REG_7_ <= n1738;
    DATAO_REG_8_ <= n1742;
    DATAO_REG_9_ <= n1746;
    DATAO_REG_10_ <= n1750;
    DATAO_REG_11_ <= n1754;
    DATAO_REG_12_ <= n1758;
    DATAO_REG_13_ <= n1762;
    DATAO_REG_14_ <= n1766;
    DATAO_REG_15_ <= n1770;
    DATAO_REG_16_ <= n1774;
    DATAO_REG_17_ <= n1778;
    DATAO_REG_18_ <= n1782;
    DATAO_REG_19_ <= n1786;
    DATAO_REG_20_ <= n1790;
    DATAO_REG_21_ <= n1794;
    DATAO_REG_22_ <= n1798;
    DATAO_REG_23_ <= n1802;
    DATAO_REG_24_ <= n1806;
    DATAO_REG_25_ <= n1810;
    DATAO_REG_26_ <= n1814;
    DATAO_REG_27_ <= n1818;
    DATAO_REG_28_ <= n1822;
    DATAO_REG_29_ <= n1826;
    DATAO_REG_30_ <= n1830;
    DATAO_REG_31_ <= n1834;
    EAX_REG_0_ <= n1838;
    EAX_REG_1_ <= n1843;
    EAX_REG_2_ <= n1848;
    EAX_REG_3_ <= n1853;
    EAX_REG_4_ <= n1858;
    EAX_REG_5_ <= n1863;
    EAX_REG_6_ <= n1868;
    EAX_REG_7_ <= n1873;
    EAX_REG_8_ <= n1878;
    EAX_REG_9_ <= n1883;
    EAX_REG_10_ <= n1888;
    EAX_REG_11_ <= n1893;
    EAX_REG_12_ <= n1898;
    EAX_REG_13_ <= n1903;
    EAX_REG_14_ <= n1908;
    EAX_REG_15_ <= n1913;
    EAX_REG_16_ <= n1918;
    EAX_REG_17_ <= n1923;
    EAX_REG_18_ <= n1928;
    EAX_REG_19_ <= n1933;
    EAX_REG_20_ <= n1938;
    EAX_REG_21_ <= n1943;
    EAX_REG_22_ <= n1948;
    EAX_REG_23_ <= n1953;
    EAX_REG_24_ <= n1958;
    EAX_REG_25_ <= n1963;
    EAX_REG_26_ <= n1968;
    EAX_REG_27_ <= n1973;
    EAX_REG_28_ <= n1978;
    EAX_REG_29_ <= n1983;
    EAX_REG_30_ <= n1988;
    EAX_REG_31_ <= n1993;
    EBX_REG_0_ <= n1998;
    EBX_REG_1_ <= n2003;
    EBX_REG_2_ <= n2008;
    EBX_REG_3_ <= n2013;
    EBX_REG_4_ <= n2018;
    EBX_REG_5_ <= n2023;
    EBX_REG_6_ <= n2028;
    EBX_REG_7_ <= n2033;
    EBX_REG_8_ <= n2038;
    EBX_REG_9_ <= n2043;
    EBX_REG_10_ <= n2048;
    EBX_REG_11_ <= n2053;
    EBX_REG_12_ <= n2058;
    EBX_REG_13_ <= n2063;
    EBX_REG_14_ <= n2068;
    EBX_REG_15_ <= n2073;
    EBX_REG_16_ <= n2078;
    EBX_REG_17_ <= n2083;
    EBX_REG_18_ <= n2088;
    EBX_REG_19_ <= n2093;
    EBX_REG_20_ <= n2098;
    EBX_REG_21_ <= n2103;
    EBX_REG_22_ <= n2108;
    EBX_REG_23_ <= n2113;
    EBX_REG_24_ <= n2118;
    EBX_REG_25_ <= n2123;
    EBX_REG_26_ <= n2128;
    EBX_REG_27_ <= n2133;
    EBX_REG_28_ <= n2138;
    EBX_REG_29_ <= n2143;
    EBX_REG_30_ <= n2148;
    EBX_REG_31_ <= n2153;
    REIP_REG_0_ <= n2158;
    REIP_REG_1_ <= n2163;
    REIP_REG_2_ <= n2168;
    REIP_REG_3_ <= n2173;
    REIP_REG_4_ <= n2178;
    REIP_REG_5_ <= n2183;
    REIP_REG_6_ <= n2188;
    REIP_REG_7_ <= n2193;
    REIP_REG_8_ <= n2198;
    REIP_REG_9_ <= n2203;
    REIP_REG_10_ <= n2208;
    REIP_REG_11_ <= n2213;
    REIP_REG_12_ <= n2218;
    REIP_REG_13_ <= n2223;
    REIP_REG_14_ <= n2228;
    REIP_REG_15_ <= n2233;
    REIP_REG_16_ <= n2238;
    REIP_REG_17_ <= n2243;
    REIP_REG_18_ <= n2248;
    REIP_REG_19_ <= n2253;
    REIP_REG_20_ <= n2258;
    REIP_REG_21_ <= n2263;
    REIP_REG_22_ <= n2268;
    REIP_REG_23_ <= n2273;
    REIP_REG_24_ <= n2278;
    REIP_REG_25_ <= n2283;
    REIP_REG_26_ <= n2288;
    REIP_REG_27_ <= n2293;
    REIP_REG_28_ <= n2298;
    REIP_REG_29_ <= n2303;
    REIP_REG_30_ <= n2308;
    REIP_REG_31_ <= n2313;
    BYTEENABLE_REG_3_ <= n2318;
    BYTEENABLE_REG_2_ <= n2323;
    BYTEENABLE_REG_1_ <= n2328;
    BYTEENABLE_REG_0_ <= n2333;
    W_R_N_REG <= n2338;
    FLUSH_REG <= n2342;
    MORE_REG <= n2347;
    STATEBS16_REG <= n2352;
    REQUESTPENDING_REG <= n2357;
    D_C_N_REG <= n2362;
    M_IO_N_REG <= n2366;
    CODEFETCH_REG <= n2370;
    ADS_N_REG <= n2375;
    READREQUEST_REG <= n2379;
    MEMORYFETCH_REG <= n2384;
  end
endmodule


