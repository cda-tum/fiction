// Benchmark "top" written by ABC on Mon Nov 27 17:06:31 2023

module top ( 
    in00, in01, in02, in03, in04, in05, in06, in07, in08, in09, in010,
    in011, in012, in013, in014, in015, in016, in017, in018, in019, in020,
    in021, in022, in023, in024, in025, in026, in027, in028, in029, in030,
    in031, in032, in033, in034, in035, in036, in037, in038, in039, in040,
    in041, in042, in043, in044, in045, in046, in047, in048, in049, in050,
    in051, in052, in053, in054, in055, in056, in057, in058, in059, in060,
    in061, in062, in063, in064, in065, in066, in067, in068, in069, in070,
    in071, in072, in073, in074, in075, in076, in077, in078, in079, in080,
    in081, in082, in083, in084, in085, in086, in087, in088, in089, in090,
    in091, in092, in093, in094, in095, in096, in097, in098, in099, in0100,
    in0101, in0102, in0103, in0104, in0105, in0106, in0107, in0108, in0109,
    in0110, in0111, in0112, in0113, in0114, in0115, in0116, in0117, in0118,
    in0119, in0120, in0121, in0122, in0123, in0124, in0125, in0126, in0127,
    in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in110,
    in111, in112, in113, in114, in115, in116, in117, in118, in119, in120,
    in121, in122, in123, in124, in125, in126, in127, in128, in129, in130,
    in131, in132, in133, in134, in135, in136, in137, in138, in139, in140,
    in141, in142, in143, in144, in145, in146, in147, in148, in149, in150,
    in151, in152, in153, in154, in155, in156, in157, in158, in159, in160,
    in161, in162, in163, in164, in165, in166, in167, in168, in169, in170,
    in171, in172, in173, in174, in175, in176, in177, in178, in179, in180,
    in181, in182, in183, in184, in185, in186, in187, in188, in189, in190,
    in191, in192, in193, in194, in195, in196, in197, in198, in199, in1100,
    in1101, in1102, in1103, in1104, in1105, in1106, in1107, in1108, in1109,
    in1110, in1111, in1112, in1113, in1114, in1115, in1116, in1117, in1118,
    in1119, in1120, in1121, in1122, in1123, in1124, in1125, in1126, in1127,
    in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in210,
    in211, in212, in213, in214, in215, in216, in217, in218, in219, in220,
    in221, in222, in223, in224, in225, in226, in227, in228, in229, in230,
    in231, in232, in233, in234, in235, in236, in237, in238, in239, in240,
    in241, in242, in243, in244, in245, in246, in247, in248, in249, in250,
    in251, in252, in253, in254, in255, in256, in257, in258, in259, in260,
    in261, in262, in263, in264, in265, in266, in267, in268, in269, in270,
    in271, in272, in273, in274, in275, in276, in277, in278, in279, in280,
    in281, in282, in283, in284, in285, in286, in287, in288, in289, in290,
    in291, in292, in293, in294, in295, in296, in297, in298, in299, in2100,
    in2101, in2102, in2103, in2104, in2105, in2106, in2107, in2108, in2109,
    in2110, in2111, in2112, in2113, in2114, in2115, in2116, in2117, in2118,
    in2119, in2120, in2121, in2122, in2123, in2124, in2125, in2126, in2127,
    in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in310,
    in311, in312, in313, in314, in315, in316, in317, in318, in319, in320,
    in321, in322, in323, in324, in325, in326, in327, in328, in329, in330,
    in331, in332, in333, in334, in335, in336, in337, in338, in339, in340,
    in341, in342, in343, in344, in345, in346, in347, in348, in349, in350,
    in351, in352, in353, in354, in355, in356, in357, in358, in359, in360,
    in361, in362, in363, in364, in365, in366, in367, in368, in369, in370,
    in371, in372, in373, in374, in375, in376, in377, in378, in379, in380,
    in381, in382, in383, in384, in385, in386, in387, in388, in389, in390,
    in391, in392, in393, in394, in395, in396, in397, in398, in399, in3100,
    in3101, in3102, in3103, in3104, in3105, in3106, in3107, in3108, in3109,
    in3110, in3111, in3112, in3113, in3114, in3115, in3116, in3117, in3118,
    in3119, in3120, in3121, in3122, in3123, in3124, in3125, in3126, in3127,
    result0, result1, result2, result3, result4, result5, result6, result7,
    result8, result9, result10, result11, result12, result13, result14,
    result15, result16, result17, result18, result19, result20, result21,
    result22, result23, result24, result25, result26, result27, result28,
    result29, result30, result31, result32, result33, result34, result35,
    result36, result37, result38, result39, result40, result41, result42,
    result43, result44, result45, result46, result47, result48, result49,
    result50, result51, result52, result53, result54, result55, result56,
    result57, result58, result59, result60, result61, result62, result63,
    result64, result65, result66, result67, result68, result69, result70,
    result71, result72, result73, result74, result75, result76, result77,
    result78, result79, result80, result81, result82, result83, result84,
    result85, result86, result87, result88, result89, result90, result91,
    result92, result93, result94, result95, result96, result97, result98,
    result99, result100, result101, result102, result103, result104,
    result105, result106, result107, result108, result109, result110,
    result111, result112, result113, result114, result115, result116,
    result117, result118, result119, result120, result121, result122,
    result123, result124, result125, result126, result127, address0,
    address1  );
  input  in00, in01, in02, in03, in04, in05, in06, in07, in08, in09,
    in010, in011, in012, in013, in014, in015, in016, in017, in018, in019,
    in020, in021, in022, in023, in024, in025, in026, in027, in028, in029,
    in030, in031, in032, in033, in034, in035, in036, in037, in038, in039,
    in040, in041, in042, in043, in044, in045, in046, in047, in048, in049,
    in050, in051, in052, in053, in054, in055, in056, in057, in058, in059,
    in060, in061, in062, in063, in064, in065, in066, in067, in068, in069,
    in070, in071, in072, in073, in074, in075, in076, in077, in078, in079,
    in080, in081, in082, in083, in084, in085, in086, in087, in088, in089,
    in090, in091, in092, in093, in094, in095, in096, in097, in098, in099,
    in0100, in0101, in0102, in0103, in0104, in0105, in0106, in0107, in0108,
    in0109, in0110, in0111, in0112, in0113, in0114, in0115, in0116, in0117,
    in0118, in0119, in0120, in0121, in0122, in0123, in0124, in0125, in0126,
    in0127, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19,
    in110, in111, in112, in113, in114, in115, in116, in117, in118, in119,
    in120, in121, in122, in123, in124, in125, in126, in127, in128, in129,
    in130, in131, in132, in133, in134, in135, in136, in137, in138, in139,
    in140, in141, in142, in143, in144, in145, in146, in147, in148, in149,
    in150, in151, in152, in153, in154, in155, in156, in157, in158, in159,
    in160, in161, in162, in163, in164, in165, in166, in167, in168, in169,
    in170, in171, in172, in173, in174, in175, in176, in177, in178, in179,
    in180, in181, in182, in183, in184, in185, in186, in187, in188, in189,
    in190, in191, in192, in193, in194, in195, in196, in197, in198, in199,
    in1100, in1101, in1102, in1103, in1104, in1105, in1106, in1107, in1108,
    in1109, in1110, in1111, in1112, in1113, in1114, in1115, in1116, in1117,
    in1118, in1119, in1120, in1121, in1122, in1123, in1124, in1125, in1126,
    in1127, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29,
    in210, in211, in212, in213, in214, in215, in216, in217, in218, in219,
    in220, in221, in222, in223, in224, in225, in226, in227, in228, in229,
    in230, in231, in232, in233, in234, in235, in236, in237, in238, in239,
    in240, in241, in242, in243, in244, in245, in246, in247, in248, in249,
    in250, in251, in252, in253, in254, in255, in256, in257, in258, in259,
    in260, in261, in262, in263, in264, in265, in266, in267, in268, in269,
    in270, in271, in272, in273, in274, in275, in276, in277, in278, in279,
    in280, in281, in282, in283, in284, in285, in286, in287, in288, in289,
    in290, in291, in292, in293, in294, in295, in296, in297, in298, in299,
    in2100, in2101, in2102, in2103, in2104, in2105, in2106, in2107, in2108,
    in2109, in2110, in2111, in2112, in2113, in2114, in2115, in2116, in2117,
    in2118, in2119, in2120, in2121, in2122, in2123, in2124, in2125, in2126,
    in2127, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39,
    in310, in311, in312, in313, in314, in315, in316, in317, in318, in319,
    in320, in321, in322, in323, in324, in325, in326, in327, in328, in329,
    in330, in331, in332, in333, in334, in335, in336, in337, in338, in339,
    in340, in341, in342, in343, in344, in345, in346, in347, in348, in349,
    in350, in351, in352, in353, in354, in355, in356, in357, in358, in359,
    in360, in361, in362, in363, in364, in365, in366, in367, in368, in369,
    in370, in371, in372, in373, in374, in375, in376, in377, in378, in379,
    in380, in381, in382, in383, in384, in385, in386, in387, in388, in389,
    in390, in391, in392, in393, in394, in395, in396, in397, in398, in399,
    in3100, in3101, in3102, in3103, in3104, in3105, in3106, in3107, in3108,
    in3109, in3110, in3111, in3112, in3113, in3114, in3115, in3116, in3117,
    in3118, in3119, in3120, in3121, in3122, in3123, in3124, in3125, in3126,
    in3127;
  output result0, result1, result2, result3, result4, result5, result6,
    result7, result8, result9, result10, result11, result12, result13,
    result14, result15, result16, result17, result18, result19, result20,
    result21, result22, result23, result24, result25, result26, result27,
    result28, result29, result30, result31, result32, result33, result34,
    result35, result36, result37, result38, result39, result40, result41,
    result42, result43, result44, result45, result46, result47, result48,
    result49, result50, result51, result52, result53, result54, result55,
    result56, result57, result58, result59, result60, result61, result62,
    result63, result64, result65, result66, result67, result68, result69,
    result70, result71, result72, result73, result74, result75, result76,
    result77, result78, result79, result80, result81, result82, result83,
    result84, result85, result86, result87, result88, result89, result90,
    result91, result92, result93, result94, result95, result96, result97,
    result98, result99, result100, result101, result102, result103,
    result104, result105, result106, result107, result108, result109,
    result110, result111, result112, result113, result114, result115,
    result116, result117, result118, result119, result120, result121,
    result122, result123, result124, result125, result126, result127,
    address0, address1;
  wire new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1454, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2715,
    new_n2716, new_n2717, new_n2718, new_n2719, new_n2720, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2830, new_n2831, new_n2832, new_n2833, new_n2834, new_n2835,
    new_n2836, new_n2837, new_n2838, new_n2839, new_n2840, new_n2841,
    new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847,
    new_n2848, new_n2849, new_n2850, new_n2851, new_n2852, new_n2853,
    new_n2854, new_n2855, new_n2856, new_n2857, new_n2858, new_n2859,
    new_n2860, new_n2861, new_n2862, new_n2863, new_n2864, new_n2865,
    new_n2866, new_n2867, new_n2868, new_n2869, new_n2870, new_n2871,
    new_n2872, new_n2873, new_n2874, new_n2875, new_n2876, new_n2877,
    new_n2878, new_n2879, new_n2880, new_n2881, new_n2882, new_n2883,
    new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889,
    new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2896, new_n2897, new_n2898, new_n2899, new_n2900, new_n2901,
    new_n2902, new_n2903, new_n2904, new_n2905, new_n2906, new_n2907,
    new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913,
    new_n2914, new_n2915, new_n2916, new_n2917, new_n2918, new_n2919,
    new_n2920, new_n2921, new_n2922, new_n2923, new_n2924, new_n2925,
    new_n2926, new_n2927, new_n2928, new_n2929, new_n2930, new_n2931,
    new_n2932, new_n2933, new_n2934, new_n2935, new_n2936, new_n2937,
    new_n2938, new_n2939, new_n2940, new_n2941, new_n2942, new_n2943,
    new_n2944, new_n2945, new_n2946, new_n2947, new_n2948, new_n2949,
    new_n2950, new_n2951, new_n2952, new_n2953, new_n2954, new_n2955,
    new_n2956, new_n2957, new_n2958, new_n2959, new_n2960, new_n2961,
    new_n2962, new_n2963, new_n2964, new_n2965, new_n2966, new_n2967,
    new_n2968, new_n2969, new_n2970, new_n2971, new_n2972, new_n2973,
    new_n2974, new_n2975, new_n2977, new_n2978, new_n2980, new_n2981,
    new_n2983, new_n2984, new_n2986, new_n2987, new_n2989, new_n2990,
    new_n2992, new_n2993, new_n2995, new_n2996, new_n2998, new_n2999,
    new_n3001, new_n3002, new_n3004, new_n3005, new_n3007, new_n3008,
    new_n3010, new_n3011, new_n3013, new_n3014, new_n3016, new_n3017,
    new_n3019, new_n3020, new_n3022, new_n3023, new_n3025, new_n3026,
    new_n3028, new_n3029, new_n3031, new_n3032, new_n3034, new_n3035,
    new_n3037, new_n3038, new_n3040, new_n3041, new_n3043, new_n3044,
    new_n3046, new_n3047, new_n3049, new_n3050, new_n3052, new_n3053,
    new_n3055, new_n3056, new_n3058, new_n3059, new_n3061, new_n3062,
    new_n3064, new_n3065, new_n3067, new_n3068, new_n3070, new_n3071,
    new_n3073, new_n3074, new_n3076, new_n3077, new_n3079, new_n3080,
    new_n3082, new_n3083, new_n3085, new_n3086, new_n3088, new_n3089,
    new_n3091, new_n3092, new_n3094, new_n3095, new_n3097, new_n3098,
    new_n3100, new_n3101, new_n3103, new_n3104, new_n3106, new_n3107,
    new_n3109, new_n3110, new_n3112, new_n3113, new_n3115, new_n3116,
    new_n3118, new_n3119, new_n3121, new_n3122, new_n3124, new_n3125,
    new_n3127, new_n3128, new_n3130, new_n3131, new_n3133, new_n3134,
    new_n3136, new_n3137, new_n3139, new_n3140, new_n3142, new_n3143,
    new_n3145, new_n3146, new_n3148, new_n3149, new_n3151, new_n3152,
    new_n3154, new_n3155, new_n3157, new_n3158, new_n3160, new_n3161,
    new_n3163, new_n3164, new_n3166, new_n3167, new_n3169, new_n3170,
    new_n3172, new_n3173, new_n3175, new_n3176, new_n3178, new_n3179,
    new_n3181, new_n3182, new_n3184, new_n3185, new_n3187, new_n3188,
    new_n3190, new_n3191, new_n3193, new_n3194, new_n3196, new_n3197,
    new_n3199, new_n3200, new_n3202, new_n3203, new_n3205, new_n3206,
    new_n3208, new_n3209, new_n3211, new_n3212, new_n3214, new_n3215,
    new_n3217, new_n3218, new_n3220, new_n3221, new_n3223, new_n3224,
    new_n3226, new_n3227, new_n3229, new_n3230, new_n3232, new_n3233,
    new_n3235, new_n3236, new_n3238, new_n3239, new_n3241, new_n3242,
    new_n3244, new_n3245, new_n3247, new_n3248, new_n3250, new_n3251,
    new_n3253, new_n3254, new_n3256, new_n3257, new_n3259, new_n3260,
    new_n3262, new_n3263, new_n3265, new_n3266, new_n3268, new_n3269,
    new_n3271, new_n3272, new_n3274, new_n3275, new_n3277, new_n3278,
    new_n3280, new_n3281, new_n3283, new_n3284, new_n3286, new_n3287,
    new_n3289, new_n3290, new_n3292, new_n3293, new_n3295, new_n3296,
    new_n3298, new_n3299, new_n3301, new_n3302, new_n3304, new_n3305,
    new_n3307, new_n3308, new_n3310, new_n3311, new_n3313, new_n3314,
    new_n3316, new_n3317, new_n3319, new_n3320, new_n3322, new_n3323,
    new_n3325, new_n3326, new_n3328, new_n3329, new_n3331, new_n3332,
    new_n3334, new_n3335, new_n3337, new_n3338, new_n3340, new_n3341,
    new_n3343, new_n3344, new_n3346, new_n3347, new_n3349, new_n3350,
    new_n3352, new_n3353, new_n3355, new_n3356, new_n3359, new_n3360;
  assign new_n643 = in0126 & ~in1126;
  assign new_n644 = ~in0125 & in1125;
  assign new_n645 = ~in0126 & in1126;
  assign new_n646 = ~new_n644 & ~new_n645;
  assign new_n647 = in0125 & ~in1125;
  assign new_n648 = in0124 & ~in1124;
  assign new_n649 = ~new_n647 & ~new_n648;
  assign new_n650 = new_n646 & ~new_n649;
  assign new_n651 = ~in0124 & in1124;
  assign new_n652 = in0123 & ~in1123;
  assign new_n653 = in0122 & ~in1122;
  assign new_n654 = ~in0122 & in1122;
  assign new_n655 = ~in0121 & in1121;
  assign new_n656 = in0120 & ~in1120;
  assign new_n657 = in0121 & ~in1121;
  assign new_n658 = ~in0120 & in1120;
  assign new_n659 = in0119 & ~in1119;
  assign new_n660 = ~in0119 & in1119;
  assign new_n661 = in0118 & ~in1118;
  assign new_n662 = ~in0118 & in1118;
  assign new_n663 = in0117 & ~in1117;
  assign new_n664 = ~in0117 & in1117;
  assign new_n665 = in0116 & ~in1116;
  assign new_n666 = ~in0116 & in1116;
  assign new_n667 = in0115 & ~in1115;
  assign new_n668 = ~in0115 & in1115;
  assign new_n669 = in0114 & ~in1114;
  assign new_n670 = ~in0114 & in1114;
  assign new_n671 = in0113 & ~in1113;
  assign new_n672 = ~in0113 & in1113;
  assign new_n673 = in0112 & ~in1112;
  assign new_n674 = ~in0112 & in1112;
  assign new_n675 = in0111 & ~in1111;
  assign new_n676 = ~in0111 & in1111;
  assign new_n677 = in0110 & ~in1110;
  assign new_n678 = ~in0109 & in1109;
  assign new_n679 = ~in0110 & in1110;
  assign new_n680 = in0109 & ~in1109;
  assign new_n681 = ~in0108 & in1108;
  assign new_n682 = in0108 & ~in1108;
  assign new_n683 = ~in0107 & in1107;
  assign new_n684 = in0107 & ~in1107;
  assign new_n685 = ~in0106 & in1106;
  assign new_n686 = in0105 & ~in1105;
  assign new_n687 = in0106 & ~in1106;
  assign new_n688 = ~in0105 & in1105;
  assign new_n689 = in0104 & ~in1104;
  assign new_n690 = ~in0104 & in1104;
  assign new_n691 = in0103 & ~in1103;
  assign new_n692 = ~in0103 & in1103;
  assign new_n693 = in0102 & ~in1102;
  assign new_n694 = ~in0101 & in1101;
  assign new_n695 = ~in0102 & in1102;
  assign new_n696 = in0101 & ~in1101;
  assign new_n697 = ~in0100 & in1100;
  assign new_n698 = in0100 & ~in1100;
  assign new_n699 = ~in099 & in199;
  assign new_n700 = in099 & ~in199;
  assign new_n701 = ~in098 & in198;
  assign new_n702 = in097 & ~in197;
  assign new_n703 = in098 & ~in198;
  assign new_n704 = ~in097 & in197;
  assign new_n705 = in096 & ~in196;
  assign new_n706 = ~in096 & in196;
  assign new_n707 = in095 & ~in195;
  assign new_n708 = ~in095 & in195;
  assign new_n709 = in094 & ~in194;
  assign new_n710 = ~in093 & in193;
  assign new_n711 = ~in094 & in194;
  assign new_n712 = in093 & ~in193;
  assign new_n713 = ~in092 & in192;
  assign new_n714 = in092 & ~in192;
  assign new_n715 = ~in091 & in191;
  assign new_n716 = in091 & ~in191;
  assign new_n717 = ~in090 & in190;
  assign new_n718 = in089 & ~in189;
  assign new_n719 = in090 & ~in190;
  assign new_n720 = ~in089 & in189;
  assign new_n721 = in088 & ~in188;
  assign new_n722 = ~in088 & in188;
  assign new_n723 = in087 & ~in187;
  assign new_n724 = ~in087 & in187;
  assign new_n725 = in086 & ~in186;
  assign new_n726 = ~in085 & in185;
  assign new_n727 = ~in086 & in186;
  assign new_n728 = in085 & ~in185;
  assign new_n729 = ~in084 & in184;
  assign new_n730 = in084 & ~in184;
  assign new_n731 = ~in083 & in183;
  assign new_n732 = in083 & ~in183;
  assign new_n733 = ~in082 & in182;
  assign new_n734 = in077 & ~in177;
  assign new_n735 = in076 & ~in176;
  assign new_n736 = ~new_n734 & ~new_n735;
  assign new_n737 = ~in079 & in179;
  assign new_n738 = ~in078 & in178;
  assign new_n739 = ~in077 & in177;
  assign new_n740 = ~new_n737 & ~new_n738;
  assign new_n741 = ~new_n739 & new_n740;
  assign new_n742 = ~new_n736 & new_n741;
  assign new_n743 = in080 & ~in180;
  assign new_n744 = in079 & ~in179;
  assign new_n745 = in078 & ~in178;
  assign new_n746 = ~new_n737 & new_n745;
  assign new_n747 = ~in076 & in176;
  assign new_n748 = ~in073 & in173;
  assign new_n749 = in071 & ~in171;
  assign new_n750 = in070 & ~in170;
  assign new_n751 = ~in069 & in169;
  assign new_n752 = ~in070 & in170;
  assign new_n753 = in069 & ~in169;
  assign new_n754 = ~in068 & in168;
  assign new_n755 = in068 & ~in168;
  assign new_n756 = ~in067 & in167;
  assign new_n757 = in067 & ~in167;
  assign new_n758 = ~in066 & in166;
  assign new_n759 = in066 & ~in166;
  assign new_n760 = ~in065 & in165;
  assign new_n761 = in064 & ~in164;
  assign new_n762 = in065 & ~in165;
  assign new_n763 = ~in064 & in164;
  assign new_n764 = ~in056 & in156;
  assign new_n765 = in055 & ~in155;
  assign new_n766 = in046 & ~in146;
  assign new_n767 = in047 & ~in147;
  assign new_n768 = ~in046 & in146;
  assign new_n769 = in045 & ~in145;
  assign new_n770 = ~in045 & in145;
  assign new_n771 = in044 & ~in144;
  assign new_n772 = ~in044 & in144;
  assign new_n773 = ~in039 & in139;
  assign new_n774 = in038 & ~in138;
  assign new_n775 = in039 & ~in139;
  assign new_n776 = ~in038 & in138;
  assign new_n777 = in037 & ~in137;
  assign new_n778 = ~in037 & in137;
  assign new_n779 = in031 & ~in131;
  assign new_n780 = in030 & ~in130;
  assign new_n781 = ~in029 & in129;
  assign new_n782 = ~in030 & in130;
  assign new_n783 = in029 & ~in129;
  assign new_n784 = ~in028 & in128;
  assign new_n785 = in028 & ~in128;
  assign new_n786 = ~in027 & in127;
  assign new_n787 = in027 & ~in127;
  assign new_n788 = ~in026 & in126;
  assign new_n789 = in026 & ~in126;
  assign new_n790 = ~in025 & in125;
  assign new_n791 = in025 & ~in125;
  assign new_n792 = ~in024 & in124;
  assign new_n793 = in024 & ~in124;
  assign new_n794 = ~in023 & in123;
  assign new_n795 = in023 & ~in123;
  assign new_n796 = ~in022 & in122;
  assign new_n797 = in022 & ~in122;
  assign new_n798 = ~in021 & in121;
  assign new_n799 = in021 & ~in121;
  assign new_n800 = ~in020 & in120;
  assign new_n801 = in020 & ~in120;
  assign new_n802 = ~in019 & in119;
  assign new_n803 = in019 & ~in119;
  assign new_n804 = ~in018 & in118;
  assign new_n805 = in018 & ~in118;
  assign new_n806 = ~in017 & in117;
  assign new_n807 = in017 & ~in117;
  assign new_n808 = ~in016 & in116;
  assign new_n809 = in016 & ~in116;
  assign new_n810 = ~in015 & in115;
  assign new_n811 = in015 & ~in115;
  assign new_n812 = ~in014 & in114;
  assign new_n813 = in014 & ~in114;
  assign new_n814 = ~in013 & in113;
  assign new_n815 = in013 & ~in113;
  assign new_n816 = ~in012 & in112;
  assign new_n817 = in012 & ~in112;
  assign new_n818 = ~in011 & in111;
  assign new_n819 = in010 & ~in110;
  assign new_n820 = in011 & ~in111;
  assign new_n821 = ~in010 & in110;
  assign new_n822 = in09 & ~in19;
  assign new_n823 = ~in09 & in19;
  assign new_n824 = in08 & ~in18;
  assign new_n825 = ~in08 & in18;
  assign new_n826 = in07 & ~in17;
  assign new_n827 = ~in07 & in17;
  assign new_n828 = in06 & ~in16;
  assign new_n829 = ~in05 & in15;
  assign new_n830 = ~in06 & in16;
  assign new_n831 = in05 & ~in15;
  assign new_n832 = ~in04 & in14;
  assign new_n833 = in04 & ~in14;
  assign new_n834 = in03 & ~in13;
  assign new_n835 = ~in02 & in12;
  assign new_n836 = ~in03 & in13;
  assign new_n837 = in02 & ~in12;
  assign new_n838 = in00 & ~in10;
  assign new_n839 = in01 & new_n838;
  assign new_n840 = in11 & ~new_n839;
  assign new_n841 = ~in01 & ~new_n838;
  assign new_n842 = ~new_n840 & ~new_n841;
  assign new_n843 = ~new_n837 & ~new_n842;
  assign new_n844 = ~new_n835 & ~new_n836;
  assign new_n845 = ~new_n843 & new_n844;
  assign new_n846 = ~new_n833 & ~new_n834;
  assign new_n847 = ~new_n845 & new_n846;
  assign new_n848 = ~new_n832 & ~new_n847;
  assign new_n849 = ~new_n831 & ~new_n848;
  assign new_n850 = ~new_n829 & ~new_n830;
  assign new_n851 = ~new_n849 & new_n850;
  assign new_n852 = ~new_n828 & ~new_n851;
  assign new_n853 = ~new_n827 & ~new_n852;
  assign new_n854 = ~new_n826 & ~new_n853;
  assign new_n855 = ~new_n825 & ~new_n854;
  assign new_n856 = ~new_n824 & ~new_n855;
  assign new_n857 = ~new_n823 & ~new_n856;
  assign new_n858 = ~new_n822 & ~new_n857;
  assign new_n859 = ~new_n821 & ~new_n858;
  assign new_n860 = ~new_n819 & ~new_n820;
  assign new_n861 = ~new_n859 & new_n860;
  assign new_n862 = ~new_n818 & ~new_n861;
  assign new_n863 = ~new_n817 & ~new_n862;
  assign new_n864 = ~new_n816 & ~new_n863;
  assign new_n865 = ~new_n815 & ~new_n864;
  assign new_n866 = ~new_n814 & ~new_n865;
  assign new_n867 = ~new_n813 & ~new_n866;
  assign new_n868 = ~new_n812 & ~new_n867;
  assign new_n869 = ~new_n811 & ~new_n868;
  assign new_n870 = ~new_n810 & ~new_n869;
  assign new_n871 = ~new_n809 & ~new_n870;
  assign new_n872 = ~new_n808 & ~new_n871;
  assign new_n873 = ~new_n807 & ~new_n872;
  assign new_n874 = ~new_n806 & ~new_n873;
  assign new_n875 = ~new_n805 & ~new_n874;
  assign new_n876 = ~new_n804 & ~new_n875;
  assign new_n877 = ~new_n803 & ~new_n876;
  assign new_n878 = ~new_n802 & ~new_n877;
  assign new_n879 = ~new_n801 & ~new_n878;
  assign new_n880 = ~new_n800 & ~new_n879;
  assign new_n881 = ~new_n799 & ~new_n880;
  assign new_n882 = ~new_n798 & ~new_n881;
  assign new_n883 = ~new_n797 & ~new_n882;
  assign new_n884 = ~new_n796 & ~new_n883;
  assign new_n885 = ~new_n795 & ~new_n884;
  assign new_n886 = ~new_n794 & ~new_n885;
  assign new_n887 = ~new_n793 & ~new_n886;
  assign new_n888 = ~new_n792 & ~new_n887;
  assign new_n889 = ~new_n791 & ~new_n888;
  assign new_n890 = ~new_n790 & ~new_n889;
  assign new_n891 = ~new_n789 & ~new_n890;
  assign new_n892 = ~new_n788 & ~new_n891;
  assign new_n893 = ~new_n787 & ~new_n892;
  assign new_n894 = ~new_n786 & ~new_n893;
  assign new_n895 = ~new_n785 & ~new_n894;
  assign new_n896 = ~new_n784 & ~new_n895;
  assign new_n897 = ~new_n783 & ~new_n896;
  assign new_n898 = ~new_n781 & ~new_n782;
  assign new_n899 = ~new_n897 & new_n898;
  assign new_n900 = ~new_n779 & ~new_n780;
  assign new_n901 = ~new_n899 & new_n900;
  assign new_n902 = ~in036 & in136;
  assign new_n903 = ~in032 & in132;
  assign new_n904 = ~in033 & in133;
  assign new_n905 = ~in035 & in135;
  assign new_n906 = ~in034 & in134;
  assign new_n907 = ~new_n905 & ~new_n906;
  assign new_n908 = ~in031 & in131;
  assign new_n909 = ~new_n902 & ~new_n903;
  assign new_n910 = ~new_n904 & ~new_n908;
  assign new_n911 = new_n909 & new_n910;
  assign new_n912 = new_n907 & new_n911;
  assign new_n913 = ~new_n901 & new_n912;
  assign new_n914 = in036 & ~in136;
  assign new_n915 = in035 & ~in135;
  assign new_n916 = in033 & ~in133;
  assign new_n917 = in034 & ~in134;
  assign new_n918 = in032 & ~in132;
  assign new_n919 = ~new_n904 & new_n918;
  assign new_n920 = ~new_n916 & ~new_n917;
  assign new_n921 = ~new_n919 & new_n920;
  assign new_n922 = new_n907 & ~new_n921;
  assign new_n923 = ~new_n915 & ~new_n922;
  assign new_n924 = ~new_n902 & ~new_n923;
  assign new_n925 = ~new_n914 & ~new_n924;
  assign new_n926 = ~new_n913 & new_n925;
  assign new_n927 = ~new_n778 & ~new_n926;
  assign new_n928 = ~new_n777 & ~new_n927;
  assign new_n929 = ~new_n776 & ~new_n928;
  assign new_n930 = ~new_n774 & ~new_n775;
  assign new_n931 = ~new_n929 & new_n930;
  assign new_n932 = ~in041 & in141;
  assign new_n933 = ~in040 & in140;
  assign new_n934 = ~new_n773 & ~new_n932;
  assign new_n935 = ~new_n933 & new_n934;
  assign new_n936 = ~new_n931 & new_n935;
  assign new_n937 = in042 & ~in142;
  assign new_n938 = in041 & ~in141;
  assign new_n939 = in040 & ~in140;
  assign new_n940 = ~new_n932 & new_n939;
  assign new_n941 = ~new_n937 & ~new_n938;
  assign new_n942 = ~new_n940 & new_n941;
  assign new_n943 = ~new_n936 & new_n942;
  assign new_n944 = ~in042 & in142;
  assign new_n945 = ~in043 & in143;
  assign new_n946 = ~new_n944 & ~new_n945;
  assign new_n947 = ~new_n943 & new_n946;
  assign new_n948 = in043 & ~in143;
  assign new_n949 = ~new_n947 & ~new_n948;
  assign new_n950 = ~new_n772 & ~new_n949;
  assign new_n951 = ~new_n771 & ~new_n950;
  assign new_n952 = ~new_n770 & ~new_n951;
  assign new_n953 = ~new_n769 & ~new_n952;
  assign new_n954 = ~new_n768 & ~new_n953;
  assign new_n955 = ~new_n766 & ~new_n767;
  assign new_n956 = ~new_n954 & new_n955;
  assign new_n957 = ~in055 & in155;
  assign new_n958 = ~in054 & in154;
  assign new_n959 = ~new_n957 & ~new_n958;
  assign new_n960 = ~in053 & in153;
  assign new_n961 = ~in052 & in152;
  assign new_n962 = ~new_n960 & ~new_n961;
  assign new_n963 = ~in049 & in149;
  assign new_n964 = ~in051 & in151;
  assign new_n965 = ~in050 & in150;
  assign new_n966 = ~new_n964 & ~new_n965;
  assign new_n967 = ~in048 & in148;
  assign new_n968 = ~in047 & in147;
  assign new_n969 = ~new_n963 & ~new_n967;
  assign new_n970 = ~new_n968 & new_n969;
  assign new_n971 = new_n959 & new_n962;
  assign new_n972 = new_n966 & new_n971;
  assign new_n973 = new_n970 & new_n972;
  assign new_n974 = ~new_n956 & new_n973;
  assign new_n975 = in053 & ~in153;
  assign new_n976 = in054 & ~in154;
  assign new_n977 = in052 & ~in152;
  assign new_n978 = in051 & ~in151;
  assign new_n979 = in050 & ~in150;
  assign new_n980 = in049 & ~in149;
  assign new_n981 = in048 & ~in148;
  assign new_n982 = ~new_n963 & new_n981;
  assign new_n983 = ~new_n979 & ~new_n980;
  assign new_n984 = ~new_n982 & new_n983;
  assign new_n985 = new_n966 & ~new_n984;
  assign new_n986 = ~new_n977 & ~new_n978;
  assign new_n987 = ~new_n985 & new_n986;
  assign new_n988 = new_n962 & ~new_n987;
  assign new_n989 = ~new_n975 & ~new_n976;
  assign new_n990 = ~new_n988 & new_n989;
  assign new_n991 = new_n959 & ~new_n990;
  assign new_n992 = ~new_n765 & ~new_n991;
  assign new_n993 = ~new_n974 & new_n992;
  assign new_n994 = ~in057 & in157;
  assign new_n995 = ~in059 & in159;
  assign new_n996 = ~in058 & in158;
  assign new_n997 = ~in063 & in163;
  assign new_n998 = ~in062 & in162;
  assign new_n999 = ~new_n997 & ~new_n998;
  assign new_n1000 = ~in061 & in161;
  assign new_n1001 = ~in060 & in160;
  assign new_n1002 = ~new_n1000 & ~new_n1001;
  assign new_n1003 = new_n999 & new_n1002;
  assign new_n1004 = ~new_n995 & ~new_n996;
  assign new_n1005 = new_n1003 & new_n1004;
  assign new_n1006 = ~new_n764 & ~new_n994;
  assign new_n1007 = new_n1005 & new_n1006;
  assign new_n1008 = ~new_n993 & new_n1007;
  assign new_n1009 = in058 & ~in158;
  assign new_n1010 = in057 & ~in157;
  assign new_n1011 = in056 & ~in156;
  assign new_n1012 = ~new_n994 & new_n1011;
  assign new_n1013 = ~new_n1009 & ~new_n1010;
  assign new_n1014 = ~new_n1012 & new_n1013;
  assign new_n1015 = new_n1005 & ~new_n1014;
  assign new_n1016 = in062 & ~in162;
  assign new_n1017 = in061 & ~in161;
  assign new_n1018 = ~new_n1016 & ~new_n1017;
  assign new_n1019 = new_n999 & ~new_n1018;
  assign new_n1020 = in060 & ~in160;
  assign new_n1021 = in059 & ~in159;
  assign new_n1022 = ~new_n1020 & ~new_n1021;
  assign new_n1023 = new_n1003 & ~new_n1022;
  assign new_n1024 = in063 & ~in163;
  assign new_n1025 = ~new_n1019 & ~new_n1024;
  assign new_n1026 = ~new_n1023 & new_n1025;
  assign new_n1027 = ~new_n1015 & new_n1026;
  assign new_n1028 = ~new_n1008 & new_n1027;
  assign new_n1029 = ~new_n763 & ~new_n1028;
  assign new_n1030 = ~new_n761 & ~new_n762;
  assign new_n1031 = ~new_n1029 & new_n1030;
  assign new_n1032 = ~new_n760 & ~new_n1031;
  assign new_n1033 = ~new_n759 & ~new_n1032;
  assign new_n1034 = ~new_n758 & ~new_n1033;
  assign new_n1035 = ~new_n757 & ~new_n1034;
  assign new_n1036 = ~new_n756 & ~new_n1035;
  assign new_n1037 = ~new_n755 & ~new_n1036;
  assign new_n1038 = ~new_n754 & ~new_n1037;
  assign new_n1039 = ~new_n753 & ~new_n1038;
  assign new_n1040 = ~new_n751 & ~new_n752;
  assign new_n1041 = ~new_n1039 & new_n1040;
  assign new_n1042 = ~new_n749 & ~new_n750;
  assign new_n1043 = ~new_n1041 & new_n1042;
  assign new_n1044 = ~in072 & in172;
  assign new_n1045 = ~in071 & in171;
  assign new_n1046 = ~new_n748 & ~new_n1044;
  assign new_n1047 = ~new_n1045 & new_n1046;
  assign new_n1048 = ~new_n1043 & new_n1047;
  assign new_n1049 = in074 & ~in174;
  assign new_n1050 = in073 & ~in173;
  assign new_n1051 = in072 & ~in172;
  assign new_n1052 = ~new_n748 & new_n1051;
  assign new_n1053 = ~new_n1049 & ~new_n1050;
  assign new_n1054 = ~new_n1052 & new_n1053;
  assign new_n1055 = ~new_n1048 & new_n1054;
  assign new_n1056 = ~in074 & in174;
  assign new_n1057 = ~new_n1055 & ~new_n1056;
  assign new_n1058 = in075 & ~in175;
  assign new_n1059 = ~new_n1057 & ~new_n1058;
  assign new_n1060 = ~in075 & in175;
  assign new_n1061 = ~new_n747 & ~new_n1060;
  assign new_n1062 = new_n741 & new_n1061;
  assign new_n1063 = ~new_n1059 & new_n1062;
  assign new_n1064 = ~new_n743 & ~new_n744;
  assign new_n1065 = ~new_n746 & new_n1064;
  assign new_n1066 = ~new_n742 & new_n1065;
  assign new_n1067 = ~new_n1063 & new_n1066;
  assign new_n1068 = ~in080 & in180;
  assign new_n1069 = ~in081 & in181;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = ~new_n1067 & new_n1070;
  assign new_n1072 = in082 & ~in182;
  assign new_n1073 = in081 & ~in181;
  assign new_n1074 = ~new_n1072 & ~new_n1073;
  assign new_n1075 = ~new_n1071 & new_n1074;
  assign new_n1076 = ~new_n733 & ~new_n1075;
  assign new_n1077 = ~new_n732 & ~new_n1076;
  assign new_n1078 = ~new_n731 & ~new_n1077;
  assign new_n1079 = ~new_n730 & ~new_n1078;
  assign new_n1080 = ~new_n729 & ~new_n1079;
  assign new_n1081 = ~new_n728 & ~new_n1080;
  assign new_n1082 = ~new_n726 & ~new_n727;
  assign new_n1083 = ~new_n1081 & new_n1082;
  assign new_n1084 = ~new_n725 & ~new_n1083;
  assign new_n1085 = ~new_n724 & ~new_n1084;
  assign new_n1086 = ~new_n723 & ~new_n1085;
  assign new_n1087 = ~new_n722 & ~new_n1086;
  assign new_n1088 = ~new_n721 & ~new_n1087;
  assign new_n1089 = ~new_n720 & ~new_n1088;
  assign new_n1090 = ~new_n718 & ~new_n719;
  assign new_n1091 = ~new_n1089 & new_n1090;
  assign new_n1092 = ~new_n717 & ~new_n1091;
  assign new_n1093 = ~new_n716 & ~new_n1092;
  assign new_n1094 = ~new_n715 & ~new_n1093;
  assign new_n1095 = ~new_n714 & ~new_n1094;
  assign new_n1096 = ~new_n713 & ~new_n1095;
  assign new_n1097 = ~new_n712 & ~new_n1096;
  assign new_n1098 = ~new_n710 & ~new_n711;
  assign new_n1099 = ~new_n1097 & new_n1098;
  assign new_n1100 = ~new_n709 & ~new_n1099;
  assign new_n1101 = ~new_n708 & ~new_n1100;
  assign new_n1102 = ~new_n707 & ~new_n1101;
  assign new_n1103 = ~new_n706 & ~new_n1102;
  assign new_n1104 = ~new_n705 & ~new_n1103;
  assign new_n1105 = ~new_n704 & ~new_n1104;
  assign new_n1106 = ~new_n702 & ~new_n703;
  assign new_n1107 = ~new_n1105 & new_n1106;
  assign new_n1108 = ~new_n701 & ~new_n1107;
  assign new_n1109 = ~new_n700 & ~new_n1108;
  assign new_n1110 = ~new_n699 & ~new_n1109;
  assign new_n1111 = ~new_n698 & ~new_n1110;
  assign new_n1112 = ~new_n697 & ~new_n1111;
  assign new_n1113 = ~new_n696 & ~new_n1112;
  assign new_n1114 = ~new_n694 & ~new_n695;
  assign new_n1115 = ~new_n1113 & new_n1114;
  assign new_n1116 = ~new_n693 & ~new_n1115;
  assign new_n1117 = ~new_n692 & ~new_n1116;
  assign new_n1118 = ~new_n691 & ~new_n1117;
  assign new_n1119 = ~new_n690 & ~new_n1118;
  assign new_n1120 = ~new_n689 & ~new_n1119;
  assign new_n1121 = ~new_n688 & ~new_n1120;
  assign new_n1122 = ~new_n686 & ~new_n687;
  assign new_n1123 = ~new_n1121 & new_n1122;
  assign new_n1124 = ~new_n685 & ~new_n1123;
  assign new_n1125 = ~new_n684 & ~new_n1124;
  assign new_n1126 = ~new_n683 & ~new_n1125;
  assign new_n1127 = ~new_n682 & ~new_n1126;
  assign new_n1128 = ~new_n681 & ~new_n1127;
  assign new_n1129 = ~new_n680 & ~new_n1128;
  assign new_n1130 = ~new_n678 & ~new_n679;
  assign new_n1131 = ~new_n1129 & new_n1130;
  assign new_n1132 = ~new_n677 & ~new_n1131;
  assign new_n1133 = ~new_n676 & ~new_n1132;
  assign new_n1134 = ~new_n675 & ~new_n1133;
  assign new_n1135 = ~new_n674 & ~new_n1134;
  assign new_n1136 = ~new_n673 & ~new_n1135;
  assign new_n1137 = ~new_n672 & ~new_n1136;
  assign new_n1138 = ~new_n671 & ~new_n1137;
  assign new_n1139 = ~new_n670 & ~new_n1138;
  assign new_n1140 = ~new_n669 & ~new_n1139;
  assign new_n1141 = ~new_n668 & ~new_n1140;
  assign new_n1142 = ~new_n667 & ~new_n1141;
  assign new_n1143 = ~new_n666 & ~new_n1142;
  assign new_n1144 = ~new_n665 & ~new_n1143;
  assign new_n1145 = ~new_n664 & ~new_n1144;
  assign new_n1146 = ~new_n663 & ~new_n1145;
  assign new_n1147 = ~new_n662 & ~new_n1146;
  assign new_n1148 = ~new_n661 & ~new_n1147;
  assign new_n1149 = ~new_n660 & ~new_n1148;
  assign new_n1150 = ~new_n659 & ~new_n1149;
  assign new_n1151 = ~new_n658 & ~new_n1150;
  assign new_n1152 = ~new_n656 & ~new_n657;
  assign new_n1153 = ~new_n1151 & new_n1152;
  assign new_n1154 = ~new_n654 & ~new_n655;
  assign new_n1155 = ~new_n1153 & new_n1154;
  assign new_n1156 = ~new_n652 & ~new_n653;
  assign new_n1157 = ~new_n1155 & new_n1156;
  assign new_n1158 = ~in0123 & in1123;
  assign new_n1159 = ~new_n651 & ~new_n1158;
  assign new_n1160 = new_n646 & new_n1159;
  assign new_n1161 = ~new_n1157 & new_n1160;
  assign new_n1162 = ~new_n643 & ~new_n650;
  assign new_n1163 = ~new_n1161 & new_n1162;
  assign new_n1164 = in0127 & new_n1163;
  assign new_n1165 = in1127 & ~new_n1164;
  assign new_n1166 = ~in0127 & ~new_n1163;
  assign new_n1167 = ~new_n1165 & ~new_n1166;
  assign new_n1168 = in00 & ~new_n1167;
  assign new_n1169 = in10 & new_n1167;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = in2127 & in3127;
  assign new_n1172 = in0127 & in1127;
  assign new_n1173 = in2126 & ~in3126;
  assign new_n1174 = ~in2125 & in3125;
  assign new_n1175 = ~in2126 & in3126;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = in2125 & ~in3125;
  assign new_n1178 = in2124 & ~in3124;
  assign new_n1179 = ~new_n1177 & ~new_n1178;
  assign new_n1180 = new_n1176 & ~new_n1179;
  assign new_n1181 = ~in2124 & in3124;
  assign new_n1182 = in2123 & ~in3123;
  assign new_n1183 = in2122 & ~in3122;
  assign new_n1184 = ~in2122 & in3122;
  assign new_n1185 = ~in2121 & in3121;
  assign new_n1186 = in2120 & ~in3120;
  assign new_n1187 = in2121 & ~in3121;
  assign new_n1188 = ~in2120 & in3120;
  assign new_n1189 = in2119 & ~in3119;
  assign new_n1190 = ~in2119 & in3119;
  assign new_n1191 = in2118 & ~in3118;
  assign new_n1192 = ~in2118 & in3118;
  assign new_n1193 = in2117 & ~in3117;
  assign new_n1194 = ~in2117 & in3117;
  assign new_n1195 = in2116 & ~in3116;
  assign new_n1196 = ~in2116 & in3116;
  assign new_n1197 = in2115 & ~in3115;
  assign new_n1198 = ~in2115 & in3115;
  assign new_n1199 = in2114 & ~in3114;
  assign new_n1200 = ~in2114 & in3114;
  assign new_n1201 = in2113 & ~in3113;
  assign new_n1202 = ~in2113 & in3113;
  assign new_n1203 = in2112 & ~in3112;
  assign new_n1204 = ~in2112 & in3112;
  assign new_n1205 = in2111 & ~in3111;
  assign new_n1206 = ~in2111 & in3111;
  assign new_n1207 = in2110 & ~in3110;
  assign new_n1208 = ~in2109 & in3109;
  assign new_n1209 = ~in2110 & in3110;
  assign new_n1210 = in2109 & ~in3109;
  assign new_n1211 = ~in2108 & in3108;
  assign new_n1212 = in2108 & ~in3108;
  assign new_n1213 = ~in2107 & in3107;
  assign new_n1214 = in2107 & ~in3107;
  assign new_n1215 = ~in2106 & in3106;
  assign new_n1216 = in2105 & ~in3105;
  assign new_n1217 = in2106 & ~in3106;
  assign new_n1218 = ~in2105 & in3105;
  assign new_n1219 = in2104 & ~in3104;
  assign new_n1220 = ~in2104 & in3104;
  assign new_n1221 = in2103 & ~in3103;
  assign new_n1222 = ~in2103 & in3103;
  assign new_n1223 = in2102 & ~in3102;
  assign new_n1224 = ~in2101 & in3101;
  assign new_n1225 = ~in2102 & in3102;
  assign new_n1226 = in2101 & ~in3101;
  assign new_n1227 = ~in2100 & in3100;
  assign new_n1228 = in2100 & ~in3100;
  assign new_n1229 = ~in299 & in399;
  assign new_n1230 = in299 & ~in399;
  assign new_n1231 = ~in298 & in398;
  assign new_n1232 = in297 & ~in397;
  assign new_n1233 = in298 & ~in398;
  assign new_n1234 = ~in297 & in397;
  assign new_n1235 = in296 & ~in396;
  assign new_n1236 = ~in296 & in396;
  assign new_n1237 = in295 & ~in395;
  assign new_n1238 = ~in295 & in395;
  assign new_n1239 = in294 & ~in394;
  assign new_n1240 = ~in293 & in393;
  assign new_n1241 = ~in294 & in394;
  assign new_n1242 = in293 & ~in393;
  assign new_n1243 = ~in292 & in392;
  assign new_n1244 = in292 & ~in392;
  assign new_n1245 = ~in291 & in391;
  assign new_n1246 = in291 & ~in391;
  assign new_n1247 = ~in290 & in390;
  assign new_n1248 = in289 & ~in389;
  assign new_n1249 = in290 & ~in390;
  assign new_n1250 = ~in289 & in389;
  assign new_n1251 = in288 & ~in388;
  assign new_n1252 = ~in288 & in388;
  assign new_n1253 = in287 & ~in387;
  assign new_n1254 = ~in287 & in387;
  assign new_n1255 = in286 & ~in386;
  assign new_n1256 = ~in285 & in385;
  assign new_n1257 = ~in286 & in386;
  assign new_n1258 = in285 & ~in385;
  assign new_n1259 = ~in284 & in384;
  assign new_n1260 = in284 & ~in384;
  assign new_n1261 = ~in283 & in383;
  assign new_n1262 = in283 & ~in383;
  assign new_n1263 = ~in282 & in382;
  assign new_n1264 = in281 & ~in381;
  assign new_n1265 = in282 & ~in382;
  assign new_n1266 = ~in281 & in381;
  assign new_n1267 = in280 & ~in380;
  assign new_n1268 = ~in280 & in380;
  assign new_n1269 = in279 & ~in379;
  assign new_n1270 = ~in279 & in379;
  assign new_n1271 = in278 & ~in378;
  assign new_n1272 = ~in277 & in377;
  assign new_n1273 = ~in278 & in378;
  assign new_n1274 = in277 & ~in377;
  assign new_n1275 = ~in276 & in376;
  assign new_n1276 = in276 & ~in376;
  assign new_n1277 = ~in275 & in375;
  assign new_n1278 = in275 & ~in375;
  assign new_n1279 = ~in274 & in374;
  assign new_n1280 = in273 & ~in373;
  assign new_n1281 = in274 & ~in374;
  assign new_n1282 = ~in273 & in373;
  assign new_n1283 = in272 & ~in372;
  assign new_n1284 = ~in272 & in372;
  assign new_n1285 = in271 & ~in371;
  assign new_n1286 = ~in271 & in371;
  assign new_n1287 = in270 & ~in370;
  assign new_n1288 = ~in269 & in369;
  assign new_n1289 = ~in270 & in370;
  assign new_n1290 = in269 & ~in369;
  assign new_n1291 = ~in268 & in368;
  assign new_n1292 = ~in263 & in363;
  assign new_n1293 = ~in258 & in358;
  assign new_n1294 = in257 & ~in357;
  assign new_n1295 = in258 & ~in358;
  assign new_n1296 = ~in257 & in357;
  assign new_n1297 = in256 & ~in356;
  assign new_n1298 = ~in256 & in356;
  assign new_n1299 = in247 & ~in347;
  assign new_n1300 = in246 & ~in346;
  assign new_n1301 = ~in246 & in346;
  assign new_n1302 = ~in245 & in345;
  assign new_n1303 = in245 & ~in345;
  assign new_n1304 = in239 & ~in339;
  assign new_n1305 = in238 & ~in338;
  assign new_n1306 = ~in238 & in338;
  assign new_n1307 = ~in237 & in337;
  assign new_n1308 = in237 & ~in337;
  assign new_n1309 = in231 & ~in331;
  assign new_n1310 = in230 & ~in330;
  assign new_n1311 = ~in229 & in329;
  assign new_n1312 = ~in230 & in330;
  assign new_n1313 = in229 & ~in329;
  assign new_n1314 = ~in228 & in328;
  assign new_n1315 = in228 & ~in328;
  assign new_n1316 = ~in227 & in327;
  assign new_n1317 = in227 & ~in327;
  assign new_n1318 = ~in226 & in326;
  assign new_n1319 = in226 & ~in326;
  assign new_n1320 = ~in225 & in325;
  assign new_n1321 = in225 & ~in325;
  assign new_n1322 = ~in224 & in324;
  assign new_n1323 = in224 & ~in324;
  assign new_n1324 = ~in223 & in323;
  assign new_n1325 = in223 & ~in323;
  assign new_n1326 = ~in222 & in322;
  assign new_n1327 = in222 & ~in322;
  assign new_n1328 = ~in221 & in321;
  assign new_n1329 = in220 & ~in320;
  assign new_n1330 = in221 & ~in321;
  assign new_n1331 = ~in220 & in320;
  assign new_n1332 = in219 & ~in319;
  assign new_n1333 = ~in219 & in319;
  assign new_n1334 = in218 & ~in318;
  assign new_n1335 = ~in218 & in318;
  assign new_n1336 = in217 & ~in317;
  assign new_n1337 = ~in217 & in317;
  assign new_n1338 = in216 & ~in316;
  assign new_n1339 = ~in216 & in316;
  assign new_n1340 = in215 & ~in315;
  assign new_n1341 = ~in214 & in314;
  assign new_n1342 = ~in215 & in315;
  assign new_n1343 = in214 & ~in314;
  assign new_n1344 = ~in213 & in313;
  assign new_n1345 = in213 & ~in313;
  assign new_n1346 = ~in212 & in312;
  assign new_n1347 = in212 & ~in312;
  assign new_n1348 = ~in211 & in311;
  assign new_n1349 = in210 & ~in310;
  assign new_n1350 = in211 & ~in311;
  assign new_n1351 = ~in210 & in310;
  assign new_n1352 = in29 & ~in39;
  assign new_n1353 = ~in29 & in39;
  assign new_n1354 = in28 & ~in38;
  assign new_n1355 = ~in28 & in38;
  assign new_n1356 = in27 & ~in37;
  assign new_n1357 = ~in26 & in36;
  assign new_n1358 = ~in27 & in37;
  assign new_n1359 = in26 & ~in36;
  assign new_n1360 = ~in25 & in35;
  assign new_n1361 = in25 & ~in35;
  assign new_n1362 = in24 & ~in34;
  assign new_n1363 = ~in23 & in33;
  assign new_n1364 = ~in24 & in34;
  assign new_n1365 = in23 & ~in33;
  assign new_n1366 = ~in22 & in32;
  assign new_n1367 = in22 & ~in32;
  assign new_n1368 = ~in21 & in31;
  assign new_n1369 = in21 & ~in31;
  assign new_n1370 = in20 & ~in30;
  assign new_n1371 = ~new_n1369 & ~new_n1370;
  assign new_n1372 = ~new_n1368 & ~new_n1371;
  assign new_n1373 = ~new_n1367 & ~new_n1372;
  assign new_n1374 = ~new_n1366 & ~new_n1373;
  assign new_n1375 = ~new_n1365 & ~new_n1374;
  assign new_n1376 = ~new_n1363 & ~new_n1364;
  assign new_n1377 = ~new_n1375 & new_n1376;
  assign new_n1378 = ~new_n1361 & ~new_n1362;
  assign new_n1379 = ~new_n1377 & new_n1378;
  assign new_n1380 = ~new_n1360 & ~new_n1379;
  assign new_n1381 = ~new_n1359 & ~new_n1380;
  assign new_n1382 = ~new_n1357 & ~new_n1358;
  assign new_n1383 = ~new_n1381 & new_n1382;
  assign new_n1384 = ~new_n1356 & ~new_n1383;
  assign new_n1385 = ~new_n1355 & ~new_n1384;
  assign new_n1386 = ~new_n1354 & ~new_n1385;
  assign new_n1387 = ~new_n1353 & ~new_n1386;
  assign new_n1388 = ~new_n1352 & ~new_n1387;
  assign new_n1389 = ~new_n1351 & ~new_n1388;
  assign new_n1390 = ~new_n1349 & ~new_n1350;
  assign new_n1391 = ~new_n1389 & new_n1390;
  assign new_n1392 = ~new_n1348 & ~new_n1391;
  assign new_n1393 = ~new_n1347 & ~new_n1392;
  assign new_n1394 = ~new_n1346 & ~new_n1393;
  assign new_n1395 = ~new_n1345 & ~new_n1394;
  assign new_n1396 = ~new_n1344 & ~new_n1395;
  assign new_n1397 = ~new_n1343 & ~new_n1396;
  assign new_n1398 = ~new_n1341 & ~new_n1342;
  assign new_n1399 = ~new_n1397 & new_n1398;
  assign new_n1400 = ~new_n1340 & ~new_n1399;
  assign new_n1401 = ~new_n1339 & ~new_n1400;
  assign new_n1402 = ~new_n1338 & ~new_n1401;
  assign new_n1403 = ~new_n1337 & ~new_n1402;
  assign new_n1404 = ~new_n1336 & ~new_n1403;
  assign new_n1405 = ~new_n1335 & ~new_n1404;
  assign new_n1406 = ~new_n1334 & ~new_n1405;
  assign new_n1407 = ~new_n1333 & ~new_n1406;
  assign new_n1408 = ~new_n1332 & ~new_n1407;
  assign new_n1409 = ~new_n1331 & ~new_n1408;
  assign new_n1410 = ~new_n1329 & ~new_n1330;
  assign new_n1411 = ~new_n1409 & new_n1410;
  assign new_n1412 = ~new_n1328 & ~new_n1411;
  assign new_n1413 = ~new_n1327 & ~new_n1412;
  assign new_n1414 = ~new_n1326 & ~new_n1413;
  assign new_n1415 = ~new_n1325 & ~new_n1414;
  assign new_n1416 = ~new_n1324 & ~new_n1415;
  assign new_n1417 = ~new_n1323 & ~new_n1416;
  assign new_n1418 = ~new_n1322 & ~new_n1417;
  assign new_n1419 = ~new_n1321 & ~new_n1418;
  assign new_n1420 = ~new_n1320 & ~new_n1419;
  assign new_n1421 = ~new_n1319 & ~new_n1420;
  assign new_n1422 = ~new_n1318 & ~new_n1421;
  assign new_n1423 = ~new_n1317 & ~new_n1422;
  assign new_n1424 = ~new_n1316 & ~new_n1423;
  assign new_n1425 = ~new_n1315 & ~new_n1424;
  assign new_n1426 = ~new_n1314 & ~new_n1425;
  assign new_n1427 = ~new_n1313 & ~new_n1426;
  assign new_n1428 = ~new_n1311 & ~new_n1312;
  assign new_n1429 = ~new_n1427 & new_n1428;
  assign new_n1430 = ~new_n1309 & ~new_n1310;
  assign new_n1431 = ~new_n1429 & new_n1430;
  assign new_n1432 = ~in236 & in336;
  assign new_n1433 = ~in232 & in332;
  assign new_n1434 = ~in233 & in333;
  assign new_n1435 = ~in235 & in335;
  assign new_n1436 = ~in234 & in334;
  assign new_n1437 = ~new_n1435 & ~new_n1436;
  assign new_n1438 = ~in231 & in331;
  assign new_n1439 = ~new_n1432 & ~new_n1433;
  assign new_n1440 = ~new_n1434 & ~new_n1438;
  assign new_n1441 = new_n1439 & new_n1440;
  assign new_n1442 = new_n1437 & new_n1441;
  assign new_n1443 = ~new_n1431 & new_n1442;
  assign new_n1444 = in236 & ~in336;
  assign new_n1445 = in235 & ~in335;
  assign new_n1446 = in233 & ~in333;
  assign new_n1447 = in234 & ~in334;
  assign new_n1448 = in232 & ~in332;
  assign new_n1449 = ~new_n1434 & new_n1448;
  assign new_n1450 = ~new_n1446 & ~new_n1447;
  assign new_n1451 = ~new_n1449 & new_n1450;
  assign new_n1452 = new_n1437 & ~new_n1451;
  assign new_n1453 = ~new_n1445 & ~new_n1452;
  assign new_n1454 = ~new_n1432 & ~new_n1453;
  assign new_n1455 = ~new_n1308 & ~new_n1444;
  assign new_n1456 = ~new_n1454 & new_n1455;
  assign new_n1457 = ~new_n1443 & new_n1456;
  assign new_n1458 = ~new_n1306 & ~new_n1307;
  assign new_n1459 = ~new_n1457 & new_n1458;
  assign new_n1460 = ~new_n1304 & ~new_n1305;
  assign new_n1461 = ~new_n1459 & new_n1460;
  assign new_n1462 = ~in241 & in341;
  assign new_n1463 = ~in239 & in339;
  assign new_n1464 = ~in244 & in344;
  assign new_n1465 = ~in243 & in343;
  assign new_n1466 = ~in242 & in342;
  assign new_n1467 = ~new_n1465 & ~new_n1466;
  assign new_n1468 = ~in240 & in340;
  assign new_n1469 = ~new_n1462 & ~new_n1463;
  assign new_n1470 = ~new_n1464 & ~new_n1468;
  assign new_n1471 = new_n1469 & new_n1470;
  assign new_n1472 = new_n1467 & new_n1471;
  assign new_n1473 = ~new_n1461 & new_n1472;
  assign new_n1474 = in244 & ~in344;
  assign new_n1475 = in243 & ~in343;
  assign new_n1476 = in241 & ~in341;
  assign new_n1477 = in242 & ~in342;
  assign new_n1478 = in240 & ~in340;
  assign new_n1479 = ~new_n1462 & new_n1478;
  assign new_n1480 = ~new_n1476 & ~new_n1477;
  assign new_n1481 = ~new_n1479 & new_n1480;
  assign new_n1482 = new_n1467 & ~new_n1481;
  assign new_n1483 = ~new_n1475 & ~new_n1482;
  assign new_n1484 = ~new_n1464 & ~new_n1483;
  assign new_n1485 = ~new_n1303 & ~new_n1474;
  assign new_n1486 = ~new_n1484 & new_n1485;
  assign new_n1487 = ~new_n1473 & new_n1486;
  assign new_n1488 = ~new_n1301 & ~new_n1302;
  assign new_n1489 = ~new_n1487 & new_n1488;
  assign new_n1490 = ~new_n1299 & ~new_n1300;
  assign new_n1491 = ~new_n1489 & new_n1490;
  assign new_n1492 = ~in251 & in351;
  assign new_n1493 = ~in250 & in350;
  assign new_n1494 = ~new_n1492 & ~new_n1493;
  assign new_n1495 = ~in248 & in348;
  assign new_n1496 = ~in255 & in355;
  assign new_n1497 = ~in254 & in354;
  assign new_n1498 = ~new_n1496 & ~new_n1497;
  assign new_n1499 = ~in253 & in353;
  assign new_n1500 = ~in252 & in352;
  assign new_n1501 = ~new_n1499 & ~new_n1500;
  assign new_n1502 = new_n1498 & new_n1501;
  assign new_n1503 = ~in247 & in347;
  assign new_n1504 = ~in249 & in349;
  assign new_n1505 = ~new_n1495 & ~new_n1503;
  assign new_n1506 = ~new_n1504 & new_n1505;
  assign new_n1507 = new_n1494 & new_n1506;
  assign new_n1508 = new_n1502 & new_n1507;
  assign new_n1509 = ~new_n1491 & new_n1508;
  assign new_n1510 = in252 & ~in352;
  assign new_n1511 = in250 & ~in350;
  assign new_n1512 = in249 & ~in349;
  assign new_n1513 = in248 & ~in348;
  assign new_n1514 = ~new_n1504 & new_n1513;
  assign new_n1515 = ~new_n1511 & ~new_n1512;
  assign new_n1516 = ~new_n1514 & new_n1515;
  assign new_n1517 = new_n1494 & ~new_n1516;
  assign new_n1518 = in251 & ~in351;
  assign new_n1519 = ~new_n1510 & ~new_n1518;
  assign new_n1520 = ~new_n1517 & new_n1519;
  assign new_n1521 = new_n1502 & ~new_n1520;
  assign new_n1522 = in255 & ~in355;
  assign new_n1523 = in254 & ~in354;
  assign new_n1524 = in253 & ~in353;
  assign new_n1525 = ~new_n1523 & ~new_n1524;
  assign new_n1526 = new_n1498 & ~new_n1525;
  assign new_n1527 = ~new_n1522 & ~new_n1526;
  assign new_n1528 = ~new_n1521 & new_n1527;
  assign new_n1529 = ~new_n1509 & new_n1528;
  assign new_n1530 = ~new_n1298 & ~new_n1529;
  assign new_n1531 = ~new_n1297 & ~new_n1530;
  assign new_n1532 = ~new_n1296 & ~new_n1531;
  assign new_n1533 = ~new_n1294 & ~new_n1295;
  assign new_n1534 = ~new_n1532 & new_n1533;
  assign new_n1535 = ~in260 & in360;
  assign new_n1536 = ~in259 & in359;
  assign new_n1537 = ~new_n1293 & ~new_n1535;
  assign new_n1538 = ~new_n1536 & new_n1537;
  assign new_n1539 = ~new_n1534 & new_n1538;
  assign new_n1540 = in261 & ~in361;
  assign new_n1541 = in260 & ~in360;
  assign new_n1542 = in259 & ~in359;
  assign new_n1543 = ~new_n1535 & new_n1542;
  assign new_n1544 = ~new_n1540 & ~new_n1541;
  assign new_n1545 = ~new_n1543 & new_n1544;
  assign new_n1546 = ~new_n1539 & new_n1545;
  assign new_n1547 = ~in261 & in361;
  assign new_n1548 = ~in262 & in362;
  assign new_n1549 = ~new_n1547 & ~new_n1548;
  assign new_n1550 = ~new_n1546 & new_n1549;
  assign new_n1551 = in263 & ~in363;
  assign new_n1552 = in262 & ~in362;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = ~new_n1550 & new_n1553;
  assign new_n1555 = ~in265 & in365;
  assign new_n1556 = ~in264 & in364;
  assign new_n1557 = ~new_n1292 & ~new_n1555;
  assign new_n1558 = ~new_n1556 & new_n1557;
  assign new_n1559 = ~new_n1554 & new_n1558;
  assign new_n1560 = in266 & ~in366;
  assign new_n1561 = in265 & ~in365;
  assign new_n1562 = in264 & ~in364;
  assign new_n1563 = ~new_n1555 & new_n1562;
  assign new_n1564 = ~new_n1560 & ~new_n1561;
  assign new_n1565 = ~new_n1563 & new_n1564;
  assign new_n1566 = ~new_n1559 & new_n1565;
  assign new_n1567 = ~in266 & in366;
  assign new_n1568 = ~in267 & in367;
  assign new_n1569 = ~new_n1567 & ~new_n1568;
  assign new_n1570 = ~new_n1566 & new_n1569;
  assign new_n1571 = in268 & ~in368;
  assign new_n1572 = in267 & ~in367;
  assign new_n1573 = ~new_n1571 & ~new_n1572;
  assign new_n1574 = ~new_n1570 & new_n1573;
  assign new_n1575 = ~new_n1291 & ~new_n1574;
  assign new_n1576 = ~new_n1290 & ~new_n1575;
  assign new_n1577 = ~new_n1288 & ~new_n1289;
  assign new_n1578 = ~new_n1576 & new_n1577;
  assign new_n1579 = ~new_n1287 & ~new_n1578;
  assign new_n1580 = ~new_n1286 & ~new_n1579;
  assign new_n1581 = ~new_n1285 & ~new_n1580;
  assign new_n1582 = ~new_n1284 & ~new_n1581;
  assign new_n1583 = ~new_n1283 & ~new_n1582;
  assign new_n1584 = ~new_n1282 & ~new_n1583;
  assign new_n1585 = ~new_n1280 & ~new_n1281;
  assign new_n1586 = ~new_n1584 & new_n1585;
  assign new_n1587 = ~new_n1279 & ~new_n1586;
  assign new_n1588 = ~new_n1278 & ~new_n1587;
  assign new_n1589 = ~new_n1277 & ~new_n1588;
  assign new_n1590 = ~new_n1276 & ~new_n1589;
  assign new_n1591 = ~new_n1275 & ~new_n1590;
  assign new_n1592 = ~new_n1274 & ~new_n1591;
  assign new_n1593 = ~new_n1272 & ~new_n1273;
  assign new_n1594 = ~new_n1592 & new_n1593;
  assign new_n1595 = ~new_n1271 & ~new_n1594;
  assign new_n1596 = ~new_n1270 & ~new_n1595;
  assign new_n1597 = ~new_n1269 & ~new_n1596;
  assign new_n1598 = ~new_n1268 & ~new_n1597;
  assign new_n1599 = ~new_n1267 & ~new_n1598;
  assign new_n1600 = ~new_n1266 & ~new_n1599;
  assign new_n1601 = ~new_n1264 & ~new_n1265;
  assign new_n1602 = ~new_n1600 & new_n1601;
  assign new_n1603 = ~new_n1263 & ~new_n1602;
  assign new_n1604 = ~new_n1262 & ~new_n1603;
  assign new_n1605 = ~new_n1261 & ~new_n1604;
  assign new_n1606 = ~new_n1260 & ~new_n1605;
  assign new_n1607 = ~new_n1259 & ~new_n1606;
  assign new_n1608 = ~new_n1258 & ~new_n1607;
  assign new_n1609 = ~new_n1256 & ~new_n1257;
  assign new_n1610 = ~new_n1608 & new_n1609;
  assign new_n1611 = ~new_n1255 & ~new_n1610;
  assign new_n1612 = ~new_n1254 & ~new_n1611;
  assign new_n1613 = ~new_n1253 & ~new_n1612;
  assign new_n1614 = ~new_n1252 & ~new_n1613;
  assign new_n1615 = ~new_n1251 & ~new_n1614;
  assign new_n1616 = ~new_n1250 & ~new_n1615;
  assign new_n1617 = ~new_n1248 & ~new_n1249;
  assign new_n1618 = ~new_n1616 & new_n1617;
  assign new_n1619 = ~new_n1247 & ~new_n1618;
  assign new_n1620 = ~new_n1246 & ~new_n1619;
  assign new_n1621 = ~new_n1245 & ~new_n1620;
  assign new_n1622 = ~new_n1244 & ~new_n1621;
  assign new_n1623 = ~new_n1243 & ~new_n1622;
  assign new_n1624 = ~new_n1242 & ~new_n1623;
  assign new_n1625 = ~new_n1240 & ~new_n1241;
  assign new_n1626 = ~new_n1624 & new_n1625;
  assign new_n1627 = ~new_n1239 & ~new_n1626;
  assign new_n1628 = ~new_n1238 & ~new_n1627;
  assign new_n1629 = ~new_n1237 & ~new_n1628;
  assign new_n1630 = ~new_n1236 & ~new_n1629;
  assign new_n1631 = ~new_n1235 & ~new_n1630;
  assign new_n1632 = ~new_n1234 & ~new_n1631;
  assign new_n1633 = ~new_n1232 & ~new_n1233;
  assign new_n1634 = ~new_n1632 & new_n1633;
  assign new_n1635 = ~new_n1231 & ~new_n1634;
  assign new_n1636 = ~new_n1230 & ~new_n1635;
  assign new_n1637 = ~new_n1229 & ~new_n1636;
  assign new_n1638 = ~new_n1228 & ~new_n1637;
  assign new_n1639 = ~new_n1227 & ~new_n1638;
  assign new_n1640 = ~new_n1226 & ~new_n1639;
  assign new_n1641 = ~new_n1224 & ~new_n1225;
  assign new_n1642 = ~new_n1640 & new_n1641;
  assign new_n1643 = ~new_n1223 & ~new_n1642;
  assign new_n1644 = ~new_n1222 & ~new_n1643;
  assign new_n1645 = ~new_n1221 & ~new_n1644;
  assign new_n1646 = ~new_n1220 & ~new_n1645;
  assign new_n1647 = ~new_n1219 & ~new_n1646;
  assign new_n1648 = ~new_n1218 & ~new_n1647;
  assign new_n1649 = ~new_n1216 & ~new_n1217;
  assign new_n1650 = ~new_n1648 & new_n1649;
  assign new_n1651 = ~new_n1215 & ~new_n1650;
  assign new_n1652 = ~new_n1214 & ~new_n1651;
  assign new_n1653 = ~new_n1213 & ~new_n1652;
  assign new_n1654 = ~new_n1212 & ~new_n1653;
  assign new_n1655 = ~new_n1211 & ~new_n1654;
  assign new_n1656 = ~new_n1210 & ~new_n1655;
  assign new_n1657 = ~new_n1208 & ~new_n1209;
  assign new_n1658 = ~new_n1656 & new_n1657;
  assign new_n1659 = ~new_n1207 & ~new_n1658;
  assign new_n1660 = ~new_n1206 & ~new_n1659;
  assign new_n1661 = ~new_n1205 & ~new_n1660;
  assign new_n1662 = ~new_n1204 & ~new_n1661;
  assign new_n1663 = ~new_n1203 & ~new_n1662;
  assign new_n1664 = ~new_n1202 & ~new_n1663;
  assign new_n1665 = ~new_n1201 & ~new_n1664;
  assign new_n1666 = ~new_n1200 & ~new_n1665;
  assign new_n1667 = ~new_n1199 & ~new_n1666;
  assign new_n1668 = ~new_n1198 & ~new_n1667;
  assign new_n1669 = ~new_n1197 & ~new_n1668;
  assign new_n1670 = ~new_n1196 & ~new_n1669;
  assign new_n1671 = ~new_n1195 & ~new_n1670;
  assign new_n1672 = ~new_n1194 & ~new_n1671;
  assign new_n1673 = ~new_n1193 & ~new_n1672;
  assign new_n1674 = ~new_n1192 & ~new_n1673;
  assign new_n1675 = ~new_n1191 & ~new_n1674;
  assign new_n1676 = ~new_n1190 & ~new_n1675;
  assign new_n1677 = ~new_n1189 & ~new_n1676;
  assign new_n1678 = ~new_n1188 & ~new_n1677;
  assign new_n1679 = ~new_n1186 & ~new_n1187;
  assign new_n1680 = ~new_n1678 & new_n1679;
  assign new_n1681 = ~new_n1184 & ~new_n1185;
  assign new_n1682 = ~new_n1680 & new_n1681;
  assign new_n1683 = ~new_n1182 & ~new_n1183;
  assign new_n1684 = ~new_n1682 & new_n1683;
  assign new_n1685 = ~in2123 & in3123;
  assign new_n1686 = ~new_n1181 & ~new_n1685;
  assign new_n1687 = new_n1176 & new_n1686;
  assign new_n1688 = ~new_n1684 & new_n1687;
  assign new_n1689 = ~new_n1173 & ~new_n1180;
  assign new_n1690 = ~new_n1688 & new_n1689;
  assign new_n1691 = in2127 & new_n1690;
  assign new_n1692 = in3127 & ~new_n1691;
  assign new_n1693 = ~in2127 & ~new_n1690;
  assign new_n1694 = ~new_n1692 & ~new_n1693;
  assign new_n1695 = in2126 & ~new_n1694;
  assign new_n1696 = in3126 & new_n1694;
  assign new_n1697 = ~new_n1695 & ~new_n1696;
  assign new_n1698 = in0126 & ~new_n1167;
  assign new_n1699 = in1126 & new_n1167;
  assign new_n1700 = ~new_n1698 & ~new_n1699;
  assign new_n1701 = new_n1697 & ~new_n1700;
  assign new_n1702 = ~new_n1697 & new_n1700;
  assign new_n1703 = in2125 & ~new_n1694;
  assign new_n1704 = in3125 & new_n1694;
  assign new_n1705 = ~new_n1703 & ~new_n1704;
  assign new_n1706 = in0125 & ~new_n1167;
  assign new_n1707 = in1125 & new_n1167;
  assign new_n1708 = ~new_n1706 & ~new_n1707;
  assign new_n1709 = ~new_n1705 & new_n1708;
  assign new_n1710 = ~new_n1702 & ~new_n1709;
  assign new_n1711 = in2124 & ~new_n1694;
  assign new_n1712 = in3124 & new_n1694;
  assign new_n1713 = ~new_n1711 & ~new_n1712;
  assign new_n1714 = in0124 & ~new_n1167;
  assign new_n1715 = in1124 & new_n1167;
  assign new_n1716 = ~new_n1714 & ~new_n1715;
  assign new_n1717 = new_n1713 & ~new_n1716;
  assign new_n1718 = new_n1705 & ~new_n1708;
  assign new_n1719 = ~new_n1717 & ~new_n1718;
  assign new_n1720 = new_n1710 & ~new_n1719;
  assign new_n1721 = ~new_n1713 & new_n1716;
  assign new_n1722 = in2123 & ~new_n1694;
  assign new_n1723 = in3123 & new_n1694;
  assign new_n1724 = ~new_n1722 & ~new_n1723;
  assign new_n1725 = in0123 & ~new_n1167;
  assign new_n1726 = in1123 & new_n1167;
  assign new_n1727 = ~new_n1725 & ~new_n1726;
  assign new_n1728 = new_n1724 & ~new_n1727;
  assign new_n1729 = in2122 & ~new_n1694;
  assign new_n1730 = in3122 & new_n1694;
  assign new_n1731 = ~new_n1729 & ~new_n1730;
  assign new_n1732 = in0122 & ~new_n1167;
  assign new_n1733 = in1122 & new_n1167;
  assign new_n1734 = ~new_n1732 & ~new_n1733;
  assign new_n1735 = new_n1731 & ~new_n1734;
  assign new_n1736 = in2121 & ~new_n1694;
  assign new_n1737 = in3121 & new_n1694;
  assign new_n1738 = ~new_n1736 & ~new_n1737;
  assign new_n1739 = in0121 & ~new_n1167;
  assign new_n1740 = in1121 & new_n1167;
  assign new_n1741 = ~new_n1739 & ~new_n1740;
  assign new_n1742 = ~new_n1738 & new_n1741;
  assign new_n1743 = new_n1738 & ~new_n1741;
  assign new_n1744 = in0117 & ~new_n1167;
  assign new_n1745 = in1117 & new_n1167;
  assign new_n1746 = ~new_n1744 & ~new_n1745;
  assign new_n1747 = in2117 & ~new_n1694;
  assign new_n1748 = in3117 & new_n1694;
  assign new_n1749 = ~new_n1747 & ~new_n1748;
  assign new_n1750 = new_n1746 & ~new_n1749;
  assign new_n1751 = in2116 & ~new_n1694;
  assign new_n1752 = in3116 & new_n1694;
  assign new_n1753 = ~new_n1751 & ~new_n1752;
  assign new_n1754 = in0116 & ~new_n1167;
  assign new_n1755 = in1116 & new_n1167;
  assign new_n1756 = ~new_n1754 & ~new_n1755;
  assign new_n1757 = new_n1753 & ~new_n1756;
  assign new_n1758 = ~new_n1746 & new_n1749;
  assign new_n1759 = ~new_n1753 & new_n1756;
  assign new_n1760 = in2115 & ~new_n1694;
  assign new_n1761 = in3115 & new_n1694;
  assign new_n1762 = ~new_n1760 & ~new_n1761;
  assign new_n1763 = in0115 & ~new_n1167;
  assign new_n1764 = in1115 & new_n1167;
  assign new_n1765 = ~new_n1763 & ~new_n1764;
  assign new_n1766 = ~new_n1762 & new_n1765;
  assign new_n1767 = in2114 & ~new_n1694;
  assign new_n1768 = in3114 & new_n1694;
  assign new_n1769 = ~new_n1767 & ~new_n1768;
  assign new_n1770 = in0114 & ~new_n1167;
  assign new_n1771 = in1114 & new_n1167;
  assign new_n1772 = ~new_n1770 & ~new_n1771;
  assign new_n1773 = new_n1769 & ~new_n1772;
  assign new_n1774 = new_n1762 & ~new_n1765;
  assign new_n1775 = ~new_n1769 & new_n1772;
  assign new_n1776 = in2113 & ~new_n1694;
  assign new_n1777 = in3113 & new_n1694;
  assign new_n1778 = ~new_n1776 & ~new_n1777;
  assign new_n1779 = in0113 & ~new_n1167;
  assign new_n1780 = in1113 & new_n1167;
  assign new_n1781 = ~new_n1779 & ~new_n1780;
  assign new_n1782 = new_n1778 & ~new_n1781;
  assign new_n1783 = in0109 & ~new_n1167;
  assign new_n1784 = in1109 & new_n1167;
  assign new_n1785 = ~new_n1783 & ~new_n1784;
  assign new_n1786 = in2109 & ~new_n1694;
  assign new_n1787 = in3109 & new_n1694;
  assign new_n1788 = ~new_n1786 & ~new_n1787;
  assign new_n1789 = new_n1785 & ~new_n1788;
  assign new_n1790 = in2108 & ~new_n1694;
  assign new_n1791 = in3108 & new_n1694;
  assign new_n1792 = ~new_n1790 & ~new_n1791;
  assign new_n1793 = in0108 & ~new_n1167;
  assign new_n1794 = in1108 & new_n1167;
  assign new_n1795 = ~new_n1793 & ~new_n1794;
  assign new_n1796 = new_n1792 & ~new_n1795;
  assign new_n1797 = ~new_n1785 & new_n1788;
  assign new_n1798 = ~new_n1792 & new_n1795;
  assign new_n1799 = in0107 & ~new_n1167;
  assign new_n1800 = in1107 & new_n1167;
  assign new_n1801 = ~new_n1799 & ~new_n1800;
  assign new_n1802 = in2107 & ~new_n1694;
  assign new_n1803 = in3107 & new_n1694;
  assign new_n1804 = ~new_n1802 & ~new_n1803;
  assign new_n1805 = new_n1801 & ~new_n1804;
  assign new_n1806 = in2106 & ~new_n1694;
  assign new_n1807 = in3106 & new_n1694;
  assign new_n1808 = ~new_n1806 & ~new_n1807;
  assign new_n1809 = in0106 & ~new_n1167;
  assign new_n1810 = in1106 & new_n1167;
  assign new_n1811 = ~new_n1809 & ~new_n1810;
  assign new_n1812 = new_n1808 & ~new_n1811;
  assign new_n1813 = ~new_n1801 & new_n1804;
  assign new_n1814 = ~new_n1808 & new_n1811;
  assign new_n1815 = in0105 & ~new_n1167;
  assign new_n1816 = in1105 & new_n1167;
  assign new_n1817 = ~new_n1815 & ~new_n1816;
  assign new_n1818 = in2105 & ~new_n1694;
  assign new_n1819 = in3105 & new_n1694;
  assign new_n1820 = ~new_n1818 & ~new_n1819;
  assign new_n1821 = new_n1817 & ~new_n1820;
  assign new_n1822 = in2104 & ~new_n1694;
  assign new_n1823 = in3104 & new_n1694;
  assign new_n1824 = ~new_n1822 & ~new_n1823;
  assign new_n1825 = in0104 & ~new_n1167;
  assign new_n1826 = in1104 & new_n1167;
  assign new_n1827 = ~new_n1825 & ~new_n1826;
  assign new_n1828 = new_n1824 & ~new_n1827;
  assign new_n1829 = ~new_n1817 & new_n1820;
  assign new_n1830 = ~new_n1824 & new_n1827;
  assign new_n1831 = in0103 & ~new_n1167;
  assign new_n1832 = in1103 & new_n1167;
  assign new_n1833 = ~new_n1831 & ~new_n1832;
  assign new_n1834 = in2103 & ~new_n1694;
  assign new_n1835 = in3103 & new_n1694;
  assign new_n1836 = ~new_n1834 & ~new_n1835;
  assign new_n1837 = new_n1833 & ~new_n1836;
  assign new_n1838 = in2102 & ~new_n1694;
  assign new_n1839 = in3102 & new_n1694;
  assign new_n1840 = ~new_n1838 & ~new_n1839;
  assign new_n1841 = in0102 & ~new_n1167;
  assign new_n1842 = in1102 & new_n1167;
  assign new_n1843 = ~new_n1841 & ~new_n1842;
  assign new_n1844 = new_n1840 & ~new_n1843;
  assign new_n1845 = ~new_n1833 & new_n1836;
  assign new_n1846 = ~new_n1840 & new_n1843;
  assign new_n1847 = in2101 & ~new_n1694;
  assign new_n1848 = in3101 & new_n1694;
  assign new_n1849 = ~new_n1847 & ~new_n1848;
  assign new_n1850 = in0101 & ~new_n1167;
  assign new_n1851 = in1101 & new_n1167;
  assign new_n1852 = ~new_n1850 & ~new_n1851;
  assign new_n1853 = ~new_n1849 & new_n1852;
  assign new_n1854 = in0100 & ~new_n1167;
  assign new_n1855 = in1100 & new_n1167;
  assign new_n1856 = ~new_n1854 & ~new_n1855;
  assign new_n1857 = in2100 & ~new_n1694;
  assign new_n1858 = in3100 & new_n1694;
  assign new_n1859 = ~new_n1857 & ~new_n1858;
  assign new_n1860 = ~new_n1856 & new_n1859;
  assign new_n1861 = new_n1849 & ~new_n1852;
  assign new_n1862 = new_n1856 & ~new_n1859;
  assign new_n1863 = in099 & ~new_n1167;
  assign new_n1864 = in199 & new_n1167;
  assign new_n1865 = ~new_n1863 & ~new_n1864;
  assign new_n1866 = in299 & ~new_n1694;
  assign new_n1867 = in399 & new_n1694;
  assign new_n1868 = ~new_n1866 & ~new_n1867;
  assign new_n1869 = ~new_n1865 & new_n1868;
  assign new_n1870 = new_n1865 & ~new_n1868;
  assign new_n1871 = in298 & ~new_n1694;
  assign new_n1872 = in398 & new_n1694;
  assign new_n1873 = ~new_n1871 & ~new_n1872;
  assign new_n1874 = in098 & ~new_n1167;
  assign new_n1875 = in198 & new_n1167;
  assign new_n1876 = ~new_n1874 & ~new_n1875;
  assign new_n1877 = new_n1873 & ~new_n1876;
  assign new_n1878 = in297 & ~new_n1694;
  assign new_n1879 = in397 & new_n1694;
  assign new_n1880 = ~new_n1878 & ~new_n1879;
  assign new_n1881 = in097 & ~new_n1167;
  assign new_n1882 = in197 & new_n1167;
  assign new_n1883 = ~new_n1881 & ~new_n1882;
  assign new_n1884 = ~new_n1880 & new_n1883;
  assign new_n1885 = ~new_n1873 & new_n1876;
  assign new_n1886 = new_n1880 & ~new_n1883;
  assign new_n1887 = in296 & ~new_n1694;
  assign new_n1888 = in396 & new_n1694;
  assign new_n1889 = ~new_n1887 & ~new_n1888;
  assign new_n1890 = in096 & ~new_n1167;
  assign new_n1891 = in196 & new_n1167;
  assign new_n1892 = ~new_n1890 & ~new_n1891;
  assign new_n1893 = ~new_n1889 & new_n1892;
  assign new_n1894 = new_n1889 & ~new_n1892;
  assign new_n1895 = in295 & ~new_n1694;
  assign new_n1896 = in395 & new_n1694;
  assign new_n1897 = ~new_n1895 & ~new_n1896;
  assign new_n1898 = in095 & ~new_n1167;
  assign new_n1899 = in195 & new_n1167;
  assign new_n1900 = ~new_n1898 & ~new_n1899;
  assign new_n1901 = ~new_n1897 & new_n1900;
  assign new_n1902 = new_n1897 & ~new_n1900;
  assign new_n1903 = in094 & ~new_n1167;
  assign new_n1904 = in194 & new_n1167;
  assign new_n1905 = ~new_n1903 & ~new_n1904;
  assign new_n1906 = in294 & ~new_n1694;
  assign new_n1907 = in394 & new_n1694;
  assign new_n1908 = ~new_n1906 & ~new_n1907;
  assign new_n1909 = new_n1905 & ~new_n1908;
  assign new_n1910 = ~new_n1905 & new_n1908;
  assign new_n1911 = in093 & ~new_n1167;
  assign new_n1912 = in193 & new_n1167;
  assign new_n1913 = ~new_n1911 & ~new_n1912;
  assign new_n1914 = in293 & ~new_n1694;
  assign new_n1915 = in393 & new_n1694;
  assign new_n1916 = ~new_n1914 & ~new_n1915;
  assign new_n1917 = new_n1913 & ~new_n1916;
  assign new_n1918 = ~new_n1913 & new_n1916;
  assign new_n1919 = in292 & ~new_n1694;
  assign new_n1920 = in392 & new_n1694;
  assign new_n1921 = ~new_n1919 & ~new_n1920;
  assign new_n1922 = in092 & ~new_n1167;
  assign new_n1923 = in192 & new_n1167;
  assign new_n1924 = ~new_n1922 & ~new_n1923;
  assign new_n1925 = ~new_n1921 & new_n1924;
  assign new_n1926 = in291 & ~new_n1694;
  assign new_n1927 = in391 & new_n1694;
  assign new_n1928 = ~new_n1926 & ~new_n1927;
  assign new_n1929 = in091 & ~new_n1167;
  assign new_n1930 = in191 & new_n1167;
  assign new_n1931 = ~new_n1929 & ~new_n1930;
  assign new_n1932 = new_n1928 & ~new_n1931;
  assign new_n1933 = new_n1921 & ~new_n1924;
  assign new_n1934 = ~new_n1928 & new_n1931;
  assign new_n1935 = in290 & ~new_n1694;
  assign new_n1936 = in390 & new_n1694;
  assign new_n1937 = ~new_n1935 & ~new_n1936;
  assign new_n1938 = in090 & ~new_n1167;
  assign new_n1939 = in190 & new_n1167;
  assign new_n1940 = ~new_n1938 & ~new_n1939;
  assign new_n1941 = new_n1937 & ~new_n1940;
  assign new_n1942 = ~new_n1937 & new_n1940;
  assign new_n1943 = in089 & ~new_n1167;
  assign new_n1944 = in189 & new_n1167;
  assign new_n1945 = ~new_n1943 & ~new_n1944;
  assign new_n1946 = in289 & ~new_n1694;
  assign new_n1947 = in389 & new_n1694;
  assign new_n1948 = ~new_n1946 & ~new_n1947;
  assign new_n1949 = ~new_n1945 & new_n1948;
  assign new_n1950 = new_n1945 & ~new_n1948;
  assign new_n1951 = in088 & ~new_n1167;
  assign new_n1952 = in188 & new_n1167;
  assign new_n1953 = ~new_n1951 & ~new_n1952;
  assign new_n1954 = in288 & ~new_n1694;
  assign new_n1955 = in388 & new_n1694;
  assign new_n1956 = ~new_n1954 & ~new_n1955;
  assign new_n1957 = ~new_n1953 & new_n1956;
  assign new_n1958 = new_n1953 & ~new_n1956;
  assign new_n1959 = in087 & ~new_n1167;
  assign new_n1960 = in187 & new_n1167;
  assign new_n1961 = ~new_n1959 & ~new_n1960;
  assign new_n1962 = in287 & ~new_n1694;
  assign new_n1963 = in387 & new_n1694;
  assign new_n1964 = ~new_n1962 & ~new_n1963;
  assign new_n1965 = ~new_n1961 & new_n1964;
  assign new_n1966 = new_n1961 & ~new_n1964;
  assign new_n1967 = in086 & ~new_n1167;
  assign new_n1968 = in186 & new_n1167;
  assign new_n1969 = ~new_n1967 & ~new_n1968;
  assign new_n1970 = in286 & ~new_n1694;
  assign new_n1971 = in386 & new_n1694;
  assign new_n1972 = ~new_n1970 & ~new_n1971;
  assign new_n1973 = ~new_n1969 & new_n1972;
  assign new_n1974 = in085 & ~new_n1167;
  assign new_n1975 = in185 & new_n1167;
  assign new_n1976 = ~new_n1974 & ~new_n1975;
  assign new_n1977 = in285 & ~new_n1694;
  assign new_n1978 = in385 & new_n1694;
  assign new_n1979 = ~new_n1977 & ~new_n1978;
  assign new_n1980 = new_n1976 & ~new_n1979;
  assign new_n1981 = new_n1969 & ~new_n1972;
  assign new_n1982 = ~new_n1976 & new_n1979;
  assign new_n1983 = in084 & ~new_n1167;
  assign new_n1984 = in184 & new_n1167;
  assign new_n1985 = ~new_n1983 & ~new_n1984;
  assign new_n1986 = in284 & ~new_n1694;
  assign new_n1987 = in384 & new_n1694;
  assign new_n1988 = ~new_n1986 & ~new_n1987;
  assign new_n1989 = new_n1985 & ~new_n1988;
  assign new_n1990 = in083 & ~new_n1167;
  assign new_n1991 = in183 & new_n1167;
  assign new_n1992 = ~new_n1990 & ~new_n1991;
  assign new_n1993 = in283 & ~new_n1694;
  assign new_n1994 = in383 & new_n1694;
  assign new_n1995 = ~new_n1993 & ~new_n1994;
  assign new_n1996 = ~new_n1992 & new_n1995;
  assign new_n1997 = ~new_n1985 & new_n1988;
  assign new_n1998 = in282 & ~new_n1694;
  assign new_n1999 = in382 & new_n1694;
  assign new_n2000 = ~new_n1998 & ~new_n1999;
  assign new_n2001 = in082 & ~new_n1167;
  assign new_n2002 = in182 & new_n1167;
  assign new_n2003 = ~new_n2001 & ~new_n2002;
  assign new_n2004 = ~new_n2000 & new_n2003;
  assign new_n2005 = new_n1992 & ~new_n1995;
  assign new_n2006 = new_n2000 & ~new_n2003;
  assign new_n2007 = in281 & ~new_n1694;
  assign new_n2008 = in381 & new_n1694;
  assign new_n2009 = ~new_n2007 & ~new_n2008;
  assign new_n2010 = in081 & ~new_n1167;
  assign new_n2011 = in181 & new_n1167;
  assign new_n2012 = ~new_n2010 & ~new_n2011;
  assign new_n2013 = new_n2009 & ~new_n2012;
  assign new_n2014 = ~new_n2009 & new_n2012;
  assign new_n2015 = in080 & ~new_n1167;
  assign new_n2016 = in180 & new_n1167;
  assign new_n2017 = ~new_n2015 & ~new_n2016;
  assign new_n2018 = in280 & ~new_n1694;
  assign new_n2019 = in380 & new_n1694;
  assign new_n2020 = ~new_n2018 & ~new_n2019;
  assign new_n2021 = new_n2017 & ~new_n2020;
  assign new_n2022 = ~new_n2017 & new_n2020;
  assign new_n2023 = in279 & ~new_n1694;
  assign new_n2024 = in379 & new_n1694;
  assign new_n2025 = ~new_n2023 & ~new_n2024;
  assign new_n2026 = in079 & ~new_n1167;
  assign new_n2027 = in179 & new_n1167;
  assign new_n2028 = ~new_n2026 & ~new_n2027;
  assign new_n2029 = new_n2025 & ~new_n2028;
  assign new_n2030 = in278 & ~new_n1694;
  assign new_n2031 = in378 & new_n1694;
  assign new_n2032 = ~new_n2030 & ~new_n2031;
  assign new_n2033 = in078 & ~new_n1167;
  assign new_n2034 = in178 & new_n1167;
  assign new_n2035 = ~new_n2033 & ~new_n2034;
  assign new_n2036 = ~new_n2032 & new_n2035;
  assign new_n2037 = ~new_n2025 & new_n2028;
  assign new_n2038 = new_n2032 & ~new_n2035;
  assign new_n2039 = in077 & ~new_n1167;
  assign new_n2040 = in177 & new_n1167;
  assign new_n2041 = ~new_n2039 & ~new_n2040;
  assign new_n2042 = in277 & ~new_n1694;
  assign new_n2043 = in377 & new_n1694;
  assign new_n2044 = ~new_n2042 & ~new_n2043;
  assign new_n2045 = new_n2041 & ~new_n2044;
  assign new_n2046 = ~new_n2041 & new_n2044;
  assign new_n2047 = in276 & ~new_n1694;
  assign new_n2048 = in376 & new_n1694;
  assign new_n2049 = ~new_n2047 & ~new_n2048;
  assign new_n2050 = in076 & ~new_n1167;
  assign new_n2051 = in176 & new_n1167;
  assign new_n2052 = ~new_n2050 & ~new_n2051;
  assign new_n2053 = ~new_n2049 & new_n2052;
  assign new_n2054 = new_n2049 & ~new_n2052;
  assign new_n2055 = in075 & ~new_n1167;
  assign new_n2056 = in175 & new_n1167;
  assign new_n2057 = ~new_n2055 & ~new_n2056;
  assign new_n2058 = in275 & ~new_n1694;
  assign new_n2059 = in375 & new_n1694;
  assign new_n2060 = ~new_n2058 & ~new_n2059;
  assign new_n2061 = ~new_n2057 & new_n2060;
  assign new_n2062 = in274 & ~new_n1694;
  assign new_n2063 = in374 & new_n1694;
  assign new_n2064 = ~new_n2062 & ~new_n2063;
  assign new_n2065 = in074 & ~new_n1167;
  assign new_n2066 = in174 & new_n1167;
  assign new_n2067 = ~new_n2065 & ~new_n2066;
  assign new_n2068 = ~new_n2064 & new_n2067;
  assign new_n2069 = new_n2057 & ~new_n2060;
  assign new_n2070 = new_n2064 & ~new_n2067;
  assign new_n2071 = in273 & ~new_n1694;
  assign new_n2072 = in373 & new_n1694;
  assign new_n2073 = ~new_n2071 & ~new_n2072;
  assign new_n2074 = in073 & ~new_n1167;
  assign new_n2075 = in173 & new_n1167;
  assign new_n2076 = ~new_n2074 & ~new_n2075;
  assign new_n2077 = new_n2073 & ~new_n2076;
  assign new_n2078 = ~new_n2073 & new_n2076;
  assign new_n2079 = in072 & ~new_n1167;
  assign new_n2080 = in172 & new_n1167;
  assign new_n2081 = ~new_n2079 & ~new_n2080;
  assign new_n2082 = in272 & ~new_n1694;
  assign new_n2083 = in372 & new_n1694;
  assign new_n2084 = ~new_n2082 & ~new_n2083;
  assign new_n2085 = new_n2081 & ~new_n2084;
  assign new_n2086 = ~new_n2081 & new_n2084;
  assign new_n2087 = in271 & ~new_n1694;
  assign new_n2088 = in371 & new_n1694;
  assign new_n2089 = ~new_n2087 & ~new_n2088;
  assign new_n2090 = in071 & ~new_n1167;
  assign new_n2091 = in171 & new_n1167;
  assign new_n2092 = ~new_n2090 & ~new_n2091;
  assign new_n2093 = new_n2089 & ~new_n2092;
  assign new_n2094 = in270 & ~new_n1694;
  assign new_n2095 = in370 & new_n1694;
  assign new_n2096 = ~new_n2094 & ~new_n2095;
  assign new_n2097 = in070 & ~new_n1167;
  assign new_n2098 = in170 & new_n1167;
  assign new_n2099 = ~new_n2097 & ~new_n2098;
  assign new_n2100 = ~new_n2096 & new_n2099;
  assign new_n2101 = ~new_n2089 & new_n2092;
  assign new_n2102 = new_n2096 & ~new_n2099;
  assign new_n2103 = in069 & ~new_n1167;
  assign new_n2104 = in169 & new_n1167;
  assign new_n2105 = ~new_n2103 & ~new_n2104;
  assign new_n2106 = in269 & ~new_n1694;
  assign new_n2107 = in369 & new_n1694;
  assign new_n2108 = ~new_n2106 & ~new_n2107;
  assign new_n2109 = new_n2105 & ~new_n2108;
  assign new_n2110 = ~new_n2105 & new_n2108;
  assign new_n2111 = in068 & ~new_n1167;
  assign new_n2112 = in168 & new_n1167;
  assign new_n2113 = ~new_n2111 & ~new_n2112;
  assign new_n2114 = in268 & ~new_n1694;
  assign new_n2115 = in368 & new_n1694;
  assign new_n2116 = ~new_n2114 & ~new_n2115;
  assign new_n2117 = new_n2113 & ~new_n2116;
  assign new_n2118 = ~new_n2113 & new_n2116;
  assign new_n2119 = in067 & ~new_n1167;
  assign new_n2120 = in167 & new_n1167;
  assign new_n2121 = ~new_n2119 & ~new_n2120;
  assign new_n2122 = in267 & ~new_n1694;
  assign new_n2123 = in367 & new_n1694;
  assign new_n2124 = ~new_n2122 & ~new_n2123;
  assign new_n2125 = new_n2121 & ~new_n2124;
  assign new_n2126 = in066 & ~new_n1167;
  assign new_n2127 = in166 & new_n1167;
  assign new_n2128 = ~new_n2126 & ~new_n2127;
  assign new_n2129 = in266 & ~new_n1694;
  assign new_n2130 = in366 & new_n1694;
  assign new_n2131 = ~new_n2129 & ~new_n2130;
  assign new_n2132 = ~new_n2128 & new_n2131;
  assign new_n2133 = ~new_n2121 & new_n2124;
  assign new_n2134 = new_n2128 & ~new_n2131;
  assign new_n2135 = in065 & ~new_n1167;
  assign new_n2136 = in165 & new_n1167;
  assign new_n2137 = ~new_n2135 & ~new_n2136;
  assign new_n2138 = in265 & ~new_n1694;
  assign new_n2139 = in365 & new_n1694;
  assign new_n2140 = ~new_n2138 & ~new_n2139;
  assign new_n2141 = ~new_n2137 & new_n2140;
  assign new_n2142 = new_n2137 & ~new_n2140;
  assign new_n2143 = in064 & ~new_n1167;
  assign new_n2144 = in164 & new_n1167;
  assign new_n2145 = ~new_n2143 & ~new_n2144;
  assign new_n2146 = in264 & ~new_n1694;
  assign new_n2147 = in364 & new_n1694;
  assign new_n2148 = ~new_n2146 & ~new_n2147;
  assign new_n2149 = ~new_n2145 & new_n2148;
  assign new_n2150 = new_n2145 & ~new_n2148;
  assign new_n2151 = in263 & ~new_n1694;
  assign new_n2152 = in363 & new_n1694;
  assign new_n2153 = ~new_n2151 & ~new_n2152;
  assign new_n2154 = in063 & ~new_n1167;
  assign new_n2155 = in163 & new_n1167;
  assign new_n2156 = ~new_n2154 & ~new_n2155;
  assign new_n2157 = new_n2153 & ~new_n2156;
  assign new_n2158 = in262 & ~new_n1694;
  assign new_n2159 = in362 & new_n1694;
  assign new_n2160 = ~new_n2158 & ~new_n2159;
  assign new_n2161 = in062 & ~new_n1167;
  assign new_n2162 = in162 & new_n1167;
  assign new_n2163 = ~new_n2161 & ~new_n2162;
  assign new_n2164 = ~new_n2160 & new_n2163;
  assign new_n2165 = ~new_n2153 & new_n2156;
  assign new_n2166 = new_n2160 & ~new_n2163;
  assign new_n2167 = in261 & ~new_n1694;
  assign new_n2168 = in361 & new_n1694;
  assign new_n2169 = ~new_n2167 & ~new_n2168;
  assign new_n2170 = in061 & ~new_n1167;
  assign new_n2171 = in161 & new_n1167;
  assign new_n2172 = ~new_n2170 & ~new_n2171;
  assign new_n2173 = ~new_n2169 & new_n2172;
  assign new_n2174 = new_n2169 & ~new_n2172;
  assign new_n2175 = in256 & ~new_n1694;
  assign new_n2176 = in356 & new_n1694;
  assign new_n2177 = ~new_n2175 & ~new_n2176;
  assign new_n2178 = in056 & ~new_n1167;
  assign new_n2179 = in156 & new_n1167;
  assign new_n2180 = ~new_n2178 & ~new_n2179;
  assign new_n2181 = ~new_n2177 & new_n2180;
  assign new_n2182 = in254 & ~new_n1694;
  assign new_n2183 = in354 & new_n1694;
  assign new_n2184 = ~new_n2182 & ~new_n2183;
  assign new_n2185 = in054 & ~new_n1167;
  assign new_n2186 = in154 & new_n1167;
  assign new_n2187 = ~new_n2185 & ~new_n2186;
  assign new_n2188 = new_n2184 & ~new_n2187;
  assign new_n2189 = in055 & ~new_n1167;
  assign new_n2190 = in155 & new_n1167;
  assign new_n2191 = ~new_n2189 & ~new_n2190;
  assign new_n2192 = in255 & ~new_n1694;
  assign new_n2193 = in355 & new_n1694;
  assign new_n2194 = ~new_n2192 & ~new_n2193;
  assign new_n2195 = ~new_n2191 & new_n2194;
  assign new_n2196 = ~new_n2184 & new_n2187;
  assign new_n2197 = in253 & ~new_n1694;
  assign new_n2198 = in353 & new_n1694;
  assign new_n2199 = ~new_n2197 & ~new_n2198;
  assign new_n2200 = in053 & ~new_n1167;
  assign new_n2201 = in153 & new_n1167;
  assign new_n2202 = ~new_n2200 & ~new_n2201;
  assign new_n2203 = ~new_n2199 & new_n2202;
  assign new_n2204 = in052 & ~new_n1167;
  assign new_n2205 = in152 & new_n1167;
  assign new_n2206 = ~new_n2204 & ~new_n2205;
  assign new_n2207 = in252 & ~new_n1694;
  assign new_n2208 = in352 & new_n1694;
  assign new_n2209 = ~new_n2207 & ~new_n2208;
  assign new_n2210 = ~new_n2206 & new_n2209;
  assign new_n2211 = in247 & ~new_n1694;
  assign new_n2212 = in347 & new_n1694;
  assign new_n2213 = ~new_n2211 & ~new_n2212;
  assign new_n2214 = in047 & ~new_n1167;
  assign new_n2215 = in147 & new_n1167;
  assign new_n2216 = ~new_n2214 & ~new_n2215;
  assign new_n2217 = new_n2213 & ~new_n2216;
  assign new_n2218 = in046 & ~new_n1167;
  assign new_n2219 = in146 & new_n1167;
  assign new_n2220 = ~new_n2218 & ~new_n2219;
  assign new_n2221 = in246 & ~new_n1694;
  assign new_n2222 = in346 & new_n1694;
  assign new_n2223 = ~new_n2221 & ~new_n2222;
  assign new_n2224 = ~new_n2220 & new_n2223;
  assign new_n2225 = in045 & ~new_n1167;
  assign new_n2226 = in145 & new_n1167;
  assign new_n2227 = ~new_n2225 & ~new_n2226;
  assign new_n2228 = in245 & ~new_n1694;
  assign new_n2229 = in345 & new_n1694;
  assign new_n2230 = ~new_n2228 & ~new_n2229;
  assign new_n2231 = new_n2227 & ~new_n2230;
  assign new_n2232 = new_n2220 & ~new_n2223;
  assign new_n2233 = ~new_n2227 & new_n2230;
  assign new_n2234 = in240 & ~new_n1694;
  assign new_n2235 = in340 & new_n1694;
  assign new_n2236 = ~new_n2234 & ~new_n2235;
  assign new_n2237 = in040 & ~new_n1167;
  assign new_n2238 = in140 & new_n1167;
  assign new_n2239 = ~new_n2237 & ~new_n2238;
  assign new_n2240 = ~new_n2236 & new_n2239;
  assign new_n2241 = in038 & ~new_n1167;
  assign new_n2242 = in138 & new_n1167;
  assign new_n2243 = ~new_n2241 & ~new_n2242;
  assign new_n2244 = in238 & ~new_n1694;
  assign new_n2245 = in338 & new_n1694;
  assign new_n2246 = ~new_n2244 & ~new_n2245;
  assign new_n2247 = ~new_n2243 & new_n2246;
  assign new_n2248 = in232 & ~new_n1694;
  assign new_n2249 = in332 & new_n1694;
  assign new_n2250 = ~new_n2248 & ~new_n2249;
  assign new_n2251 = in032 & ~new_n1167;
  assign new_n2252 = in132 & new_n1167;
  assign new_n2253 = ~new_n2251 & ~new_n2252;
  assign new_n2254 = ~new_n2250 & new_n2253;
  assign new_n2255 = in031 & ~new_n1167;
  assign new_n2256 = in131 & new_n1167;
  assign new_n2257 = ~new_n2255 & ~new_n2256;
  assign new_n2258 = in231 & ~new_n1694;
  assign new_n2259 = in331 & new_n1694;
  assign new_n2260 = ~new_n2258 & ~new_n2259;
  assign new_n2261 = ~new_n2257 & new_n2260;
  assign new_n2262 = in030 & ~new_n1167;
  assign new_n2263 = in130 & new_n1167;
  assign new_n2264 = ~new_n2262 & ~new_n2263;
  assign new_n2265 = in230 & ~new_n1694;
  assign new_n2266 = in330 & new_n1694;
  assign new_n2267 = ~new_n2265 & ~new_n2266;
  assign new_n2268 = ~new_n2264 & new_n2267;
  assign new_n2269 = in229 & ~new_n1694;
  assign new_n2270 = in329 & new_n1694;
  assign new_n2271 = ~new_n2269 & ~new_n2270;
  assign new_n2272 = in029 & ~new_n1167;
  assign new_n2273 = in129 & new_n1167;
  assign new_n2274 = ~new_n2272 & ~new_n2273;
  assign new_n2275 = ~new_n2271 & new_n2274;
  assign new_n2276 = new_n2264 & ~new_n2267;
  assign new_n2277 = new_n2271 & ~new_n2274;
  assign new_n2278 = in028 & ~new_n1167;
  assign new_n2279 = in128 & new_n1167;
  assign new_n2280 = ~new_n2278 & ~new_n2279;
  assign new_n2281 = in228 & ~new_n1694;
  assign new_n2282 = in328 & new_n1694;
  assign new_n2283 = ~new_n2281 & ~new_n2282;
  assign new_n2284 = ~new_n2280 & new_n2283;
  assign new_n2285 = in227 & ~new_n1694;
  assign new_n2286 = in327 & new_n1694;
  assign new_n2287 = ~new_n2285 & ~new_n2286;
  assign new_n2288 = in027 & ~new_n1167;
  assign new_n2289 = in127 & new_n1167;
  assign new_n2290 = ~new_n2288 & ~new_n2289;
  assign new_n2291 = ~new_n2287 & new_n2290;
  assign new_n2292 = new_n2280 & ~new_n2283;
  assign new_n2293 = new_n2287 & ~new_n2290;
  assign new_n2294 = in026 & ~new_n1167;
  assign new_n2295 = in126 & new_n1167;
  assign new_n2296 = ~new_n2294 & ~new_n2295;
  assign new_n2297 = in226 & ~new_n1694;
  assign new_n2298 = in326 & new_n1694;
  assign new_n2299 = ~new_n2297 & ~new_n2298;
  assign new_n2300 = ~new_n2296 & new_n2299;
  assign new_n2301 = in225 & ~new_n1694;
  assign new_n2302 = in325 & new_n1694;
  assign new_n2303 = ~new_n2301 & ~new_n2302;
  assign new_n2304 = in025 & ~new_n1167;
  assign new_n2305 = in125 & new_n1167;
  assign new_n2306 = ~new_n2304 & ~new_n2305;
  assign new_n2307 = ~new_n2303 & new_n2306;
  assign new_n2308 = new_n2296 & ~new_n2299;
  assign new_n2309 = new_n2303 & ~new_n2306;
  assign new_n2310 = in024 & ~new_n1167;
  assign new_n2311 = in124 & new_n1167;
  assign new_n2312 = ~new_n2310 & ~new_n2311;
  assign new_n2313 = in224 & ~new_n1694;
  assign new_n2314 = in324 & new_n1694;
  assign new_n2315 = ~new_n2313 & ~new_n2314;
  assign new_n2316 = ~new_n2312 & new_n2315;
  assign new_n2317 = in223 & ~new_n1694;
  assign new_n2318 = in323 & new_n1694;
  assign new_n2319 = ~new_n2317 & ~new_n2318;
  assign new_n2320 = in023 & ~new_n1167;
  assign new_n2321 = in123 & new_n1167;
  assign new_n2322 = ~new_n2320 & ~new_n2321;
  assign new_n2323 = ~new_n2319 & new_n2322;
  assign new_n2324 = new_n2312 & ~new_n2315;
  assign new_n2325 = new_n2319 & ~new_n2322;
  assign new_n2326 = in222 & ~new_n1694;
  assign new_n2327 = in322 & new_n1694;
  assign new_n2328 = ~new_n2326 & ~new_n2327;
  assign new_n2329 = in022 & ~new_n1167;
  assign new_n2330 = in122 & new_n1167;
  assign new_n2331 = ~new_n2329 & ~new_n2330;
  assign new_n2332 = new_n2328 & ~new_n2331;
  assign new_n2333 = ~new_n2328 & new_n2331;
  assign new_n2334 = in221 & ~new_n1694;
  assign new_n2335 = in321 & new_n1694;
  assign new_n2336 = ~new_n2334 & ~new_n2335;
  assign new_n2337 = in021 & ~new_n1167;
  assign new_n2338 = in121 & new_n1167;
  assign new_n2339 = ~new_n2337 & ~new_n2338;
  assign new_n2340 = ~new_n2336 & new_n2339;
  assign new_n2341 = in220 & ~new_n1694;
  assign new_n2342 = in320 & new_n1694;
  assign new_n2343 = ~new_n2341 & ~new_n2342;
  assign new_n2344 = in020 & ~new_n1167;
  assign new_n2345 = in120 & new_n1167;
  assign new_n2346 = ~new_n2344 & ~new_n2345;
  assign new_n2347 = new_n2343 & ~new_n2346;
  assign new_n2348 = new_n2336 & ~new_n2339;
  assign new_n2349 = ~new_n2343 & new_n2346;
  assign new_n2350 = in219 & ~new_n1694;
  assign new_n2351 = in319 & new_n1694;
  assign new_n2352 = ~new_n2350 & ~new_n2351;
  assign new_n2353 = in019 & ~new_n1167;
  assign new_n2354 = in119 & new_n1167;
  assign new_n2355 = ~new_n2353 & ~new_n2354;
  assign new_n2356 = new_n2352 & ~new_n2355;
  assign new_n2357 = ~new_n2352 & new_n2355;
  assign new_n2358 = in218 & ~new_n1694;
  assign new_n2359 = in318 & new_n1694;
  assign new_n2360 = ~new_n2358 & ~new_n2359;
  assign new_n2361 = in018 & ~new_n1167;
  assign new_n2362 = in118 & new_n1167;
  assign new_n2363 = ~new_n2361 & ~new_n2362;
  assign new_n2364 = new_n2360 & ~new_n2363;
  assign new_n2365 = in017 & ~new_n1167;
  assign new_n2366 = in117 & new_n1167;
  assign new_n2367 = ~new_n2365 & ~new_n2366;
  assign new_n2368 = in217 & ~new_n1694;
  assign new_n2369 = in317 & new_n1694;
  assign new_n2370 = ~new_n2368 & ~new_n2369;
  assign new_n2371 = new_n2367 & ~new_n2370;
  assign new_n2372 = ~new_n2360 & new_n2363;
  assign new_n2373 = ~new_n2367 & new_n2370;
  assign new_n2374 = in216 & ~new_n1694;
  assign new_n2375 = in316 & new_n1694;
  assign new_n2376 = ~new_n2374 & ~new_n2375;
  assign new_n2377 = in016 & ~new_n1167;
  assign new_n2378 = in116 & new_n1167;
  assign new_n2379 = ~new_n2377 & ~new_n2378;
  assign new_n2380 = ~new_n2376 & new_n2379;
  assign new_n2381 = new_n2376 & ~new_n2379;
  assign new_n2382 = in015 & ~new_n1167;
  assign new_n2383 = in115 & new_n1167;
  assign new_n2384 = ~new_n2382 & ~new_n2383;
  assign new_n2385 = in215 & ~new_n1694;
  assign new_n2386 = in315 & new_n1694;
  assign new_n2387 = ~new_n2385 & ~new_n2386;
  assign new_n2388 = ~new_n2384 & new_n2387;
  assign new_n2389 = in214 & ~new_n1694;
  assign new_n2390 = in314 & new_n1694;
  assign new_n2391 = ~new_n2389 & ~new_n2390;
  assign new_n2392 = in014 & ~new_n1167;
  assign new_n2393 = in114 & new_n1167;
  assign new_n2394 = ~new_n2392 & ~new_n2393;
  assign new_n2395 = ~new_n2391 & new_n2394;
  assign new_n2396 = new_n2384 & ~new_n2387;
  assign new_n2397 = new_n2391 & ~new_n2394;
  assign new_n2398 = in213 & ~new_n1694;
  assign new_n2399 = in313 & new_n1694;
  assign new_n2400 = ~new_n2398 & ~new_n2399;
  assign new_n2401 = in013 & ~new_n1167;
  assign new_n2402 = in113 & new_n1167;
  assign new_n2403 = ~new_n2401 & ~new_n2402;
  assign new_n2404 = new_n2400 & ~new_n2403;
  assign new_n2405 = ~new_n2400 & new_n2403;
  assign new_n2406 = in212 & ~new_n1694;
  assign new_n2407 = in312 & new_n1694;
  assign new_n2408 = ~new_n2406 & ~new_n2407;
  assign new_n2409 = in012 & ~new_n1167;
  assign new_n2410 = in112 & new_n1167;
  assign new_n2411 = ~new_n2409 & ~new_n2410;
  assign new_n2412 = ~new_n2408 & new_n2411;
  assign new_n2413 = in211 & ~new_n1694;
  assign new_n2414 = in311 & new_n1694;
  assign new_n2415 = ~new_n2413 & ~new_n2414;
  assign new_n2416 = in011 & ~new_n1167;
  assign new_n2417 = in111 & new_n1167;
  assign new_n2418 = ~new_n2416 & ~new_n2417;
  assign new_n2419 = new_n2415 & ~new_n2418;
  assign new_n2420 = new_n2408 & ~new_n2411;
  assign new_n2421 = ~new_n2415 & new_n2418;
  assign new_n2422 = in210 & ~new_n1694;
  assign new_n2423 = in310 & new_n1694;
  assign new_n2424 = ~new_n2422 & ~new_n2423;
  assign new_n2425 = in010 & ~new_n1167;
  assign new_n2426 = in110 & new_n1167;
  assign new_n2427 = ~new_n2425 & ~new_n2426;
  assign new_n2428 = new_n2424 & ~new_n2427;
  assign new_n2429 = ~new_n2424 & new_n2427;
  assign new_n2430 = in29 & ~new_n1694;
  assign new_n2431 = in39 & new_n1694;
  assign new_n2432 = ~new_n2430 & ~new_n2431;
  assign new_n2433 = in09 & ~new_n1167;
  assign new_n2434 = in19 & new_n1167;
  assign new_n2435 = ~new_n2433 & ~new_n2434;
  assign new_n2436 = new_n2432 & ~new_n2435;
  assign new_n2437 = in28 & ~new_n1694;
  assign new_n2438 = in38 & new_n1694;
  assign new_n2439 = ~new_n2437 & ~new_n2438;
  assign new_n2440 = in08 & ~new_n1167;
  assign new_n2441 = in18 & new_n1167;
  assign new_n2442 = ~new_n2440 & ~new_n2441;
  assign new_n2443 = ~new_n2439 & new_n2442;
  assign new_n2444 = ~new_n2432 & new_n2435;
  assign new_n2445 = new_n2439 & ~new_n2442;
  assign new_n2446 = in07 & ~new_n1167;
  assign new_n2447 = in17 & new_n1167;
  assign new_n2448 = ~new_n2446 & ~new_n2447;
  assign new_n2449 = in27 & ~new_n1694;
  assign new_n2450 = in37 & new_n1694;
  assign new_n2451 = ~new_n2449 & ~new_n2450;
  assign new_n2452 = new_n2448 & ~new_n2451;
  assign new_n2453 = ~new_n2448 & new_n2451;
  assign new_n2454 = in26 & ~new_n1694;
  assign new_n2455 = in36 & new_n1694;
  assign new_n2456 = ~new_n2454 & ~new_n2455;
  assign new_n2457 = in06 & ~new_n1167;
  assign new_n2458 = in16 & new_n1167;
  assign new_n2459 = ~new_n2457 & ~new_n2458;
  assign new_n2460 = new_n2456 & ~new_n2459;
  assign new_n2461 = in05 & ~new_n1167;
  assign new_n2462 = in15 & new_n1167;
  assign new_n2463 = ~new_n2461 & ~new_n2462;
  assign new_n2464 = in25 & ~new_n1694;
  assign new_n2465 = in35 & new_n1694;
  assign new_n2466 = ~new_n2464 & ~new_n2465;
  assign new_n2467 = new_n2463 & ~new_n2466;
  assign new_n2468 = ~new_n2456 & new_n2459;
  assign new_n2469 = ~new_n2463 & new_n2466;
  assign new_n2470 = in24 & ~new_n1694;
  assign new_n2471 = in34 & new_n1694;
  assign new_n2472 = ~new_n2470 & ~new_n2471;
  assign new_n2473 = in04 & ~new_n1167;
  assign new_n2474 = in14 & new_n1167;
  assign new_n2475 = ~new_n2473 & ~new_n2474;
  assign new_n2476 = new_n2472 & ~new_n2475;
  assign new_n2477 = in23 & ~new_n1694;
  assign new_n2478 = in33 & new_n1694;
  assign new_n2479 = ~new_n2477 & ~new_n2478;
  assign new_n2480 = in03 & ~new_n1167;
  assign new_n2481 = in13 & new_n1167;
  assign new_n2482 = ~new_n2480 & ~new_n2481;
  assign new_n2483 = ~new_n2479 & new_n2482;
  assign new_n2484 = ~new_n2472 & new_n2475;
  assign new_n2485 = new_n2479 & ~new_n2482;
  assign new_n2486 = in02 & ~new_n1167;
  assign new_n2487 = in12 & new_n1167;
  assign new_n2488 = ~new_n2486 & ~new_n2487;
  assign new_n2489 = in22 & ~new_n1694;
  assign new_n2490 = in32 & new_n1694;
  assign new_n2491 = ~new_n2489 & ~new_n2490;
  assign new_n2492 = in01 & ~new_n1167;
  assign new_n2493 = in11 & new_n1167;
  assign new_n2494 = ~new_n2492 & ~new_n2493;
  assign new_n2495 = in21 & ~new_n1694;
  assign new_n2496 = in31 & new_n1694;
  assign new_n2497 = ~new_n2495 & ~new_n2496;
  assign new_n2498 = ~new_n2494 & new_n2497;
  assign new_n2499 = in20 & ~new_n1694;
  assign new_n2500 = in30 & new_n1694;
  assign new_n2501 = ~new_n2499 & ~new_n2500;
  assign new_n2502 = new_n2494 & ~new_n2497;
  assign new_n2503 = ~new_n1170 & new_n2501;
  assign new_n2504 = ~new_n2502 & new_n2503;
  assign new_n2505 = ~new_n2498 & ~new_n2504;
  assign new_n2506 = new_n2491 & ~new_n2505;
  assign new_n2507 = new_n2488 & ~new_n2506;
  assign new_n2508 = ~new_n2491 & new_n2505;
  assign new_n2509 = ~new_n2507 & ~new_n2508;
  assign new_n2510 = ~new_n2485 & ~new_n2509;
  assign new_n2511 = ~new_n2483 & ~new_n2484;
  assign new_n2512 = ~new_n2510 & new_n2511;
  assign new_n2513 = ~new_n2469 & ~new_n2476;
  assign new_n2514 = ~new_n2512 & new_n2513;
  assign new_n2515 = ~new_n2467 & ~new_n2468;
  assign new_n2516 = ~new_n2514 & new_n2515;
  assign new_n2517 = ~new_n2453 & ~new_n2460;
  assign new_n2518 = ~new_n2516 & new_n2517;
  assign new_n2519 = ~new_n2452 & ~new_n2518;
  assign new_n2520 = ~new_n2445 & ~new_n2519;
  assign new_n2521 = ~new_n2443 & ~new_n2444;
  assign new_n2522 = ~new_n2520 & new_n2521;
  assign new_n2523 = ~new_n2436 & ~new_n2522;
  assign new_n2524 = ~new_n2429 & ~new_n2523;
  assign new_n2525 = ~new_n2428 & ~new_n2524;
  assign new_n2526 = ~new_n2421 & ~new_n2525;
  assign new_n2527 = ~new_n2419 & ~new_n2420;
  assign new_n2528 = ~new_n2526 & new_n2527;
  assign new_n2529 = ~new_n2405 & ~new_n2412;
  assign new_n2530 = ~new_n2528 & new_n2529;
  assign new_n2531 = ~new_n2397 & ~new_n2404;
  assign new_n2532 = ~new_n2530 & new_n2531;
  assign new_n2533 = ~new_n2395 & ~new_n2396;
  assign new_n2534 = ~new_n2532 & new_n2533;
  assign new_n2535 = ~new_n2381 & ~new_n2388;
  assign new_n2536 = ~new_n2534 & new_n2535;
  assign new_n2537 = ~new_n2380 & ~new_n2536;
  assign new_n2538 = ~new_n2373 & ~new_n2537;
  assign new_n2539 = ~new_n2371 & ~new_n2372;
  assign new_n2540 = ~new_n2538 & new_n2539;
  assign new_n2541 = ~new_n2364 & ~new_n2540;
  assign new_n2542 = ~new_n2357 & ~new_n2541;
  assign new_n2543 = ~new_n2356 & ~new_n2542;
  assign new_n2544 = ~new_n2349 & ~new_n2543;
  assign new_n2545 = ~new_n2347 & ~new_n2348;
  assign new_n2546 = ~new_n2544 & new_n2545;
  assign new_n2547 = ~new_n2333 & ~new_n2340;
  assign new_n2548 = ~new_n2546 & new_n2547;
  assign new_n2549 = ~new_n2325 & ~new_n2332;
  assign new_n2550 = ~new_n2548 & new_n2549;
  assign new_n2551 = ~new_n2323 & ~new_n2324;
  assign new_n2552 = ~new_n2550 & new_n2551;
  assign new_n2553 = ~new_n2309 & ~new_n2316;
  assign new_n2554 = ~new_n2552 & new_n2553;
  assign new_n2555 = ~new_n2307 & ~new_n2308;
  assign new_n2556 = ~new_n2554 & new_n2555;
  assign new_n2557 = ~new_n2293 & ~new_n2300;
  assign new_n2558 = ~new_n2556 & new_n2557;
  assign new_n2559 = ~new_n2291 & ~new_n2292;
  assign new_n2560 = ~new_n2558 & new_n2559;
  assign new_n2561 = ~new_n2277 & ~new_n2284;
  assign new_n2562 = ~new_n2560 & new_n2561;
  assign new_n2563 = ~new_n2275 & ~new_n2276;
  assign new_n2564 = ~new_n2562 & new_n2563;
  assign new_n2565 = ~new_n2261 & ~new_n2268;
  assign new_n2566 = ~new_n2564 & new_n2565;
  assign new_n2567 = in233 & ~new_n1694;
  assign new_n2568 = in333 & new_n1694;
  assign new_n2569 = ~new_n2567 & ~new_n2568;
  assign new_n2570 = in033 & ~new_n1167;
  assign new_n2571 = in133 & new_n1167;
  assign new_n2572 = ~new_n2570 & ~new_n2571;
  assign new_n2573 = ~new_n2569 & new_n2572;
  assign new_n2574 = in234 & ~new_n1694;
  assign new_n2575 = in334 & new_n1694;
  assign new_n2576 = ~new_n2574 & ~new_n2575;
  assign new_n2577 = in034 & ~new_n1167;
  assign new_n2578 = in134 & new_n1167;
  assign new_n2579 = ~new_n2577 & ~new_n2578;
  assign new_n2580 = ~new_n2576 & new_n2579;
  assign new_n2581 = ~new_n2573 & ~new_n2580;
  assign new_n2582 = in237 & ~new_n1694;
  assign new_n2583 = in337 & new_n1694;
  assign new_n2584 = ~new_n2582 & ~new_n2583;
  assign new_n2585 = in037 & ~new_n1167;
  assign new_n2586 = in137 & new_n1167;
  assign new_n2587 = ~new_n2585 & ~new_n2586;
  assign new_n2588 = ~new_n2584 & new_n2587;
  assign new_n2589 = new_n2243 & ~new_n2246;
  assign new_n2590 = ~new_n2588 & ~new_n2589;
  assign new_n2591 = in235 & ~new_n1694;
  assign new_n2592 = in335 & new_n1694;
  assign new_n2593 = ~new_n2591 & ~new_n2592;
  assign new_n2594 = in035 & ~new_n1167;
  assign new_n2595 = in135 & new_n1167;
  assign new_n2596 = ~new_n2594 & ~new_n2595;
  assign new_n2597 = ~new_n2593 & new_n2596;
  assign new_n2598 = in036 & ~new_n1167;
  assign new_n2599 = in136 & new_n1167;
  assign new_n2600 = ~new_n2598 & ~new_n2599;
  assign new_n2601 = in236 & ~new_n1694;
  assign new_n2602 = in336 & new_n1694;
  assign new_n2603 = ~new_n2601 & ~new_n2602;
  assign new_n2604 = new_n2600 & ~new_n2603;
  assign new_n2605 = ~new_n2597 & ~new_n2604;
  assign new_n2606 = new_n2257 & ~new_n2260;
  assign new_n2607 = ~new_n2254 & ~new_n2606;
  assign new_n2608 = new_n2581 & new_n2607;
  assign new_n2609 = new_n2590 & new_n2605;
  assign new_n2610 = new_n2608 & new_n2609;
  assign new_n2611 = ~new_n2566 & new_n2610;
  assign new_n2612 = in039 & ~new_n1167;
  assign new_n2613 = in139 & new_n1167;
  assign new_n2614 = ~new_n2612 & ~new_n2613;
  assign new_n2615 = in239 & ~new_n1694;
  assign new_n2616 = in339 & new_n1694;
  assign new_n2617 = ~new_n2615 & ~new_n2616;
  assign new_n2618 = ~new_n2614 & new_n2617;
  assign new_n2619 = new_n2584 & ~new_n2587;
  assign new_n2620 = ~new_n2600 & new_n2603;
  assign new_n2621 = new_n2593 & ~new_n2596;
  assign new_n2622 = new_n2576 & ~new_n2579;
  assign new_n2623 = new_n2569 & ~new_n2572;
  assign new_n2624 = new_n2250 & ~new_n2253;
  assign new_n2625 = ~new_n2623 & ~new_n2624;
  assign new_n2626 = new_n2581 & ~new_n2625;
  assign new_n2627 = ~new_n2621 & ~new_n2622;
  assign new_n2628 = ~new_n2626 & new_n2627;
  assign new_n2629 = new_n2605 & ~new_n2628;
  assign new_n2630 = ~new_n2619 & ~new_n2620;
  assign new_n2631 = ~new_n2629 & new_n2630;
  assign new_n2632 = new_n2590 & ~new_n2631;
  assign new_n2633 = ~new_n2247 & ~new_n2618;
  assign new_n2634 = ~new_n2632 & new_n2633;
  assign new_n2635 = ~new_n2611 & new_n2634;
  assign new_n2636 = in242 & ~new_n1694;
  assign new_n2637 = in342 & new_n1694;
  assign new_n2638 = ~new_n2636 & ~new_n2637;
  assign new_n2639 = in042 & ~new_n1167;
  assign new_n2640 = in142 & new_n1167;
  assign new_n2641 = ~new_n2639 & ~new_n2640;
  assign new_n2642 = ~new_n2638 & new_n2641;
  assign new_n2643 = in043 & ~new_n1167;
  assign new_n2644 = in143 & new_n1167;
  assign new_n2645 = ~new_n2643 & ~new_n2644;
  assign new_n2646 = in243 & ~new_n1694;
  assign new_n2647 = in343 & new_n1694;
  assign new_n2648 = ~new_n2646 & ~new_n2647;
  assign new_n2649 = new_n2645 & ~new_n2648;
  assign new_n2650 = ~new_n2642 & ~new_n2649;
  assign new_n2651 = in044 & ~new_n1167;
  assign new_n2652 = in144 & new_n1167;
  assign new_n2653 = ~new_n2651 & ~new_n2652;
  assign new_n2654 = in244 & ~new_n1694;
  assign new_n2655 = in344 & new_n1694;
  assign new_n2656 = ~new_n2654 & ~new_n2655;
  assign new_n2657 = new_n2653 & ~new_n2656;
  assign new_n2658 = new_n2614 & ~new_n2617;
  assign new_n2659 = in241 & ~new_n1694;
  assign new_n2660 = in341 & new_n1694;
  assign new_n2661 = ~new_n2659 & ~new_n2660;
  assign new_n2662 = in041 & ~new_n1167;
  assign new_n2663 = in141 & new_n1167;
  assign new_n2664 = ~new_n2662 & ~new_n2663;
  assign new_n2665 = ~new_n2661 & new_n2664;
  assign new_n2666 = ~new_n2240 & ~new_n2657;
  assign new_n2667 = ~new_n2658 & ~new_n2665;
  assign new_n2668 = new_n2666 & new_n2667;
  assign new_n2669 = new_n2650 & new_n2668;
  assign new_n2670 = ~new_n2635 & new_n2669;
  assign new_n2671 = ~new_n2653 & new_n2656;
  assign new_n2672 = ~new_n2645 & new_n2648;
  assign new_n2673 = new_n2661 & ~new_n2664;
  assign new_n2674 = new_n2638 & ~new_n2641;
  assign new_n2675 = new_n2236 & ~new_n2239;
  assign new_n2676 = ~new_n2665 & new_n2675;
  assign new_n2677 = ~new_n2673 & ~new_n2674;
  assign new_n2678 = ~new_n2676 & new_n2677;
  assign new_n2679 = new_n2650 & ~new_n2678;
  assign new_n2680 = ~new_n2672 & ~new_n2679;
  assign new_n2681 = ~new_n2657 & ~new_n2680;
  assign new_n2682 = ~new_n2233 & ~new_n2671;
  assign new_n2683 = ~new_n2681 & new_n2682;
  assign new_n2684 = ~new_n2670 & new_n2683;
  assign new_n2685 = ~new_n2231 & ~new_n2232;
  assign new_n2686 = ~new_n2684 & new_n2685;
  assign new_n2687 = ~new_n2217 & ~new_n2224;
  assign new_n2688 = ~new_n2686 & new_n2687;
  assign new_n2689 = in050 & ~new_n1167;
  assign new_n2690 = in150 & new_n1167;
  assign new_n2691 = ~new_n2689 & ~new_n2690;
  assign new_n2692 = in250 & ~new_n1694;
  assign new_n2693 = in350 & new_n1694;
  assign new_n2694 = ~new_n2692 & ~new_n2693;
  assign new_n2695 = new_n2691 & ~new_n2694;
  assign new_n2696 = in049 & ~new_n1167;
  assign new_n2697 = in149 & new_n1167;
  assign new_n2698 = ~new_n2696 & ~new_n2697;
  assign new_n2699 = in249 & ~new_n1694;
  assign new_n2700 = in349 & new_n1694;
  assign new_n2701 = ~new_n2699 & ~new_n2700;
  assign new_n2702 = new_n2698 & ~new_n2701;
  assign new_n2703 = ~new_n2695 & ~new_n2702;
  assign new_n2704 = ~new_n2213 & new_n2216;
  assign new_n2705 = in251 & ~new_n1694;
  assign new_n2706 = in351 & new_n1694;
  assign new_n2707 = ~new_n2705 & ~new_n2706;
  assign new_n2708 = in051 & ~new_n1167;
  assign new_n2709 = in151 & new_n1167;
  assign new_n2710 = ~new_n2708 & ~new_n2709;
  assign new_n2711 = ~new_n2707 & new_n2710;
  assign new_n2712 = new_n2206 & ~new_n2209;
  assign new_n2713 = ~new_n2711 & ~new_n2712;
  assign new_n2714 = in048 & ~new_n1167;
  assign new_n2715 = in148 & new_n1167;
  assign new_n2716 = ~new_n2714 & ~new_n2715;
  assign new_n2717 = in248 & ~new_n1694;
  assign new_n2718 = in348 & new_n1694;
  assign new_n2719 = ~new_n2717 & ~new_n2718;
  assign new_n2720 = new_n2716 & ~new_n2719;
  assign new_n2721 = ~new_n2704 & ~new_n2720;
  assign new_n2722 = new_n2703 & new_n2721;
  assign new_n2723 = new_n2713 & new_n2722;
  assign new_n2724 = ~new_n2688 & new_n2723;
  assign new_n2725 = new_n2199 & ~new_n2202;
  assign new_n2726 = ~new_n2691 & new_n2694;
  assign new_n2727 = new_n2707 & ~new_n2710;
  assign new_n2728 = ~new_n2698 & new_n2701;
  assign new_n2729 = ~new_n2716 & new_n2719;
  assign new_n2730 = ~new_n2728 & ~new_n2729;
  assign new_n2731 = new_n2703 & ~new_n2730;
  assign new_n2732 = ~new_n2726 & ~new_n2727;
  assign new_n2733 = ~new_n2731 & new_n2732;
  assign new_n2734 = new_n2713 & ~new_n2733;
  assign new_n2735 = ~new_n2210 & ~new_n2725;
  assign new_n2736 = ~new_n2734 & new_n2735;
  assign new_n2737 = ~new_n2724 & new_n2736;
  assign new_n2738 = ~new_n2196 & ~new_n2203;
  assign new_n2739 = ~new_n2737 & new_n2738;
  assign new_n2740 = ~new_n2188 & ~new_n2195;
  assign new_n2741 = ~new_n2739 & new_n2740;
  assign new_n2742 = in258 & ~new_n1694;
  assign new_n2743 = in358 & new_n1694;
  assign new_n2744 = ~new_n2742 & ~new_n2743;
  assign new_n2745 = in058 & ~new_n1167;
  assign new_n2746 = in158 & new_n1167;
  assign new_n2747 = ~new_n2745 & ~new_n2746;
  assign new_n2748 = ~new_n2744 & new_n2747;
  assign new_n2749 = in259 & ~new_n1694;
  assign new_n2750 = in359 & new_n1694;
  assign new_n2751 = ~new_n2749 & ~new_n2750;
  assign new_n2752 = in059 & ~new_n1167;
  assign new_n2753 = in159 & new_n1167;
  assign new_n2754 = ~new_n2752 & ~new_n2753;
  assign new_n2755 = ~new_n2751 & new_n2754;
  assign new_n2756 = ~new_n2748 & ~new_n2755;
  assign new_n2757 = new_n2191 & ~new_n2194;
  assign new_n2758 = in260 & ~new_n1694;
  assign new_n2759 = in360 & new_n1694;
  assign new_n2760 = ~new_n2758 & ~new_n2759;
  assign new_n2761 = in060 & ~new_n1167;
  assign new_n2762 = in160 & new_n1167;
  assign new_n2763 = ~new_n2761 & ~new_n2762;
  assign new_n2764 = ~new_n2760 & new_n2763;
  assign new_n2765 = in257 & ~new_n1694;
  assign new_n2766 = in357 & new_n1694;
  assign new_n2767 = ~new_n2765 & ~new_n2766;
  assign new_n2768 = in057 & ~new_n1167;
  assign new_n2769 = in157 & new_n1167;
  assign new_n2770 = ~new_n2768 & ~new_n2769;
  assign new_n2771 = ~new_n2767 & new_n2770;
  assign new_n2772 = ~new_n2181 & ~new_n2757;
  assign new_n2773 = ~new_n2764 & ~new_n2771;
  assign new_n2774 = new_n2772 & new_n2773;
  assign new_n2775 = new_n2756 & new_n2774;
  assign new_n2776 = ~new_n2741 & new_n2775;
  assign new_n2777 = new_n2760 & ~new_n2763;
  assign new_n2778 = new_n2751 & ~new_n2754;
  assign new_n2779 = new_n2744 & ~new_n2747;
  assign new_n2780 = new_n2767 & ~new_n2770;
  assign new_n2781 = new_n2177 & ~new_n2180;
  assign new_n2782 = ~new_n2771 & new_n2781;
  assign new_n2783 = ~new_n2779 & ~new_n2780;
  assign new_n2784 = ~new_n2782 & new_n2783;
  assign new_n2785 = new_n2756 & ~new_n2784;
  assign new_n2786 = ~new_n2778 & ~new_n2785;
  assign new_n2787 = ~new_n2764 & ~new_n2786;
  assign new_n2788 = ~new_n2174 & ~new_n2777;
  assign new_n2789 = ~new_n2787 & new_n2788;
  assign new_n2790 = ~new_n2776 & new_n2789;
  assign new_n2791 = ~new_n2173 & ~new_n2790;
  assign new_n2792 = ~new_n2166 & ~new_n2791;
  assign new_n2793 = ~new_n2164 & ~new_n2165;
  assign new_n2794 = ~new_n2792 & new_n2793;
  assign new_n2795 = ~new_n2157 & ~new_n2794;
  assign new_n2796 = ~new_n2150 & ~new_n2795;
  assign new_n2797 = ~new_n2149 & ~new_n2796;
  assign new_n2798 = ~new_n2142 & ~new_n2797;
  assign new_n2799 = ~new_n2141 & ~new_n2798;
  assign new_n2800 = ~new_n2134 & ~new_n2799;
  assign new_n2801 = ~new_n2132 & ~new_n2133;
  assign new_n2802 = ~new_n2800 & new_n2801;
  assign new_n2803 = ~new_n2125 & ~new_n2802;
  assign new_n2804 = ~new_n2118 & ~new_n2803;
  assign new_n2805 = ~new_n2117 & ~new_n2804;
  assign new_n2806 = ~new_n2110 & ~new_n2805;
  assign new_n2807 = ~new_n2109 & ~new_n2806;
  assign new_n2808 = ~new_n2102 & ~new_n2807;
  assign new_n2809 = ~new_n2100 & ~new_n2101;
  assign new_n2810 = ~new_n2808 & new_n2809;
  assign new_n2811 = ~new_n2086 & ~new_n2093;
  assign new_n2812 = ~new_n2810 & new_n2811;
  assign new_n2813 = ~new_n2078 & ~new_n2085;
  assign new_n2814 = ~new_n2812 & new_n2813;
  assign new_n2815 = ~new_n2070 & ~new_n2077;
  assign new_n2816 = ~new_n2814 & new_n2815;
  assign new_n2817 = ~new_n2068 & ~new_n2069;
  assign new_n2818 = ~new_n2816 & new_n2817;
  assign new_n2819 = ~new_n2054 & ~new_n2061;
  assign new_n2820 = ~new_n2818 & new_n2819;
  assign new_n2821 = ~new_n2053 & ~new_n2820;
  assign new_n2822 = ~new_n2046 & ~new_n2821;
  assign new_n2823 = ~new_n2045 & ~new_n2822;
  assign new_n2824 = ~new_n2038 & ~new_n2823;
  assign new_n2825 = ~new_n2036 & ~new_n2037;
  assign new_n2826 = ~new_n2824 & new_n2825;
  assign new_n2827 = ~new_n2022 & ~new_n2029;
  assign new_n2828 = ~new_n2826 & new_n2827;
  assign new_n2829 = ~new_n2014 & ~new_n2021;
  assign new_n2830 = ~new_n2828 & new_n2829;
  assign new_n2831 = ~new_n2006 & ~new_n2013;
  assign new_n2832 = ~new_n2830 & new_n2831;
  assign new_n2833 = ~new_n2004 & ~new_n2005;
  assign new_n2834 = ~new_n2832 & new_n2833;
  assign new_n2835 = ~new_n1996 & ~new_n1997;
  assign new_n2836 = ~new_n2834 & new_n2835;
  assign new_n2837 = ~new_n1989 & ~new_n2836;
  assign new_n2838 = ~new_n1982 & ~new_n2837;
  assign new_n2839 = ~new_n1980 & ~new_n1981;
  assign new_n2840 = ~new_n2838 & new_n2839;
  assign new_n2841 = ~new_n1973 & ~new_n2840;
  assign new_n2842 = ~new_n1966 & ~new_n2841;
  assign new_n2843 = ~new_n1965 & ~new_n2842;
  assign new_n2844 = ~new_n1958 & ~new_n2843;
  assign new_n2845 = ~new_n1957 & ~new_n2844;
  assign new_n2846 = ~new_n1950 & ~new_n2845;
  assign new_n2847 = ~new_n1949 & ~new_n2846;
  assign new_n2848 = ~new_n1942 & ~new_n2847;
  assign new_n2849 = ~new_n1941 & ~new_n2848;
  assign new_n2850 = ~new_n1934 & ~new_n2849;
  assign new_n2851 = ~new_n1932 & ~new_n1933;
  assign new_n2852 = ~new_n2850 & new_n2851;
  assign new_n2853 = ~new_n1925 & ~new_n2852;
  assign new_n2854 = ~new_n1918 & ~new_n2853;
  assign new_n2855 = ~new_n1917 & ~new_n2854;
  assign new_n2856 = ~new_n1910 & ~new_n2855;
  assign new_n2857 = ~new_n1909 & ~new_n2856;
  assign new_n2858 = ~new_n1902 & ~new_n2857;
  assign new_n2859 = ~new_n1901 & ~new_n2858;
  assign new_n2860 = ~new_n1894 & ~new_n2859;
  assign new_n2861 = ~new_n1893 & ~new_n2860;
  assign new_n2862 = ~new_n1886 & ~new_n2861;
  assign new_n2863 = ~new_n1884 & ~new_n1885;
  assign new_n2864 = ~new_n2862 & new_n2863;
  assign new_n2865 = ~new_n1877 & ~new_n2864;
  assign new_n2866 = ~new_n1870 & ~new_n2865;
  assign new_n2867 = ~new_n1869 & ~new_n2866;
  assign new_n2868 = ~new_n1862 & ~new_n2867;
  assign new_n2869 = ~new_n1860 & ~new_n1861;
  assign new_n2870 = ~new_n2868 & new_n2869;
  assign new_n2871 = ~new_n1846 & ~new_n1853;
  assign new_n2872 = ~new_n2870 & new_n2871;
  assign new_n2873 = ~new_n1844 & ~new_n1845;
  assign new_n2874 = ~new_n2872 & new_n2873;
  assign new_n2875 = ~new_n1830 & ~new_n1837;
  assign new_n2876 = ~new_n2874 & new_n2875;
  assign new_n2877 = ~new_n1828 & ~new_n1829;
  assign new_n2878 = ~new_n2876 & new_n2877;
  assign new_n2879 = ~new_n1814 & ~new_n1821;
  assign new_n2880 = ~new_n2878 & new_n2879;
  assign new_n2881 = ~new_n1812 & ~new_n1813;
  assign new_n2882 = ~new_n2880 & new_n2881;
  assign new_n2883 = ~new_n1798 & ~new_n1805;
  assign new_n2884 = ~new_n2882 & new_n2883;
  assign new_n2885 = ~new_n1796 & ~new_n1797;
  assign new_n2886 = ~new_n2884 & new_n2885;
  assign new_n2887 = in2110 & ~new_n1694;
  assign new_n2888 = in3110 & new_n1694;
  assign new_n2889 = ~new_n2887 & ~new_n2888;
  assign new_n2890 = in0110 & ~new_n1167;
  assign new_n2891 = in1110 & new_n1167;
  assign new_n2892 = ~new_n2890 & ~new_n2891;
  assign new_n2893 = ~new_n2889 & new_n2892;
  assign new_n2894 = in2111 & ~new_n1694;
  assign new_n2895 = in3111 & new_n1694;
  assign new_n2896 = ~new_n2894 & ~new_n2895;
  assign new_n2897 = in0111 & ~new_n1167;
  assign new_n2898 = in1111 & new_n1167;
  assign new_n2899 = ~new_n2897 & ~new_n2898;
  assign new_n2900 = ~new_n2896 & new_n2899;
  assign new_n2901 = ~new_n1789 & ~new_n2893;
  assign new_n2902 = ~new_n2900 & new_n2901;
  assign new_n2903 = ~new_n2886 & new_n2902;
  assign new_n2904 = in2112 & ~new_n1694;
  assign new_n2905 = in3112 & new_n1694;
  assign new_n2906 = ~new_n2904 & ~new_n2905;
  assign new_n2907 = in0112 & ~new_n1167;
  assign new_n2908 = in1112 & new_n1167;
  assign new_n2909 = ~new_n2907 & ~new_n2908;
  assign new_n2910 = new_n2906 & ~new_n2909;
  assign new_n2911 = new_n2896 & ~new_n2899;
  assign new_n2912 = new_n2889 & ~new_n2892;
  assign new_n2913 = ~new_n2900 & new_n2912;
  assign new_n2914 = ~new_n2910 & ~new_n2911;
  assign new_n2915 = ~new_n2913 & new_n2914;
  assign new_n2916 = ~new_n2903 & new_n2915;
  assign new_n2917 = ~new_n2906 & new_n2909;
  assign new_n2918 = ~new_n2916 & ~new_n2917;
  assign new_n2919 = ~new_n1782 & ~new_n2918;
  assign new_n2920 = ~new_n1778 & new_n1781;
  assign new_n2921 = ~new_n1775 & ~new_n2920;
  assign new_n2922 = ~new_n2919 & new_n2921;
  assign new_n2923 = ~new_n1773 & ~new_n1774;
  assign new_n2924 = ~new_n2922 & new_n2923;
  assign new_n2925 = ~new_n1759 & ~new_n1766;
  assign new_n2926 = ~new_n2924 & new_n2925;
  assign new_n2927 = ~new_n1757 & ~new_n1758;
  assign new_n2928 = ~new_n2926 & new_n2927;
  assign new_n2929 = in0118 & ~new_n1167;
  assign new_n2930 = in1118 & new_n1167;
  assign new_n2931 = ~new_n2929 & ~new_n2930;
  assign new_n2932 = in2118 & ~new_n1694;
  assign new_n2933 = in3118 & new_n1694;
  assign new_n2934 = ~new_n2932 & ~new_n2933;
  assign new_n2935 = new_n2931 & ~new_n2934;
  assign new_n2936 = in2119 & ~new_n1694;
  assign new_n2937 = in3119 & new_n1694;
  assign new_n2938 = ~new_n2936 & ~new_n2937;
  assign new_n2939 = in0119 & ~new_n1167;
  assign new_n2940 = in1119 & new_n1167;
  assign new_n2941 = ~new_n2939 & ~new_n2940;
  assign new_n2942 = ~new_n2938 & new_n2941;
  assign new_n2943 = ~new_n1750 & ~new_n2935;
  assign new_n2944 = ~new_n2942 & new_n2943;
  assign new_n2945 = ~new_n2928 & new_n2944;
  assign new_n2946 = in2120 & ~new_n1694;
  assign new_n2947 = in3120 & new_n1694;
  assign new_n2948 = ~new_n2946 & ~new_n2947;
  assign new_n2949 = in0120 & ~new_n1167;
  assign new_n2950 = in1120 & new_n1167;
  assign new_n2951 = ~new_n2949 & ~new_n2950;
  assign new_n2952 = new_n2948 & ~new_n2951;
  assign new_n2953 = new_n2938 & ~new_n2941;
  assign new_n2954 = ~new_n2931 & new_n2934;
  assign new_n2955 = ~new_n2942 & new_n2954;
  assign new_n2956 = ~new_n2952 & ~new_n2953;
  assign new_n2957 = ~new_n2955 & new_n2956;
  assign new_n2958 = ~new_n2945 & new_n2957;
  assign new_n2959 = ~new_n2948 & new_n2951;
  assign new_n2960 = ~new_n2958 & ~new_n2959;
  assign new_n2961 = ~new_n1743 & ~new_n2960;
  assign new_n2962 = ~new_n1731 & new_n1734;
  assign new_n2963 = ~new_n1742 & ~new_n2962;
  assign new_n2964 = ~new_n2961 & new_n2963;
  assign new_n2965 = ~new_n1728 & ~new_n1735;
  assign new_n2966 = ~new_n2964 & new_n2965;
  assign new_n2967 = ~new_n1724 & new_n1727;
  assign new_n2968 = ~new_n1721 & ~new_n2967;
  assign new_n2969 = new_n1710 & new_n2968;
  assign new_n2970 = ~new_n2966 & new_n2969;
  assign new_n2971 = ~new_n1701 & ~new_n1720;
  assign new_n2972 = ~new_n2970 & new_n2971;
  assign new_n2973 = new_n1172 & new_n2972;
  assign new_n2974 = new_n1171 & ~new_n2973;
  assign new_n2975 = ~new_n1172 & ~new_n2972;
  assign address1 = ~new_n2974 & ~new_n2975;
  assign new_n2977 = ~new_n1170 & ~address1;
  assign new_n2978 = ~new_n2501 & address1;
  assign result0 = new_n2977 | new_n2978;
  assign new_n2980 = ~new_n2497 & address1;
  assign new_n2981 = ~new_n2494 & ~address1;
  assign result1 = new_n2980 | new_n2981;
  assign new_n2983 = ~new_n2488 & ~address1;
  assign new_n2984 = ~new_n2491 & address1;
  assign result2 = new_n2983 | new_n2984;
  assign new_n2986 = ~new_n2482 & ~address1;
  assign new_n2987 = ~new_n2479 & address1;
  assign result3 = new_n2986 | new_n2987;
  assign new_n2989 = ~new_n2475 & ~address1;
  assign new_n2990 = ~new_n2472 & address1;
  assign result4 = new_n2989 | new_n2990;
  assign new_n2992 = ~new_n2463 & ~address1;
  assign new_n2993 = ~new_n2466 & address1;
  assign result5 = new_n2992 | new_n2993;
  assign new_n2995 = ~new_n2459 & ~address1;
  assign new_n2996 = ~new_n2456 & address1;
  assign result6 = new_n2995 | new_n2996;
  assign new_n2998 = ~new_n2448 & ~address1;
  assign new_n2999 = ~new_n2451 & address1;
  assign result7 = new_n2998 | new_n2999;
  assign new_n3001 = ~new_n2442 & ~address1;
  assign new_n3002 = ~new_n2439 & address1;
  assign result8 = new_n3001 | new_n3002;
  assign new_n3004 = ~new_n2435 & ~address1;
  assign new_n3005 = ~new_n2432 & address1;
  assign result9 = new_n3004 | new_n3005;
  assign new_n3007 = ~new_n2427 & ~address1;
  assign new_n3008 = ~new_n2424 & address1;
  assign result10 = new_n3007 | new_n3008;
  assign new_n3010 = ~new_n2418 & ~address1;
  assign new_n3011 = ~new_n2415 & address1;
  assign result11 = new_n3010 | new_n3011;
  assign new_n3013 = ~new_n2411 & ~address1;
  assign new_n3014 = ~new_n2408 & address1;
  assign result12 = new_n3013 | new_n3014;
  assign new_n3016 = ~new_n2403 & ~address1;
  assign new_n3017 = ~new_n2400 & address1;
  assign result13 = new_n3016 | new_n3017;
  assign new_n3019 = ~new_n2394 & ~address1;
  assign new_n3020 = ~new_n2391 & address1;
  assign result14 = new_n3019 | new_n3020;
  assign new_n3022 = ~new_n2384 & ~address1;
  assign new_n3023 = ~new_n2387 & address1;
  assign result15 = new_n3022 | new_n3023;
  assign new_n3025 = ~new_n2379 & ~address1;
  assign new_n3026 = ~new_n2376 & address1;
  assign result16 = new_n3025 | new_n3026;
  assign new_n3028 = ~new_n2367 & ~address1;
  assign new_n3029 = ~new_n2370 & address1;
  assign result17 = new_n3028 | new_n3029;
  assign new_n3031 = ~new_n2363 & ~address1;
  assign new_n3032 = ~new_n2360 & address1;
  assign result18 = new_n3031 | new_n3032;
  assign new_n3034 = ~new_n2355 & ~address1;
  assign new_n3035 = ~new_n2352 & address1;
  assign result19 = new_n3034 | new_n3035;
  assign new_n3037 = ~new_n2346 & ~address1;
  assign new_n3038 = ~new_n2343 & address1;
  assign result20 = new_n3037 | new_n3038;
  assign new_n3040 = ~new_n2339 & ~address1;
  assign new_n3041 = ~new_n2336 & address1;
  assign result21 = new_n3040 | new_n3041;
  assign new_n3043 = ~new_n2331 & ~address1;
  assign new_n3044 = ~new_n2328 & address1;
  assign result22 = new_n3043 | new_n3044;
  assign new_n3046 = ~new_n2322 & ~address1;
  assign new_n3047 = ~new_n2319 & address1;
  assign result23 = new_n3046 | new_n3047;
  assign new_n3049 = ~new_n2312 & ~address1;
  assign new_n3050 = ~new_n2315 & address1;
  assign result24 = new_n3049 | new_n3050;
  assign new_n3052 = ~new_n2306 & ~address1;
  assign new_n3053 = ~new_n2303 & address1;
  assign result25 = new_n3052 | new_n3053;
  assign new_n3055 = ~new_n2296 & ~address1;
  assign new_n3056 = ~new_n2299 & address1;
  assign result26 = new_n3055 | new_n3056;
  assign new_n3058 = ~new_n2290 & ~address1;
  assign new_n3059 = ~new_n2287 & address1;
  assign result27 = new_n3058 | new_n3059;
  assign new_n3061 = ~new_n2280 & ~address1;
  assign new_n3062 = ~new_n2283 & address1;
  assign result28 = new_n3061 | new_n3062;
  assign new_n3064 = ~new_n2274 & ~address1;
  assign new_n3065 = ~new_n2271 & address1;
  assign result29 = new_n3064 | new_n3065;
  assign new_n3067 = ~new_n2264 & ~address1;
  assign new_n3068 = ~new_n2267 & address1;
  assign result30 = new_n3067 | new_n3068;
  assign new_n3070 = ~new_n2260 & address1;
  assign new_n3071 = ~new_n2257 & ~address1;
  assign result31 = new_n3070 | new_n3071;
  assign new_n3073 = ~new_n2253 & ~address1;
  assign new_n3074 = ~new_n2250 & address1;
  assign result32 = new_n3073 | new_n3074;
  assign new_n3076 = ~new_n2572 & ~address1;
  assign new_n3077 = ~new_n2569 & address1;
  assign result33 = new_n3076 | new_n3077;
  assign new_n3079 = ~new_n2579 & ~address1;
  assign new_n3080 = ~new_n2576 & address1;
  assign result34 = new_n3079 | new_n3080;
  assign new_n3082 = ~new_n2596 & ~address1;
  assign new_n3083 = ~new_n2593 & address1;
  assign result35 = new_n3082 | new_n3083;
  assign new_n3085 = ~new_n2600 & ~address1;
  assign new_n3086 = ~new_n2603 & address1;
  assign result36 = new_n3085 | new_n3086;
  assign new_n3088 = ~new_n2587 & ~address1;
  assign new_n3089 = ~new_n2584 & address1;
  assign result37 = new_n3088 | new_n3089;
  assign new_n3091 = ~new_n2243 & ~address1;
  assign new_n3092 = ~new_n2246 & address1;
  assign result38 = new_n3091 | new_n3092;
  assign new_n3094 = ~new_n2614 & ~address1;
  assign new_n3095 = ~new_n2617 & address1;
  assign result39 = new_n3094 | new_n3095;
  assign new_n3097 = ~new_n2239 & ~address1;
  assign new_n3098 = ~new_n2236 & address1;
  assign result40 = new_n3097 | new_n3098;
  assign new_n3100 = ~new_n2664 & ~address1;
  assign new_n3101 = ~new_n2661 & address1;
  assign result41 = new_n3100 | new_n3101;
  assign new_n3103 = ~new_n2641 & ~address1;
  assign new_n3104 = ~new_n2638 & address1;
  assign result42 = new_n3103 | new_n3104;
  assign new_n3106 = ~new_n2645 & ~address1;
  assign new_n3107 = ~new_n2648 & address1;
  assign result43 = new_n3106 | new_n3107;
  assign new_n3109 = ~new_n2653 & ~address1;
  assign new_n3110 = ~new_n2656 & address1;
  assign result44 = new_n3109 | new_n3110;
  assign new_n3112 = ~new_n2227 & ~address1;
  assign new_n3113 = ~new_n2230 & address1;
  assign result45 = new_n3112 | new_n3113;
  assign new_n3115 = ~new_n2220 & ~address1;
  assign new_n3116 = ~new_n2223 & address1;
  assign result46 = new_n3115 | new_n3116;
  assign new_n3118 = ~new_n2216 & ~address1;
  assign new_n3119 = ~new_n2213 & address1;
  assign result47 = new_n3118 | new_n3119;
  assign new_n3121 = ~new_n2716 & ~address1;
  assign new_n3122 = ~new_n2719 & address1;
  assign result48 = new_n3121 | new_n3122;
  assign new_n3124 = ~new_n2698 & ~address1;
  assign new_n3125 = ~new_n2701 & address1;
  assign result49 = new_n3124 | new_n3125;
  assign new_n3127 = ~new_n2694 & address1;
  assign new_n3128 = ~new_n2691 & ~address1;
  assign result50 = new_n3127 | new_n3128;
  assign new_n3130 = ~new_n2710 & ~address1;
  assign new_n3131 = ~new_n2707 & address1;
  assign result51 = new_n3130 | new_n3131;
  assign new_n3133 = ~new_n2206 & ~address1;
  assign new_n3134 = ~new_n2209 & address1;
  assign result52 = new_n3133 | new_n3134;
  assign new_n3136 = ~new_n2202 & ~address1;
  assign new_n3137 = ~new_n2199 & address1;
  assign result53 = new_n3136 | new_n3137;
  assign new_n3139 = ~new_n2187 & ~address1;
  assign new_n3140 = ~new_n2184 & address1;
  assign result54 = new_n3139 | new_n3140;
  assign new_n3142 = ~new_n2191 & ~address1;
  assign new_n3143 = ~new_n2194 & address1;
  assign result55 = new_n3142 | new_n3143;
  assign new_n3145 = ~new_n2180 & ~address1;
  assign new_n3146 = ~new_n2177 & address1;
  assign result56 = new_n3145 | new_n3146;
  assign new_n3148 = ~new_n2770 & ~address1;
  assign new_n3149 = ~new_n2767 & address1;
  assign result57 = new_n3148 | new_n3149;
  assign new_n3151 = ~new_n2747 & ~address1;
  assign new_n3152 = ~new_n2744 & address1;
  assign result58 = new_n3151 | new_n3152;
  assign new_n3154 = ~new_n2754 & ~address1;
  assign new_n3155 = ~new_n2751 & address1;
  assign result59 = new_n3154 | new_n3155;
  assign new_n3157 = ~new_n2763 & ~address1;
  assign new_n3158 = ~new_n2760 & address1;
  assign result60 = new_n3157 | new_n3158;
  assign new_n3160 = ~new_n2172 & ~address1;
  assign new_n3161 = ~new_n2169 & address1;
  assign result61 = new_n3160 | new_n3161;
  assign new_n3163 = ~new_n2163 & ~address1;
  assign new_n3164 = ~new_n2160 & address1;
  assign result62 = new_n3163 | new_n3164;
  assign new_n3166 = ~new_n2156 & ~address1;
  assign new_n3167 = ~new_n2153 & address1;
  assign result63 = new_n3166 | new_n3167;
  assign new_n3169 = ~new_n2145 & ~address1;
  assign new_n3170 = ~new_n2148 & address1;
  assign result64 = new_n3169 | new_n3170;
  assign new_n3172 = ~new_n2137 & ~address1;
  assign new_n3173 = ~new_n2140 & address1;
  assign result65 = new_n3172 | new_n3173;
  assign new_n3175 = ~new_n2131 & address1;
  assign new_n3176 = ~new_n2128 & ~address1;
  assign result66 = new_n3175 | new_n3176;
  assign new_n3178 = ~new_n2124 & address1;
  assign new_n3179 = ~new_n2121 & ~address1;
  assign result67 = new_n3178 | new_n3179;
  assign new_n3181 = ~new_n2113 & ~address1;
  assign new_n3182 = ~new_n2116 & address1;
  assign result68 = new_n3181 | new_n3182;
  assign new_n3184 = ~new_n2105 & ~address1;
  assign new_n3185 = ~new_n2108 & address1;
  assign result69 = new_n3184 | new_n3185;
  assign new_n3187 = ~new_n2099 & ~address1;
  assign new_n3188 = ~new_n2096 & address1;
  assign result70 = new_n3187 | new_n3188;
  assign new_n3190 = ~new_n2092 & ~address1;
  assign new_n3191 = ~new_n2089 & address1;
  assign result71 = new_n3190 | new_n3191;
  assign new_n3193 = ~new_n2081 & ~address1;
  assign new_n3194 = ~new_n2084 & address1;
  assign result72 = new_n3193 | new_n3194;
  assign new_n3196 = ~new_n2076 & ~address1;
  assign new_n3197 = ~new_n2073 & address1;
  assign result73 = new_n3196 | new_n3197;
  assign new_n3199 = ~new_n2067 & ~address1;
  assign new_n3200 = ~new_n2064 & address1;
  assign result74 = new_n3199 | new_n3200;
  assign new_n3202 = ~new_n2057 & ~address1;
  assign new_n3203 = ~new_n2060 & address1;
  assign result75 = new_n3202 | new_n3203;
  assign new_n3205 = ~new_n2052 & ~address1;
  assign new_n3206 = ~new_n2049 & address1;
  assign result76 = new_n3205 | new_n3206;
  assign new_n3208 = ~new_n2041 & ~address1;
  assign new_n3209 = ~new_n2044 & address1;
  assign result77 = new_n3208 | new_n3209;
  assign new_n3211 = ~new_n2035 & ~address1;
  assign new_n3212 = ~new_n2032 & address1;
  assign result78 = new_n3211 | new_n3212;
  assign new_n3214 = ~new_n2028 & ~address1;
  assign new_n3215 = ~new_n2025 & address1;
  assign result79 = new_n3214 | new_n3215;
  assign new_n3217 = ~new_n2017 & ~address1;
  assign new_n3218 = ~new_n2020 & address1;
  assign result80 = new_n3217 | new_n3218;
  assign new_n3220 = ~new_n2012 & ~address1;
  assign new_n3221 = ~new_n2009 & address1;
  assign result81 = new_n3220 | new_n3221;
  assign new_n3223 = ~new_n2003 & ~address1;
  assign new_n3224 = ~new_n2000 & address1;
  assign result82 = new_n3223 | new_n3224;
  assign new_n3226 = ~new_n1992 & ~address1;
  assign new_n3227 = ~new_n1995 & address1;
  assign result83 = new_n3226 | new_n3227;
  assign new_n3229 = ~new_n1985 & ~address1;
  assign new_n3230 = ~new_n1988 & address1;
  assign result84 = new_n3229 | new_n3230;
  assign new_n3232 = ~new_n1976 & ~address1;
  assign new_n3233 = ~new_n1979 & address1;
  assign result85 = new_n3232 | new_n3233;
  assign new_n3235 = ~new_n1969 & ~address1;
  assign new_n3236 = ~new_n1972 & address1;
  assign result86 = new_n3235 | new_n3236;
  assign new_n3238 = ~new_n1961 & ~address1;
  assign new_n3239 = ~new_n1964 & address1;
  assign result87 = new_n3238 | new_n3239;
  assign new_n3241 = ~new_n1953 & ~address1;
  assign new_n3242 = ~new_n1956 & address1;
  assign result88 = new_n3241 | new_n3242;
  assign new_n3244 = ~new_n1948 & address1;
  assign new_n3245 = ~new_n1945 & ~address1;
  assign result89 = new_n3244 | new_n3245;
  assign new_n3247 = ~new_n1940 & ~address1;
  assign new_n3248 = ~new_n1937 & address1;
  assign result90 = new_n3247 | new_n3248;
  assign new_n3250 = ~new_n1931 & ~address1;
  assign new_n3251 = ~new_n1928 & address1;
  assign result91 = new_n3250 | new_n3251;
  assign new_n3253 = ~new_n1924 & ~address1;
  assign new_n3254 = ~new_n1921 & address1;
  assign result92 = new_n3253 | new_n3254;
  assign new_n3256 = ~new_n1913 & ~address1;
  assign new_n3257 = ~new_n1916 & address1;
  assign result93 = new_n3256 | new_n3257;
  assign new_n3259 = ~new_n1905 & ~address1;
  assign new_n3260 = ~new_n1908 & address1;
  assign result94 = new_n3259 | new_n3260;
  assign new_n3262 = ~new_n1900 & ~address1;
  assign new_n3263 = ~new_n1897 & address1;
  assign result95 = new_n3262 | new_n3263;
  assign new_n3265 = ~new_n1892 & ~address1;
  assign new_n3266 = ~new_n1889 & address1;
  assign result96 = new_n3265 | new_n3266;
  assign new_n3268 = ~new_n1883 & ~address1;
  assign new_n3269 = ~new_n1880 & address1;
  assign result97 = new_n3268 | new_n3269;
  assign new_n3271 = ~new_n1876 & ~address1;
  assign new_n3272 = ~new_n1873 & address1;
  assign result98 = new_n3271 | new_n3272;
  assign new_n3274 = ~new_n1865 & ~address1;
  assign new_n3275 = ~new_n1868 & address1;
  assign result99 = new_n3274 | new_n3275;
  assign new_n3277 = ~new_n1856 & ~address1;
  assign new_n3278 = ~new_n1859 & address1;
  assign result100 = new_n3277 | new_n3278;
  assign new_n3280 = ~new_n1852 & ~address1;
  assign new_n3281 = ~new_n1849 & address1;
  assign result101 = new_n3280 | new_n3281;
  assign new_n3283 = ~new_n1843 & ~address1;
  assign new_n3284 = ~new_n1840 & address1;
  assign result102 = new_n3283 | new_n3284;
  assign new_n3286 = ~new_n1833 & ~address1;
  assign new_n3287 = ~new_n1836 & address1;
  assign result103 = new_n3286 | new_n3287;
  assign new_n3289 = ~new_n1827 & ~address1;
  assign new_n3290 = ~new_n1824 & address1;
  assign result104 = new_n3289 | new_n3290;
  assign new_n3292 = ~new_n1817 & ~address1;
  assign new_n3293 = ~new_n1820 & address1;
  assign result105 = new_n3292 | new_n3293;
  assign new_n3295 = ~new_n1811 & ~address1;
  assign new_n3296 = ~new_n1808 & address1;
  assign result106 = new_n3295 | new_n3296;
  assign new_n3298 = ~new_n1801 & ~address1;
  assign new_n3299 = ~new_n1804 & address1;
  assign result107 = new_n3298 | new_n3299;
  assign new_n3301 = ~new_n1795 & ~address1;
  assign new_n3302 = ~new_n1792 & address1;
  assign result108 = new_n3301 | new_n3302;
  assign new_n3304 = ~new_n1785 & ~address1;
  assign new_n3305 = ~new_n1788 & address1;
  assign result109 = new_n3304 | new_n3305;
  assign new_n3307 = ~new_n2892 & ~address1;
  assign new_n3308 = ~new_n2889 & address1;
  assign result110 = new_n3307 | new_n3308;
  assign new_n3310 = ~new_n2899 & ~address1;
  assign new_n3311 = ~new_n2896 & address1;
  assign result111 = new_n3310 | new_n3311;
  assign new_n3313 = ~new_n2909 & ~address1;
  assign new_n3314 = ~new_n2906 & address1;
  assign result112 = new_n3313 | new_n3314;
  assign new_n3316 = ~new_n1781 & ~address1;
  assign new_n3317 = ~new_n1778 & address1;
  assign result113 = new_n3316 | new_n3317;
  assign new_n3319 = ~new_n1772 & ~address1;
  assign new_n3320 = ~new_n1769 & address1;
  assign result114 = new_n3319 | new_n3320;
  assign new_n3322 = ~new_n1765 & ~address1;
  assign new_n3323 = ~new_n1762 & address1;
  assign result115 = new_n3322 | new_n3323;
  assign new_n3325 = ~new_n1756 & ~address1;
  assign new_n3326 = ~new_n1753 & address1;
  assign result116 = new_n3325 | new_n3326;
  assign new_n3328 = ~new_n1746 & ~address1;
  assign new_n3329 = ~new_n1749 & address1;
  assign result117 = new_n3328 | new_n3329;
  assign new_n3331 = ~new_n2934 & address1;
  assign new_n3332 = ~new_n2931 & ~address1;
  assign result118 = new_n3331 | new_n3332;
  assign new_n3334 = ~new_n2941 & ~address1;
  assign new_n3335 = ~new_n2938 & address1;
  assign result119 = new_n3334 | new_n3335;
  assign new_n3337 = ~new_n2951 & ~address1;
  assign new_n3338 = ~new_n2948 & address1;
  assign result120 = new_n3337 | new_n3338;
  assign new_n3340 = ~new_n1741 & ~address1;
  assign new_n3341 = ~new_n1738 & address1;
  assign result121 = new_n3340 | new_n3341;
  assign new_n3343 = ~new_n1734 & ~address1;
  assign new_n3344 = ~new_n1731 & address1;
  assign result122 = new_n3343 | new_n3344;
  assign new_n3346 = ~new_n1727 & ~address1;
  assign new_n3347 = ~new_n1724 & address1;
  assign result123 = new_n3346 | new_n3347;
  assign new_n3349 = ~new_n1716 & ~address1;
  assign new_n3350 = ~new_n1713 & address1;
  assign result124 = new_n3349 | new_n3350;
  assign new_n3352 = ~new_n1708 & ~address1;
  assign new_n3353 = ~new_n1705 & address1;
  assign result125 = new_n3352 | new_n3353;
  assign new_n3355 = ~new_n1700 & ~address1;
  assign new_n3356 = ~new_n1697 & address1;
  assign result126 = new_n3355 | new_n3356;
  assign result127 = new_n1171 & new_n1172;
  assign new_n3359 = new_n1167 & ~address1;
  assign new_n3360 = new_n1694 & address1;
  assign address0 = new_n3359 | new_n3360;
endmodule


