module c7552 ( 
    \1 , 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50, 53, 54,
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74, 75, 76,
    77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97, 100, 103,
    106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127, 130, 133,
    134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155, 156, 157,
    158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171,
    172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185,
    186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199,
    200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213,
    214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227,
    228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241,
    242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277, 280, 283,
    286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322, 325, 328,
    331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364, 367, 382,
    387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342  );
  input  \1 , 5, 9, 12, 15, 18, 23, 26, 29, 32, 35, 38, 41, 44, 47, 50,
    53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 69, 70, 73, 74,
    75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 94, 97,
    100, 103, 106, 109, 110, 111, 112, 113, 114, 115, 118, 121, 124, 127,
    130, 133, 134, 135, 138, 141, 144, 147, 150, 151, 152, 153, 154, 155,
    156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169,
    170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183,
    184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197,
    198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211,
    212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225,
    226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239,
    240, 241, 242, 245, 248, 251, 254, 257, 260, 263, 267, 271, 274, 277,
    280, 283, 286, 289, 293, 296, 299, 303, 307, 310, 313, 316, 319, 322,
    325, 328, 331, 334, 337, 340, 343, 346, 349, 352, 355, 358, 361, 364,
    367, 382;
  output 387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342;
  wire n317, n318, n320, n321, n323, n324, n326, n327, n330, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1218, n1219,
    n1220, n1221, n1222, n1224, n1225, n1226, n1227, n1228, n1229, n1231,
    n1232, n1233, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1273, n1274, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1710,
    n1711, n1712, n1713, n1715, n1716, n1717, n1718, n1719, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766,
    n1767, n1768, n1769, n1771, n1772, n1773, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1791, n1792, n1793, n1794, n1795, n1797, n1798, n1799, n1800,
    n1801, n1802, n1804, n1805, n1806, n1808, n1809, n1810, n1811, n1812,
    n1814, n1815, n1816, n1817, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1857,
    n1858, n1860, n1861, n1862, n1863, n1864, n1865, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1877, n1878, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1896, n1897, n1898, n1899, n1900, n1902, n1903,
    n1904, n1905, n1906, n1907, n1909, n1910, n1911, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1951, n1952, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388;
  assign 881 = 5 | 57;
  assign n317 = 150 & 184;
  assign n318 = 228 & n317;
  assign 882 = ~240 | ~n318;
  assign n320 = 152 & 210;
  assign n321 = 218 & n320;
  assign 883 = ~230 | ~n321;
  assign n323 = 182 & 183;
  assign n324 = 185 & n323;
  assign 884 = ~186 | ~n324;
  assign n326 = 162 & 172;
  assign n327 = 188 & n326;
  assign 885 = ~199 | ~n327;
  assign 1110 = 5 | ~242;
  assign n330 = 133 & 134;
  assign 1113 = 5 | ~n330;
  assign 1781 = \1  & 163;
  assign n333 = 18 & 229;
  assign n334 = ~18 & 41;
  assign n335 = ~n333 & ~n334;
  assign n336 = ~18 & ~n335;
  assign n337 = ~18 & ~310;
  assign n338 = ~18 & ~n337;
  assign n339 = n336 & n338;
  assign n340 = ~n336 & ~n338;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~367 & ~n341;
  assign n343 = 367 & n341;
  assign 10025 = n342 | n343;
  assign n345 = 267 & 382;
  assign n346 = 38 & ~n345;
  assign n347 = 38 & n345;
  assign n348 = ~38 & ~n345;
  assign n349 = ~n347 & ~n348;
  assign n350 = 263 & 382;
  assign n351 = 38 & ~n350;
  assign n352 = ~n349 & n351;
  assign n353 = ~n346 & ~n352;
  assign n354 = 18 & 213;
  assign n355 = 18 & ~n354;
  assign n356 = 9 & 12;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~260 & n357;
  assign n359 = 260 & n357;
  assign n360 = ~260 & ~n357;
  assign n361 = ~n359 & ~n360;
  assign n362 = 18 & 214;
  assign n363 = 18 & ~n362;
  assign n364 = ~n356 & ~n363;
  assign n365 = ~257 & n364;
  assign n366 = ~n361 & n365;
  assign n367 = 257 & n364;
  assign n368 = ~257 & ~n364;
  assign n369 = ~n367 & ~n368;
  assign n370 = 18 & 215;
  assign n371 = 18 & ~n370;
  assign n372 = ~n356 & ~n371;
  assign n373 = ~106 & n372;
  assign n374 = ~n361 & ~n369;
  assign n375 = n373 & n374;
  assign n376 = 106 & n372;
  assign n377 = ~106 & ~n372;
  assign n378 = ~n376 & ~n377;
  assign n379 = 18 & 216;
  assign n380 = 18 & ~n379;
  assign n381 = ~n356 & ~n380;
  assign n382 = ~254 & n381;
  assign n383 = ~n361 & ~n378;
  assign n384 = n382 & n383;
  assign n385 = ~n369 & n384;
  assign n386 = 254 & n381;
  assign n387 = ~254 & ~n381;
  assign n388 = ~n386 & ~n387;
  assign n389 = 18 & 209;
  assign n390 = 18 & ~n389;
  assign n391 = ~n356 & ~n390;
  assign n392 = ~251 & n391;
  assign n393 = ~n378 & ~n388;
  assign n394 = ~n361 & n393;
  assign n395 = n392 & n394;
  assign n396 = ~n369 & n395;
  assign n397 = ~n358 & ~n366;
  assign n398 = ~n375 & n397;
  assign n399 = ~n385 & n398;
  assign n400 = ~n396 & n399;
  assign n401 = 38 & n350;
  assign n402 = ~38 & ~n350;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n349 & ~n403;
  assign n405 = ~n400 & n404;
  assign n406 = n353 & ~n405;
  assign n407 = 18 & 153;
  assign n408 = 18 & ~n407;
  assign n409 = ~n356 & ~n408;
  assign n410 = ~303 & n409;
  assign n411 = 303 & n409;
  assign n412 = ~303 & ~n409;
  assign n413 = ~n411 & ~n412;
  assign n414 = 18 & 154;
  assign n415 = 18 & ~n414;
  assign n416 = ~n356 & ~n415;
  assign n417 = ~299 & n416;
  assign n418 = ~n413 & n417;
  assign n419 = 299 & n416;
  assign n420 = ~299 & ~n416;
  assign n421 = ~n419 & ~n420;
  assign n422 = 18 & 155;
  assign n423 = 18 & ~n422;
  assign n424 = ~n356 & ~n423;
  assign n425 = ~296 & n424;
  assign n426 = ~n413 & ~n421;
  assign n427 = n425 & n426;
  assign n428 = 296 & n424;
  assign n429 = ~296 & ~n424;
  assign n430 = ~n428 & ~n429;
  assign n431 = 18 & 156;
  assign n432 = 18 & ~n431;
  assign n433 = ~n356 & ~n432;
  assign n434 = ~293 & n433;
  assign n435 = ~n413 & ~n430;
  assign n436 = n434 & n435;
  assign n437 = ~n421 & n436;
  assign n438 = ~n410 & ~n418;
  assign n439 = ~n427 & n438;
  assign n440 = ~n437 & n439;
  assign n441 = 18 & 157;
  assign n442 = 18 & ~n441;
  assign n443 = ~n356 & ~n442;
  assign n444 = ~289 & n443;
  assign n445 = 289 & n443;
  assign n446 = ~289 & ~n443;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~18 & 135;
  assign n449 = 18 & 158;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~286 & ~n450;
  assign n452 = ~n447 & n451;
  assign n453 = 286 & ~n450;
  assign n454 = ~286 & n450;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~18 & 144;
  assign n457 = 18 & 159;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~283 & ~n458;
  assign n460 = ~n447 & ~n455;
  assign n461 = n459 & n460;
  assign n462 = 283 & ~n458;
  assign n463 = ~283 & n458;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~18 & 138;
  assign n466 = 18 & 160;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~280 & ~n467;
  assign n469 = ~n447 & ~n464;
  assign n470 = n468 & n469;
  assign n471 = ~n455 & n470;
  assign n472 = 280 & ~n467;
  assign n473 = ~280 & n467;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~18 & 147;
  assign n476 = 18 & 151;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~277 & ~n477;
  assign n479 = ~n464 & ~n474;
  assign n480 = ~n447 & n479;
  assign n481 = n478 & n480;
  assign n482 = ~n455 & n481;
  assign n483 = ~n444 & ~n452;
  assign n484 = ~n461 & n483;
  assign n485 = ~n471 & n484;
  assign n486 = ~n482 & n485;
  assign n487 = 293 & n433;
  assign n488 = ~293 & ~n433;
  assign n489 = ~n487 & ~n488;
  assign n490 = ~n421 & ~n489;
  assign n491 = ~n430 & n490;
  assign n492 = ~n413 & n491;
  assign n493 = ~n486 & n492;
  assign n494 = n440 & ~n493;
  assign n495 = 251 & n391;
  assign n496 = ~251 & ~n391;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n369 & ~n497;
  assign n499 = ~n378 & n498;
  assign n500 = ~n361 & n499;
  assign n501 = ~n388 & n500;
  assign n502 = n404 & n501;
  assign n503 = ~n494 & n502;
  assign n504 = 18 & 219;
  assign n505 = ~18 & 66;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~364 & ~n506;
  assign n508 = 364 & ~n506;
  assign n509 = ~364 & n506;
  assign n510 = ~n508 & ~n509;
  assign n511 = 18 & 220;
  assign n512 = ~18 & 50;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~361 & ~n513;
  assign n515 = ~n510 & n514;
  assign n516 = 361 & ~n513;
  assign n517 = ~361 & n513;
  assign n518 = ~n516 & ~n517;
  assign n519 = 18 & 221;
  assign n520 = ~18 & 32;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~358 & ~n521;
  assign n523 = ~n510 & ~n518;
  assign n524 = n522 & n523;
  assign n525 = 358 & ~n521;
  assign n526 = ~358 & n521;
  assign n527 = ~n525 & ~n526;
  assign n528 = 18 & 222;
  assign n529 = ~18 & 35;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~355 & ~n530;
  assign n532 = ~n510 & ~n527;
  assign n533 = n531 & n532;
  assign n534 = ~n518 & n533;
  assign n535 = ~n507 & ~n515;
  assign n536 = ~n524 & n535;
  assign n537 = ~n534 & n536;
  assign n538 = 18 & 223;
  assign n539 = ~18 & 47;
  assign n540 = ~n538 & ~n539;
  assign n541 = ~352 & ~n540;
  assign n542 = 352 & ~n540;
  assign n543 = ~352 & n540;
  assign n544 = ~n542 & ~n543;
  assign n545 = 18 & 224;
  assign n546 = ~18 & 121;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~349 & ~n547;
  assign n549 = ~n544 & n548;
  assign n550 = 349 & ~n547;
  assign n551 = ~349 & n547;
  assign n552 = ~n550 & ~n551;
  assign n553 = 18 & 225;
  assign n554 = ~18 & 94;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~346 & ~n555;
  assign n557 = ~n544 & ~n552;
  assign n558 = n556 & n557;
  assign n559 = 346 & ~n555;
  assign n560 = ~346 & n555;
  assign n561 = ~n559 & ~n560;
  assign n562 = 18 & 226;
  assign n563 = ~18 & 97;
  assign n564 = ~n562 & ~n563;
  assign n565 = ~343 & ~n564;
  assign n566 = ~n544 & ~n561;
  assign n567 = n565 & n566;
  assign n568 = ~n552 & n567;
  assign n569 = 343 & ~n564;
  assign n570 = ~343 & n564;
  assign n571 = ~n569 & ~n570;
  assign n572 = 18 & 217;
  assign n573 = ~18 & 118;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~340 & ~n574;
  assign n576 = ~n561 & ~n571;
  assign n577 = ~n544 & n576;
  assign n578 = n575 & n577;
  assign n579 = ~n552 & n578;
  assign n580 = ~n541 & ~n549;
  assign n581 = ~n558 & n580;
  assign n582 = ~n568 & n581;
  assign n583 = ~n579 & n582;
  assign n584 = 355 & ~n530;
  assign n585 = ~355 & n530;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n518 & ~n586;
  assign n588 = ~n527 & n587;
  assign n589 = ~n510 & n588;
  assign n590 = ~n583 & n589;
  assign n591 = n537 & ~n590;
  assign n592 = 277 & ~n477;
  assign n593 = ~277 & n477;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n455 & ~n594;
  assign n596 = ~n464 & n595;
  assign n597 = ~n447 & n596;
  assign n598 = ~n474 & n597;
  assign n599 = n492 & n598;
  assign n600 = ~n591 & n599;
  assign n601 = n502 & n600;
  assign n602 = 18 & 231;
  assign n603 = ~18 & 100;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~334 & ~n604;
  assign n606 = 334 & ~n604;
  assign n607 = ~334 & n604;
  assign n608 = ~n606 & ~n607;
  assign n609 = 18 & 232;
  assign n610 = ~18 & 124;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~331 & ~n611;
  assign n613 = ~n608 & n612;
  assign n614 = 331 & ~n611;
  assign n615 = ~331 & n611;
  assign n616 = ~n614 & ~n615;
  assign n617 = 18 & 233;
  assign n618 = ~18 & 127;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~328 & ~n619;
  assign n621 = ~n608 & ~n616;
  assign n622 = n620 & n621;
  assign n623 = 328 & ~n619;
  assign n624 = ~328 & n619;
  assign n625 = ~n623 & ~n624;
  assign n626 = 18 & 234;
  assign n627 = ~18 & 130;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~325 & ~n628;
  assign n630 = ~n608 & ~n625;
  assign n631 = n629 & n630;
  assign n632 = ~n616 & n631;
  assign n633 = ~n605 & ~n613;
  assign n634 = ~n622 & n633;
  assign n635 = ~n632 & n634;
  assign n636 = 18 & 235;
  assign n637 = ~18 & 103;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~322 & ~n638;
  assign n640 = 322 & ~n638;
  assign n641 = ~322 & n638;
  assign n642 = ~n640 & ~n641;
  assign n643 = 18 & 236;
  assign n644 = ~18 & 23;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~319 & ~n645;
  assign n647 = ~n642 & n646;
  assign n648 = 319 & ~n645;
  assign n649 = ~319 & n645;
  assign n650 = ~n648 & ~n649;
  assign n651 = 18 & 237;
  assign n652 = ~18 & 26;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~316 & ~n653;
  assign n655 = ~n642 & ~n650;
  assign n656 = n654 & n655;
  assign n657 = 316 & ~n653;
  assign n658 = ~316 & n653;
  assign n659 = ~n657 & ~n658;
  assign n660 = 18 & 238;
  assign n661 = ~18 & 29;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~313 & ~n662;
  assign n664 = ~n642 & ~n659;
  assign n665 = n663 & n664;
  assign n666 = ~n650 & n665;
  assign n667 = 313 & ~n662;
  assign n668 = ~313 & n662;
  assign n669 = ~n667 & ~n668;
  assign n670 = n336 & ~n338;
  assign n671 = ~n659 & ~n669;
  assign n672 = ~n642 & n671;
  assign n673 = n670 & n672;
  assign n674 = ~n650 & n673;
  assign n675 = ~n639 & ~n647;
  assign n676 = ~n656 & n675;
  assign n677 = ~n666 & n676;
  assign n678 = ~n674 & n677;
  assign n679 = 325 & ~n628;
  assign n680 = ~325 & n628;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~n616 & ~n681;
  assign n683 = ~n625 & n682;
  assign n684 = ~n608 & n683;
  assign n685 = ~n678 & n684;
  assign n686 = n635 & ~n685;
  assign n687 = 340 & ~n574;
  assign n688 = ~340 & n574;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~n552 & ~n689;
  assign n691 = ~n561 & n690;
  assign n692 = ~n544 & n691;
  assign n693 = ~n571 & n692;
  assign n694 = n589 & n693;
  assign n695 = ~n686 & n694;
  assign n696 = n599 & n695;
  assign n697 = n502 & n696;
  assign n698 = ~n341 & ~n650;
  assign n699 = ~n659 & n698;
  assign n700 = ~n642 & n699;
  assign n701 = ~n669 & n700;
  assign n702 = n684 & n701;
  assign n703 = 367 & n702;
  assign n704 = n694 & n703;
  assign n705 = n599 & n704;
  assign n706 = n502 & n705;
  assign n707 = n406 & ~n503;
  assign n708 = ~n601 & n707;
  assign n709 = ~n697 & n708;
  assign 10101 = n706 | ~n709;
  assign n711 = ~271 & 382;
  assign n712 = 38 & ~n711;
  assign n713 = 38 & n711;
  assign n714 = ~38 & ~n711;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~245 & 382;
  assign n717 = 38 & ~n716;
  assign n718 = ~n715 & n717;
  assign n719 = ~n712 & ~n718;
  assign n720 = 38 & n716;
  assign n721 = ~38 & ~n716;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~n715 & ~n722;
  assign n724 = ~18 & 88;
  assign n725 = 18 & ~260;
  assign n726 = ~n724 & ~n725;
  assign n727 = 18 & 166;
  assign n728 = 18 & ~n727;
  assign n729 = ~n356 & ~n728;
  assign n730 = ~n726 & n729;
  assign n731 = n726 & n729;
  assign n732 = ~n726 & ~n729;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~18 & 112;
  assign n735 = 18 & ~257;
  assign n736 = ~n734 & ~n735;
  assign n737 = 18 & 167;
  assign n738 = 18 & ~n737;
  assign n739 = ~n356 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = ~n733 & n740;
  assign n742 = n736 & n739;
  assign n743 = ~n736 & ~n739;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~18 & 87;
  assign n746 = 18 & ~106;
  assign n747 = ~n745 & ~n746;
  assign n748 = 18 & 168;
  assign n749 = 18 & ~n748;
  assign n750 = ~n356 & ~n749;
  assign n751 = ~n747 & n750;
  assign n752 = ~n733 & ~n744;
  assign n753 = n751 & n752;
  assign n754 = n747 & n750;
  assign n755 = ~n747 & ~n750;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~18 & 111;
  assign n758 = 18 & ~254;
  assign n759 = ~n757 & ~n758;
  assign n760 = 18 & 169;
  assign n761 = 18 & ~n760;
  assign n762 = ~n356 & ~n761;
  assign n763 = ~n759 & n762;
  assign n764 = ~n733 & ~n756;
  assign n765 = n763 & n764;
  assign n766 = ~n744 & n765;
  assign n767 = n759 & n762;
  assign n768 = ~n759 & ~n762;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~18 & 113;
  assign n771 = 18 & ~251;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n356 & ~n772;
  assign n774 = ~n756 & ~n769;
  assign n775 = ~n733 & n774;
  assign n776 = n773 & n775;
  assign n777 = ~n744 & n776;
  assign n778 = ~n730 & ~n741;
  assign n779 = ~n753 & n778;
  assign n780 = ~n766 & n779;
  assign n781 = ~n777 & n780;
  assign n782 = n723 & ~n781;
  assign n783 = n719 & ~n782;
  assign n784 = ~18 & 110;
  assign n785 = 18 & ~303;
  assign n786 = ~n784 & ~n785;
  assign n787 = 18 & 173;
  assign n788 = 18 & ~n787;
  assign n789 = ~n356 & ~n788;
  assign n790 = ~n786 & n789;
  assign n791 = n786 & n789;
  assign n792 = ~n786 & ~n789;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~18 & 109;
  assign n795 = 18 & ~299;
  assign n796 = ~n794 & ~n795;
  assign n797 = 18 & 174;
  assign n798 = 18 & ~n797;
  assign n799 = ~n356 & ~n798;
  assign n800 = ~n796 & n799;
  assign n801 = ~n793 & n800;
  assign n802 = n796 & n799;
  assign n803 = ~n796 & ~n799;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~18 & 86;
  assign n806 = 18 & ~296;
  assign n807 = ~n805 & ~n806;
  assign n808 = 18 & 175;
  assign n809 = 18 & ~n808;
  assign n810 = ~n356 & ~n809;
  assign n811 = ~n807 & n810;
  assign n812 = ~n793 & ~n804;
  assign n813 = n811 & n812;
  assign n814 = n807 & n810;
  assign n815 = ~n807 & ~n810;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~18 & 63;
  assign n818 = 18 & ~293;
  assign n819 = ~n817 & ~n818;
  assign n820 = 18 & 176;
  assign n821 = 18 & ~n820;
  assign n822 = ~n356 & ~n821;
  assign n823 = ~n819 & n822;
  assign n824 = ~n793 & ~n816;
  assign n825 = n823 & n824;
  assign n826 = ~n804 & n825;
  assign n827 = ~n790 & ~n801;
  assign n828 = ~n813 & n827;
  assign n829 = ~n826 & n828;
  assign n830 = n819 & n822;
  assign n831 = ~n819 & ~n822;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n816 & ~n832;
  assign n834 = ~n804 & n833;
  assign n835 = ~n793 & n834;
  assign n836 = ~18 & 64;
  assign n837 = 18 & ~289;
  assign n838 = ~n836 & ~n837;
  assign n839 = 18 & 177;
  assign n840 = 18 & ~n839;
  assign n841 = ~n356 & ~n840;
  assign n842 = ~n838 & n841;
  assign n843 = n838 & n841;
  assign n844 = ~n838 & ~n841;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~18 & 85;
  assign n847 = 18 & ~286;
  assign n848 = ~n846 & ~n847;
  assign n849 = 18 & 178;
  assign n850 = ~n448 & ~n849;
  assign n851 = ~n848 & ~n850;
  assign n852 = ~n845 & n851;
  assign n853 = n848 & ~n850;
  assign n854 = ~n848 & n850;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~18 & 84;
  assign n857 = 18 & ~283;
  assign n858 = ~n856 & ~n857;
  assign n859 = 18 & 179;
  assign n860 = ~n456 & ~n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = ~n845 & ~n855;
  assign n863 = n861 & n862;
  assign n864 = n858 & ~n860;
  assign n865 = ~n858 & n860;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~18 & 83;
  assign n868 = 18 & ~280;
  assign n869 = ~n867 & ~n868;
  assign n870 = 18 & 180;
  assign n871 = ~n465 & ~n870;
  assign n872 = ~n869 & ~n871;
  assign n873 = ~n845 & ~n866;
  assign n874 = n872 & n873;
  assign n875 = ~n855 & n874;
  assign n876 = n869 & ~n871;
  assign n877 = ~n869 & n871;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~18 & 65;
  assign n880 = 18 & ~277;
  assign n881 = ~n879 & ~n880;
  assign n882 = 18 & 171;
  assign n883 = ~n475 & ~n882;
  assign n884 = ~n881 & ~n883;
  assign n885 = ~n866 & ~n878;
  assign n886 = ~n845 & n885;
  assign n887 = n884 & n886;
  assign n888 = ~n855 & n887;
  assign n889 = ~n842 & ~n852;
  assign n890 = ~n863 & n889;
  assign n891 = ~n875 & n890;
  assign n892 = ~n888 & n891;
  assign n893 = n835 & ~n892;
  assign n894 = n829 & ~n893;
  assign n895 = ~n356 & n772;
  assign n896 = n356 & ~n772;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n769 & ~n897;
  assign n899 = ~n756 & n898;
  assign n900 = ~n744 & n899;
  assign n901 = ~n733 & n900;
  assign n902 = n723 & n901;
  assign n903 = ~n894 & n902;
  assign n904 = 18 & ~364;
  assign n905 = ~18 & 62;
  assign n906 = ~n904 & ~n905;
  assign n907 = 18 & 189;
  assign n908 = ~n505 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = n906 & ~n908;
  assign n911 = ~n906 & n908;
  assign n912 = ~n910 & ~n911;
  assign n913 = 18 & ~361;
  assign n914 = ~18 & 61;
  assign n915 = ~n913 & ~n914;
  assign n916 = 18 & 190;
  assign n917 = ~n512 & ~n916;
  assign n918 = ~n915 & ~n917;
  assign n919 = ~n912 & n918;
  assign n920 = n915 & ~n917;
  assign n921 = ~n915 & n917;
  assign n922 = ~n920 & ~n921;
  assign n923 = 18 & ~358;
  assign n924 = ~18 & 60;
  assign n925 = ~n923 & ~n924;
  assign n926 = 18 & 191;
  assign n927 = ~n520 & ~n926;
  assign n928 = ~n925 & ~n927;
  assign n929 = ~n912 & ~n922;
  assign n930 = n928 & n929;
  assign n931 = n925 & ~n927;
  assign n932 = ~n925 & n927;
  assign n933 = ~n931 & ~n932;
  assign n934 = 18 & ~355;
  assign n935 = ~18 & 79;
  assign n936 = ~n934 & ~n935;
  assign n937 = 18 & 192;
  assign n938 = ~n529 & ~n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~n912 & ~n933;
  assign n941 = n939 & n940;
  assign n942 = ~n922 & n941;
  assign n943 = ~n909 & ~n919;
  assign n944 = ~n930 & n943;
  assign n945 = ~n942 & n944;
  assign n946 = n936 & ~n938;
  assign n947 = ~n936 & n938;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~n933 & ~n948;
  assign n950 = ~n922 & n949;
  assign n951 = ~n912 & n950;
  assign n952 = 18 & ~352;
  assign n953 = ~18 & 80;
  assign n954 = ~n952 & ~n953;
  assign n955 = 18 & 193;
  assign n956 = ~n539 & ~n955;
  assign n957 = ~n954 & ~n956;
  assign n958 = n954 & ~n956;
  assign n959 = ~n954 & n956;
  assign n960 = ~n958 & ~n959;
  assign n961 = 18 & ~349;
  assign n962 = ~18 & 81;
  assign n963 = ~n961 & ~n962;
  assign n964 = 18 & 194;
  assign n965 = ~n546 & ~n964;
  assign n966 = ~n963 & ~n965;
  assign n967 = ~n960 & n966;
  assign n968 = n963 & ~n965;
  assign n969 = ~n963 & n965;
  assign n970 = ~n968 & ~n969;
  assign n971 = 18 & ~346;
  assign n972 = ~18 & 59;
  assign n973 = ~n971 & ~n972;
  assign n974 = 18 & 195;
  assign n975 = ~n554 & ~n974;
  assign n976 = ~n973 & ~n975;
  assign n977 = ~n960 & ~n970;
  assign n978 = n976 & n977;
  assign n979 = n973 & ~n975;
  assign n980 = ~n973 & n975;
  assign n981 = ~n979 & ~n980;
  assign n982 = 18 & ~343;
  assign n983 = ~18 & 78;
  assign n984 = ~n982 & ~n983;
  assign n985 = 18 & 196;
  assign n986 = ~n563 & ~n985;
  assign n987 = ~n984 & ~n986;
  assign n988 = ~n960 & ~n981;
  assign n989 = n987 & n988;
  assign n990 = ~n970 & n989;
  assign n991 = n984 & ~n986;
  assign n992 = ~n984 & n986;
  assign n993 = ~n991 & ~n992;
  assign n994 = 18 & ~340;
  assign n995 = ~18 & 77;
  assign n996 = ~n994 & ~n995;
  assign n997 = 18 & 187;
  assign n998 = ~n573 & ~n997;
  assign n999 = ~n996 & ~n998;
  assign n1000 = ~n981 & ~n993;
  assign n1001 = ~n960 & n1000;
  assign n1002 = n999 & n1001;
  assign n1003 = ~n970 & n1002;
  assign n1004 = ~n957 & ~n967;
  assign n1005 = ~n978 & n1004;
  assign n1006 = ~n990 & n1005;
  assign n1007 = ~n1003 & n1006;
  assign n1008 = n951 & ~n1007;
  assign n1009 = n945 & ~n1008;
  assign n1010 = n881 & ~n883;
  assign n1011 = ~n881 & n883;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n878 & ~n1012;
  assign n1014 = ~n866 & n1013;
  assign n1015 = ~n855 & n1014;
  assign n1016 = ~n845 & n1015;
  assign n1017 = n835 & n1016;
  assign n1018 = ~n1009 & n1017;
  assign n1019 = n902 & n1018;
  assign n1020 = 18 & ~334;
  assign n1021 = ~18 & 56;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = 18 & 200;
  assign n1024 = ~n603 & ~n1023;
  assign n1025 = ~n1022 & ~n1024;
  assign n1026 = n1022 & ~n1024;
  assign n1027 = ~n1022 & n1024;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = 18 & ~331;
  assign n1030 = ~18 & 55;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = 18 & 201;
  assign n1033 = ~n610 & ~n1032;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = ~n1028 & n1034;
  assign n1036 = n1031 & ~n1033;
  assign n1037 = ~n1031 & n1033;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = 18 & ~328;
  assign n1040 = ~18 & 54;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = 18 & 202;
  assign n1043 = ~n618 & ~n1042;
  assign n1044 = ~n1041 & ~n1043;
  assign n1045 = ~n1028 & ~n1038;
  assign n1046 = n1044 & n1045;
  assign n1047 = n1041 & ~n1043;
  assign n1048 = ~n1041 & n1043;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = 18 & ~325;
  assign n1051 = ~18 & 53;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = 18 & 203;
  assign n1054 = ~n627 & ~n1053;
  assign n1055 = ~n1052 & ~n1054;
  assign n1056 = ~n1028 & ~n1049;
  assign n1057 = n1055 & n1056;
  assign n1058 = ~n1038 & n1057;
  assign n1059 = ~n1025 & ~n1035;
  assign n1060 = ~n1046 & n1059;
  assign n1061 = ~n1058 & n1060;
  assign n1062 = n1052 & ~n1054;
  assign n1063 = ~n1052 & n1054;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n1049 & ~n1064;
  assign n1066 = ~n1038 & n1065;
  assign n1067 = ~n1028 & n1066;
  assign n1068 = 18 & ~322;
  assign n1069 = ~18 & 73;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = 18 & 204;
  assign n1072 = ~n637 & ~n1071;
  assign n1073 = ~n1070 & ~n1072;
  assign n1074 = n1070 & ~n1072;
  assign n1075 = ~n1070 & n1072;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = 18 & ~319;
  assign n1078 = ~18 & 75;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = 18 & 205;
  assign n1081 = ~n644 & ~n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign n1083 = ~n1076 & n1082;
  assign n1084 = n1079 & ~n1081;
  assign n1085 = ~n1079 & n1081;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = 18 & ~316;
  assign n1088 = ~18 & 76;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = 18 & 206;
  assign n1091 = ~n652 & ~n1090;
  assign n1092 = ~n1089 & ~n1091;
  assign n1093 = ~n1076 & ~n1086;
  assign n1094 = n1092 & n1093;
  assign n1095 = n1089 & ~n1091;
  assign n1096 = ~n1089 & n1091;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = 18 & ~313;
  assign n1099 = ~18 & 74;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = 18 & 207;
  assign n1102 = ~n661 & ~n1101;
  assign n1103 = ~n1100 & ~n1102;
  assign n1104 = ~n1076 & ~n1097;
  assign n1105 = n1103 & n1104;
  assign n1106 = ~n1086 & n1105;
  assign n1107 = n1100 & ~n1102;
  assign n1108 = ~n1100 & n1102;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~18 & 70;
  assign n1111 = ~18 & ~n1110;
  assign n1112 = 18 & 198;
  assign n1113 = ~n334 & ~n1112;
  assign n1114 = ~18 & ~n1113;
  assign n1115 = ~n1111 & n1114;
  assign n1116 = ~n1097 & ~n1109;
  assign n1117 = ~n1076 & n1116;
  assign n1118 = n1115 & n1117;
  assign n1119 = ~n1086 & n1118;
  assign n1120 = ~n1073 & ~n1083;
  assign n1121 = ~n1094 & n1120;
  assign n1122 = ~n1106 & n1121;
  assign n1123 = ~n1119 & n1122;
  assign n1124 = n1067 & ~n1123;
  assign n1125 = n1061 & ~n1124;
  assign n1126 = n996 & ~n998;
  assign n1127 = ~n996 & n998;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n993 & ~n1128;
  assign n1130 = ~n981 & n1129;
  assign n1131 = ~n970 & n1130;
  assign n1132 = ~n960 & n1131;
  assign n1133 = n951 & n1132;
  assign n1134 = ~n1125 & n1133;
  assign n1135 = n1017 & n1134;
  assign n1136 = n902 & n1135;
  assign n1137 = n1111 & n1114;
  assign n1138 = ~n1111 & ~n1114;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1109 & ~n1139;
  assign n1141 = ~n1097 & n1140;
  assign n1142 = ~n1086 & n1141;
  assign n1143 = ~n1076 & n1142;
  assign n1144 = n1067 & n1143;
  assign n1145 = 89 & n1144;
  assign n1146 = n1133 & n1145;
  assign n1147 = n1017 & n1146;
  assign n1148 = n902 & n1147;
  assign n1149 = n783 & ~n903;
  assign n1150 = ~n1019 & n1149;
  assign n1151 = ~n1136 & n1150;
  assign 10102 = n1148 | ~n1151;
  assign n1153 = ~n430 & ~n489;
  assign n1154 = ~n421 & n1153;
  assign n1155 = ~n413 & n1154;
  assign n1156 = ~n486 & n1155;
  assign n1157 = n440 & ~n1156;
  assign n1158 = ~n388 & ~n497;
  assign n1159 = ~n378 & n1158;
  assign n1160 = ~n369 & n1159;
  assign n1161 = ~n361 & n1160;
  assign n1162 = n404 & n1161;
  assign n1163 = ~n1157 & n1162;
  assign n1164 = ~n527 & ~n586;
  assign n1165 = ~n518 & n1164;
  assign n1166 = ~n510 & n1165;
  assign n1167 = ~n583 & n1166;
  assign n1168 = n537 & ~n1167;
  assign n1169 = ~n474 & ~n594;
  assign n1170 = ~n464 & n1169;
  assign n1171 = ~n455 & n1170;
  assign n1172 = ~n447 & n1171;
  assign n1173 = n1155 & n1172;
  assign n1174 = ~n1168 & n1173;
  assign n1175 = n1162 & n1174;
  assign n1176 = ~n625 & ~n681;
  assign n1177 = ~n616 & n1176;
  assign n1178 = ~n608 & n1177;
  assign n1179 = ~n678 & n1178;
  assign n1180 = n635 & ~n1179;
  assign n1181 = ~n571 & ~n689;
  assign n1182 = ~n561 & n1181;
  assign n1183 = ~n552 & n1182;
  assign n1184 = ~n544 & n1183;
  assign n1185 = n1166 & n1184;
  assign n1186 = ~n1180 & n1185;
  assign n1187 = n1173 & n1186;
  assign n1188 = n1162 & n1187;
  assign n1189 = ~n341 & ~n669;
  assign n1190 = ~n659 & n1189;
  assign n1191 = ~n650 & n1190;
  assign n1192 = ~n642 & n1191;
  assign n1193 = n1178 & n1192;
  assign n1194 = 367 & n1193;
  assign n1195 = n1185 & n1194;
  assign n1196 = n1173 & n1195;
  assign n1197 = n1162 & n1196;
  assign n1198 = n406 & ~n1163;
  assign n1199 = ~n1175 & n1198;
  assign n1200 = ~n1188 & n1199;
  assign 10104 = n1197 | ~n1200;
  assign n1202 = ~n650 & n654;
  assign n1203 = ~n659 & n663;
  assign n1204 = ~n650 & n1203;
  assign n1205 = n670 & n671;
  assign n1206 = ~n650 & n1205;
  assign n1207 = 367 & ~n341;
  assign n1208 = ~n659 & n1207;
  assign n1209 = ~n669 & n1208;
  assign n1210 = ~n650 & n1209;
  assign n1211 = ~n646 & ~n1202;
  assign n1212 = ~n1204 & n1211;
  assign n1213 = ~n1206 & n1212;
  assign n1214 = ~n1210 & n1213;
  assign n1215 = ~n642 & n1214;
  assign n1216 = n642 & ~n1214;
  assign 10109 = n1215 | n1216;
  assign n1218 = ~n654 & ~n1203;
  assign n1219 = ~n1205 & n1218;
  assign n1220 = ~n1209 & n1219;
  assign n1221 = ~n650 & n1220;
  assign n1222 = n650 & ~n1220;
  assign 10110 = n1221 | n1222;
  assign n1224 = ~n669 & n670;
  assign n1225 = ~n669 & n1207;
  assign n1226 = ~n663 & ~n1224;
  assign n1227 = ~n1225 & n1226;
  assign n1228 = ~n659 & n1227;
  assign n1229 = n659 & ~n1227;
  assign 10111 = n1228 | n1229;
  assign n1231 = ~n670 & ~n1207;
  assign n1232 = ~n669 & n1231;
  assign n1233 = n669 & ~n1231;
  assign 10112 = n1232 | n1233;
  assign n1235 = ~n616 & n620;
  assign n1236 = ~n625 & n629;
  assign n1237 = ~n616 & n1236;
  assign n1238 = ~n612 & ~n1235;
  assign n1239 = ~n1237 & n1238;
  assign n1240 = ~n608 & ~n1239;
  assign n1241 = n608 & n1239;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = 367 & n701;
  assign n1244 = n678 & ~n1243;
  assign n1245 = n1242 & n1244;
  assign n1246 = ~n1177 & n1239;
  assign n1247 = ~n608 & n1246;
  assign n1248 = n608 & ~n1246;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~n1244 & ~n1249;
  assign 10350 = n1245 | n1250;
  assign n1252 = ~n620 & ~n1236;
  assign n1253 = ~n616 & ~n1252;
  assign n1254 = n616 & n1252;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = n1244 & n1255;
  assign n1257 = ~n1176 & n1252;
  assign n1258 = ~n616 & n1257;
  assign n1259 = n616 & ~n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1244 & ~n1260;
  assign 10351 = n1256 | n1261;
  assign n1263 = ~n625 & ~n629;
  assign n1264 = n625 & n629;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = n1244 & ~n1265;
  assign n1267 = 325 & n628;
  assign n1268 = ~n625 & ~n1267;
  assign n1269 = n625 & n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1244 & n1270;
  assign 10352 = n1266 | n1271;
  assign n1273 = ~n681 & n1244;
  assign n1274 = n681 & ~n1244;
  assign 10353 = n1273 | n1274;
  assign n1276 = 18 & 212;
  assign n1277 = 18 & ~n1276;
  assign n1278 = ~n356 & ~n1277;
  assign n1279 = 18 & 211;
  assign n1280 = 18 & ~n1279;
  assign n1281 = ~n356 & ~n1280;
  assign n1282 = n1278 & ~n1281;
  assign n1283 = ~n1278 & n1281;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = n356 & ~n391;
  assign n1286 = ~n356 & n391;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~n372 & n381;
  assign n1289 = n372 & ~n381;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n357 & n364;
  assign n1292 = n357 & ~n364;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1287 & n1290;
  assign n1295 = n1293 & n1294;
  assign n1296 = n1287 & n1290;
  assign n1297 = ~n1293 & n1296;
  assign n1298 = ~n1295 & ~n1297;
  assign n1299 = n1287 & ~n1290;
  assign n1300 = n1293 & n1299;
  assign n1301 = ~n1287 & ~n1290;
  assign n1302 = ~n1293 & n1301;
  assign n1303 = ~n1300 & ~n1302;
  assign n1304 = n1298 & n1303;
  assign n1305 = ~n1284 & n1304;
  assign n1306 = n1284 & ~n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n424 & n433;
  assign n1309 = n424 & ~n433;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n409 & n416;
  assign n1312 = n409 & ~n416;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1310 & n1313;
  assign n1315 = n1310 & ~n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = ~18 & 141;
  assign n1318 = 18 & 161;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n477 & ~n1319;
  assign n1321 = ~n477 & n1319;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = n458 & ~n467;
  assign n1324 = ~n458 & n467;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = ~n443 & ~n450;
  assign n1327 = n443 & n450;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1322 & n1325;
  assign n1330 = n1328 & n1329;
  assign n1331 = n1322 & n1325;
  assign n1332 = ~n1328 & n1331;
  assign n1333 = ~n1330 & ~n1332;
  assign n1334 = n1322 & ~n1325;
  assign n1335 = n1328 & n1334;
  assign n1336 = ~n1322 & ~n1325;
  assign n1337 = ~n1328 & n1336;
  assign n1338 = ~n1335 & ~n1337;
  assign n1339 = n1333 & n1338;
  assign n1340 = ~n1316 & n1339;
  assign n1341 = n1316 & ~n1339;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n521 & ~n530;
  assign n1344 = ~n521 & n530;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = n506 & ~n513;
  assign n1347 = ~n506 & n513;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1345 & n1348;
  assign n1350 = n1345 & ~n1348;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = 18 & 227;
  assign n1353 = ~18 & 115;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = n574 & ~n1354;
  assign n1356 = ~n574 & n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = n555 & ~n564;
  assign n1359 = ~n555 & n564;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = n540 & ~n547;
  assign n1362 = ~n540 & n547;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = ~n1357 & n1360;
  assign n1365 = n1363 & n1364;
  assign n1366 = n1357 & n1360;
  assign n1367 = ~n1363 & n1366;
  assign n1368 = ~n1365 & ~n1367;
  assign n1369 = n1357 & ~n1360;
  assign n1370 = n1363 & n1369;
  assign n1371 = ~n1357 & ~n1360;
  assign n1372 = ~n1363 & n1371;
  assign n1373 = ~n1370 & ~n1372;
  assign n1374 = n1368 & n1373;
  assign n1375 = ~n1351 & n1374;
  assign n1376 = n1351 & ~n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = n619 & ~n628;
  assign n1379 = ~n619 & n628;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n604 & ~n611;
  assign n1382 = ~n604 & n611;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n1380 & n1383;
  assign n1385 = n1380 & ~n1383;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = 18 & 239;
  assign n1388 = ~18 & 44;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = n335 & ~n1389;
  assign n1391 = ~n335 & n1389;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = n653 & ~n662;
  assign n1394 = ~n653 & n662;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = n638 & ~n645;
  assign n1397 = ~n638 & n645;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1392 & n1395;
  assign n1400 = n1398 & n1399;
  assign n1401 = n1392 & n1395;
  assign n1402 = ~n1398 & n1401;
  assign n1403 = ~n1400 & ~n1402;
  assign n1404 = n1392 & ~n1395;
  assign n1405 = n1398 & n1404;
  assign n1406 = ~n1392 & ~n1395;
  assign n1407 = ~n1398 & n1406;
  assign n1408 = ~n1405 & ~n1407;
  assign n1409 = n1403 & n1408;
  assign n1410 = ~n1386 & n1409;
  assign n1411 = n1386 & ~n1409;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~n1307 & ~n1342;
  assign n1414 = ~n1377 & n1413;
  assign 10574 = n1412 | ~n1414;
  assign n1416 = ~18 & 245;
  assign n1417 = 18 & ~263;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~18 & 271;
  assign n1420 = 18 & ~267;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~n1418 & n1421;
  assign n1423 = n1418 & ~n1421;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~18 & 114;
  assign n1426 = 18 & ~248;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = n772 & ~n1427;
  assign n1429 = ~n772 & n1427;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = n747 & ~n759;
  assign n1432 = ~n747 & n759;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = n726 & ~n736;
  assign n1435 = ~n726 & n736;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1430 & n1433;
  assign n1438 = n1436 & n1437;
  assign n1439 = n1430 & n1433;
  assign n1440 = ~n1436 & n1439;
  assign n1441 = ~n1438 & ~n1440;
  assign n1442 = n1430 & ~n1433;
  assign n1443 = n1436 & n1442;
  assign n1444 = ~n1430 & ~n1433;
  assign n1445 = ~n1436 & n1444;
  assign n1446 = ~n1443 & ~n1445;
  assign n1447 = n1441 & n1446;
  assign n1448 = ~n1424 & n1447;
  assign n1449 = n1424 & ~n1447;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n807 & ~n819;
  assign n1452 = ~n807 & n819;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = n786 & ~n796;
  assign n1455 = ~n786 & n796;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1453 & n1456;
  assign n1458 = n1453 & ~n1456;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~18 & 82;
  assign n1461 = 18 & ~274;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = n881 & ~n1462;
  assign n1464 = ~n881 & n1462;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = n858 & ~n869;
  assign n1467 = ~n858 & n869;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = n838 & ~n848;
  assign n1470 = ~n838 & n848;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = ~n1465 & n1468;
  assign n1473 = n1471 & n1472;
  assign n1474 = n1465 & n1468;
  assign n1475 = ~n1471 & n1474;
  assign n1476 = ~n1473 & ~n1475;
  assign n1477 = n1465 & ~n1468;
  assign n1478 = n1471 & n1477;
  assign n1479 = ~n1465 & ~n1468;
  assign n1480 = ~n1471 & n1479;
  assign n1481 = ~n1478 & ~n1480;
  assign n1482 = n1476 & n1481;
  assign n1483 = ~n1459 & n1482;
  assign n1484 = n1459 & ~n1482;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = n925 & ~n936;
  assign n1487 = ~n925 & n936;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = n906 & ~n915;
  assign n1490 = ~n906 & n915;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n1488 & n1491;
  assign n1493 = n1488 & ~n1491;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = 18 & ~337;
  assign n1496 = ~18 & 58;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = n996 & ~n1497;
  assign n1499 = ~n996 & n1497;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = n973 & ~n984;
  assign n1502 = ~n973 & n984;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = n954 & ~n963;
  assign n1505 = ~n954 & n963;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = ~n1500 & n1503;
  assign n1508 = n1506 & n1507;
  assign n1509 = n1500 & n1503;
  assign n1510 = ~n1506 & n1509;
  assign n1511 = ~n1508 & ~n1510;
  assign n1512 = n1500 & ~n1503;
  assign n1513 = n1506 & n1512;
  assign n1514 = ~n1500 & ~n1503;
  assign n1515 = ~n1506 & n1514;
  assign n1516 = ~n1513 & ~n1515;
  assign n1517 = n1511 & n1516;
  assign n1518 = ~n1494 & n1517;
  assign n1519 = n1494 & ~n1517;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = n1041 & ~n1052;
  assign n1522 = ~n1041 & n1052;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = n1022 & ~n1031;
  assign n1525 = ~n1022 & n1031;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = ~n1523 & n1526;
  assign n1528 = n1523 & ~n1526;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = 18 & ~307;
  assign n1531 = ~18 & 69;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = 18 & ~310;
  assign n1534 = ~n1110 & ~n1533;
  assign n1535 = ~n1532 & n1534;
  assign n1536 = n1532 & ~n1534;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = n1089 & ~n1100;
  assign n1539 = ~n1089 & n1100;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = n1070 & ~n1079;
  assign n1542 = ~n1070 & n1079;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1537 & n1540;
  assign n1545 = n1543 & n1544;
  assign n1546 = n1537 & n1540;
  assign n1547 = ~n1543 & n1546;
  assign n1548 = ~n1545 & ~n1547;
  assign n1549 = n1537 & ~n1540;
  assign n1550 = n1543 & n1549;
  assign n1551 = ~n1537 & ~n1540;
  assign n1552 = ~n1543 & n1551;
  assign n1553 = ~n1550 & ~n1552;
  assign n1554 = n1548 & n1553;
  assign n1555 = ~n1529 & n1554;
  assign n1556 = n1529 & ~n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1450 & ~n1485;
  assign n1559 = ~n1520 & n1558;
  assign 10575 = n1557 | ~n1559;
  assign n1561 = 18 & 165;
  assign n1562 = 18 & ~n1561;
  assign n1563 = ~n356 & ~n1562;
  assign n1564 = 18 & 164;
  assign n1565 = 18 & ~n1564;
  assign n1566 = ~n356 & ~n1565;
  assign n1567 = n1563 & ~n1566;
  assign n1568 = ~n1563 & n1566;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = 18 & 170;
  assign n1571 = 18 & ~n1570;
  assign n1572 = ~n356 & ~n1571;
  assign n1573 = n356 & ~n1572;
  assign n1574 = ~n356 & n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n750 & n762;
  assign n1577 = n750 & ~n762;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = ~n729 & n739;
  assign n1580 = n729 & ~n739;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1575 & n1578;
  assign n1583 = n1581 & n1582;
  assign n1584 = n1575 & n1578;
  assign n1585 = ~n1581 & n1584;
  assign n1586 = ~n1583 & ~n1585;
  assign n1587 = n1575 & ~n1578;
  assign n1588 = n1581 & n1587;
  assign n1589 = ~n1575 & ~n1578;
  assign n1590 = ~n1581 & n1589;
  assign n1591 = ~n1588 & ~n1590;
  assign n1592 = n1586 & n1591;
  assign n1593 = ~n1569 & n1592;
  assign n1594 = n1569 & ~n1592;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = ~n810 & n822;
  assign n1597 = n810 & ~n822;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n789 & n799;
  assign n1600 = n789 & ~n799;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = ~n1598 & n1601;
  assign n1603 = n1598 & ~n1601;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = 18 & 181;
  assign n1606 = ~n1317 & ~n1605;
  assign n1607 = n883 & ~n1606;
  assign n1608 = ~n883 & n1606;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = n860 & ~n871;
  assign n1611 = ~n860 & n871;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~n841 & ~n850;
  assign n1614 = n841 & n850;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1609 & n1612;
  assign n1617 = n1615 & n1616;
  assign n1618 = n1609 & n1612;
  assign n1619 = ~n1615 & n1618;
  assign n1620 = ~n1617 & ~n1619;
  assign n1621 = n1609 & ~n1612;
  assign n1622 = n1615 & n1621;
  assign n1623 = ~n1609 & ~n1612;
  assign n1624 = ~n1615 & n1623;
  assign n1625 = ~n1622 & ~n1624;
  assign n1626 = n1620 & n1625;
  assign n1627 = ~n1604 & n1626;
  assign n1628 = n1604 & ~n1626;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = n927 & ~n938;
  assign n1631 = ~n927 & n938;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = n908 & ~n917;
  assign n1634 = ~n908 & n917;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n1632 & n1635;
  assign n1637 = n1632 & ~n1635;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = 18 & 197;
  assign n1640 = ~n1353 & ~n1639;
  assign n1641 = n998 & ~n1640;
  assign n1642 = ~n998 & n1640;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = n975 & ~n986;
  assign n1645 = ~n975 & n986;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = n956 & ~n965;
  assign n1648 = ~n956 & n965;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = ~n1643 & n1646;
  assign n1651 = n1649 & n1650;
  assign n1652 = n1643 & n1646;
  assign n1653 = ~n1649 & n1652;
  assign n1654 = ~n1651 & ~n1653;
  assign n1655 = n1643 & ~n1646;
  assign n1656 = n1649 & n1655;
  assign n1657 = ~n1643 & ~n1646;
  assign n1658 = ~n1649 & n1657;
  assign n1659 = ~n1656 & ~n1658;
  assign n1660 = n1654 & n1659;
  assign n1661 = ~n1638 & n1660;
  assign n1662 = n1638 & ~n1660;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = n1043 & ~n1054;
  assign n1665 = ~n1043 & n1054;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = n1024 & ~n1033;
  assign n1668 = ~n1024 & n1033;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = ~n1666 & n1669;
  assign n1671 = n1666 & ~n1669;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = 18 & 208;
  assign n1674 = ~n1388 & ~n1673;
  assign n1675 = n1113 & ~n1674;
  assign n1676 = ~n1113 & n1674;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n1091 & ~n1102;
  assign n1679 = ~n1091 & n1102;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n1072 & ~n1081;
  assign n1682 = ~n1072 & n1081;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1677 & n1680;
  assign n1685 = n1683 & n1684;
  assign n1686 = n1677 & n1680;
  assign n1687 = ~n1683 & n1686;
  assign n1688 = ~n1685 & ~n1687;
  assign n1689 = n1677 & ~n1680;
  assign n1690 = n1683 & n1689;
  assign n1691 = ~n1677 & ~n1680;
  assign n1692 = ~n1683 & n1691;
  assign n1693 = ~n1690 & ~n1692;
  assign n1694 = n1688 & n1693;
  assign n1695 = ~n1672 & n1694;
  assign n1696 = n1672 & ~n1694;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~n1595 & ~n1629;
  assign n1699 = ~n1663 & n1698;
  assign 10576 = n1697 | ~n1699;
  assign n1701 = n719 & ~n723;
  assign n1702 = n894 & ~n1018;
  assign n1703 = ~n1135 & n1702;
  assign n1704 = ~n1147 & n1703;
  assign n1705 = n901 & ~n1704;
  assign n1706 = n781 & ~n1705;
  assign n1707 = ~n1701 & ~n1706;
  assign n1708 = ~n719 & n1706;
  assign 10628 = n1707 | n1708;
  assign n1710 = n591 & ~n695;
  assign n1711 = ~n704 & n1710;
  assign n1712 = ~n594 & n1711;
  assign n1713 = n594 & ~n1711;
  assign 10632 = n1712 | n1713;
  assign n1715 = n494 & ~n600;
  assign n1716 = ~n696 & n1715;
  assign n1717 = ~n705 & n1716;
  assign n1718 = ~n497 & n1717;
  assign n1719 = n497 & ~n1717;
  assign 10641 = n1718 | n1719;
  assign n1721 = n945 & ~n951;
  assign n1722 = n1061 & ~n1067;
  assign n1723 = 89 & n1143;
  assign n1724 = n1123 & ~n1723;
  assign n1725 = ~n1722 & ~n1724;
  assign n1726 = ~n1061 & n1724;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = n1132 & ~n1727;
  assign n1729 = n1007 & ~n1728;
  assign n1730 = ~n1721 & ~n1729;
  assign n1731 = ~n945 & n1729;
  assign 10704 = n1730 | n1731;
  assign n1733 = n353 & ~n404;
  assign n1734 = n1157 & ~n1174;
  assign n1735 = ~n1187 & n1734;
  assign n1736 = ~n1196 & n1735;
  assign n1737 = n1161 & ~n1736;
  assign n1738 = n400 & ~n1737;
  assign n1739 = ~n1733 & ~n1738;
  assign n1740 = ~n353 & n1738;
  assign 10706 = n1739 | n1740;
  assign n1742 = ~n455 & n459;
  assign n1743 = ~n464 & n468;
  assign n1744 = ~n455 & n1743;
  assign n1745 = n478 & n479;
  assign n1746 = ~n455 & n1745;
  assign n1747 = ~n594 & ~n1711;
  assign n1748 = ~n464 & n1747;
  assign n1749 = ~n474 & n1748;
  assign n1750 = ~n455 & n1749;
  assign n1751 = ~n451 & ~n1742;
  assign n1752 = ~n1744 & n1751;
  assign n1753 = ~n1746 & n1752;
  assign n1754 = ~n1750 & n1753;
  assign n1755 = ~n447 & n1754;
  assign n1756 = n447 & ~n1754;
  assign 10711 = n1755 | n1756;
  assign n1758 = ~n459 & ~n1743;
  assign n1759 = ~n1745 & n1758;
  assign n1760 = ~n1749 & n1759;
  assign n1761 = ~n455 & n1760;
  assign n1762 = n455 & ~n1760;
  assign 10712 = n1761 | n1762;
  assign n1764 = ~n474 & n478;
  assign n1765 = ~n474 & n1747;
  assign n1766 = ~n468 & ~n1764;
  assign n1767 = ~n1765 & n1766;
  assign n1768 = ~n464 & n1767;
  assign n1769 = n464 & ~n1767;
  assign 10713 = n1768 | n1769;
  assign n1771 = ~n478 & ~n1747;
  assign n1772 = ~n474 & n1771;
  assign n1773 = n474 & ~n1771;
  assign 10714 = n1772 | n1773;
  assign n1775 = ~n369 & n373;
  assign n1776 = ~n378 & n382;
  assign n1777 = ~n369 & n1776;
  assign n1778 = n392 & n393;
  assign n1779 = ~n369 & n1778;
  assign n1780 = ~n497 & ~n1717;
  assign n1781 = ~n378 & n1780;
  assign n1782 = ~n388 & n1781;
  assign n1783 = ~n369 & n1782;
  assign n1784 = ~n365 & ~n1775;
  assign n1785 = ~n1777 & n1784;
  assign n1786 = ~n1779 & n1785;
  assign n1787 = ~n1783 & n1786;
  assign n1788 = ~n361 & n1787;
  assign n1789 = n361 & ~n1787;
  assign 10715 = n1788 | n1789;
  assign n1791 = ~n373 & ~n1776;
  assign n1792 = ~n1778 & n1791;
  assign n1793 = ~n1782 & n1792;
  assign n1794 = ~n369 & n1793;
  assign n1795 = n369 & ~n1793;
  assign 10716 = n1794 | n1795;
  assign n1797 = ~n388 & n392;
  assign n1798 = ~n388 & n1780;
  assign n1799 = ~n382 & ~n1797;
  assign n1800 = ~n1798 & n1799;
  assign n1801 = ~n378 & n1800;
  assign n1802 = n378 & ~n1800;
  assign 10717 = n1801 | n1802;
  assign n1804 = ~n392 & ~n1780;
  assign n1805 = ~n388 & n1804;
  assign n1806 = n388 & ~n1804;
  assign 10718 = n1805 | n1806;
  assign n1808 = ~882 & ~883;
  assign n1809 = ~884 & ~885;
  assign n1810 = ~10574 & ~10575;
  assign n1811 = ~10576 & n1810;
  assign n1812 = n1808 & n1809;
  assign 10729 = ~n1811 | ~n1812;
  assign n1814 = n501 & ~n1717;
  assign n1815 = n400 & ~n1814;
  assign n1816 = ~n353 & n1815;
  assign n1817 = ~n1733 & ~n1815;
  assign 10759 = n1816 | n1817;
  assign n1819 = ~n421 & n425;
  assign n1820 = ~n430 & n434;
  assign n1821 = ~n421 & n1820;
  assign n1822 = ~n417 & ~n1819;
  assign n1823 = ~n1821 & n1822;
  assign n1824 = ~n413 & ~n1823;
  assign n1825 = n413 & n1823;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = n598 & ~n1711;
  assign n1828 = n486 & ~n1827;
  assign n1829 = n1826 & n1828;
  assign n1830 = ~n1154 & n1823;
  assign n1831 = ~n413 & n1830;
  assign n1832 = n413 & ~n1830;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1828 & ~n1833;
  assign 10760 = n1829 | n1834;
  assign n1836 = ~n425 & ~n1820;
  assign n1837 = ~n421 & ~n1836;
  assign n1838 = n421 & n1836;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = n1828 & n1839;
  assign n1841 = ~n1153 & n1836;
  assign n1842 = ~n421 & n1841;
  assign n1843 = n421 & ~n1841;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1828 & ~n1844;
  assign 10761 = n1840 | n1845;
  assign n1847 = ~n430 & ~n434;
  assign n1848 = n430 & n434;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = n1828 & ~n1849;
  assign n1851 = 293 & ~n433;
  assign n1852 = ~n430 & ~n1851;
  assign n1853 = n430 & n1851;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1828 & n1854;
  assign 10762 = n1850 | n1855;
  assign n1857 = ~n489 & n1828;
  assign n1858 = n489 & ~n1828;
  assign 10763 = n1857 | n1858;
  assign n1860 = ~n635 & n1244;
  assign n1861 = n635 & ~n684;
  assign n1862 = ~n1244 & ~n1861;
  assign n1863 = ~n1860 & ~n1862;
  assign n1864 = ~n689 & n1863;
  assign n1865 = n689 & ~n1863;
  assign 10827 = n1864 | n1865;
  assign n1867 = ~n349 & ~n351;
  assign n1868 = n349 & n351;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = n1815 & ~n1869;
  assign n1871 = ~38 & n350;
  assign n1872 = ~n349 & ~n1871;
  assign n1873 = n349 & n1871;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1815 & n1874;
  assign 10837 = n1870 | n1875;
  assign n1877 = ~n403 & n1815;
  assign n1878 = n403 & ~n1815;
  assign 10839 = n1877 | n1878;
  assign n1880 = ~n552 & n556;
  assign n1881 = ~n561 & n565;
  assign n1882 = ~n552 & n1881;
  assign n1883 = n575 & n576;
  assign n1884 = ~n552 & n1883;
  assign n1885 = ~n689 & ~n1863;
  assign n1886 = ~n561 & n1885;
  assign n1887 = ~n571 & n1886;
  assign n1888 = ~n552 & n1887;
  assign n1889 = ~n548 & ~n1880;
  assign n1890 = ~n1882 & n1889;
  assign n1891 = ~n1884 & n1890;
  assign n1892 = ~n1888 & n1891;
  assign n1893 = ~n544 & n1892;
  assign n1894 = n544 & ~n1892;
  assign 10868 = n1893 | n1894;
  assign n1896 = ~n556 & ~n1881;
  assign n1897 = ~n1883 & n1896;
  assign n1898 = ~n1887 & n1897;
  assign n1899 = ~n552 & n1898;
  assign n1900 = n552 & ~n1898;
  assign 10869 = n1899 | n1900;
  assign n1902 = ~n571 & n575;
  assign n1903 = ~n571 & n1885;
  assign n1904 = ~n565 & ~n1902;
  assign n1905 = ~n1903 & n1904;
  assign n1906 = ~n561 & n1905;
  assign n1907 = n561 & ~n1905;
  assign 10870 = n1906 | n1907;
  assign n1909 = ~n575 & ~n1885;
  assign n1910 = ~n571 & n1909;
  assign n1911 = n571 & ~n1909;
  assign 10871 = n1910 | n1911;
  assign n1913 = ~n518 & n522;
  assign n1914 = ~n527 & n531;
  assign n1915 = ~n518 & n1914;
  assign n1916 = ~n514 & ~n1913;
  assign n1917 = ~n1915 & n1916;
  assign n1918 = ~n510 & ~n1917;
  assign n1919 = n510 & n1917;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = n693 & ~n1863;
  assign n1922 = n583 & ~n1921;
  assign n1923 = n1920 & n1922;
  assign n1924 = ~n1165 & n1917;
  assign n1925 = ~n510 & n1924;
  assign n1926 = n510 & ~n1924;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1922 & ~n1927;
  assign 10905 = n1923 | n1928;
  assign n1930 = ~n522 & ~n1914;
  assign n1931 = ~n518 & ~n1930;
  assign n1932 = n518 & n1930;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = n1922 & n1933;
  assign n1935 = ~n1164 & n1930;
  assign n1936 = ~n518 & n1935;
  assign n1937 = n518 & ~n1935;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1922 & ~n1938;
  assign 10906 = n1934 | n1939;
  assign n1941 = ~n527 & ~n531;
  assign n1942 = n527 & n531;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = n1922 & ~n1943;
  assign n1945 = 355 & n530;
  assign n1946 = ~n527 & ~n1945;
  assign n1947 = n527 & n1945;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~n1922 & n1948;
  assign 10907 = n1944 | n1949;
  assign n1951 = ~n586 & n1922;
  assign n1952 = n586 & ~n1922;
  assign 10908 = n1951 | n1952;
  assign n1954 = ~n478 & n1759;
  assign n1955 = n478 & ~n1759;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = n1766 & n1956;
  assign n1958 = ~n1766 & ~n1956;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960 = n1753 & n1959;
  assign n1961 = ~n1753 & ~n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n594 & n1962;
  assign n1964 = n594 & ~n1962;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n474 & n1965;
  assign n1967 = n474 & ~n1965;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n447 & n1968;
  assign n1970 = n447 & ~n1968;
  assign n1971 = ~n1969 & ~n1970;
  assign n1972 = ~n464 & n1971;
  assign n1973 = n464 & ~n1971;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = ~n455 & n1974;
  assign n1976 = n455 & ~n1974;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = n1168 & ~n1186;
  assign n1979 = ~n1195 & n1978;
  assign n1980 = n1977 & n1979;
  assign n1981 = ~n464 & ~n594;
  assign n1982 = ~n455 & n1981;
  assign n1983 = ~n474 & n1982;
  assign n1984 = n1753 & ~n1983;
  assign n1985 = ~n1169 & n1766;
  assign n1986 = ~n474 & n1981;
  assign n1987 = n1759 & ~n1986;
  assign n1988 = 277 & n477;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n1987 & n1988;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = ~n1985 & n1991;
  assign n1993 = n1985 & ~n1991;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~n1984 & n1994;
  assign n1996 = n1984 & ~n1994;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n594 & n1997;
  assign n1999 = n594 & ~n1997;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~n474 & n2000;
  assign n2002 = n474 & ~n2000;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = ~n447 & n2003;
  assign n2005 = n447 & ~n2003;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~n464 & n2006;
  assign n2008 = n464 & ~n2006;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n455 & n2009;
  assign n2011 = n455 & ~n2009;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n1979 & ~n2012;
  assign n2014 = ~n1980 & ~n2013;
  assign n2015 = ~n434 & n1836;
  assign n2016 = n434 & ~n1836;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n1823 & n2017;
  assign n2019 = ~n1823 & ~n2017;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n489 & n2020;
  assign n2022 = n489 & ~n2020;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = ~n430 & n2023;
  assign n2025 = n430 & ~n2023;
  assign n2026 = ~n2024 & ~n2025;
  assign n2027 = ~n413 & n2026;
  assign n2028 = n413 & ~n2026;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~n421 & n2029;
  assign n2031 = n421 & ~n2029;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = n486 & ~n2032;
  assign n2034 = n1979 & n2033;
  assign n2035 = ~n1841 & ~n1851;
  assign n2036 = n1841 & n1851;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = ~n1830 & n2037;
  assign n2039 = n1830 & ~n2037;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~n489 & n2040;
  assign n2042 = n489 & ~n2040;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = ~n430 & n2043;
  assign n2045 = n430 & ~n2043;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~n413 & n2046;
  assign n2048 = n413 & ~n2046;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = ~n421 & n2049;
  assign n2051 = n421 & ~n2049;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = ~n486 & ~n2052;
  assign n2054 = n1979 & n2053;
  assign n2055 = n486 & ~n1172;
  assign n2056 = ~n2032 & n2055;
  assign n2057 = ~n1979 & n2056;
  assign n2058 = ~n2052 & ~n2055;
  assign n2059 = ~n1979 & n2058;
  assign n2060 = ~n2034 & ~n2054;
  assign n2061 = ~n2057 & n2060;
  assign n2062 = ~n2059 & n2061;
  assign n2063 = ~n2014 & n2062;
  assign n2064 = n2014 & ~n2062;
  assign 11333 = ~n2063 & ~n2064;
  assign n2066 = ~n392 & n1792;
  assign n2067 = n392 & ~n1792;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = n1799 & n2068;
  assign n2070 = ~n1799 & ~n2068;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = n1786 & n2071;
  assign n2073 = ~n1786 & ~n2071;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = ~n497 & n2074;
  assign n2076 = n497 & ~n2074;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = ~n388 & n2077;
  assign n2079 = n388 & ~n2077;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n361 & n2080;
  assign n2082 = n361 & ~n2080;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n378 & n2083;
  assign n2085 = n378 & ~n2083;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = ~n369 & n2086;
  assign n2088 = n369 & ~n2086;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n1736 & n2089;
  assign n2091 = ~n378 & ~n497;
  assign n2092 = ~n369 & n2091;
  assign n2093 = ~n388 & n2092;
  assign n2094 = n1786 & ~n2093;
  assign n2095 = ~n1158 & n1799;
  assign n2096 = ~n388 & n2091;
  assign n2097 = n1792 & ~n2096;
  assign n2098 = 251 & ~n391;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = n2097 & n2098;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = ~n2095 & n2101;
  assign n2103 = n2095 & ~n2101;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n2094 & n2104;
  assign n2106 = n2094 & ~n2104;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = ~n497 & n2107;
  assign n2109 = n497 & ~n2107;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n388 & n2110;
  assign n2112 = n388 & ~n2110;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n361 & n2113;
  assign n2115 = n361 & ~n2113;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = ~n378 & n2116;
  assign n2118 = n378 & ~n2116;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~n369 & n2119;
  assign n2121 = n369 & ~n2119;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n1736 & ~n2122;
  assign n2124 = ~n2090 & ~n2123;
  assign n2125 = ~n351 & n353;
  assign n2126 = n351 & ~n353;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = n353 & n2127;
  assign n2129 = ~n353 & ~n2127;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n403 & n2130;
  assign n2132 = n403 & ~n2130;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = ~n349 & n2133;
  assign n2135 = n349 & ~n2133;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = n400 & ~n2136;
  assign n2138 = n1736 & n2137;
  assign n2139 = ~n1733 & ~n1871;
  assign n2140 = n1733 & n1871;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~n1733 & n2141;
  assign n2143 = n1733 & ~n2141;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~n403 & n2144;
  assign n2146 = n403 & ~n2144;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n349 & n2147;
  assign n2149 = n349 & ~n2147;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = ~n400 & ~n2150;
  assign n2152 = n1736 & n2151;
  assign n2153 = n400 & ~n1161;
  assign n2154 = ~n2136 & n2153;
  assign n2155 = ~n1736 & n2154;
  assign n2156 = ~n2150 & ~n2153;
  assign n2157 = ~n1736 & n2156;
  assign n2158 = ~n2138 & ~n2152;
  assign n2159 = ~n2155 & n2158;
  assign n2160 = ~n2157 & n2159;
  assign n2161 = ~n2124 & n2160;
  assign n2162 = n2124 & ~n2160;
  assign 11334 = ~n2161 & ~n2162;
  assign n2164 = ~n575 & n1897;
  assign n2165 = n575 & ~n1897;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = n1904 & n2166;
  assign n2168 = ~n1904 & ~n2166;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = n1891 & n2169;
  assign n2171 = ~n1891 & ~n2169;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n689 & n2172;
  assign n2174 = n689 & ~n2172;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = ~n571 & n2175;
  assign n2177 = n571 & ~n2175;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = ~n544 & n2178;
  assign n2180 = n544 & ~n2178;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n561 & n2181;
  assign n2183 = n561 & ~n2181;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~n552 & n2184;
  assign n2186 = n552 & ~n2184;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = n635 & ~n1178;
  assign n2189 = 367 & n1192;
  assign n2190 = n678 & ~n2189;
  assign n2191 = ~n2188 & ~n2190;
  assign n2192 = ~n635 & n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = n2187 & n2193;
  assign n2195 = ~n561 & ~n689;
  assign n2196 = ~n552 & n2195;
  assign n2197 = ~n571 & n2196;
  assign n2198 = n1891 & ~n2197;
  assign n2199 = ~n1181 & n1904;
  assign n2200 = ~n571 & n2195;
  assign n2201 = n1897 & ~n2200;
  assign n2202 = 340 & n574;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = n2201 & n2202;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = ~n2199 & n2205;
  assign n2207 = n2199 & ~n2205;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~n2198 & n2208;
  assign n2210 = n2198 & ~n2208;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n689 & n2211;
  assign n2213 = n689 & ~n2211;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n571 & n2214;
  assign n2216 = n571 & ~n2214;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n544 & n2217;
  assign n2219 = n544 & ~n2217;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~n561 & n2220;
  assign n2222 = n561 & ~n2220;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = ~n552 & n2223;
  assign n2225 = n552 & ~n2223;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = ~n2193 & ~n2226;
  assign n2228 = ~n2194 & ~n2227;
  assign n2229 = ~n531 & n1930;
  assign n2230 = n531 & ~n1930;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = n1917 & n2231;
  assign n2233 = ~n1917 & ~n2231;
  assign n2234 = ~n2232 & ~n2233;
  assign n2235 = ~n586 & n2234;
  assign n2236 = n586 & ~n2234;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n527 & n2237;
  assign n2239 = n527 & ~n2237;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n510 & n2240;
  assign n2242 = n510 & ~n2240;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = ~n518 & n2243;
  assign n2245 = n518 & ~n2243;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n583 & ~n2246;
  assign n2248 = n2193 & n2247;
  assign n2249 = ~n1935 & ~n1945;
  assign n2250 = n1935 & n1945;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = ~n1924 & n2251;
  assign n2253 = n1924 & ~n2251;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = ~n586 & n2254;
  assign n2256 = n586 & ~n2254;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = ~n527 & n2257;
  assign n2259 = n527 & ~n2257;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = ~n510 & n2260;
  assign n2262 = n510 & ~n2260;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~n518 & n2263;
  assign n2265 = n518 & ~n2263;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n583 & ~n2266;
  assign n2268 = n2193 & n2267;
  assign n2269 = n583 & ~n1184;
  assign n2270 = ~n2246 & n2269;
  assign n2271 = ~n2193 & n2270;
  assign n2272 = ~n2266 & ~n2269;
  assign n2273 = ~n2193 & n2272;
  assign n2274 = ~n2248 & ~n2268;
  assign n2275 = ~n2271 & n2274;
  assign n2276 = ~n2273 & n2275;
  assign n2277 = ~n2228 & n2276;
  assign n2278 = n2228 & ~n2276;
  assign 11340 = ~n2277 & ~n2278;
  assign n2280 = ~n670 & n1219;
  assign n2281 = n670 & ~n1219;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = n1226 & n2282;
  assign n2284 = ~n1226 & ~n2282;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = n1213 & n2285;
  assign n2287 = ~n1213 & ~n2285;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n341 & n2288;
  assign n2290 = n341 & ~n2288;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n669 & n2291;
  assign n2293 = n669 & ~n2291;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n642 & n2294;
  assign n2296 = n642 & ~n2294;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = ~n659 & n2297;
  assign n2299 = n659 & ~n2297;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = ~n650 & n2300;
  assign n2302 = n650 & ~n2300;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~367 & n2303;
  assign n2305 = ~n341 & ~n659;
  assign n2306 = ~n650 & n2305;
  assign n2307 = ~n669 & n2306;
  assign n2308 = n1213 & ~n2307;
  assign n2309 = ~n1189 & n1226;
  assign n2310 = ~n669 & n2305;
  assign n2311 = n1219 & ~n2310;
  assign n2312 = ~n336 & n338;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = n2311 & n2312;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n2309 & n2315;
  assign n2317 = n2309 & ~n2315;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = ~n2308 & n2318;
  assign n2320 = n2308 & ~n2318;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = ~n341 & n2321;
  assign n2323 = n341 & ~n2321;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n669 & n2324;
  assign n2326 = n669 & ~n2324;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = ~n642 & n2327;
  assign n2329 = n642 & ~n2327;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = ~n659 & n2330;
  assign n2332 = n659 & ~n2330;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = ~n650 & n2333;
  assign n2335 = n650 & ~n2333;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = 367 & ~n2336;
  assign n2338 = ~n2304 & ~n2337;
  assign n2339 = ~n629 & n1252;
  assign n2340 = n629 & ~n1252;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = n1239 & n2341;
  assign n2343 = ~n1239 & ~n2341;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~n681 & n2344;
  assign n2346 = n681 & ~n2344;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n625 & n2347;
  assign n2349 = n625 & ~n2347;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~n608 & n2350;
  assign n2352 = n608 & ~n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n616 & n2353;
  assign n2355 = n616 & ~n2353;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = n678 & ~n2356;
  assign n2358 = ~367 & n2357;
  assign n2359 = ~n1257 & ~n1267;
  assign n2360 = n1257 & n1267;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n1246 & n2361;
  assign n2363 = n1246 & ~n2361;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = ~n681 & n2364;
  assign n2366 = n681 & ~n2364;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n625 & n2367;
  assign n2369 = n625 & ~n2367;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = ~n608 & n2370;
  assign n2372 = n608 & ~n2370;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~n616 & n2373;
  assign n2375 = n616 & ~n2373;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n678 & ~n2376;
  assign n2378 = ~367 & n2377;
  assign n2379 = n678 & ~n1192;
  assign n2380 = ~n2356 & n2379;
  assign n2381 = 367 & n2380;
  assign n2382 = ~n2376 & ~n2379;
  assign n2383 = 367 & n2382;
  assign n2384 = ~n2358 & ~n2378;
  assign n2385 = ~n2381 & n2384;
  assign n2386 = ~n2383 & n2385;
  assign n2387 = ~n2338 & n2386;
  assign n2388 = n2338 & ~n2386;
  assign 11342 = ~n2387 & ~n2388;
  assign 582 = ~15;
  assign 387 = \1 ;
  assign 388 = \1 ;
  assign 478 = 248;
  assign 482 = 254;
  assign 484 = 257;
  assign 486 = 260;
  assign 489 = 263;
  assign 492 = 267;
  assign 501 = 274;
  assign 505 = 280;
  assign 507 = 283;
  assign 509 = 286;
  assign 511 = 289;
  assign 513 = 293;
  assign 515 = 296;
  assign 517 = 299;
  assign 519 = 303;
  assign 535 = 307;
  assign 537 = 310;
  assign 539 = 313;
  assign 541 = 316;
  assign 543 = 319;
  assign 545 = 322;
  assign 547 = 325;
  assign 549 = 328;
  assign 551 = 331;
  assign 553 = 334;
  assign 556 = 337;
  assign 559 = 343;
  assign 561 = 346;
  assign 563 = 349;
  assign 565 = 352;
  assign 567 = 355;
  assign 569 = 358;
  assign 571 = 361;
  assign 573 = 364;
  assign 643 = 251;
  assign 707 = 277;
  assign 813 = 340;
  assign 889 = \1 ;
  assign 945 = 106;
  assign 1111 = 582;
  assign 1112 = 1110;
  assign 1114 = 582;
  assign 1489 = 1113;
  assign 1490 = \1 ;
  assign 10103 = 10102;
  assign 10838 = 10837;
  assign 10840 = 10839;
endmodule


