// Benchmark "top" written by ABC on Mon Feb 19 11:52:42 2024

module top ( 
    p_127gat_18_, p_155gat_22_, p_120gat_17_, p_64gat_9_, p_106gat_15_,
    p_204gat_29_, p_1gat_0_, p_43gat_6_, p_85gat_12_, p_141gat_20_,
    p_183gat_26_, p_57gat_8_, p_148gat_21_, p_169gat_24_, p_225gat_32_,
    p_99gat_14_, p_230gat_37_, p_134gat_19_, p_162gat_23_, p_29gat_4_,
    p_78gat_11_, p_226gat_33_, p_22gat_3_, p_231gat_38_, p_36gat_5_,
    p_113gat_16_, p_8gat_1_, p_50gat_7_, p_227gat_34_, p_92gat_13_,
    p_197gat_28_, p_232gat_39_, p_233gat_40_, p_71gat_10_, p_190gat_27_,
    p_15gat_2_, p_228gat_35_, p_176gat_25_, p_218gat_31_, p_211gat_30_,
    p_229gat_36_,
    p_1332gat_585_, p_1331gat_572_, p_1334gat_577_, p_1354gat_562_,
    p_1352gat_570_, p_1336gat_586_, p_1330gat_576_, p_1335gat_573_,
    p_1353gat_566_, p_1329gat_580_, p_1328gat_584_, p_1342gat_559_,
    p_1351gat_557_, p_1333gat_581_, p_1349gat_565_, p_1350gat_561_,
    p_1348gat_569_, p_1347gat_556_, p_1341gat_563_, p_1325gat_579_,
    p_1326gat_575_, p_1344gat_568_, p_1324gat_583_, p_1343gat_555_,
    p_1345gat_564_, p_1337gat_582_, p_1327gat_571_, p_1340gat_567_,
    p_1346gat_560_, p_1339gat_574_, p_1355gat_558_, p_1338gat_578_  );
  input  p_127gat_18_, p_155gat_22_, p_120gat_17_, p_64gat_9_,
    p_106gat_15_, p_204gat_29_, p_1gat_0_, p_43gat_6_, p_85gat_12_,
    p_141gat_20_, p_183gat_26_, p_57gat_8_, p_148gat_21_, p_169gat_24_,
    p_225gat_32_, p_99gat_14_, p_230gat_37_, p_134gat_19_, p_162gat_23_,
    p_29gat_4_, p_78gat_11_, p_226gat_33_, p_22gat_3_, p_231gat_38_,
    p_36gat_5_, p_113gat_16_, p_8gat_1_, p_50gat_7_, p_227gat_34_,
    p_92gat_13_, p_197gat_28_, p_232gat_39_, p_233gat_40_, p_71gat_10_,
    p_190gat_27_, p_15gat_2_, p_228gat_35_, p_176gat_25_, p_218gat_31_,
    p_211gat_30_, p_229gat_36_;
  output p_1332gat_585_, p_1331gat_572_, p_1334gat_577_, p_1354gat_562_,
    p_1352gat_570_, p_1336gat_586_, p_1330gat_576_, p_1335gat_573_,
    p_1353gat_566_, p_1329gat_580_, p_1328gat_584_, p_1342gat_559_,
    p_1351gat_557_, p_1333gat_581_, p_1349gat_565_, p_1350gat_561_,
    p_1348gat_569_, p_1347gat_556_, p_1341gat_563_, p_1325gat_579_,
    p_1326gat_575_, p_1344gat_568_, p_1324gat_583_, p_1343gat_555_,
    p_1345gat_564_, p_1337gat_582_, p_1327gat_571_, p_1340gat_567_,
    p_1346gat_560_, p_1339gat_574_, p_1355gat_558_, p_1338gat_578_;
  wire new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n393, new_n394, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n402, new_n403, new_n404, new_n405, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n430, new_n431, new_n432, new_n433, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n443, new_n444, new_n445,
    new_n446, new_n448, new_n449, new_n450, new_n451, new_n453, new_n454,
    new_n455, new_n456, new_n458, new_n459, new_n460, new_n461, new_n463,
    new_n464, new_n465, new_n466, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n500, new_n501, new_n502, new_n503, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n513,
    new_n514, new_n515, new_n516, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n526, new_n527, new_n528, new_n529,
    new_n531, new_n532, new_n533, new_n534, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584;
  assign new_n74 = p_106gat_15_ & p_99gat_14_;
  assign new_n75 = p_106gat_15_ & ~new_n74;
  assign new_n76 = p_99gat_14_ & ~new_n74;
  assign new_n77 = ~new_n75 & ~new_n76;
  assign new_n78 = p_85gat_12_ & p_92gat_13_;
  assign new_n79 = p_92gat_13_ & ~new_n78;
  assign new_n80 = p_85gat_12_ & ~new_n78;
  assign new_n81 = ~new_n79 & ~new_n80;
  assign new_n82 = ~new_n77 & ~new_n81;
  assign new_n83 = ~new_n77 & ~new_n82;
  assign new_n84 = ~new_n81 & ~new_n82;
  assign new_n85 = ~new_n83 & ~new_n84;
  assign new_n86 = p_43gat_6_ & p_50gat_7_;
  assign new_n87 = p_50gat_7_ & ~new_n86;
  assign new_n88 = p_43gat_6_ & ~new_n86;
  assign new_n89 = ~new_n87 & ~new_n88;
  assign new_n90 = p_29gat_4_ & p_36gat_5_;
  assign new_n91 = p_36gat_5_ & ~new_n90;
  assign new_n92 = p_29gat_4_ & ~new_n90;
  assign new_n93 = ~new_n91 & ~new_n92;
  assign new_n94 = ~new_n89 & ~new_n93;
  assign new_n95 = ~new_n89 & ~new_n94;
  assign new_n96 = ~new_n93 & ~new_n94;
  assign new_n97 = ~new_n95 & ~new_n96;
  assign new_n98 = ~new_n85 & ~new_n97;
  assign new_n99 = ~new_n85 & ~new_n98;
  assign new_n100 = ~new_n97 & ~new_n98;
  assign new_n101 = ~new_n99 & ~new_n100;
  assign new_n102 = p_232gat_39_ & p_233gat_40_;
  assign new_n103 = ~new_n101 & new_n102;
  assign new_n104 = ~new_n101 & ~new_n103;
  assign new_n105 = new_n102 & ~new_n103;
  assign new_n106 = ~new_n104 & ~new_n105;
  assign new_n107 = p_190gat_27_ & p_218gat_31_;
  assign new_n108 = p_218gat_31_ & ~new_n107;
  assign new_n109 = p_190gat_27_ & ~new_n107;
  assign new_n110 = ~new_n108 & ~new_n109;
  assign new_n111 = p_134gat_19_ & p_162gat_23_;
  assign new_n112 = p_162gat_23_ & ~new_n111;
  assign new_n113 = p_134gat_19_ & ~new_n111;
  assign new_n114 = ~new_n112 & ~new_n113;
  assign new_n115 = ~new_n110 & ~new_n114;
  assign new_n116 = ~new_n110 & ~new_n115;
  assign new_n117 = ~new_n114 & ~new_n115;
  assign new_n118 = ~new_n116 & ~new_n117;
  assign new_n119 = ~new_n106 & ~new_n118;
  assign new_n120 = ~new_n106 & ~new_n119;
  assign new_n121 = ~new_n118 & ~new_n119;
  assign new_n122 = ~new_n120 & ~new_n121;
  assign new_n123 = p_218gat_31_ & p_211gat_30_;
  assign new_n124 = p_218gat_31_ & ~new_n123;
  assign new_n125 = p_211gat_30_ & ~new_n123;
  assign new_n126 = ~new_n124 & ~new_n125;
  assign new_n127 = p_204gat_29_ & p_197gat_28_;
  assign new_n128 = p_204gat_29_ & ~new_n127;
  assign new_n129 = p_197gat_28_ & ~new_n127;
  assign new_n130 = ~new_n128 & ~new_n129;
  assign new_n131 = ~new_n126 & ~new_n130;
  assign new_n132 = ~new_n126 & ~new_n131;
  assign new_n133 = ~new_n130 & ~new_n131;
  assign new_n134 = ~new_n132 & ~new_n133;
  assign new_n135 = p_155gat_22_ & p_162gat_23_;
  assign new_n136 = p_162gat_23_ & ~new_n135;
  assign new_n137 = p_155gat_22_ & ~new_n135;
  assign new_n138 = ~new_n136 & ~new_n137;
  assign new_n139 = p_141gat_20_ & p_148gat_21_;
  assign new_n140 = p_148gat_21_ & ~new_n139;
  assign new_n141 = p_141gat_20_ & ~new_n139;
  assign new_n142 = ~new_n140 & ~new_n141;
  assign new_n143 = ~new_n138 & ~new_n142;
  assign new_n144 = ~new_n138 & ~new_n143;
  assign new_n145 = ~new_n142 & ~new_n143;
  assign new_n146 = ~new_n144 & ~new_n145;
  assign new_n147 = ~new_n134 & ~new_n146;
  assign new_n148 = ~new_n134 & ~new_n147;
  assign new_n149 = ~new_n146 & ~new_n147;
  assign new_n150 = ~new_n148 & ~new_n149;
  assign new_n151 = p_233gat_40_ & p_228gat_35_;
  assign new_n152 = ~new_n150 & new_n151;
  assign new_n153 = ~new_n150 & ~new_n152;
  assign new_n154 = new_n151 & ~new_n152;
  assign new_n155 = ~new_n153 & ~new_n154;
  assign new_n156 = p_106gat_15_ & p_78gat_11_;
  assign new_n157 = p_106gat_15_ & ~new_n156;
  assign new_n158 = p_78gat_11_ & ~new_n156;
  assign new_n159 = ~new_n157 & ~new_n158;
  assign new_n160 = p_22gat_3_ & p_50gat_7_;
  assign new_n161 = p_50gat_7_ & ~new_n160;
  assign new_n162 = p_22gat_3_ & ~new_n160;
  assign new_n163 = ~new_n161 & ~new_n162;
  assign new_n164 = ~new_n159 & ~new_n163;
  assign new_n165 = ~new_n159 & ~new_n164;
  assign new_n166 = ~new_n163 & ~new_n164;
  assign new_n167 = ~new_n165 & ~new_n166;
  assign new_n168 = ~new_n155 & ~new_n167;
  assign new_n169 = ~new_n155 & ~new_n168;
  assign new_n170 = ~new_n167 & ~new_n168;
  assign new_n171 = ~new_n169 & ~new_n170;
  assign new_n172 = p_183gat_26_ & p_190gat_27_;
  assign new_n173 = p_190gat_27_ & ~new_n172;
  assign new_n174 = p_183gat_26_ & ~new_n172;
  assign new_n175 = ~new_n173 & ~new_n174;
  assign new_n176 = p_169gat_24_ & p_176gat_25_;
  assign new_n177 = p_176gat_25_ & ~new_n176;
  assign new_n178 = p_169gat_24_ & ~new_n176;
  assign new_n179 = ~new_n177 & ~new_n178;
  assign new_n180 = ~new_n175 & ~new_n179;
  assign new_n181 = ~new_n175 & ~new_n180;
  assign new_n182 = ~new_n179 & ~new_n180;
  assign new_n183 = ~new_n181 & ~new_n182;
  assign new_n184 = ~new_n134 & ~new_n183;
  assign new_n185 = ~new_n134 & ~new_n184;
  assign new_n186 = ~new_n183 & ~new_n184;
  assign new_n187 = ~new_n185 & ~new_n186;
  assign new_n188 = p_226gat_33_ & p_233gat_40_;
  assign new_n189 = ~new_n187 & new_n188;
  assign new_n190 = ~new_n187 & ~new_n189;
  assign new_n191 = new_n188 & ~new_n189;
  assign new_n192 = ~new_n190 & ~new_n191;
  assign new_n193 = p_64gat_9_ & p_92gat_13_;
  assign new_n194 = p_92gat_13_ & ~new_n193;
  assign new_n195 = p_64gat_9_ & ~new_n193;
  assign new_n196 = ~new_n194 & ~new_n195;
  assign new_n197 = p_36gat_5_ & p_8gat_1_;
  assign new_n198 = p_36gat_5_ & ~new_n197;
  assign new_n199 = p_8gat_1_ & ~new_n197;
  assign new_n200 = ~new_n198 & ~new_n199;
  assign new_n201 = ~new_n196 & ~new_n200;
  assign new_n202 = ~new_n196 & ~new_n201;
  assign new_n203 = ~new_n200 & ~new_n201;
  assign new_n204 = ~new_n202 & ~new_n203;
  assign new_n205 = ~new_n192 & ~new_n204;
  assign new_n206 = ~new_n192 & ~new_n205;
  assign new_n207 = ~new_n204 & ~new_n205;
  assign new_n208 = ~new_n206 & ~new_n207;
  assign new_n209 = p_127gat_18_ & p_134gat_19_;
  assign new_n210 = p_134gat_19_ & ~new_n209;
  assign new_n211 = p_127gat_18_ & ~new_n209;
  assign new_n212 = ~new_n210 & ~new_n211;
  assign new_n213 = p_120gat_17_ & p_113gat_16_;
  assign new_n214 = p_120gat_17_ & ~new_n213;
  assign new_n215 = p_113gat_16_ & ~new_n213;
  assign new_n216 = ~new_n214 & ~new_n215;
  assign new_n217 = ~new_n212 & ~new_n216;
  assign new_n218 = ~new_n212 & ~new_n217;
  assign new_n219 = ~new_n216 & ~new_n217;
  assign new_n220 = ~new_n218 & ~new_n219;
  assign new_n221 = ~new_n183 & ~new_n220;
  assign new_n222 = ~new_n183 & ~new_n221;
  assign new_n223 = ~new_n220 & ~new_n221;
  assign new_n224 = ~new_n222 & ~new_n223;
  assign new_n225 = p_227gat_34_ & p_233gat_40_;
  assign new_n226 = ~new_n224 & new_n225;
  assign new_n227 = ~new_n224 & ~new_n226;
  assign new_n228 = new_n225 & ~new_n226;
  assign new_n229 = ~new_n227 & ~new_n228;
  assign new_n230 = p_99gat_14_ & p_71gat_10_;
  assign new_n231 = p_99gat_14_ & ~new_n230;
  assign new_n232 = p_71gat_10_ & ~new_n230;
  assign new_n233 = ~new_n231 & ~new_n232;
  assign new_n234 = p_43gat_6_ & p_15gat_2_;
  assign new_n235 = p_43gat_6_ & ~new_n234;
  assign new_n236 = p_15gat_2_ & ~new_n234;
  assign new_n237 = ~new_n235 & ~new_n236;
  assign new_n238 = ~new_n233 & ~new_n237;
  assign new_n239 = ~new_n233 & ~new_n238;
  assign new_n240 = ~new_n237 & ~new_n238;
  assign new_n241 = ~new_n239 & ~new_n240;
  assign new_n242 = ~new_n229 & ~new_n241;
  assign new_n243 = ~new_n229 & ~new_n242;
  assign new_n244 = ~new_n241 & ~new_n242;
  assign new_n245 = ~new_n243 & ~new_n244;
  assign new_n246 = ~new_n146 & ~new_n220;
  assign new_n247 = ~new_n146 & ~new_n246;
  assign new_n248 = ~new_n220 & ~new_n246;
  assign new_n249 = ~new_n247 & ~new_n248;
  assign new_n250 = p_225gat_32_ & p_233gat_40_;
  assign new_n251 = ~new_n249 & new_n250;
  assign new_n252 = ~new_n249 & ~new_n251;
  assign new_n253 = new_n250 & ~new_n251;
  assign new_n254 = ~new_n252 & ~new_n253;
  assign new_n255 = p_85gat_12_ & p_57gat_8_;
  assign new_n256 = p_85gat_12_ & ~new_n255;
  assign new_n257 = p_57gat_8_ & ~new_n255;
  assign new_n258 = ~new_n256 & ~new_n257;
  assign new_n259 = p_1gat_0_ & p_29gat_4_;
  assign new_n260 = p_29gat_4_ & ~new_n259;
  assign new_n261 = p_1gat_0_ & ~new_n259;
  assign new_n262 = ~new_n260 & ~new_n261;
  assign new_n263 = ~new_n258 & ~new_n262;
  assign new_n264 = ~new_n258 & ~new_n263;
  assign new_n265 = ~new_n262 & ~new_n263;
  assign new_n266 = ~new_n264 & ~new_n265;
  assign new_n267 = ~new_n254 & ~new_n266;
  assign new_n268 = ~new_n254 & ~new_n267;
  assign new_n269 = ~new_n266 & ~new_n267;
  assign new_n270 = ~new_n268 & ~new_n269;
  assign new_n271 = new_n171 & new_n208;
  assign new_n272 = new_n245 & new_n271;
  assign new_n273 = ~new_n270 & new_n272;
  assign new_n274 = ~new_n245 & new_n271;
  assign new_n275 = new_n270 & new_n274;
  assign new_n276 = new_n171 & ~new_n208;
  assign new_n277 = new_n245 & new_n276;
  assign new_n278 = new_n270 & new_n277;
  assign new_n279 = ~new_n171 & new_n208;
  assign new_n280 = new_n245 & new_n279;
  assign new_n281 = new_n270 & new_n280;
  assign new_n282 = ~new_n273 & ~new_n275;
  assign new_n283 = ~new_n278 & new_n282;
  assign new_n284 = ~new_n281 & new_n283;
  assign new_n285 = p_78gat_11_ & p_71gat_10_;
  assign new_n286 = p_78gat_11_ & ~new_n285;
  assign new_n287 = p_71gat_10_ & ~new_n285;
  assign new_n288 = ~new_n286 & ~new_n287;
  assign new_n289 = p_64gat_9_ & p_57gat_8_;
  assign new_n290 = p_64gat_9_ & ~new_n289;
  assign new_n291 = p_57gat_8_ & ~new_n289;
  assign new_n292 = ~new_n290 & ~new_n291;
  assign new_n293 = ~new_n288 & ~new_n292;
  assign new_n294 = ~new_n288 & ~new_n293;
  assign new_n295 = ~new_n292 & ~new_n293;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = ~new_n85 & ~new_n296;
  assign new_n298 = ~new_n85 & ~new_n297;
  assign new_n299 = ~new_n296 & ~new_n297;
  assign new_n300 = ~new_n298 & ~new_n299;
  assign new_n301 = p_230gat_37_ & p_233gat_40_;
  assign new_n302 = ~new_n300 & new_n301;
  assign new_n303 = ~new_n300 & ~new_n302;
  assign new_n304 = new_n301 & ~new_n302;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = p_204gat_29_ & p_176gat_25_;
  assign new_n307 = p_204gat_29_ & ~new_n306;
  assign new_n308 = p_176gat_25_ & ~new_n306;
  assign new_n309 = ~new_n307 & ~new_n308;
  assign new_n310 = p_120gat_17_ & p_148gat_21_;
  assign new_n311 = p_148gat_21_ & ~new_n310;
  assign new_n312 = p_120gat_17_ & ~new_n310;
  assign new_n313 = ~new_n311 & ~new_n312;
  assign new_n314 = ~new_n309 & ~new_n313;
  assign new_n315 = ~new_n309 & ~new_n314;
  assign new_n316 = ~new_n313 & ~new_n314;
  assign new_n317 = ~new_n315 & ~new_n316;
  assign new_n318 = ~new_n305 & ~new_n317;
  assign new_n319 = ~new_n305 & ~new_n318;
  assign new_n320 = ~new_n317 & ~new_n318;
  assign new_n321 = ~new_n319 & ~new_n320;
  assign new_n322 = p_22gat_3_ & p_15gat_2_;
  assign new_n323 = p_22gat_3_ & ~new_n322;
  assign new_n324 = p_15gat_2_ & ~new_n322;
  assign new_n325 = ~new_n323 & ~new_n324;
  assign new_n326 = p_1gat_0_ & p_8gat_1_;
  assign new_n327 = p_8gat_1_ & ~new_n326;
  assign new_n328 = p_1gat_0_ & ~new_n326;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = ~new_n325 & ~new_n329;
  assign new_n331 = ~new_n325 & ~new_n330;
  assign new_n332 = ~new_n329 & ~new_n330;
  assign new_n333 = ~new_n331 & ~new_n332;
  assign new_n334 = ~new_n296 & ~new_n333;
  assign new_n335 = ~new_n296 & ~new_n334;
  assign new_n336 = ~new_n333 & ~new_n334;
  assign new_n337 = ~new_n335 & ~new_n336;
  assign new_n338 = p_231gat_38_ & p_233gat_40_;
  assign new_n339 = ~new_n337 & new_n338;
  assign new_n340 = ~new_n337 & ~new_n339;
  assign new_n341 = new_n338 & ~new_n339;
  assign new_n342 = ~new_n340 & ~new_n341;
  assign new_n343 = p_183gat_26_ & p_211gat_30_;
  assign new_n344 = p_211gat_30_ & ~new_n343;
  assign new_n345 = p_183gat_26_ & ~new_n343;
  assign new_n346 = ~new_n344 & ~new_n345;
  assign new_n347 = p_127gat_18_ & p_155gat_22_;
  assign new_n348 = p_155gat_22_ & ~new_n347;
  assign new_n349 = p_127gat_18_ & ~new_n347;
  assign new_n350 = ~new_n348 & ~new_n349;
  assign new_n351 = ~new_n346 & ~new_n350;
  assign new_n352 = ~new_n346 & ~new_n351;
  assign new_n353 = ~new_n350 & ~new_n351;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = ~new_n342 & ~new_n354;
  assign new_n356 = ~new_n342 & ~new_n355;
  assign new_n357 = ~new_n354 & ~new_n355;
  assign new_n358 = ~new_n356 & ~new_n357;
  assign new_n359 = ~new_n97 & ~new_n333;
  assign new_n360 = ~new_n97 & ~new_n359;
  assign new_n361 = ~new_n333 & ~new_n359;
  assign new_n362 = ~new_n360 & ~new_n361;
  assign new_n363 = p_233gat_40_ & p_229gat_36_;
  assign new_n364 = ~new_n362 & new_n363;
  assign new_n365 = ~new_n362 & ~new_n364;
  assign new_n366 = new_n363 & ~new_n364;
  assign new_n367 = ~new_n365 & ~new_n366;
  assign new_n368 = p_169gat_24_ & p_197gat_28_;
  assign new_n369 = p_197gat_28_ & ~new_n368;
  assign new_n370 = p_169gat_24_ & ~new_n368;
  assign new_n371 = ~new_n369 & ~new_n370;
  assign new_n372 = p_141gat_20_ & p_113gat_16_;
  assign new_n373 = p_141gat_20_ & ~new_n372;
  assign new_n374 = p_113gat_16_ & ~new_n372;
  assign new_n375 = ~new_n373 & ~new_n374;
  assign new_n376 = ~new_n371 & ~new_n375;
  assign new_n377 = ~new_n371 & ~new_n376;
  assign new_n378 = ~new_n375 & ~new_n376;
  assign new_n379 = ~new_n377 & ~new_n378;
  assign new_n380 = ~new_n367 & ~new_n379;
  assign new_n381 = ~new_n367 & ~new_n380;
  assign new_n382 = ~new_n379 & ~new_n380;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = new_n122 & ~new_n284;
  assign new_n385 = ~new_n321 & new_n384;
  assign new_n386 = ~new_n358 & new_n385;
  assign new_n387 = new_n383 & new_n386;
  assign new_n388 = ~new_n270 & new_n387;
  assign new_n389 = p_57gat_8_ & new_n388;
  assign new_n390 = new_n388 & ~new_n389;
  assign new_n391 = p_57gat_8_ & ~new_n389;
  assign p_1332gat_585_ = new_n390 | new_n391;
  assign new_n393 = ~new_n122 & ~new_n284;
  assign new_n394 = new_n321 & new_n393;
  assign new_n395 = new_n358 & new_n394;
  assign new_n396 = ~new_n383 & new_n395;
  assign new_n397 = ~new_n171 & new_n396;
  assign new_n398 = p_50gat_7_ & new_n397;
  assign new_n399 = new_n397 & ~new_n398;
  assign new_n400 = p_50gat_7_ & ~new_n398;
  assign p_1331gat_572_ = new_n399 | new_n400;
  assign new_n402 = ~new_n245 & new_n387;
  assign new_n403 = p_71gat_10_ & new_n402;
  assign new_n404 = new_n402 & ~new_n403;
  assign new_n405 = p_71gat_10_ & ~new_n403;
  assign p_1334gat_577_ = new_n404 | new_n405;
  assign new_n407 = new_n122 & new_n321;
  assign new_n408 = new_n358 & new_n407;
  assign new_n409 = ~new_n383 & new_n408;
  assign new_n410 = ~new_n358 & new_n407;
  assign new_n411 = new_n383 & new_n410;
  assign new_n412 = new_n122 & ~new_n321;
  assign new_n413 = new_n358 & new_n412;
  assign new_n414 = new_n383 & new_n413;
  assign new_n415 = ~new_n122 & new_n321;
  assign new_n416 = new_n358 & new_n415;
  assign new_n417 = new_n383 & new_n416;
  assign new_n418 = ~new_n409 & ~new_n411;
  assign new_n419 = ~new_n414 & new_n418;
  assign new_n420 = ~new_n417 & new_n419;
  assign new_n421 = ~new_n171 & ~new_n420;
  assign new_n422 = ~new_n208 & new_n421;
  assign new_n423 = new_n245 & new_n422;
  assign new_n424 = new_n270 & new_n423;
  assign new_n425 = ~new_n358 & new_n424;
  assign new_n426 = p_211gat_30_ & new_n425;
  assign new_n427 = new_n425 & ~new_n426;
  assign new_n428 = p_211gat_30_ & ~new_n426;
  assign p_1354gat_562_ = new_n427 | new_n428;
  assign new_n430 = ~new_n383 & new_n424;
  assign new_n431 = p_197gat_28_ & new_n430;
  assign new_n432 = new_n430 & ~new_n431;
  assign new_n433 = p_197gat_28_ & ~new_n431;
  assign p_1352gat_570_ = new_n432 | new_n433;
  assign new_n435 = ~new_n321 & new_n393;
  assign new_n436 = new_n358 & new_n435;
  assign new_n437 = new_n383 & new_n436;
  assign new_n438 = ~new_n270 & new_n437;
  assign new_n439 = p_85gat_12_ & new_n438;
  assign new_n440 = new_n438 & ~new_n439;
  assign new_n441 = p_85gat_12_ & ~new_n439;
  assign p_1336gat_586_ = new_n440 | new_n441;
  assign new_n443 = ~new_n245 & new_n396;
  assign new_n444 = p_43gat_6_ & new_n443;
  assign new_n445 = new_n443 & ~new_n444;
  assign new_n446 = p_43gat_6_ & ~new_n444;
  assign p_1330gat_576_ = new_n445 | new_n446;
  assign new_n448 = ~new_n171 & new_n387;
  assign new_n449 = p_78gat_11_ & new_n448;
  assign new_n450 = new_n448 & ~new_n449;
  assign new_n451 = p_78gat_11_ & ~new_n449;
  assign p_1335gat_573_ = new_n450 | new_n451;
  assign new_n453 = ~new_n321 & new_n424;
  assign new_n454 = p_204gat_29_ & new_n453;
  assign new_n455 = new_n453 & ~new_n454;
  assign new_n456 = p_204gat_29_ & ~new_n454;
  assign p_1353gat_566_ = new_n455 | new_n456;
  assign new_n458 = ~new_n208 & new_n396;
  assign new_n459 = p_36gat_5_ & new_n458;
  assign new_n460 = new_n458 & ~new_n459;
  assign new_n461 = p_36gat_5_ & ~new_n459;
  assign p_1329gat_580_ = new_n460 | new_n461;
  assign new_n463 = ~new_n270 & new_n396;
  assign new_n464 = p_29gat_4_ & new_n463;
  assign new_n465 = new_n463 & ~new_n464;
  assign new_n466 = p_29gat_4_ & ~new_n464;
  assign p_1328gat_584_ = new_n465 | new_n466;
  assign new_n468 = new_n171 & ~new_n420;
  assign new_n469 = new_n208 & new_n468;
  assign new_n470 = ~new_n245 & new_n469;
  assign new_n471 = ~new_n270 & new_n470;
  assign new_n472 = ~new_n358 & new_n471;
  assign new_n473 = p_127gat_18_ & new_n472;
  assign new_n474 = new_n472 & ~new_n473;
  assign new_n475 = p_127gat_18_ & ~new_n473;
  assign p_1342gat_559_ = new_n474 | new_n475;
  assign new_n477 = ~new_n208 & new_n468;
  assign new_n478 = ~new_n245 & new_n477;
  assign new_n479 = new_n270 & new_n478;
  assign new_n480 = ~new_n122 & new_n479;
  assign new_n481 = p_190gat_27_ & new_n480;
  assign new_n482 = new_n480 & ~new_n481;
  assign new_n483 = p_190gat_27_ & ~new_n481;
  assign p_1351gat_557_ = new_n482 | new_n483;
  assign new_n485 = ~new_n208 & new_n387;
  assign new_n486 = p_64gat_9_ & new_n485;
  assign new_n487 = new_n485 & ~new_n486;
  assign new_n488 = p_64gat_9_ & ~new_n486;
  assign p_1333gat_581_ = new_n487 | new_n488;
  assign new_n490 = ~new_n321 & new_n479;
  assign new_n491 = p_176gat_25_ & new_n490;
  assign new_n492 = new_n490 & ~new_n491;
  assign new_n493 = p_176gat_25_ & ~new_n491;
  assign p_1349gat_565_ = new_n492 | new_n493;
  assign new_n495 = ~new_n358 & new_n479;
  assign new_n496 = p_183gat_26_ & new_n495;
  assign new_n497 = new_n495 & ~new_n496;
  assign new_n498 = p_183gat_26_ & ~new_n496;
  assign p_1350gat_561_ = new_n497 | new_n498;
  assign new_n500 = ~new_n383 & new_n479;
  assign new_n501 = p_169gat_24_ & new_n500;
  assign new_n502 = new_n500 & ~new_n501;
  assign new_n503 = p_169gat_24_ & ~new_n501;
  assign p_1348gat_569_ = new_n502 | new_n503;
  assign new_n505 = new_n208 & new_n421;
  assign new_n506 = new_n245 & new_n505;
  assign new_n507 = ~new_n270 & new_n506;
  assign new_n508 = ~new_n122 & new_n507;
  assign new_n509 = p_162gat_23_ & new_n508;
  assign new_n510 = new_n508 & ~new_n509;
  assign new_n511 = p_162gat_23_ & ~new_n509;
  assign p_1347gat_556_ = new_n510 | new_n511;
  assign new_n513 = ~new_n321 & new_n471;
  assign new_n514 = p_120gat_17_ & new_n513;
  assign new_n515 = new_n513 & ~new_n514;
  assign new_n516 = p_120gat_17_ & ~new_n514;
  assign p_1341gat_563_ = new_n515 | new_n516;
  assign new_n518 = new_n321 & new_n384;
  assign new_n519 = ~new_n358 & new_n518;
  assign new_n520 = ~new_n383 & new_n519;
  assign new_n521 = ~new_n208 & new_n520;
  assign new_n522 = p_8gat_1_ & new_n521;
  assign new_n523 = new_n521 & ~new_n522;
  assign new_n524 = p_8gat_1_ & ~new_n522;
  assign p_1325gat_579_ = new_n523 | new_n524;
  assign new_n526 = ~new_n245 & new_n520;
  assign new_n527 = p_15gat_2_ & new_n526;
  assign new_n528 = new_n526 & ~new_n527;
  assign new_n529 = p_15gat_2_ & ~new_n527;
  assign p_1326gat_575_ = new_n528 | new_n529;
  assign new_n531 = ~new_n383 & new_n507;
  assign new_n532 = p_141gat_20_ & new_n531;
  assign new_n533 = new_n531 & ~new_n532;
  assign new_n534 = p_141gat_20_ & ~new_n532;
  assign p_1344gat_568_ = new_n533 | new_n534;
  assign new_n536 = ~new_n270 & new_n520;
  assign new_n537 = p_1gat_0_ & new_n536;
  assign new_n538 = new_n536 & ~new_n537;
  assign new_n539 = p_1gat_0_ & ~new_n537;
  assign p_1324gat_583_ = new_n538 | new_n539;
  assign new_n541 = ~new_n122 & new_n471;
  assign new_n542 = p_134gat_19_ & new_n541;
  assign new_n543 = new_n541 & ~new_n542;
  assign new_n544 = p_134gat_19_ & ~new_n542;
  assign p_1343gat_555_ = new_n543 | new_n544;
  assign new_n546 = ~new_n321 & new_n507;
  assign new_n547 = p_148gat_21_ & new_n546;
  assign new_n548 = new_n546 & ~new_n547;
  assign new_n549 = p_148gat_21_ & ~new_n547;
  assign p_1345gat_564_ = new_n548 | new_n549;
  assign new_n551 = ~new_n208 & new_n437;
  assign new_n552 = p_92gat_13_ & new_n551;
  assign new_n553 = new_n551 & ~new_n552;
  assign new_n554 = p_92gat_13_ & ~new_n552;
  assign p_1337gat_582_ = new_n553 | new_n554;
  assign new_n556 = ~new_n171 & new_n520;
  assign new_n557 = p_22gat_3_ & new_n556;
  assign new_n558 = new_n556 & ~new_n557;
  assign new_n559 = p_22gat_3_ & ~new_n557;
  assign p_1327gat_571_ = new_n558 | new_n559;
  assign new_n561 = ~new_n383 & new_n471;
  assign new_n562 = p_113gat_16_ & new_n561;
  assign new_n563 = new_n561 & ~new_n562;
  assign new_n564 = p_113gat_16_ & ~new_n562;
  assign p_1340gat_567_ = new_n563 | new_n564;
  assign new_n566 = ~new_n358 & new_n507;
  assign new_n567 = p_155gat_22_ & new_n566;
  assign new_n568 = new_n566 & ~new_n567;
  assign new_n569 = p_155gat_22_ & ~new_n567;
  assign p_1346gat_560_ = new_n568 | new_n569;
  assign new_n571 = ~new_n171 & new_n437;
  assign new_n572 = p_106gat_15_ & new_n571;
  assign new_n573 = new_n571 & ~new_n572;
  assign new_n574 = p_106gat_15_ & ~new_n572;
  assign p_1339gat_574_ = new_n573 | new_n574;
  assign new_n576 = ~new_n122 & new_n424;
  assign new_n577 = p_218gat_31_ & new_n576;
  assign new_n578 = new_n576 & ~new_n577;
  assign new_n579 = p_218gat_31_ & ~new_n577;
  assign p_1355gat_558_ = new_n578 | new_n579;
  assign new_n581 = ~new_n245 & new_n437;
  assign new_n582 = p_99gat_14_ & new_n581;
  assign new_n583 = new_n581 & ~new_n582;
  assign new_n584 = p_99gat_14_ & ~new_n582;
  assign p_1338gat_578_ = new_n583 | new_n584;
endmodule


