// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pv108_3_, pv109_0_, pv118_4_, pv149_4_, pv257_2_, pv268_0_, pv288_2_,
    pv108_4_, pv118_3_, pv149_5_, pv216_0_, pv257_1_, pv268_1_, pv278_0_,
    pv288_3_, pv289_0_, pv2_0_, pv108_5_, pv118_6_, pv149_6_, pv248_0_,
    pv257_4_, pv288_4_, pv118_5_, pv149_7_, pv207_0_, pv257_3_, pv258_0_,
    pv288_5_, pv60_0_, pv78_1_, pv88_2_, pv118_0_, pv172_0_, pv189_4_,
    pv215_0_, pv257_6_, pv259_0_, pv268_4_, pv78_0_, pv88_3_, pv108_0_,
    pv189_5_, pv199_4_, pv205_0_, pv213_5_, pv234_4_, pv249_0_, pv257_5_,
    pv268_5_, pv302_0_, pv108_1_, pv118_2_, pv223_5_, pv234_3_, pv268_2_,
    pv279_0_, pv288_0_, pv1_0_, pv108_2_, pv118_1_, pv171_0_, pv234_2_,
    pv257_7_, pv268_3_, pv269_0_, pv288_1_, pv4_0_, pv32_7_, pv39_0_,
    pv100_3_, pv101_0_, pv132_0_, pv189_0_, pv199_1_, pv229_1_, pv239_2_,
    pv32_6_, pv38_0_, pv65_0_, pv100_4_, pv189_1_, pv199_0_, pv229_2_,
    pv239_1_, pv245_0_, pv32_5_, pv37_0_, pv62_0_, pv100_5_, pv189_2_,
    pv199_3_, pv239_0_, pv275_0_, pv5_0_, pv32_4_, pv63_0_, pv102_0_,
    pv189_3_, pv199_2_, pv229_0_, pv32_3_, pv35_0_, pv68_0_, pv71_0_,
    pv110_0_, pv149_0_, pv246_0_, pv277_0_, pv295_0_, pv3_0_, pv32_2_,
    pv34_0_, pv69_0_, pv70_0_, pv100_0_, pv118_7_, pv149_1_, pv32_1_,
    pv33_0_, pv66_0_, pv100_1_, pv149_2_, pv169_0_, pv257_0_, pv32_0_,
    pv67_0_, pv100_2_, pv149_3_, pv169_1_, pv247_0_, pv32_10_, pv53_0_,
    pv124_1_, pv165_2_, pv242_0_, pv7_0_, pv32_11_, pv52_0_, pv124_2_,
    pv132_7_, pv134_1_, pv165_3_, pv11_0_, pv55_0_, pv132_6_, pv134_0_,
    pv165_0_, pv262_0_, pv10_0_, pv124_0_, pv132_5_, pv165_1_, pv175_0_,
    pv243_0_, pv272_0_, pv294_0_, pv57_0_, pv132_4_, pv165_6_, pv194_4_,
    pv229_5_, pv56_0_, pv91_1_, pv132_3_, pv165_7_, pv177_0_, pv194_3_,
    pv274_0_, pv292_0_, pv6_0_, pv32_9_, pv40_0_, pv59_0_, pv94_1_,
    pv132_2_, pv165_4_, pv229_3_, pv239_4_, pv244_0_, pv293_0_, pv32_8_,
    pv41_0_, pv94_0_, pv132_1_, pv165_5_, pv229_4_, pv239_3_, pv42_0_,
    pv78_5_, pv84_2_, pv183_2_, pv194_0_, pv213_2_, pv223_3_, pv234_1_,
    pv260_0_, pv291_0_, pv16_0_, pv43_0_, pv78_4_, pv84_3_, pv183_3_,
    pv213_1_, pv223_4_, pv234_0_, pv270_0_, pv44_0_, pv78_3_, pv84_4_,
    pv88_0_, pv91_0_, pv183_4_, pv194_2_, pv204_0_, pv213_4_, pv223_1_,
    pv240_0_, pv301_0_, pv45_0_, pv78_2_, pv84_5_, pv88_1_, pv183_5_,
    pv194_1_, pv213_3_, pv214_0_, pv223_2_, pv8_0_, pv13_0_, pv46_0_,
    pv124_5_, pv202_0_, pv288_6_, pv12_0_, pv223_0_, pv241_0_, pv288_7_,
    pv15_0_, pv48_0_, pv51_0_, pv84_0_, pv124_3_, pv174_0_, pv183_0_,
    pv213_0_, pv271_0_, pv280_0_, pv9_0_, pv14_0_, pv50_0_, pv84_1_,
    pv124_4_, pv183_1_, pv203_0_, pv261_0_, pv290_0_,
    pv778, pv789, pv1213_5_, pv1243_0_, pv1261, pv1371, pv1382, pv1470,
    pv1512_3_, pv1613_1_, pv1757_0_, pv1781_1_, pv1829_2_, pv1953_2_,
    pv375_0_, pv410_0_, pv508_0_, pv539, pv1213_6_, pv1260, pv1372,
    pv1440_0_, pv1758_0_, pv1781_0_, pv1829_1_, pv1953_3_, pv657, pv787,
    pv1213_7_, pv1263, pv1380, pv1759_0_, pv1829_4_, pv1953_4_, pv656,
    pv779, pv1213_8_, pv1262, pv1370, pv1829_3_, pv1953_5_, pv763,
    pv1213_9_, pv1243_4_, pv1265, pv1375, pv1386, pv1481_0_, pv1717_0_,
    pv1829_6_, pv634_0_, pv1243_3_, pv1264, pv1480_0_, pv1741_0_,
    pv1829_5_, pv321_2_, pv512, pv783, pv1243_2_, pv1256, pv1267,
    pv1281_0_, pv1373, pv1384, pv1829_8_, pv1953_0_, pv775, pv784,
    pv1243_1_, pv1257, pv1266, pv1365, pv1374, pv1459_0_, pv1829_7_,
    pv1953_1_, pv543, pv587, pv651, pv781, pv1297_1_, pv1423, pv1771_0_,
    pv1900_0_, pv1921_1_, pv393_0_, pv500_0_, pv544, pv650, pv782,
    pv1213_11_, pv1297_2_, pv1771_1_, pv1921_0_, pv1992_0_, pv541, pv620,
    pv707, pv802_0_, pv1213_10_, pv1274_0_, pv1297_3_, pv1432, pv1726_0_,
    pv1921_3_, pv1968_0_, pv1992_1_, pv357, pv423_0_, pv542, pv621, pv630,
    pv780, pv1297_4_, pv1671_0_, pv1921_2_, pv547, pv655, pv1467_0_,
    pv1629_0_, pv1863_0_, pv1896_0_, pv1921_5_, pv1953_6_, pv377, pv548,
    pv654, pv821_0_, pv1431, pv1897_0_, pv1921_4_, pv1953_7_, pv1960_1_,
    pv527, pv538, pv545, pv653, pv1829_0_, pv1898_0_, pv537, pv546,
    pv597_0_, pv652, pv801, pv1864_0_, pv1899_0_, pv572_8_, pv585_0_,
    pv1709_1_, pv1760_0_, pv373, pv572_7_, pv1439_0_, pv1709_0_, pv572_6_,
    pv1539, pv1719, pv1960_0_, pv572_5_, pv1392_0_, pv1536_0_, pv1679_0_,
    pv1833_0_, pv356, pv435_0_, pv1492_0_, pv1537, pv511_0_, pv540,
    pv609_0_, pv1426, pv1620_0_, pv1736, pv1429, pv1832, pv432, pv572_9_,
    pv1297_0_, pv1428, pv1495_0_, pv1693_0_, pv1901_0_, pv572_0_,
    pv1243_8_, pv1258, pv1243_7_, pv1259, pv1552_0_, pv1745_0_, pv1829_9_,
    pv798_0_, pv1243_6_, pv1552_1_, pv1645_0_, pv1652_0_, pv603_0_,
    pv1213_0_, pv1243_5_, pv1378, pv1387, pv572_4_, pv826_0_, pv1213_1_,
    pv1669, pv572_3_, pv591_0_, pv966, pv1213_2_, pv1709_4_, pv398_0_,
    pv572_2_, pv640_0_, pv1213_3_, pv1512_1_, pv1709_3_, pv572_1_, pv986,
    pv1213_4_, pv1243_9_, pv1451_0_, pv1512_2_, pv1613_0_, pv1709_2_  );
  input  pv108_3_, pv109_0_, pv118_4_, pv149_4_, pv257_2_, pv268_0_,
    pv288_2_, pv108_4_, pv118_3_, pv149_5_, pv216_0_, pv257_1_, pv268_1_,
    pv278_0_, pv288_3_, pv289_0_, pv2_0_, pv108_5_, pv118_6_, pv149_6_,
    pv248_0_, pv257_4_, pv288_4_, pv118_5_, pv149_7_, pv207_0_, pv257_3_,
    pv258_0_, pv288_5_, pv60_0_, pv78_1_, pv88_2_, pv118_0_, pv172_0_,
    pv189_4_, pv215_0_, pv257_6_, pv259_0_, pv268_4_, pv78_0_, pv88_3_,
    pv108_0_, pv189_5_, pv199_4_, pv205_0_, pv213_5_, pv234_4_, pv249_0_,
    pv257_5_, pv268_5_, pv302_0_, pv108_1_, pv118_2_, pv223_5_, pv234_3_,
    pv268_2_, pv279_0_, pv288_0_, pv1_0_, pv108_2_, pv118_1_, pv171_0_,
    pv234_2_, pv257_7_, pv268_3_, pv269_0_, pv288_1_, pv4_0_, pv32_7_,
    pv39_0_, pv100_3_, pv101_0_, pv132_0_, pv189_0_, pv199_1_, pv229_1_,
    pv239_2_, pv32_6_, pv38_0_, pv65_0_, pv100_4_, pv189_1_, pv199_0_,
    pv229_2_, pv239_1_, pv245_0_, pv32_5_, pv37_0_, pv62_0_, pv100_5_,
    pv189_2_, pv199_3_, pv239_0_, pv275_0_, pv5_0_, pv32_4_, pv63_0_,
    pv102_0_, pv189_3_, pv199_2_, pv229_0_, pv32_3_, pv35_0_, pv68_0_,
    pv71_0_, pv110_0_, pv149_0_, pv246_0_, pv277_0_, pv295_0_, pv3_0_,
    pv32_2_, pv34_0_, pv69_0_, pv70_0_, pv100_0_, pv118_7_, pv149_1_,
    pv32_1_, pv33_0_, pv66_0_, pv100_1_, pv149_2_, pv169_0_, pv257_0_,
    pv32_0_, pv67_0_, pv100_2_, pv149_3_, pv169_1_, pv247_0_, pv32_10_,
    pv53_0_, pv124_1_, pv165_2_, pv242_0_, pv7_0_, pv32_11_, pv52_0_,
    pv124_2_, pv132_7_, pv134_1_, pv165_3_, pv11_0_, pv55_0_, pv132_6_,
    pv134_0_, pv165_0_, pv262_0_, pv10_0_, pv124_0_, pv132_5_, pv165_1_,
    pv175_0_, pv243_0_, pv272_0_, pv294_0_, pv57_0_, pv132_4_, pv165_6_,
    pv194_4_, pv229_5_, pv56_0_, pv91_1_, pv132_3_, pv165_7_, pv177_0_,
    pv194_3_, pv274_0_, pv292_0_, pv6_0_, pv32_9_, pv40_0_, pv59_0_,
    pv94_1_, pv132_2_, pv165_4_, pv229_3_, pv239_4_, pv244_0_, pv293_0_,
    pv32_8_, pv41_0_, pv94_0_, pv132_1_, pv165_5_, pv229_4_, pv239_3_,
    pv42_0_, pv78_5_, pv84_2_, pv183_2_, pv194_0_, pv213_2_, pv223_3_,
    pv234_1_, pv260_0_, pv291_0_, pv16_0_, pv43_0_, pv78_4_, pv84_3_,
    pv183_3_, pv213_1_, pv223_4_, pv234_0_, pv270_0_, pv44_0_, pv78_3_,
    pv84_4_, pv88_0_, pv91_0_, pv183_4_, pv194_2_, pv204_0_, pv213_4_,
    pv223_1_, pv240_0_, pv301_0_, pv45_0_, pv78_2_, pv84_5_, pv88_1_,
    pv183_5_, pv194_1_, pv213_3_, pv214_0_, pv223_2_, pv8_0_, pv13_0_,
    pv46_0_, pv124_5_, pv202_0_, pv288_6_, pv12_0_, pv223_0_, pv241_0_,
    pv288_7_, pv15_0_, pv48_0_, pv51_0_, pv84_0_, pv124_3_, pv174_0_,
    pv183_0_, pv213_0_, pv271_0_, pv280_0_, pv9_0_, pv14_0_, pv50_0_,
    pv84_1_, pv124_4_, pv183_1_, pv203_0_, pv261_0_, pv290_0_;
  output pv778, pv789, pv1213_5_, pv1243_0_, pv1261, pv1371, pv1382, pv1470,
    pv1512_3_, pv1613_1_, pv1757_0_, pv1781_1_, pv1829_2_, pv1953_2_,
    pv375_0_, pv410_0_, pv508_0_, pv539, pv1213_6_, pv1260, pv1372,
    pv1440_0_, pv1758_0_, pv1781_0_, pv1829_1_, pv1953_3_, pv657, pv787,
    pv1213_7_, pv1263, pv1380, pv1759_0_, pv1829_4_, pv1953_4_, pv656,
    pv779, pv1213_8_, pv1262, pv1370, pv1829_3_, pv1953_5_, pv763,
    pv1213_9_, pv1243_4_, pv1265, pv1375, pv1386, pv1481_0_, pv1717_0_,
    pv1829_6_, pv634_0_, pv1243_3_, pv1264, pv1480_0_, pv1741_0_,
    pv1829_5_, pv321_2_, pv512, pv783, pv1243_2_, pv1256, pv1267,
    pv1281_0_, pv1373, pv1384, pv1829_8_, pv1953_0_, pv775, pv784,
    pv1243_1_, pv1257, pv1266, pv1365, pv1374, pv1459_0_, pv1829_7_,
    pv1953_1_, pv543, pv587, pv651, pv781, pv1297_1_, pv1423, pv1771_0_,
    pv1900_0_, pv1921_1_, pv393_0_, pv500_0_, pv544, pv650, pv782,
    pv1213_11_, pv1297_2_, pv1771_1_, pv1921_0_, pv1992_0_, pv541, pv620,
    pv707, pv802_0_, pv1213_10_, pv1274_0_, pv1297_3_, pv1432, pv1726_0_,
    pv1921_3_, pv1968_0_, pv1992_1_, pv357, pv423_0_, pv542, pv621, pv630,
    pv780, pv1297_4_, pv1671_0_, pv1921_2_, pv547, pv655, pv1467_0_,
    pv1629_0_, pv1863_0_, pv1896_0_, pv1921_5_, pv1953_6_, pv377, pv548,
    pv654, pv821_0_, pv1431, pv1897_0_, pv1921_4_, pv1953_7_, pv1960_1_,
    pv527, pv538, pv545, pv653, pv1829_0_, pv1898_0_, pv537, pv546,
    pv597_0_, pv652, pv801, pv1864_0_, pv1899_0_, pv572_8_, pv585_0_,
    pv1709_1_, pv1760_0_, pv373, pv572_7_, pv1439_0_, pv1709_0_, pv572_6_,
    pv1539, pv1719, pv1960_0_, pv572_5_, pv1392_0_, pv1536_0_, pv1679_0_,
    pv1833_0_, pv356, pv435_0_, pv1492_0_, pv1537, pv511_0_, pv540,
    pv609_0_, pv1426, pv1620_0_, pv1736, pv1429, pv1832, pv432, pv572_9_,
    pv1297_0_, pv1428, pv1495_0_, pv1693_0_, pv1901_0_, pv572_0_,
    pv1243_8_, pv1258, pv1243_7_, pv1259, pv1552_0_, pv1745_0_, pv1829_9_,
    pv798_0_, pv1243_6_, pv1552_1_, pv1645_0_, pv1652_0_, pv603_0_,
    pv1213_0_, pv1243_5_, pv1378, pv1387, pv572_4_, pv826_0_, pv1213_1_,
    pv1669, pv572_3_, pv591_0_, pv966, pv1213_2_, pv1709_4_, pv398_0_,
    pv572_2_, pv640_0_, pv1213_3_, pv1512_1_, pv1709_3_, pv572_1_, pv986,
    pv1213_4_, pv1243_9_, pv1451_0_, pv1512_2_, pv1613_0_, pv1709_2_;
  wire new_n483, new_n484, new_n485, new_n487, new_n488, new_n489, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1125, new_n1126, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1170,
    new_n1171, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1303, new_n1304, new_n1305, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1355,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1425, new_n1426,
    new_n1428, new_n1429, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1454, new_n1455, new_n1456,
    new_n1457, new_n1458, new_n1459, new_n1460, new_n1461, new_n1462,
    new_n1463, new_n1464, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1470, new_n1471, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1489, new_n1490, new_n1491,
    new_n1493, new_n1494, new_n1495, new_n1496, new_n1497, new_n1498,
    new_n1499, new_n1500, new_n1501, new_n1502, new_n1503, new_n1504,
    new_n1506, new_n1507, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1521, new_n1522, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1544, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1559,
    new_n1560, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1585, new_n1586, new_n1587, new_n1588,
    new_n1589, new_n1590, new_n1591, new_n1592, new_n1593, new_n1594,
    new_n1595, new_n1596, new_n1598, new_n1599, new_n1600, new_n1602,
    new_n1603, new_n1604, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1620, new_n1621, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1628, new_n1629, new_n1630,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1658, new_n1659,
    new_n1661, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1684, new_n1685, new_n1689,
    new_n1691, new_n1692, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1699, new_n1700, new_n1701, new_n1702, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1709, new_n1710, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979,
    new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2046, new_n2047, new_n2048, new_n2050, new_n2051,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2086,
    new_n2087, new_n2088, new_n2089, new_n2090, new_n2091, new_n2092,
    new_n2093, new_n2094, new_n2095, new_n2096, new_n2097, new_n2098,
    new_n2099, new_n2100, new_n2101, new_n2102, new_n2104, new_n2105,
    new_n2106, new_n2109, new_n2110, new_n2111, new_n2112, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2131, new_n2132, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2165, new_n2166, new_n2167, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2182,
    new_n2183, new_n2184, new_n2186, new_n2187, new_n2188, new_n2189,
    new_n2190, new_n2191, new_n2194, new_n2195, new_n2196, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2214, new_n2215, new_n2217, new_n2218, new_n2219,
    new_n2220, new_n2222, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2230, new_n2231, new_n2232, new_n2234, new_n2235, new_n2237,
    new_n2238, new_n2239, new_n2240, new_n2241, new_n2242, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2265, new_n2266,
    new_n2268, new_n2269, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2286, new_n2287, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2321, new_n2322, new_n2323, new_n2325, new_n2326, new_n2327,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2337, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2359, new_n2360, new_n2361, new_n2362,
    new_n2363, new_n2365, new_n2366, new_n2367, new_n2368, new_n2369,
    new_n2370, new_n2371, new_n2372, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2440,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2455, new_n2456, new_n2457,
    new_n2460, new_n2461, new_n2462, new_n2463, new_n2465, new_n2466,
    new_n2468, new_n2469, new_n2470, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2480, new_n2482, new_n2483,
    new_n2484, new_n2485, new_n2486, new_n2487, new_n2488, new_n2489,
    new_n2490, new_n2491, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2503,
    new_n2504, new_n2506, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2559, new_n2560,
    new_n2562, new_n2563, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2571, new_n2572, new_n2573, new_n2574, new_n2576,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628,
    new_n2630, new_n2631, new_n2632, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2644, new_n2645, new_n2646, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2674, new_n2675, new_n2676, new_n2677,
    new_n2678, new_n2679, new_n2680, new_n2681, new_n2682, new_n2684,
    new_n2685, new_n2686, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2730, new_n2731,
    new_n2732, new_n2733, new_n2734, new_n2735, new_n2736, new_n2737,
    new_n2738, new_n2739, new_n2740, new_n2741, new_n2742, new_n2743,
    new_n2744, new_n2745, new_n2746, new_n2747, new_n2748, new_n2749,
    new_n2751, new_n2752, new_n2753;
  assign pv778 = pv5_0_ & pv9_0_;
  assign new_n483 = pv71_0_ & pv202_0_;
  assign new_n484 = ~pv13_0_ & new_n483;
  assign new_n485 = pv4_0_ & ~new_n484;
  assign pv789 = pv9_0_ & new_n485;
  assign new_n487 = pv149_2_ & ~pv149_3_;
  assign new_n488 = ~pv149_0_ & new_n487;
  assign new_n489 = pv149_1_ & new_n488;
  assign new_n490 = pv149_4_ & new_n489;
  assign new_n491 = ~pv174_0_ & new_n490;
  assign new_n492 = ~pv149_0_ & pv149_2_;
  assign new_n493 = ~pv149_1_ & new_n492;
  assign new_n494 = pv149_3_ & new_n493;
  assign new_n495 = ~new_n491 & ~new_n494;
  assign new_n496 = pv60_0_ & ~new_n495;
  assign new_n497 = ~pv149_4_ & ~pv149_3_;
  assign new_n498 = new_n493 & new_n497;
  assign new_n499 = ~pv149_5_ & new_n498;
  assign new_n500 = pv149_4_ & ~pv149_3_;
  assign new_n501 = new_n493 & new_n500;
  assign new_n502 = ~pv149_5_ & new_n501;
  assign new_n503 = pv149_5_ & new_n498;
  assign new_n504 = ~new_n499 & ~new_n502;
  assign new_n505 = ~new_n503 & new_n504;
  assign new_n506 = pv277_0_ & new_n491;
  assign new_n507 = pv278_0_ & ~new_n506;
  assign new_n508 = new_n491 & ~new_n507;
  assign new_n509 = ~pv149_0_ & ~pv149_1_;
  assign new_n510 = ~pv149_2_ & new_n509;
  assign new_n511 = ~pv174_0_ & new_n510;
  assign pv707 = ~pv149_3_ & new_n511;
  assign new_n513 = pv149_4_ & pv707;
  assign new_n514 = ~pv149_5_ & new_n513;
  assign new_n515 = pv149_5_ & new_n513;
  assign new_n516 = pv88_2_ & pv88_3_;
  assign new_n517 = ~pv149_4_ & new_n516;
  assign new_n518 = pv707 & new_n517;
  assign new_n519 = ~pv149_5_ & new_n518;
  assign new_n520 = ~pv88_2_ & pv88_3_;
  assign new_n521 = ~pv149_4_ & new_n520;
  assign new_n522 = pv707 & new_n521;
  assign new_n523 = ~pv149_5_ & new_n522;
  assign new_n524 = pv149_5_ & ~pv88_2_;
  assign new_n525 = ~pv149_3_ & new_n524;
  assign new_n526 = new_n511 & new_n525;
  assign new_n527 = ~pv149_4_ & new_n526;
  assign new_n528 = pv88_3_ & new_n527;
  assign new_n529 = pv149_5_ & pv88_2_;
  assign new_n530 = ~pv149_3_ & new_n529;
  assign new_n531 = new_n511 & new_n530;
  assign new_n532 = ~pv149_4_ & new_n531;
  assign new_n533 = ~pv88_3_ & new_n532;
  assign new_n534 = pv88_2_ & ~pv88_3_;
  assign new_n535 = ~pv149_4_ & new_n534;
  assign new_n536 = pv707 & new_n535;
  assign new_n537 = ~pv149_5_ & new_n536;
  assign new_n538 = ~pv88_3_ & new_n527;
  assign new_n539 = ~new_n514 & ~new_n515;
  assign new_n540 = ~new_n519 & ~new_n523;
  assign new_n541 = new_n539 & new_n540;
  assign new_n542 = ~new_n528 & ~new_n533;
  assign new_n543 = ~new_n537 & ~new_n538;
  assign new_n544 = new_n542 & new_n543;
  assign new_n545 = new_n541 & new_n544;
  assign new_n546 = pv149_3_ & new_n511;
  assign new_n547 = new_n505 & ~new_n508;
  assign new_n548 = new_n545 & new_n547;
  assign new_n549 = ~new_n494 & ~new_n546;
  assign new_n550 = new_n548 & new_n549;
  assign new_n551 = ~pv53_0_ & ~pv56_0_;
  assign new_n552 = ~pv57_0_ & new_n551;
  assign new_n553 = ~new_n493 & ~new_n510;
  assign new_n554 = pv169_1_ & ~new_n553;
  assign new_n555 = ~new_n545 & new_n554;
  assign new_n556 = pv60_0_ & new_n555;
  assign new_n557 = new_n546 & new_n554;
  assign new_n558 = pv56_0_ & new_n557;
  assign new_n559 = pv60_0_ & new_n557;
  assign new_n560 = pv56_0_ & new_n555;
  assign new_n561 = ~new_n556 & ~new_n558;
  assign new_n562 = ~new_n559 & ~new_n560;
  assign new_n563 = new_n561 & new_n562;
  assign new_n564 = ~new_n550 & ~new_n552;
  assign new_n565 = new_n563 & new_n564;
  assign new_n566 = ~pv149_0_ & pv149_1_;
  assign new_n567 = ~pv149_2_ & new_n566;
  assign new_n568 = pv149_4_ & new_n567;
  assign new_n569 = ~pv149_5_ & new_n568;
  assign new_n570 = ~pv149_3_ & new_n569;
  assign new_n571 = pv149_7_ & new_n570;
  assign new_n572 = pv149_6_ & new_n571;
  assign new_n573 = ~pv149_4_ & new_n489;
  assign new_n574 = pv149_1_ & new_n492;
  assign new_n575 = pv149_3_ & new_n574;
  assign new_n576 = ~pv165_6_ & ~pv165_4_;
  assign new_n577 = ~pv165_5_ & new_n576;
  assign new_n578 = pv165_3_ & new_n577;
  assign new_n579 = pv70_0_ & new_n578;
  assign new_n580 = pv149_5_ & new_n568;
  assign new_n581 = ~pv149_3_ & new_n580;
  assign new_n582 = pv149_7_ & new_n581;
  assign new_n583 = pv149_6_ & new_n582;
  assign new_n584 = ~pv149_7_ & new_n581;
  assign new_n585 = pv149_6_ & new_n584;
  assign new_n586 = ~new_n583 & ~new_n585;
  assign pv802_0_ = pv52_0_ | pv51_0_;
  assign new_n588 = ~new_n586 & ~pv802_0_;
  assign new_n589 = ~pv55_0_ & new_n588;
  assign new_n590 = ~new_n490 & ~new_n510;
  assign new_n591 = ~new_n589 & new_n590;
  assign new_n592 = ~pv292_0_ & ~new_n579;
  assign new_n593 = ~new_n591 & new_n592;
  assign new_n594 = ~pv291_0_ & new_n593;
  assign pv763 = pv169_0_ & new_n594;
  assign new_n596 = pv165_3_ & pv165_5_;
  assign new_n597 = pv165_7_ & new_n596;
  assign new_n598 = pv261_0_ & new_n597;
  assign new_n599 = pv70_0_ & new_n598;
  assign new_n600 = pv763 & new_n599;
  assign new_n601 = pv165_2_ & new_n600;
  assign new_n602 = pv165_0_ & new_n601;
  assign new_n603 = pv165_1_ & new_n602;
  assign new_n604 = pv165_4_ & new_n603;
  assign new_n605 = pv165_6_ & new_n604;
  assign new_n606 = pv165_3_ & pv165_4_;
  assign new_n607 = pv165_6_ & new_n606;
  assign new_n608 = pv165_5_ & new_n607;
  assign new_n609 = pv165_7_ & new_n608;
  assign new_n610 = pv165_2_ & new_n609;
  assign new_n611 = pv165_0_ & new_n610;
  assign new_n612 = pv165_1_ & new_n611;
  assign new_n613 = pv261_0_ & new_n612;
  assign new_n614 = ~pv204_0_ & new_n613;
  assign new_n615 = ~new_n605 & ~new_n614;
  assign new_n616 = ~pv262_0_ & new_n615;
  assign new_n617 = pv53_0_ & ~pv56_0_;
  assign new_n618 = ~new_n573 & new_n617;
  assign new_n619 = ~new_n575 & new_n618;
  assign new_n620 = new_n616 & new_n619;
  assign new_n621 = ~new_n565 & ~new_n572;
  assign new_n622 = ~new_n620 & new_n621;
  assign new_n623 = ~new_n496 & ~new_n622;
  assign new_n624 = pv763 & new_n616;
  assign new_n625 = new_n507 & new_n575;
  assign new_n626 = ~new_n491 & new_n553;
  assign new_n627 = ~new_n573 & new_n626;
  assign new_n628 = ~pv174_0_ & ~new_n627;
  assign new_n629 = ~pv60_0_ & ~pv59_0_;
  assign new_n630 = ~new_n507 & ~new_n629;
  assign new_n631 = new_n575 & new_n630;
  assign new_n632 = ~new_n625 & ~new_n628;
  assign new_n633 = ~new_n631 & new_n632;
  assign new_n634 = ~new_n507 & new_n575;
  assign new_n635 = ~pv59_0_ & new_n634;
  assign new_n636 = ~new_n616 & new_n633;
  assign new_n637 = ~new_n635 & new_n636;
  assign new_n638 = pv257_0_ & new_n637;
  assign new_n639 = ~new_n491 & ~new_n575;
  assign new_n640 = ~new_n573 & new_n639;
  assign new_n641 = ~new_n553 & new_n640;
  assign new_n642 = pv223_5_ & new_n641;
  assign new_n643 = new_n553 & ~new_n640;
  assign new_n644 = pv183_5_ & new_n643;
  assign new_n645 = ~new_n642 & ~new_n644;
  assign new_n646 = new_n616 & ~new_n633;
  assign new_n647 = ~new_n635 & new_n646;
  assign new_n648 = ~new_n645 & new_n647;
  assign new_n649 = ~new_n638 & ~new_n648;
  assign new_n650 = ~new_n624 & ~new_n649;
  assign new_n651 = ~pv56_0_ & ~pv59_0_;
  assign new_n652 = ~pv60_0_ & new_n651;
  assign new_n653 = pv763 & ~new_n652;
  assign new_n654 = new_n624 & ~new_n653;
  assign new_n655 = new_n624 & new_n654;
  assign new_n656 = ~new_n653 & new_n655;
  assign new_n657 = ~new_n650 & ~new_n656;
  assign new_n658 = new_n622 & ~new_n623;
  assign new_n659 = ~new_n657 & new_n658;
  assign new_n660 = ~new_n622 & new_n623;
  assign new_n661 = pv32_5_ & new_n660;
  assign pv1213_5_ = new_n659 | new_n661;
  assign new_n663 = new_n575 & new_n616;
  assign new_n664 = ~pv59_0_ & new_n663;
  assign new_n665 = ~new_n507 & new_n664;
  assign new_n666 = pv149_4_ & new_n665;
  assign new_n667 = new_n633 & new_n666;
  assign new_n668 = pv257_7_ & new_n637;
  assign new_n669 = pv234_0_ & new_n641;
  assign new_n670 = pv194_0_ & new_n643;
  assign new_n671 = ~new_n669 & ~new_n670;
  assign new_n672 = new_n647 & ~new_n671;
  assign new_n673 = ~new_n667 & ~new_n668;
  assign new_n674 = ~new_n672 & new_n673;
  assign new_n675 = ~new_n624 & ~new_n674;
  assign new_n676 = pv32_2_ & new_n653;
  assign new_n677 = pv32_5_ & ~new_n653;
  assign new_n678 = ~new_n676 & ~new_n677;
  assign new_n679 = new_n624 & ~new_n678;
  assign new_n680 = ~new_n675 & ~new_n679;
  assign new_n681 = new_n658 & ~new_n680;
  assign new_n682 = pv78_4_ & new_n660;
  assign pv321_2_ = ~new_n681 & ~new_n682;
  assign pv1260 = pv3_0_ & pv11_0_;
  assign pv1261 = ~pv62_0_ & pv1260;
  assign new_n686 = pv268_4_ & pv268_3_;
  assign new_n687 = pv268_2_ & new_n686;
  assign new_n688 = pv268_5_ & new_n687;
  assign new_n689 = pv268_1_ & ~new_n688;
  assign new_n690 = ~pv268_1_ & new_n688;
  assign pv1371 = new_n689 | new_n690;
  assign new_n692 = pv10_0_ & ~pv13_0_;
  assign new_n693 = ~new_n493 & ~new_n511;
  assign new_n694 = pv802_0_ & ~new_n693;
  assign new_n695 = ~new_n494 & ~new_n694;
  assign pv782 = pv7_0_ & new_n692;
  assign pv1382 = ~new_n695 & pv782;
  assign new_n698 = pv165_0_ & pv165_1_;
  assign new_n699 = ~pv165_2_ & new_n698;
  assign new_n700 = pv165_7_ & new_n699;
  assign new_n701 = ~pv290_0_ & new_n700;
  assign new_n702 = ~pv165_7_ & new_n699;
  assign new_n703 = pv172_0_ & pv56_0_;
  assign new_n704 = pv207_0_ & ~new_n703;
  assign new_n705 = pv59_0_ & new_n554;
  assign new_n706 = new_n704 & new_n705;
  assign new_n707 = ~new_n493 & new_n706;
  assign new_n708 = ~pv149_4_ & new_n567;
  assign new_n709 = pv149_5_ & new_n708;
  assign new_n710 = ~pv149_3_ & new_n709;
  assign new_n711 = ~pv149_7_ & new_n710;
  assign new_n712 = ~pv149_6_ & new_n711;
  assign new_n713 = ~pv174_0_ & new_n583;
  assign new_n714 = ~new_n554 & ~new_n712;
  assign new_n715 = new_n704 & new_n714;
  assign new_n716 = ~new_n713 & new_n715;
  assign new_n717 = ~new_n493 & new_n716;
  assign new_n718 = pv172_0_ & pv215_0_;
  assign new_n719 = pv67_0_ & new_n718;
  assign new_n720 = pv59_0_ & new_n713;
  assign new_n721 = new_n704 & new_n720;
  assign new_n722 = ~new_n493 & new_n721;
  assign new_n723 = pv62_0_ & new_n712;
  assign new_n724 = new_n704 & new_n723;
  assign new_n725 = ~new_n493 & new_n724;
  assign new_n726 = ~pv214_0_ & ~new_n707;
  assign new_n727 = ~new_n717 & new_n726;
  assign new_n728 = ~new_n719 & ~new_n722;
  assign new_n729 = ~new_n725 & new_n728;
  assign new_n730 = new_n727 & new_n729;
  assign new_n731 = pv241_0_ & ~new_n639;
  assign new_n732 = ~new_n573 & ~new_n731;
  assign new_n733 = ~pv275_0_ & pv272_0_;
  assign new_n734 = ~new_n732 & new_n733;
  assign new_n735 = ~pv802_0_ & new_n734;
  assign new_n736 = pv261_0_ & new_n735;
  assign new_n737 = new_n507 & new_n736;
  assign new_n738 = pv261_0_ & ~pv802_0_;
  assign new_n739 = ~new_n732 & new_n738;
  assign new_n740 = ~new_n507 & new_n739;
  assign new_n741 = pv56_0_ & ~new_n639;
  assign new_n742 = ~pv802_0_ & ~new_n640;
  assign new_n743 = ~new_n507 & new_n742;
  assign new_n744 = pv242_0_ & new_n743;
  assign new_n745 = ~new_n741 & new_n744;
  assign new_n746 = pv272_0_ & ~pv802_0_;
  assign new_n747 = pv134_0_ & new_n746;
  assign new_n748 = pv242_0_ & new_n747;
  assign new_n749 = pv134_1_ & new_n748;
  assign new_n750 = ~pv275_0_ & new_n749;
  assign new_n751 = new_n507 & new_n750;
  assign new_n752 = new_n730 & ~new_n737;
  assign new_n753 = ~new_n740 & new_n752;
  assign new_n754 = ~new_n745 & ~new_n751;
  assign new_n755 = new_n753 & new_n754;
  assign new_n756 = ~new_n701 & ~new_n702;
  assign new_n757 = ~pv302_0_ & new_n755;
  assign new_n758 = new_n756 & new_n757;
  assign new_n759 = ~pv149_5_ & new_n708;
  assign new_n760 = ~pv149_3_ & new_n759;
  assign new_n761 = pv149_7_ & new_n760;
  assign new_n762 = pv149_6_ & new_n761;
  assign new_n763 = pv67_0_ & pv14_0_;
  assign new_n764 = new_n758 & new_n763;
  assign pv1470 = ~new_n762 & new_n764;
  assign new_n766 = pv149_5_ & new_n501;
  assign new_n767 = pv88_3_ & new_n532;
  assign new_n768 = ~pv88_2_ & ~pv88_3_;
  assign new_n769 = ~pv149_4_ & new_n768;
  assign new_n770 = pv707 & new_n769;
  assign new_n771 = ~pv149_5_ & new_n770;
  assign new_n772 = ~new_n767 & ~new_n771;
  assign new_n773 = ~new_n554 & ~new_n772;
  assign new_n774 = ~new_n766 & ~new_n773;
  assign new_n775 = pv56_0_ & ~new_n774;
  assign new_n776 = ~pv172_0_ & new_n775;
  assign new_n777 = pv278_0_ & ~new_n640;
  assign new_n778 = pv171_0_ & ~new_n553;
  assign new_n779 = pv56_0_ & new_n778;
  assign new_n780 = ~pv248_0_ & ~new_n703;
  assign new_n781 = ~new_n777 & new_n780;
  assign new_n782 = pv177_0_ & new_n781;
  assign new_n783 = ~new_n779 & new_n782;
  assign new_n784 = ~pv274_0_ & ~pv271_0_;
  assign new_n785 = new_n554 & ~new_n772;
  assign new_n786 = pv59_0_ & new_n785;
  assign new_n787 = ~new_n776 & ~new_n783;
  assign new_n788 = ~new_n784 & new_n787;
  assign new_n789 = ~new_n786 & new_n788;
  assign new_n790 = new_n493 & new_n704;
  assign new_n791 = pv149_7_ & new_n493;
  assign new_n792 = pv56_0_ & new_n791;
  assign new_n793 = ~new_n790 & ~new_n792;
  assign new_n794 = ~new_n789 & new_n793;
  assign pv1536_0_ = ~new_n755 | ~new_n794;
  assign new_n796 = new_n755 & pv1536_0_;
  assign new_n797 = pv223_2_ & new_n641;
  assign new_n798 = pv183_2_ & new_n643;
  assign new_n799 = ~new_n797 & ~new_n798;
  assign new_n800 = new_n616 & ~new_n635;
  assign new_n801 = ~new_n633 & new_n800;
  assign new_n802 = ~new_n799 & new_n801;
  assign new_n803 = ~new_n624 & new_n802;
  assign new_n804 = new_n622 & new_n803;
  assign new_n805 = ~new_n624 & new_n804;
  assign new_n806 = ~new_n623 & new_n805;
  assign new_n807 = pv32_2_ & new_n660;
  assign pv1213_2_ = new_n806 | new_n807;
  assign new_n809 = pv223_3_ & new_n641;
  assign new_n810 = pv183_3_ & new_n643;
  assign new_n811 = ~new_n809 & ~new_n810;
  assign new_n812 = new_n801 & ~new_n811;
  assign new_n813 = ~new_n624 & new_n812;
  assign new_n814 = new_n622 & new_n813;
  assign new_n815 = ~new_n624 & new_n814;
  assign new_n816 = ~new_n623 & new_n815;
  assign new_n817 = pv32_3_ & new_n660;
  assign pv1213_3_ = new_n816 | new_n817;
  assign new_n819 = pv223_1_ & new_n641;
  assign new_n820 = pv183_1_ & new_n643;
  assign new_n821 = ~new_n819 & ~new_n820;
  assign new_n822 = new_n801 & ~new_n821;
  assign new_n823 = ~new_n624 & new_n822;
  assign new_n824 = new_n622 & new_n823;
  assign new_n825 = ~new_n624 & new_n824;
  assign new_n826 = ~new_n623 & new_n825;
  assign new_n827 = pv32_1_ & new_n660;
  assign pv1213_1_ = new_n826 | new_n827;
  assign new_n829 = pv223_0_ & new_n641;
  assign new_n830 = pv183_0_ & new_n643;
  assign new_n831 = ~new_n829 & ~new_n830;
  assign new_n832 = new_n801 & ~new_n831;
  assign new_n833 = ~new_n624 & new_n832;
  assign new_n834 = new_n622 & new_n833;
  assign new_n835 = ~new_n624 & new_n834;
  assign new_n836 = ~new_n623 & new_n835;
  assign new_n837 = pv32_0_ & new_n660;
  assign pv1213_0_ = new_n836 | new_n837;
  assign new_n839 = pv149_3_ & new_n759;
  assign new_n840 = ~pv149_7_ & new_n839;
  assign new_n841 = ~pv149_6_ & new_n840;
  assign new_n842 = ~pv802_0_ & new_n841;
  assign new_n843 = pv1213_2_ & pv1213_3_;
  assign new_n844 = ~pv1213_1_ & new_n843;
  assign new_n845 = ~pv1213_0_ & new_n844;
  assign new_n846 = ~new_n842 & new_n845;
  assign new_n847 = pv288_6_ & new_n846;
  assign new_n848 = pv288_7_ & new_n847;
  assign new_n849 = ~pv1213_3_ & ~pv1213_0_;
  assign new_n850 = pv1213_2_ & new_n849;
  assign new_n851 = ~pv1213_1_ & new_n850;
  assign new_n852 = ~new_n842 & new_n851;
  assign new_n853 = pv288_6_ & new_n852;
  assign new_n854 = pv288_7_ & new_n853;
  assign new_n855 = ~pv288_6_ & pv288_7_;
  assign new_n856 = ~pv288_4_ & pv288_5_;
  assign new_n857 = new_n855 & new_n856;
  assign new_n858 = ~new_n855 & ~new_n856;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = ~pv288_2_ & pv288_3_;
  assign new_n861 = ~new_n859 & new_n860;
  assign new_n862 = pv288_2_ & ~pv288_3_;
  assign new_n863 = new_n861 & new_n862;
  assign new_n864 = ~new_n855 & new_n856;
  assign new_n865 = pv288_6_ & ~pv288_7_;
  assign new_n866 = ~new_n855 & ~new_n865;
  assign new_n867 = pv288_4_ & ~pv288_5_;
  assign new_n868 = ~new_n866 & new_n867;
  assign new_n869 = new_n866 & ~new_n867;
  assign new_n870 = ~new_n868 & ~new_n869;
  assign new_n871 = ~new_n864 & ~new_n870;
  assign new_n872 = new_n864 & new_n870;
  assign new_n873 = ~new_n871 & ~new_n872;
  assign new_n874 = new_n862 & ~new_n873;
  assign new_n875 = new_n861 & ~new_n873;
  assign new_n876 = ~new_n863 & ~new_n874;
  assign new_n877 = ~new_n875 & new_n876;
  assign new_n878 = pv288_2_ & pv288_3_;
  assign new_n879 = ~new_n877 & new_n878;
  assign new_n880 = ~pv288_6_ & ~pv288_7_;
  assign new_n881 = pv288_4_ & pv288_5_;
  assign new_n882 = ~new_n880 & new_n881;
  assign new_n883 = new_n880 & ~new_n881;
  assign new_n884 = ~new_n882 & ~new_n883;
  assign new_n885 = new_n864 & new_n867;
  assign new_n886 = new_n866 & new_n867;
  assign new_n887 = new_n864 & new_n866;
  assign new_n888 = ~new_n885 & ~new_n886;
  assign new_n889 = ~new_n887 & new_n888;
  assign new_n890 = new_n884 & ~new_n889;
  assign new_n891 = ~new_n884 & new_n889;
  assign new_n892 = ~new_n890 & ~new_n891;
  assign new_n893 = new_n878 & ~new_n892;
  assign new_n894 = ~new_n877 & ~new_n892;
  assign new_n895 = ~new_n879 & ~new_n893;
  assign new_n896 = ~new_n894 & new_n895;
  assign new_n897 = new_n881 & ~new_n889;
  assign new_n898 = new_n880 & new_n881;
  assign new_n899 = new_n880 & ~new_n889;
  assign new_n900 = ~new_n897 & ~new_n898;
  assign new_n901 = ~new_n899 & new_n900;
  assign new_n902 = new_n880 & new_n901;
  assign new_n903 = ~new_n880 & ~new_n901;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = new_n896 & ~new_n904;
  assign new_n906 = ~new_n896 & new_n904;
  assign new_n907 = ~new_n905 & ~new_n906;
  assign new_n908 = ~pv1213_0_ & ~new_n907;
  assign new_n909 = pv1213_0_ & new_n907;
  assign new_n910 = ~new_n908 & ~new_n909;
  assign new_n911 = new_n862 & new_n873;
  assign new_n912 = ~new_n862 & ~new_n873;
  assign new_n913 = ~new_n911 & ~new_n912;
  assign new_n914 = ~new_n861 & ~new_n913;
  assign new_n915 = new_n861 & new_n913;
  assign new_n916 = ~new_n914 & ~new_n915;
  assign new_n917 = ~pv1213_2_ & ~new_n916;
  assign new_n918 = pv1213_2_ & new_n916;
  assign new_n919 = ~new_n917 & ~new_n918;
  assign new_n920 = new_n859 & new_n860;
  assign new_n921 = ~new_n859 & ~new_n860;
  assign new_n922 = ~new_n920 & ~new_n921;
  assign new_n923 = ~pv1213_3_ & ~new_n922;
  assign new_n924 = pv1213_3_ & new_n922;
  assign new_n925 = ~new_n923 & ~new_n924;
  assign new_n926 = new_n878 & new_n892;
  assign new_n927 = ~new_n878 & ~new_n892;
  assign new_n928 = ~new_n926 & ~new_n927;
  assign new_n929 = ~new_n877 & new_n928;
  assign new_n930 = new_n877 & ~new_n928;
  assign new_n931 = ~new_n929 & ~new_n930;
  assign new_n932 = ~pv1213_1_ & ~new_n931;
  assign new_n933 = pv1213_1_ & new_n931;
  assign new_n934 = ~new_n932 & ~new_n933;
  assign new_n935 = new_n910 & new_n919;
  assign new_n936 = new_n925 & new_n935;
  assign new_n937 = new_n934 & new_n936;
  assign new_n938 = ~new_n842 & new_n937;
  assign new_n939 = new_n878 & new_n938;
  assign new_n940 = ~pv1213_0_ & ~new_n904;
  assign new_n941 = pv1213_0_ & new_n904;
  assign new_n942 = ~new_n940 & ~new_n941;
  assign new_n943 = ~pv1213_2_ & ~new_n873;
  assign new_n944 = pv1213_2_ & new_n873;
  assign new_n945 = ~new_n943 & ~new_n944;
  assign new_n946 = ~pv1213_3_ & ~new_n859;
  assign new_n947 = pv1213_3_ & new_n859;
  assign new_n948 = ~new_n946 & ~new_n947;
  assign new_n949 = ~pv1213_1_ & ~new_n892;
  assign new_n950 = pv1213_1_ & new_n892;
  assign new_n951 = ~new_n949 & ~new_n950;
  assign new_n952 = new_n942 & new_n945;
  assign new_n953 = new_n948 & new_n952;
  assign new_n954 = new_n951 & new_n953;
  assign new_n955 = ~new_n842 & new_n954;
  assign new_n956 = new_n881 & new_n955;
  assign new_n957 = ~pv288_0_ & pv288_1_;
  assign new_n958 = ~new_n922 & new_n957;
  assign new_n959 = pv288_0_ & ~pv288_1_;
  assign new_n960 = new_n958 & new_n959;
  assign new_n961 = ~new_n916 & new_n959;
  assign new_n962 = ~new_n916 & new_n958;
  assign new_n963 = ~new_n960 & ~new_n961;
  assign new_n964 = ~new_n962 & new_n963;
  assign new_n965 = pv288_0_ & pv288_1_;
  assign new_n966 = ~new_n964 & new_n965;
  assign new_n967 = ~new_n931 & new_n965;
  assign new_n968 = ~new_n931 & ~new_n964;
  assign new_n969 = ~new_n966 & ~new_n967;
  assign new_n970 = ~new_n968 & new_n969;
  assign new_n971 = ~new_n907 & new_n970;
  assign new_n972 = new_n907 & ~new_n970;
  assign new_n973 = ~new_n971 & ~new_n972;
  assign new_n974 = ~pv1213_0_ & ~new_n973;
  assign new_n975 = pv1213_0_ & new_n973;
  assign new_n976 = ~new_n974 & ~new_n975;
  assign new_n977 = new_n916 & new_n959;
  assign new_n978 = ~new_n916 & ~new_n959;
  assign new_n979 = ~new_n977 & ~new_n978;
  assign new_n980 = ~new_n958 & ~new_n979;
  assign new_n981 = new_n958 & new_n979;
  assign new_n982 = ~new_n980 & ~new_n981;
  assign new_n983 = ~pv1213_2_ & ~new_n982;
  assign new_n984 = pv1213_2_ & new_n982;
  assign new_n985 = ~new_n983 & ~new_n984;
  assign new_n986 = new_n922 & new_n957;
  assign new_n987 = ~new_n922 & ~new_n957;
  assign new_n988 = ~new_n986 & ~new_n987;
  assign new_n989 = ~pv1213_3_ & ~new_n988;
  assign new_n990 = pv1213_3_ & new_n988;
  assign new_n991 = ~new_n989 & ~new_n990;
  assign new_n992 = new_n931 & new_n965;
  assign new_n993 = ~new_n931 & ~new_n965;
  assign new_n994 = ~new_n992 & ~new_n993;
  assign new_n995 = ~new_n964 & new_n994;
  assign new_n996 = new_n964 & ~new_n994;
  assign new_n997 = ~new_n995 & ~new_n996;
  assign new_n998 = ~pv1213_1_ & ~new_n997;
  assign new_n999 = pv1213_1_ & new_n997;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = new_n976 & new_n985;
  assign new_n1002 = new_n991 & new_n1001;
  assign new_n1003 = new_n1000 & new_n1002;
  assign new_n1004 = ~new_n842 & new_n1003;
  assign new_n1005 = new_n965 & new_n1004;
  assign new_n1006 = new_n982 & new_n988;
  assign new_n1007 = new_n997 & new_n1006;
  assign new_n1008 = ~new_n973 & ~new_n1007;
  assign new_n1009 = new_n973 & new_n1007;
  assign new_n1010 = ~new_n1008 & ~new_n1009;
  assign new_n1011 = ~pv1213_0_ & ~new_n1010;
  assign new_n1012 = pv1213_0_ & new_n1010;
  assign new_n1013 = ~new_n1011 & ~new_n1012;
  assign new_n1014 = ~new_n982 & ~new_n988;
  assign new_n1015 = ~new_n1006 & ~new_n1014;
  assign new_n1016 = ~pv1213_2_ & ~new_n1015;
  assign new_n1017 = pv1213_2_ & new_n1015;
  assign new_n1018 = ~new_n1016 & ~new_n1017;
  assign new_n1019 = ~pv1213_3_ & new_n988;
  assign new_n1020 = pv1213_3_ & ~new_n988;
  assign new_n1021 = ~new_n1019 & ~new_n1020;
  assign new_n1022 = ~new_n997 & ~new_n1006;
  assign new_n1023 = ~new_n1007 & ~new_n1022;
  assign new_n1024 = ~pv1213_1_ & ~new_n1023;
  assign new_n1025 = pv1213_1_ & new_n1023;
  assign new_n1026 = ~new_n1024 & ~new_n1025;
  assign new_n1027 = new_n1013 & new_n1018;
  assign new_n1028 = new_n1021 & new_n1027;
  assign new_n1029 = new_n1026 & new_n1028;
  assign new_n1030 = ~new_n842 & new_n1029;
  assign new_n1031 = new_n965 & new_n1030;
  assign new_n1032 = new_n859 & new_n873;
  assign new_n1033 = new_n892 & new_n1032;
  assign new_n1034 = ~new_n904 & ~new_n1033;
  assign new_n1035 = new_n904 & new_n1033;
  assign new_n1036 = ~new_n1034 & ~new_n1035;
  assign new_n1037 = ~pv1213_0_ & ~new_n1036;
  assign new_n1038 = pv1213_0_ & new_n1036;
  assign new_n1039 = ~new_n1037 & ~new_n1038;
  assign new_n1040 = ~new_n859 & ~new_n873;
  assign new_n1041 = ~new_n1032 & ~new_n1040;
  assign new_n1042 = ~pv1213_2_ & ~new_n1041;
  assign new_n1043 = pv1213_2_ & new_n1041;
  assign new_n1044 = ~new_n1042 & ~new_n1043;
  assign new_n1045 = ~pv1213_3_ & new_n859;
  assign new_n1046 = pv1213_3_ & ~new_n859;
  assign new_n1047 = ~new_n1045 & ~new_n1046;
  assign new_n1048 = ~new_n892 & ~new_n1032;
  assign new_n1049 = ~new_n1033 & ~new_n1048;
  assign new_n1050 = ~pv1213_1_ & ~new_n1049;
  assign new_n1051 = pv1213_1_ & new_n1049;
  assign new_n1052 = ~new_n1050 & ~new_n1051;
  assign new_n1053 = new_n1039 & new_n1044;
  assign new_n1054 = new_n1047 & new_n1053;
  assign new_n1055 = new_n1052 & new_n1054;
  assign new_n1056 = ~new_n842 & new_n1055;
  assign new_n1057 = new_n881 & new_n1056;
  assign new_n1058 = new_n916 & new_n922;
  assign new_n1059 = new_n931 & new_n1058;
  assign new_n1060 = ~new_n907 & ~new_n1059;
  assign new_n1061 = new_n907 & new_n1059;
  assign new_n1062 = ~new_n1060 & ~new_n1061;
  assign new_n1063 = ~pv1213_0_ & ~new_n1062;
  assign new_n1064 = pv1213_0_ & new_n1062;
  assign new_n1065 = ~new_n1063 & ~new_n1064;
  assign new_n1066 = ~new_n916 & ~new_n922;
  assign new_n1067 = ~new_n1058 & ~new_n1066;
  assign new_n1068 = ~pv1213_2_ & ~new_n1067;
  assign new_n1069 = pv1213_2_ & new_n1067;
  assign new_n1070 = ~new_n1068 & ~new_n1069;
  assign new_n1071 = ~pv1213_3_ & new_n922;
  assign new_n1072 = pv1213_3_ & ~new_n922;
  assign new_n1073 = ~new_n1071 & ~new_n1072;
  assign new_n1074 = ~new_n931 & ~new_n1058;
  assign new_n1075 = ~new_n1059 & ~new_n1074;
  assign new_n1076 = ~pv1213_1_ & ~new_n1075;
  assign new_n1077 = pv1213_1_ & new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = new_n1065 & new_n1070;
  assign new_n1080 = new_n1073 & new_n1079;
  assign new_n1081 = new_n1078 & new_n1080;
  assign new_n1082 = ~new_n842 & new_n1081;
  assign new_n1083 = new_n878 & new_n1082;
  assign new_n1084 = ~new_n848 & ~new_n854;
  assign new_n1085 = ~new_n939 & new_n1084;
  assign new_n1086 = ~new_n956 & new_n1085;
  assign new_n1087 = ~new_n1005 & new_n1086;
  assign new_n1088 = ~new_n1031 & new_n1087;
  assign new_n1089 = ~new_n1057 & new_n1088;
  assign new_n1090 = ~new_n1083 & new_n1089;
  assign new_n1091 = ~pv1536_0_ & ~new_n1090;
  assign pv1512_3_ = new_n796 | new_n1091;
  assign new_n1093 = pv149_6_ & new_n840;
  assign new_n1094 = ~pv149_7_ & new_n570;
  assign new_n1095 = ~pv149_6_ & new_n1094;
  assign new_n1096 = ~pv149_6_ & new_n571;
  assign new_n1097 = ~new_n1093 & new_n1095;
  assign new_n1098 = ~new_n1096 & new_n1097;
  assign new_n1099 = pv132_2_ & new_n1098;
  assign new_n1100 = ~new_n1093 & ~new_n1095;
  assign new_n1101 = new_n1096 & new_n1100;
  assign new_n1102 = pv118_0_ & new_n1101;
  assign pv1953_2_ = new_n1099 | new_n1102;
  assign new_n1104 = pv132_3_ & new_n1098;
  assign new_n1105 = pv118_1_ & new_n1101;
  assign pv1953_3_ = new_n1104 | new_n1105;
  assign new_n1107 = ~pv1953_2_ & pv1953_3_;
  assign new_n1108 = pv1953_2_ & ~pv1953_3_;
  assign new_n1109 = ~new_n1107 & ~new_n1108;
  assign new_n1110 = pv132_4_ & new_n1098;
  assign new_n1111 = pv118_2_ & new_n1101;
  assign pv1953_4_ = new_n1110 | new_n1111;
  assign new_n1113 = pv132_5_ & new_n1098;
  assign new_n1114 = pv118_3_ & new_n1101;
  assign pv1953_5_ = new_n1113 | new_n1114;
  assign new_n1116 = ~pv1953_4_ & pv1953_5_;
  assign new_n1117 = pv1953_4_ & ~pv1953_5_;
  assign new_n1118 = ~new_n1116 & ~new_n1117;
  assign new_n1119 = new_n1109 & ~new_n1118;
  assign new_n1120 = ~new_n1109 & new_n1118;
  assign new_n1121 = ~new_n1119 & ~new_n1120;
  assign new_n1122 = pv132_6_ & new_n1098;
  assign new_n1123 = pv118_4_ & new_n1101;
  assign pv1953_6_ = new_n1122 | new_n1123;
  assign new_n1125 = pv132_7_ & new_n1098;
  assign new_n1126 = pv118_5_ & new_n1101;
  assign pv1953_7_ = new_n1125 | new_n1126;
  assign new_n1128 = ~pv1953_6_ & pv1953_7_;
  assign new_n1129 = pv1953_6_ & ~pv1953_7_;
  assign new_n1130 = ~new_n1128 & ~new_n1129;
  assign new_n1131 = pv149_7_ & new_n710;
  assign new_n1132 = pv149_6_ & new_n1131;
  assign new_n1133 = pv149_6_ & new_n711;
  assign new_n1134 = ~new_n1132 & ~new_n1133;
  assign new_n1135 = new_n1096 & new_n1134;
  assign new_n1136 = pv118_6_ & new_n1135;
  assign new_n1137 = ~new_n1096 & ~new_n1134;
  assign new_n1138 = pv48_0_ & new_n1137;
  assign pv1960_0_ = new_n1136 | new_n1138;
  assign new_n1140 = pv118_7_ & new_n1135;
  assign new_n1141 = pv46_0_ & new_n1137;
  assign pv1960_1_ = new_n1140 | new_n1141;
  assign new_n1143 = ~pv1960_0_ & pv1960_1_;
  assign new_n1144 = pv1960_0_ & ~pv1960_1_;
  assign new_n1145 = ~new_n1143 & ~new_n1144;
  assign new_n1146 = new_n1130 & ~new_n1145;
  assign new_n1147 = ~new_n1130 & new_n1145;
  assign new_n1148 = ~new_n1146 & ~new_n1147;
  assign new_n1149 = new_n1121 & ~new_n1148;
  assign new_n1150 = ~new_n1121 & new_n1148;
  assign pv1613_1_ = ~new_n1149 & ~new_n1150;
  assign new_n1152 = ~pv16_0_ & pv15_0_;
  assign new_n1153 = pv16_0_ & pv15_0_;
  assign pv1757_0_ = new_n1152 | new_n1153;
  assign new_n1155 = pv257_6_ & new_n637;
  assign new_n1156 = pv229_5_ & new_n641;
  assign new_n1157 = pv189_5_ & new_n643;
  assign new_n1158 = ~new_n1156 & ~new_n1157;
  assign new_n1159 = new_n647 & ~new_n1158;
  assign new_n1160 = ~new_n1155 & ~new_n1159;
  assign new_n1161 = ~new_n624 & ~new_n1160;
  assign new_n1162 = pv32_1_ & new_n653;
  assign new_n1163 = pv32_4_ & ~new_n653;
  assign new_n1164 = ~new_n1162 & ~new_n1163;
  assign new_n1165 = new_n624 & ~new_n1164;
  assign new_n1166 = ~new_n1161 & ~new_n1165;
  assign new_n1167 = new_n658 & ~new_n1166;
  assign new_n1168 = pv32_11_ & new_n660;
  assign pv1213_11_ = new_n1167 | new_n1168;
  assign new_n1170 = ~new_n572 & ~pv1213_11_;
  assign new_n1171 = ~pv78_3_ & new_n572;
  assign pv1781_1_ = new_n1170 | new_n1171;
  assign new_n1173 = pv234_2_ & new_n641;
  assign new_n1174 = pv194_2_ & new_n643;
  assign new_n1175 = ~new_n1173 & ~new_n1174;
  assign new_n1176 = new_n647 & ~new_n1175;
  assign new_n1177 = pv149_6_ & new_n665;
  assign new_n1178 = new_n633 & new_n1177;
  assign new_n1179 = ~new_n1176 & ~new_n1178;
  assign new_n1180 = ~new_n624 & ~new_n1179;
  assign new_n1181 = pv32_4_ & new_n653;
  assign new_n1182 = pv32_7_ & ~new_n653;
  assign new_n1183 = ~new_n1181 & ~new_n1182;
  assign new_n1184 = new_n624 & ~new_n1183;
  assign new_n1185 = ~new_n1180 & ~new_n1184;
  assign new_n1186 = new_n658 & ~new_n1185;
  assign new_n1187 = pv84_0_ & new_n660;
  assign pv1243_2_ = new_n1186 | new_n1187;
  assign new_n1189 = pv37_0_ & ~pv1243_2_;
  assign new_n1190 = ~pv37_0_ & ~pv1213_5_;
  assign pv1829_2_ = new_n1189 | new_n1190;
  assign new_n1192 = pv109_0_ & ~pv13_0_;
  assign new_n1193 = pv1_0_ & ~new_n1192;
  assign pv1431 = pv9_0_ & new_n1193;
  assign pv787 = pv7_0_ & pv9_0_;
  assign pv1423 = pv1_0_ & pv9_0_;
  assign pv1258 = pv2_0_ & pv9_0_;
  assign pv1263 = pv4_0_ & pv9_0_;
  assign pv1387 = pv8_0_ & pv9_0_;
  assign pv1259 = pv3_0_ & pv9_0_;
  assign pv780 = pv6_0_ & pv9_0_;
  assign new_n1202 = ~pv1431 & ~pv787;
  assign new_n1203 = ~pv1423 & new_n1202;
  assign new_n1204 = ~pv1423 & ~pv1258;
  assign new_n1205 = ~pv789 & new_n1204;
  assign new_n1206 = new_n1203 & new_n1205;
  assign new_n1207 = ~pv778 & ~pv780;
  assign new_n1208 = ~pv1263 & ~pv1387;
  assign new_n1209 = ~pv1259 & new_n1208;
  assign new_n1210 = new_n1207 & new_n1209;
  assign pv375_0_ = ~new_n1206 | ~new_n1210;
  assign new_n1212 = pv62_0_ & new_n555;
  assign new_n1213 = ~new_n545 & ~new_n554;
  assign new_n1214 = new_n505 & ~new_n785;
  assign new_n1215 = ~new_n1213 & new_n1214;
  assign new_n1216 = pv59_0_ & ~new_n1215;
  assign new_n1217 = ~new_n775 & ~new_n1212;
  assign new_n1218 = ~new_n1216 & new_n1217;
  assign new_n1219 = ~new_n699 & ~pv1757_0_;
  assign pv410_0_ = new_n1218 | ~new_n1219;
  assign new_n1221 = pv59_0_ & new_n557;
  assign new_n1222 = pv62_0_ & new_n1132;
  assign new_n1223 = ~pv149_6_ & new_n1131;
  assign new_n1224 = pv149_6_ & new_n1094;
  assign new_n1225 = ~new_n572 & ~new_n1223;
  assign new_n1226 = ~new_n1224 & new_n1225;
  assign new_n1227 = pv56_0_ & ~new_n1226;
  assign new_n1228 = ~new_n491 & new_n693;
  assign new_n1229 = pv802_0_ & ~new_n1228;
  assign new_n1230 = ~new_n1227 & ~new_n1229;
  assign new_n1231 = ~pv84_2_ & pv84_3_;
  assign new_n1232 = pv84_2_ & ~pv84_3_;
  assign new_n1233 = ~new_n1231 & ~new_n1232;
  assign new_n1234 = ~pv84_4_ & pv84_5_;
  assign new_n1235 = pv84_4_ & ~pv84_5_;
  assign new_n1236 = ~new_n1234 & ~new_n1235;
  assign new_n1237 = new_n1233 & ~new_n1236;
  assign new_n1238 = ~new_n1233 & new_n1236;
  assign new_n1239 = ~new_n1237 & ~new_n1238;
  assign new_n1240 = ~pv88_0_ & pv88_1_;
  assign new_n1241 = pv88_0_ & ~pv88_1_;
  assign new_n1242 = ~new_n1240 & ~new_n1241;
  assign new_n1243 = ~new_n520 & ~new_n534;
  assign new_n1244 = new_n1242 & ~new_n1243;
  assign new_n1245 = ~new_n1242 & new_n1243;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = new_n1239 & ~new_n1246;
  assign new_n1248 = ~new_n1239 & new_n1246;
  assign new_n1249 = ~new_n1247 & ~new_n1248;
  assign new_n1250 = pv94_1_ & new_n1249;
  assign new_n1251 = ~pv94_1_ & ~new_n1249;
  assign new_n1252 = ~new_n1250 & ~new_n1251;
  assign new_n1253 = pv78_1_ & ~pv78_0_;
  assign new_n1254 = ~pv78_1_ & pv78_0_;
  assign new_n1255 = ~new_n1253 & ~new_n1254;
  assign new_n1256 = pv78_3_ & ~pv78_2_;
  assign new_n1257 = ~pv78_3_ & pv78_2_;
  assign new_n1258 = ~new_n1256 & ~new_n1257;
  assign new_n1259 = new_n1255 & ~new_n1258;
  assign new_n1260 = ~new_n1255 & new_n1258;
  assign new_n1261 = ~new_n1259 & ~new_n1260;
  assign new_n1262 = pv78_5_ & ~pv78_4_;
  assign new_n1263 = ~pv78_5_ & pv78_4_;
  assign new_n1264 = ~new_n1262 & ~new_n1263;
  assign new_n1265 = ~pv84_0_ & pv84_1_;
  assign new_n1266 = pv84_0_ & ~pv84_1_;
  assign new_n1267 = ~new_n1265 & ~new_n1266;
  assign new_n1268 = new_n1264 & ~new_n1267;
  assign new_n1269 = ~new_n1264 & new_n1267;
  assign new_n1270 = ~new_n1268 & ~new_n1269;
  assign new_n1271 = new_n1261 & ~new_n1270;
  assign new_n1272 = ~new_n1261 & new_n1270;
  assign new_n1273 = ~new_n1271 & ~new_n1272;
  assign new_n1274 = pv94_0_ & new_n1273;
  assign new_n1275 = ~pv94_0_ & ~new_n1273;
  assign new_n1276 = ~new_n1274 & ~new_n1275;
  assign new_n1277 = ~new_n1252 & ~new_n1276;
  assign new_n1278 = ~new_n1230 & ~new_n1277;
  assign new_n1279 = new_n1223 & ~new_n1278;
  assign new_n1280 = new_n546 & ~new_n554;
  assign new_n1281 = ~new_n491 & ~new_n1279;
  assign new_n1282 = ~new_n494 & new_n1281;
  assign new_n1283 = ~new_n575 & ~new_n1280;
  assign new_n1284 = new_n1282 & new_n1283;
  assign new_n1285 = pv56_0_ & ~new_n1284;
  assign new_n1286 = pv56_0_ & ~new_n1134;
  assign new_n1287 = ~new_n1221 & ~new_n1222;
  assign new_n1288 = ~new_n1285 & ~new_n1286;
  assign pv508_0_ = ~new_n1287 | ~new_n1288;
  assign pv539 = new_n491 & pv1213_2_;
  assign new_n1291 = pv257_1_ & new_n637;
  assign new_n1292 = pv229_0_ & new_n641;
  assign new_n1293 = pv189_0_ & new_n643;
  assign new_n1294 = ~new_n1292 & ~new_n1293;
  assign new_n1295 = new_n647 & ~new_n1294;
  assign new_n1296 = ~new_n1291 & ~new_n1295;
  assign new_n1297 = ~new_n624 & ~new_n1296;
  assign new_n1298 = new_n624 & new_n653;
  assign new_n1299 = ~new_n1297 & ~new_n1298;
  assign new_n1300 = new_n658 & ~new_n1299;
  assign new_n1301 = pv32_6_ & new_n660;
  assign pv1213_6_ = new_n1300 | new_n1301;
  assign new_n1303 = pv268_5_ & new_n686;
  assign new_n1304 = pv268_2_ & ~new_n1303;
  assign new_n1305 = ~pv268_2_ & new_n1303;
  assign pv1372 = new_n1304 | new_n1305;
  assign pv1440_0_ = ~pv14_0_ | new_n507;
  assign new_n1308 = pv16_0_ & ~pv15_0_;
  assign pv1758_0_ = new_n1152 | new_n1308;
  assign new_n1310 = pv257_5_ & new_n637;
  assign new_n1311 = pv229_4_ & new_n641;
  assign new_n1312 = pv189_4_ & new_n643;
  assign new_n1313 = ~new_n1311 & ~new_n1312;
  assign new_n1314 = new_n647 & ~new_n1313;
  assign new_n1315 = ~new_n1310 & ~new_n1314;
  assign new_n1316 = ~new_n624 & ~new_n1315;
  assign new_n1317 = pv32_0_ & new_n653;
  assign new_n1318 = pv32_3_ & ~new_n653;
  assign new_n1319 = ~new_n1317 & ~new_n1318;
  assign new_n1320 = new_n624 & ~new_n1319;
  assign new_n1321 = ~new_n1316 & ~new_n1320;
  assign new_n1322 = new_n658 & ~new_n1321;
  assign new_n1323 = pv32_10_ & new_n660;
  assign pv1213_10_ = new_n1322 | new_n1323;
  assign new_n1325 = ~new_n572 & ~pv1213_10_;
  assign new_n1326 = ~pv78_2_ & new_n572;
  assign pv1781_0_ = new_n1325 | new_n1326;
  assign new_n1328 = pv234_1_ & new_n641;
  assign new_n1329 = pv194_1_ & new_n643;
  assign new_n1330 = ~new_n1328 & ~new_n1329;
  assign new_n1331 = new_n647 & ~new_n1330;
  assign new_n1332 = pv149_5_ & new_n665;
  assign new_n1333 = new_n633 & new_n1332;
  assign new_n1334 = ~new_n1331 & ~new_n1333;
  assign new_n1335 = ~new_n624 & ~new_n1334;
  assign new_n1336 = pv32_3_ & new_n653;
  assign new_n1337 = pv32_6_ & ~new_n653;
  assign new_n1338 = ~new_n1336 & ~new_n1337;
  assign new_n1339 = new_n624 & ~new_n1338;
  assign new_n1340 = ~new_n1335 & ~new_n1339;
  assign new_n1341 = new_n658 & ~new_n1340;
  assign new_n1342 = pv78_5_ & new_n660;
  assign pv1243_1_ = new_n1341 | new_n1342;
  assign new_n1344 = pv37_0_ & ~pv1243_1_;
  assign new_n1345 = pv223_4_ & new_n641;
  assign new_n1346 = pv183_4_ & new_n643;
  assign new_n1347 = ~new_n1345 & ~new_n1346;
  assign new_n1348 = new_n647 & ~new_n1347;
  assign new_n1349 = ~new_n1155 & ~new_n1348;
  assign new_n1350 = new_n658 & ~new_n1349;
  assign new_n1351 = ~new_n624 & new_n1350;
  assign new_n1352 = ~new_n624 & new_n1351;
  assign new_n1353 = pv32_4_ & new_n660;
  assign pv1213_4_ = new_n1352 | new_n1353;
  assign new_n1355 = ~pv37_0_ & ~pv1213_4_;
  assign pv1829_1_ = new_n1344 | new_n1355;
  assign new_n1357 = pv257_2_ & new_n637;
  assign new_n1358 = pv229_1_ & new_n641;
  assign new_n1359 = pv189_1_ & new_n643;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = new_n647 & ~new_n1360;
  assign new_n1362 = ~new_n1357 & ~new_n1361;
  assign new_n1363 = ~new_n624 & ~new_n1362;
  assign new_n1364 = pv32_0_ & ~new_n653;
  assign new_n1365 = ~new_n653 & ~new_n1364;
  assign new_n1366 = new_n624 & ~new_n1365;
  assign new_n1367 = ~new_n1363 & ~new_n1366;
  assign new_n1368 = new_n658 & ~new_n1367;
  assign new_n1369 = pv32_7_ & new_n660;
  assign pv1213_7_ = new_n1368 | new_n1369;
  assign new_n1371 = new_n507 & ~pv802_0_;
  assign new_n1372 = pv248_0_ & ~pv802_0_;
  assign new_n1373 = pv194_3_ & pv194_1_;
  assign new_n1374 = pv199_2_ & new_n1373;
  assign new_n1375 = pv199_0_ & new_n1374;
  assign new_n1376 = pv199_4_ & new_n1375;
  assign new_n1377 = pv199_1_ & new_n1376;
  assign new_n1378 = pv199_3_ & new_n1377;
  assign new_n1379 = pv194_2_ & new_n1378;
  assign new_n1380 = pv194_4_ & new_n1379;
  assign new_n1381 = pv194_0_ & new_n1380;
  assign new_n1382 = ~pv802_0_ & new_n1381;
  assign new_n1383 = ~new_n1371 & ~new_n1372;
  assign new_n1384 = ~new_n1382 & new_n1383;
  assign new_n1385 = ~new_n639 & new_n1384;
  assign new_n1386 = ~new_n740 & new_n1385;
  assign new_n1387 = ~pv274_0_ & pv271_0_;
  assign new_n1388 = ~new_n572 & new_n1387;
  assign new_n1389 = pv134_1_ & pv134_0_;
  assign new_n1390 = new_n1388 & new_n1389;
  assign new_n1391 = new_n507 & new_n1390;
  assign new_n1392 = ~new_n1381 & new_n1391;
  assign new_n1393 = new_n573 & ~pv802_0_;
  assign new_n1394 = ~new_n1372 & new_n1393;
  assign new_n1395 = ~new_n507 & new_n1394;
  assign new_n1396 = ~new_n740 & new_n1395;
  assign new_n1397 = ~new_n1381 & new_n1396;
  assign new_n1398 = ~new_n1386 & ~new_n1392;
  assign new_n1399 = ~new_n1397 & new_n1398;
  assign new_n1400 = pv7_0_ & ~new_n1399;
  assign pv1380 = new_n692 & new_n1400;
  assign new_n1402 = new_n510 & new_n1308;
  assign new_n1403 = new_n490 & new_n1308;
  assign new_n1404 = pv56_0_ & new_n1093;
  assign new_n1405 = pv14_0_ & ~new_n1404;
  assign new_n1406 = pv101_0_ & new_n1405;
  assign new_n1407 = ~new_n1402 & ~new_n1403;
  assign pv1759_0_ = new_n1406 | ~new_n1407;
  assign new_n1409 = pv234_4_ & new_n641;
  assign new_n1410 = pv194_4_ & new_n643;
  assign new_n1411 = ~new_n1409 & ~new_n1410;
  assign new_n1412 = ~new_n624 & ~new_n635;
  assign new_n1413 = ~new_n1411 & new_n1412;
  assign new_n1414 = new_n616 & new_n1413;
  assign new_n1415 = ~new_n633 & new_n1414;
  assign new_n1416 = ~new_n624 & new_n1415;
  assign new_n1417 = pv32_6_ & new_n653;
  assign new_n1418 = pv32_9_ & ~new_n653;
  assign new_n1419 = ~new_n1417 & ~new_n1418;
  assign new_n1420 = new_n624 & ~new_n1419;
  assign new_n1421 = ~new_n1416 & ~new_n1420;
  assign new_n1422 = new_n658 & ~new_n1421;
  assign new_n1423 = pv84_2_ & new_n660;
  assign pv1243_4_ = new_n1422 | new_n1423;
  assign new_n1425 = pv37_0_ & ~pv1243_4_;
  assign new_n1426 = ~pv37_0_ & ~pv1213_7_;
  assign pv1829_4_ = new_n1425 | new_n1426;
  assign new_n1428 = pv257_6_ & ~pv257_7_;
  assign new_n1429 = ~pv257_6_ & pv257_7_;
  assign pv656 = new_n1428 | new_n1429;
  assign pv779 = pv6_0_ & new_n692;
  assign new_n1432 = pv257_3_ & new_n637;
  assign new_n1433 = pv229_2_ & new_n641;
  assign new_n1434 = pv189_2_ & new_n643;
  assign new_n1435 = ~new_n1433 & ~new_n1434;
  assign new_n1436 = new_n647 & ~new_n1435;
  assign new_n1437 = ~new_n1432 & ~new_n1436;
  assign new_n1438 = ~new_n624 & ~new_n1437;
  assign new_n1439 = pv32_1_ & ~new_n653;
  assign new_n1440 = ~new_n653 & ~new_n1439;
  assign new_n1441 = new_n624 & ~new_n1440;
  assign new_n1442 = ~new_n1438 & ~new_n1441;
  assign new_n1443 = new_n658 & ~new_n1442;
  assign new_n1444 = pv32_8_ & new_n660;
  assign pv1213_8_ = new_n1443 | new_n1444;
  assign pv1262 = pv4_0_ & new_n692;
  assign new_n1447 = pv268_4_ & pv268_2_;
  assign new_n1448 = pv268_3_ & new_n1447;
  assign new_n1449 = pv268_1_ & new_n1448;
  assign new_n1450 = pv268_5_ & new_n1449;
  assign new_n1451 = pv268_0_ & ~new_n1450;
  assign new_n1452 = ~pv268_0_ & new_n1450;
  assign pv1370 = new_n1451 | new_n1452;
  assign new_n1454 = pv234_3_ & new_n641;
  assign new_n1455 = pv194_3_ & new_n643;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = new_n647 & ~new_n1456;
  assign new_n1458 = pv149_7_ & new_n665;
  assign new_n1459 = new_n633 & new_n1458;
  assign new_n1460 = ~new_n1457 & ~new_n1459;
  assign new_n1461 = ~new_n624 & ~new_n1460;
  assign new_n1462 = pv32_5_ & new_n653;
  assign new_n1463 = pv32_8_ & ~new_n653;
  assign new_n1464 = ~new_n1462 & ~new_n1463;
  assign new_n1465 = new_n624 & ~new_n1464;
  assign new_n1466 = ~new_n1461 & ~new_n1465;
  assign new_n1467 = new_n658 & ~new_n1466;
  assign new_n1468 = pv84_1_ & new_n660;
  assign pv1243_3_ = new_n1467 | new_n1468;
  assign new_n1470 = pv37_0_ & ~pv1243_3_;
  assign new_n1471 = ~pv37_0_ & ~pv1213_6_;
  assign pv1829_3_ = new_n1470 | new_n1471;
  assign new_n1473 = pv257_4_ & new_n637;
  assign new_n1474 = pv229_3_ & new_n641;
  assign new_n1475 = pv189_3_ & new_n643;
  assign new_n1476 = ~new_n1474 & ~new_n1475;
  assign new_n1477 = new_n647 & ~new_n1476;
  assign new_n1478 = ~new_n1473 & ~new_n1477;
  assign new_n1479 = ~new_n624 & ~new_n1478;
  assign new_n1480 = pv32_2_ & ~new_n653;
  assign new_n1481 = ~new_n653 & ~new_n1480;
  assign new_n1482 = new_n624 & ~new_n1481;
  assign new_n1483 = ~new_n1479 & ~new_n1482;
  assign new_n1484 = new_n658 & ~new_n1483;
  assign new_n1485 = pv32_9_ & new_n660;
  assign pv1213_9_ = new_n1484 | new_n1485;
  assign pv1264 = pv4_0_ & pv12_0_;
  assign pv1265 = pv52_0_ & pv1264;
  assign new_n1489 = ~pv56_0_ & ~pv50_0_;
  assign new_n1490 = ~pv62_0_ & new_n1489;
  assign new_n1491 = ~new_n616 & ~new_n1490;
  assign pv1386 = pv782 & new_n1491;
  assign new_n1493 = ~pv280_0_ & new_n494;
  assign new_n1494 = pv165_2_ & pv165_1_;
  assign new_n1495 = ~pv165_0_ & new_n1494;
  assign new_n1496 = pv203_0_ & new_n1495;
  assign new_n1497 = pv240_0_ & ~new_n1493;
  assign new_n1498 = ~new_n1496 & new_n1497;
  assign new_n1499 = new_n758 & new_n1498;
  assign new_n1500 = ~new_n699 & new_n1499;
  assign new_n1501 = ~pv172_0_ & new_n1500;
  assign new_n1502 = ~new_n507 & ~new_n640;
  assign new_n1503 = ~new_n494 & ~new_n1502;
  assign new_n1504 = pv802_0_ & ~new_n1503;
  assign pv1717_0_ = new_n1501 | new_n1504;
  assign new_n1506 = pv239_1_ & new_n641;
  assign new_n1507 = pv199_1_ & new_n643;
  assign new_n1508 = ~new_n1506 & ~new_n1507;
  assign new_n1509 = new_n1412 & ~new_n1508;
  assign new_n1510 = new_n616 & new_n1509;
  assign new_n1511 = ~new_n633 & new_n1510;
  assign new_n1512 = ~new_n624 & new_n1511;
  assign new_n1513 = pv32_8_ & new_n653;
  assign new_n1514 = pv32_11_ & ~new_n653;
  assign new_n1515 = ~new_n1513 & ~new_n1514;
  assign new_n1516 = new_n624 & ~new_n1515;
  assign new_n1517 = ~new_n1512 & ~new_n1516;
  assign new_n1518 = new_n658 & ~new_n1517;
  assign new_n1519 = pv84_4_ & new_n660;
  assign pv1243_6_ = new_n1518 | new_n1519;
  assign new_n1521 = pv37_0_ & ~pv1243_6_;
  assign new_n1522 = ~pv37_0_ & ~pv1213_9_;
  assign pv1829_6_ = new_n1521 | new_n1522;
  assign new_n1524 = ~pv202_0_ & ~pv271_0_;
  assign new_n1525 = pv274_0_ & new_n1524;
  assign new_n1526 = pv274_0_ & ~new_n1525;
  assign new_n1527 = ~pv271_0_ & new_n1526;
  assign new_n1528 = pv269_0_ & ~new_n1525;
  assign new_n1529 = pv271_0_ & new_n1528;
  assign pv634_0_ = ~new_n1527 & ~new_n1529;
  assign new_n1531 = new_n493 & pv1757_0_;
  assign new_n1532 = pv802_0_ & new_n1531;
  assign new_n1533 = ~new_n493 & pv1757_0_;
  assign new_n1534 = ~new_n1278 & ~new_n1532;
  assign pv1480_0_ = new_n1533 | ~new_n1534;
  assign new_n1536 = ~new_n699 & new_n707;
  assign new_n1537 = ~new_n699 & new_n717;
  assign new_n1538 = pv290_0_ & new_n699;
  assign new_n1539 = ~new_n699 & new_n722;
  assign new_n1540 = ~new_n725 & ~new_n1536;
  assign new_n1541 = ~new_n1537 & new_n1540;
  assign new_n1542 = ~new_n1538 & ~new_n1539;
  assign pv1741_0_ = ~new_n1541 | ~new_n1542;
  assign new_n1544 = pv239_0_ & new_n641;
  assign new_n1545 = pv199_0_ & new_n643;
  assign new_n1546 = ~new_n1544 & ~new_n1545;
  assign new_n1547 = new_n1412 & ~new_n1546;
  assign new_n1548 = new_n616 & new_n1547;
  assign new_n1549 = ~new_n633 & new_n1548;
  assign new_n1550 = ~new_n624 & new_n1549;
  assign new_n1551 = pv32_7_ & new_n653;
  assign new_n1552 = pv32_10_ & ~new_n653;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = new_n624 & ~new_n1553;
  assign new_n1555 = ~new_n1550 & ~new_n1554;
  assign new_n1556 = new_n658 & ~new_n1555;
  assign new_n1557 = pv84_3_ & new_n660;
  assign pv1243_5_ = new_n1556 | new_n1557;
  assign new_n1559 = pv37_0_ & ~pv1243_5_;
  assign new_n1560 = ~pv37_0_ & ~pv1213_8_;
  assign pv1829_5_ = new_n1559 | new_n1560;
  assign new_n1562 = pv39_0_ & ~pv38_0_;
  assign new_n1563 = ~pv39_0_ & pv38_0_;
  assign new_n1564 = ~new_n1562 & ~new_n1563;
  assign new_n1565 = pv42_0_ & ~pv44_0_;
  assign new_n1566 = ~pv42_0_ & pv44_0_;
  assign new_n1567 = ~new_n1565 & ~new_n1566;
  assign pv512 = new_n1564 & new_n1567;
  assign pv783 = pv5_0_ & pv11_0_;
  assign pv1256 = pv2_0_ & new_n692;
  assign pv1267 = pv2_0_ & pv11_0_;
  assign new_n1572 = ~pv302_0_ & new_n493;
  assign new_n1573 = new_n511 & new_n554;
  assign new_n1574 = ~new_n1572 & ~new_n1573;
  assign new_n1575 = ~new_n712 & ~new_n713;
  assign new_n1576 = new_n1574 & new_n1575;
  assign new_n1577 = ~new_n699 & new_n704;
  assign new_n1578 = ~pv289_0_ & new_n1577;
  assign new_n1579 = ~new_n1576 & new_n1578;
  assign new_n1580 = pv14_0_ & new_n1579;
  assign new_n1581 = ~new_n585 & ~new_n1580;
  assign new_n1582 = ~new_n699 & new_n1581;
  assign new_n1583 = new_n704 & new_n1582;
  assign new_n1584 = new_n490 & new_n1583;
  assign new_n1585 = pv290_0_ & new_n490;
  assign new_n1586 = new_n699 & new_n1585;
  assign new_n1587 = ~new_n1584 & ~new_n1586;
  assign new_n1588 = ~pv149_6_ & new_n761;
  assign new_n1589 = pv56_0_ & new_n1588;
  assign new_n1590 = pv14_0_ & new_n1587;
  assign new_n1591 = pv213_0_ & new_n1590;
  assign new_n1592 = ~new_n1589 & new_n1591;
  assign new_n1593 = ~pv165_3_ & new_n577;
  assign new_n1594 = ~pv165_7_ & new_n1593;
  assign new_n1595 = ~new_n704 & ~new_n1594;
  assign new_n1596 = ~new_n1587 & ~new_n1595;
  assign pv1281_0_ = new_n1592 | new_n1596;
  assign new_n1598 = pv268_4_ & pv268_5_;
  assign new_n1599 = pv268_3_ & ~new_n1598;
  assign new_n1600 = ~pv268_3_ & new_n1598;
  assign pv1373 = new_n1599 | new_n1600;
  assign new_n1602 = pv56_0_ & ~new_n1278;
  assign new_n1603 = new_n1224 & new_n1602;
  assign new_n1604 = ~new_n699 & new_n1603;
  assign pv1384 = pv782 & new_n1604;
  assign new_n1606 = pv239_3_ & new_n641;
  assign new_n1607 = pv199_3_ & new_n643;
  assign new_n1608 = ~new_n1606 & ~new_n1607;
  assign new_n1609 = new_n1412 & ~new_n1608;
  assign new_n1610 = new_n616 & new_n1609;
  assign new_n1611 = ~new_n633 & new_n1610;
  assign new_n1612 = ~new_n624 & new_n1611;
  assign new_n1613 = pv32_10_ & new_n624;
  assign new_n1614 = new_n624 & new_n1613;
  assign new_n1615 = new_n653 & new_n1614;
  assign new_n1616 = ~new_n1612 & ~new_n1615;
  assign new_n1617 = new_n658 & ~new_n1616;
  assign new_n1618 = pv88_0_ & new_n660;
  assign pv1243_8_ = new_n1617 | new_n1618;
  assign new_n1620 = pv37_0_ & ~pv1243_8_;
  assign new_n1621 = ~pv37_0_ & ~pv1213_11_;
  assign pv1829_8_ = new_n1620 | new_n1621;
  assign new_n1623 = pv132_0_ & new_n1098;
  assign new_n1624 = new_n1093 & ~new_n1095;
  assign new_n1625 = ~new_n1096 & new_n1624;
  assign new_n1626 = pv108_5_ & new_n1625;
  assign pv1953_0_ = new_n1623 | new_n1626;
  assign new_n1628 = pv14_0_ & new_n758;
  assign new_n1629 = ~new_n615 & new_n1628;
  assign new_n1630 = pv763 & new_n1629;
  assign pv775 = pv70_0_ & new_n1630;
  assign pv784 = pv7_0_ & pv11_0_;
  assign new_n1633 = ~pv57_0_ & new_n1223;
  assign new_n1634 = ~new_n494 & new_n545;
  assign new_n1635 = new_n505 & new_n1634;
  assign new_n1636 = ~new_n491 & ~new_n546;
  assign new_n1637 = new_n772 & new_n1636;
  assign new_n1638 = new_n1635 & new_n1637;
  assign new_n1639 = pv57_0_ & ~new_n1638;
  assign new_n1640 = ~pv60_0_ & ~pv63_0_;
  assign new_n1641 = new_n572 & ~new_n1640;
  assign new_n1642 = ~new_n1633 & ~new_n1639;
  assign new_n1643 = pv12_0_ & new_n1642;
  assign new_n1644 = ~pv174_0_ & new_n1643;
  assign new_n1645 = pv2_0_ & new_n1644;
  assign new_n1646 = ~new_n1641 & new_n1645;
  assign pv1257 = ~pv35_0_ & new_n1646;
  assign pv1266 = pv4_0_ & pv11_0_;
  assign new_n1649 = ~new_n712 & ~new_n785;
  assign new_n1650 = new_n758 & new_n1649;
  assign new_n1651 = ~new_n1223 & new_n1650;
  assign new_n1652 = pv14_0_ & new_n1651;
  assign new_n1653 = pv62_0_ & new_n1652;
  assign new_n1654 = new_n505 & new_n1653;
  assign new_n1655 = ~new_n1133 & new_n1654;
  assign new_n1656 = new_n616 & new_n1655;
  assign pv1365 = ~new_n1213 & new_n1656;
  assign new_n1658 = pv268_4_ & ~pv268_5_;
  assign new_n1659 = ~pv268_4_ & pv268_5_;
  assign pv1374 = new_n1658 | new_n1659;
  assign new_n1661 = ~pv258_0_ & new_n1491;
  assign new_n1662 = pv268_0_ & new_n1450;
  assign new_n1663 = pv258_0_ & new_n1662;
  assign new_n1664 = ~new_n1661 & ~new_n1663;
  assign new_n1665 = pv14_0_ & new_n1664;
  assign new_n1666 = pv259_0_ & new_n1665;
  assign new_n1667 = pv14_0_ & ~new_n1664;
  assign new_n1668 = ~pv259_0_ & new_n1667;
  assign pv1459_0_ = new_n1666 | new_n1668;
  assign new_n1670 = pv239_2_ & new_n641;
  assign new_n1671 = pv199_2_ & new_n643;
  assign new_n1672 = ~new_n1670 & ~new_n1671;
  assign new_n1673 = new_n1412 & ~new_n1672;
  assign new_n1674 = new_n616 & new_n1673;
  assign new_n1675 = ~new_n633 & new_n1674;
  assign new_n1676 = ~new_n624 & new_n1675;
  assign new_n1677 = pv32_9_ & new_n624;
  assign new_n1678 = new_n624 & new_n1677;
  assign new_n1679 = new_n653 & new_n1678;
  assign new_n1680 = ~new_n1676 & ~new_n1679;
  assign new_n1681 = new_n658 & ~new_n1680;
  assign new_n1682 = pv84_5_ & new_n660;
  assign pv1243_7_ = new_n1681 | new_n1682;
  assign new_n1684 = pv37_0_ & ~pv1243_7_;
  assign new_n1685 = ~pv37_0_ & ~pv1213_10_;
  assign pv1829_7_ = new_n1684 | new_n1685;
  assign pv1953_1_ = pv132_1_ & new_n1098;
  assign pv543 = new_n491 & pv1213_6_;
  assign new_n1689 = pv802_0_ & ~new_n640;
  assign pv587 = ~pv243_0_ & ~new_n1689;
  assign new_n1691 = pv257_2_ & pv257_4_;
  assign new_n1692 = pv257_5_ & new_n1691;
  assign new_n1693 = pv257_3_ & new_n1692;
  assign new_n1694 = pv257_7_ & new_n1693;
  assign new_n1695 = pv257_6_ & new_n1694;
  assign new_n1696 = pv257_1_ & ~new_n1695;
  assign new_n1697 = ~pv257_1_ & new_n1695;
  assign pv651 = new_n1696 | new_n1697;
  assign new_n1699 = pv56_0_ & ~new_n586;
  assign new_n1700 = ~pv174_0_ & new_n1699;
  assign new_n1701 = ~pv52_0_ & ~new_n1700;
  assign new_n1702 = pv6_0_ & pv12_0_;
  assign pv781 = ~new_n1701 & new_n1702;
  assign new_n1704 = pv14_0_ & ~new_n1586;
  assign new_n1705 = pv213_2_ & new_n1704;
  assign new_n1706 = ~new_n1589 & new_n1705;
  assign new_n1707 = pv165_4_ & new_n1586;
  assign pv1297_1_ = new_n1706 | new_n1707;
  assign new_n1709 = ~pv88_2_ & new_n572;
  assign new_n1710 = ~pv134_0_ & ~new_n572;
  assign pv1771_0_ = new_n1709 | new_n1710;
  assign new_n1712 = pv149_7_ & new_n839;
  assign new_n1713 = ~pv149_6_ & new_n1712;
  assign new_n1714 = pv56_0_ & new_n1713;
  assign new_n1715 = pv108_4_ & ~new_n1714;
  assign pv1900_0_ = new_n1152 | new_n1715;
  assign new_n1717 = ~pv149_7_ & new_n760;
  assign new_n1718 = pv149_6_ & new_n1717;
  assign new_n1719 = ~new_n1095 & ~new_n1713;
  assign new_n1720 = new_n1718 & new_n1719;
  assign new_n1721 = ~new_n1588 & new_n1720;
  assign new_n1722 = pv100_1_ & new_n1721;
  assign new_n1723 = new_n1095 & ~new_n1713;
  assign new_n1724 = ~new_n1718 & new_n1723;
  assign new_n1725 = ~new_n1588 & new_n1724;
  assign new_n1726 = pv124_1_ & new_n1725;
  assign new_n1727 = ~new_n1718 & new_n1719;
  assign new_n1728 = new_n1588 & new_n1727;
  assign new_n1729 = pv213_1_ & new_n1728;
  assign new_n1730 = ~new_n1095 & new_n1713;
  assign new_n1731 = ~new_n1718 & new_n1730;
  assign new_n1732 = ~new_n1588 & new_n1731;
  assign new_n1733 = pv108_1_ & new_n1732;
  assign new_n1734 = ~new_n1722 & ~new_n1726;
  assign new_n1735 = ~new_n1729 & ~new_n1733;
  assign pv1921_1_ = ~new_n1734 | ~new_n1735;
  assign new_n1737 = pv239_4_ & new_n641;
  assign new_n1738 = pv199_4_ & new_n643;
  assign new_n1739 = ~new_n1737 & ~new_n1738;
  assign new_n1740 = new_n1412 & ~new_n1739;
  assign new_n1741 = new_n616 & new_n1740;
  assign new_n1742 = ~new_n633 & new_n1741;
  assign new_n1743 = ~new_n624 & new_n1742;
  assign new_n1744 = pv32_11_ & new_n624;
  assign new_n1745 = new_n624 & new_n1744;
  assign new_n1746 = new_n653 & new_n1745;
  assign new_n1747 = ~new_n1743 & ~new_n1746;
  assign new_n1748 = new_n658 & ~new_n1747;
  assign new_n1749 = pv88_1_ & new_n660;
  assign pv1243_9_ = new_n1748 | new_n1749;
  assign new_n1751 = ~pv1213_2_ & ~pv1213_0_;
  assign new_n1752 = ~pv1213_3_ & new_n1751;
  assign new_n1753 = ~pv1213_1_ & new_n1752;
  assign new_n1754 = ~new_n842 & new_n1753;
  assign new_n1755 = ~new_n880 & new_n1754;
  assign new_n1756 = pv1213_3_ & new_n1751;
  assign new_n1757 = ~pv1213_1_ & new_n1756;
  assign new_n1758 = ~new_n842 & new_n1757;
  assign new_n1759 = pv288_6_ & new_n1758;
  assign new_n1760 = ~new_n1755 & ~new_n1759;
  assign new_n1761 = new_n616 & new_n1760;
  assign new_n1762 = new_n616 & new_n1084;
  assign new_n1763 = new_n1761 & new_n1762;
  assign new_n1764 = pv288_6_ & pv288_7_;
  assign new_n1765 = ~new_n1763 & new_n1764;
  assign new_n1766 = new_n957 & ~new_n973;
  assign new_n1767 = new_n959 & ~new_n988;
  assign new_n1768 = ~new_n959 & ~new_n988;
  assign new_n1769 = ~new_n1767 & ~new_n1768;
  assign new_n1770 = new_n959 & ~new_n982;
  assign new_n1771 = new_n988 & ~new_n1015;
  assign new_n1772 = ~new_n988 & new_n1015;
  assign new_n1773 = ~new_n1771 & ~new_n1772;
  assign new_n1774 = ~new_n959 & ~new_n1773;
  assign new_n1775 = ~new_n1770 & ~new_n1774;
  assign new_n1776 = new_n1769 & new_n1775;
  assign new_n1777 = new_n959 & ~new_n997;
  assign new_n1778 = ~new_n1023 & ~new_n1772;
  assign new_n1779 = new_n1023 & new_n1772;
  assign new_n1780 = ~new_n1778 & ~new_n1779;
  assign new_n1781 = ~new_n959 & ~new_n1780;
  assign new_n1782 = ~new_n1777 & ~new_n1781;
  assign new_n1783 = new_n1776 & new_n1782;
  assign new_n1784 = new_n959 & ~new_n973;
  assign new_n1785 = ~new_n1010 & ~new_n1779;
  assign new_n1786 = new_n1010 & new_n1779;
  assign new_n1787 = ~new_n1785 & ~new_n1786;
  assign new_n1788 = ~new_n959 & ~new_n1787;
  assign new_n1789 = ~new_n1784 & ~new_n1788;
  assign new_n1790 = ~new_n1783 & ~new_n1789;
  assign new_n1791 = new_n1783 & new_n1789;
  assign new_n1792 = ~new_n1790 & ~new_n1791;
  assign new_n1793 = ~new_n957 & ~new_n1792;
  assign new_n1794 = ~new_n1766 & ~new_n1793;
  assign new_n1795 = ~pv1213_0_ & ~new_n1794;
  assign new_n1796 = pv1213_0_ & new_n1794;
  assign new_n1797 = ~new_n1795 & ~new_n1796;
  assign new_n1798 = new_n957 & ~new_n982;
  assign new_n1799 = ~new_n1769 & ~new_n1775;
  assign new_n1800 = ~new_n1776 & ~new_n1799;
  assign new_n1801 = ~new_n957 & ~new_n1800;
  assign new_n1802 = ~new_n1798 & ~new_n1801;
  assign new_n1803 = ~pv1213_2_ & ~new_n1802;
  assign new_n1804 = pv1213_2_ & new_n1802;
  assign new_n1805 = ~new_n1803 & ~new_n1804;
  assign new_n1806 = new_n957 & ~new_n988;
  assign new_n1807 = ~new_n957 & new_n1769;
  assign new_n1808 = ~new_n1806 & ~new_n1807;
  assign new_n1809 = ~pv1213_3_ & ~new_n1808;
  assign new_n1810 = pv1213_3_ & new_n1808;
  assign new_n1811 = ~new_n1809 & ~new_n1810;
  assign new_n1812 = new_n957 & ~new_n997;
  assign new_n1813 = ~new_n1776 & ~new_n1782;
  assign new_n1814 = ~new_n1783 & ~new_n1813;
  assign new_n1815 = ~new_n957 & ~new_n1814;
  assign new_n1816 = ~new_n1812 & ~new_n1815;
  assign new_n1817 = ~pv1213_1_ & ~new_n1816;
  assign new_n1818 = pv1213_1_ & new_n1816;
  assign new_n1819 = ~new_n1817 & ~new_n1818;
  assign new_n1820 = ~pv288_0_ & ~pv288_1_;
  assign new_n1821 = new_n1797 & new_n1805;
  assign new_n1822 = new_n1811 & new_n1821;
  assign new_n1823 = new_n1819 & new_n1822;
  assign new_n1824 = ~new_n842 & new_n1823;
  assign new_n1825 = ~new_n1820 & new_n1824;
  assign new_n1826 = ~pv1213_0_ & ~new_n1789;
  assign new_n1827 = pv1213_0_ & new_n1789;
  assign new_n1828 = ~new_n1826 & ~new_n1827;
  assign new_n1829 = ~pv1213_2_ & ~new_n1775;
  assign new_n1830 = pv1213_2_ & new_n1775;
  assign new_n1831 = ~new_n1829 & ~new_n1830;
  assign new_n1832 = ~pv1213_3_ & ~new_n1769;
  assign new_n1833 = pv1213_3_ & new_n1769;
  assign new_n1834 = ~new_n1832 & ~new_n1833;
  assign new_n1835 = ~pv1213_1_ & ~new_n1782;
  assign new_n1836 = pv1213_1_ & new_n1782;
  assign new_n1837 = ~new_n1835 & ~new_n1836;
  assign new_n1838 = new_n1828 & new_n1831;
  assign new_n1839 = new_n1834 & new_n1838;
  assign new_n1840 = new_n1837 & new_n1839;
  assign new_n1841 = ~new_n842 & new_n1840;
  assign new_n1842 = pv288_0_ & new_n1841;
  assign new_n1843 = ~new_n1825 & ~new_n1842;
  assign new_n1844 = new_n616 & new_n1843;
  assign new_n1845 = ~new_n1005 & ~new_n1031;
  assign new_n1846 = new_n616 & new_n1845;
  assign new_n1847 = new_n1844 & new_n1846;
  assign new_n1848 = new_n965 & ~new_n1847;
  assign new_n1849 = new_n860 & ~new_n907;
  assign new_n1850 = new_n862 & ~new_n922;
  assign new_n1851 = ~new_n862 & ~new_n922;
  assign new_n1852 = ~new_n1850 & ~new_n1851;
  assign new_n1853 = new_n862 & ~new_n916;
  assign new_n1854 = new_n922 & ~new_n1067;
  assign new_n1855 = ~new_n922 & new_n1067;
  assign new_n1856 = ~new_n1854 & ~new_n1855;
  assign new_n1857 = ~new_n862 & ~new_n1856;
  assign new_n1858 = ~new_n1853 & ~new_n1857;
  assign new_n1859 = new_n1852 & new_n1858;
  assign new_n1860 = new_n862 & ~new_n931;
  assign new_n1861 = ~new_n1075 & ~new_n1855;
  assign new_n1862 = new_n1075 & new_n1855;
  assign new_n1863 = ~new_n1861 & ~new_n1862;
  assign new_n1864 = ~new_n862 & ~new_n1863;
  assign new_n1865 = ~new_n1860 & ~new_n1864;
  assign new_n1866 = new_n1859 & new_n1865;
  assign new_n1867 = new_n862 & ~new_n907;
  assign new_n1868 = ~new_n1062 & ~new_n1862;
  assign new_n1869 = new_n1062 & new_n1862;
  assign new_n1870 = ~new_n1868 & ~new_n1869;
  assign new_n1871 = ~new_n862 & ~new_n1870;
  assign new_n1872 = ~new_n1867 & ~new_n1871;
  assign new_n1873 = ~new_n1866 & ~new_n1872;
  assign new_n1874 = new_n1866 & new_n1872;
  assign new_n1875 = ~new_n1873 & ~new_n1874;
  assign new_n1876 = ~new_n860 & ~new_n1875;
  assign new_n1877 = ~new_n1849 & ~new_n1876;
  assign new_n1878 = ~pv1213_0_ & ~new_n1877;
  assign new_n1879 = pv1213_0_ & new_n1877;
  assign new_n1880 = ~new_n1878 & ~new_n1879;
  assign new_n1881 = new_n860 & ~new_n916;
  assign new_n1882 = ~new_n1852 & ~new_n1858;
  assign new_n1883 = ~new_n1859 & ~new_n1882;
  assign new_n1884 = ~new_n860 & ~new_n1883;
  assign new_n1885 = ~new_n1881 & ~new_n1884;
  assign new_n1886 = ~pv1213_2_ & ~new_n1885;
  assign new_n1887 = pv1213_2_ & new_n1885;
  assign new_n1888 = ~new_n1886 & ~new_n1887;
  assign new_n1889 = new_n860 & ~new_n922;
  assign new_n1890 = ~new_n860 & new_n1852;
  assign new_n1891 = ~new_n1889 & ~new_n1890;
  assign new_n1892 = ~pv1213_3_ & ~new_n1891;
  assign new_n1893 = pv1213_3_ & new_n1891;
  assign new_n1894 = ~new_n1892 & ~new_n1893;
  assign new_n1895 = new_n860 & ~new_n931;
  assign new_n1896 = ~new_n1859 & ~new_n1865;
  assign new_n1897 = ~new_n1866 & ~new_n1896;
  assign new_n1898 = ~new_n860 & ~new_n1897;
  assign new_n1899 = ~new_n1895 & ~new_n1898;
  assign new_n1900 = ~pv1213_1_ & ~new_n1899;
  assign new_n1901 = pv1213_1_ & new_n1899;
  assign new_n1902 = ~new_n1900 & ~new_n1901;
  assign new_n1903 = ~pv288_2_ & ~pv288_3_;
  assign new_n1904 = new_n1880 & new_n1888;
  assign new_n1905 = new_n1894 & new_n1904;
  assign new_n1906 = new_n1902 & new_n1905;
  assign new_n1907 = ~new_n842 & new_n1906;
  assign new_n1908 = ~new_n1903 & new_n1907;
  assign new_n1909 = ~pv1213_0_ & ~new_n1872;
  assign new_n1910 = pv1213_0_ & new_n1872;
  assign new_n1911 = ~new_n1909 & ~new_n1910;
  assign new_n1912 = ~pv1213_2_ & ~new_n1858;
  assign new_n1913 = pv1213_2_ & new_n1858;
  assign new_n1914 = ~new_n1912 & ~new_n1913;
  assign new_n1915 = ~pv1213_3_ & ~new_n1852;
  assign new_n1916 = pv1213_3_ & new_n1852;
  assign new_n1917 = ~new_n1915 & ~new_n1916;
  assign new_n1918 = ~pv1213_1_ & ~new_n1865;
  assign new_n1919 = pv1213_1_ & new_n1865;
  assign new_n1920 = ~new_n1918 & ~new_n1919;
  assign new_n1921 = new_n1911 & new_n1914;
  assign new_n1922 = new_n1917 & new_n1921;
  assign new_n1923 = new_n1920 & new_n1922;
  assign new_n1924 = ~new_n842 & new_n1923;
  assign new_n1925 = pv288_2_ & new_n1924;
  assign new_n1926 = ~new_n1908 & ~new_n1925;
  assign new_n1927 = new_n616 & new_n1926;
  assign new_n1928 = ~new_n939 & ~new_n1083;
  assign new_n1929 = new_n616 & new_n1928;
  assign new_n1930 = new_n1927 & new_n1929;
  assign new_n1931 = new_n878 & ~new_n1930;
  assign new_n1932 = new_n856 & ~new_n904;
  assign new_n1933 = ~new_n859 & new_n867;
  assign new_n1934 = ~new_n859 & ~new_n867;
  assign new_n1935 = ~new_n1933 & ~new_n1934;
  assign new_n1936 = new_n867 & ~new_n873;
  assign new_n1937 = new_n859 & ~new_n1041;
  assign new_n1938 = ~new_n859 & new_n1041;
  assign new_n1939 = ~new_n1937 & ~new_n1938;
  assign new_n1940 = ~new_n867 & ~new_n1939;
  assign new_n1941 = ~new_n1936 & ~new_n1940;
  assign new_n1942 = new_n1935 & new_n1941;
  assign new_n1943 = new_n867 & ~new_n892;
  assign new_n1944 = ~new_n1049 & ~new_n1938;
  assign new_n1945 = new_n1049 & new_n1938;
  assign new_n1946 = ~new_n1944 & ~new_n1945;
  assign new_n1947 = ~new_n867 & ~new_n1946;
  assign new_n1948 = ~new_n1943 & ~new_n1947;
  assign new_n1949 = new_n1942 & new_n1948;
  assign new_n1950 = new_n867 & ~new_n904;
  assign new_n1951 = ~new_n1036 & ~new_n1945;
  assign new_n1952 = new_n1036 & new_n1945;
  assign new_n1953 = ~new_n1951 & ~new_n1952;
  assign new_n1954 = ~new_n867 & ~new_n1953;
  assign new_n1955 = ~new_n1950 & ~new_n1954;
  assign new_n1956 = ~new_n1949 & ~new_n1955;
  assign new_n1957 = new_n1949 & new_n1955;
  assign new_n1958 = ~new_n1956 & ~new_n1957;
  assign new_n1959 = ~new_n856 & ~new_n1958;
  assign new_n1960 = ~new_n1932 & ~new_n1959;
  assign new_n1961 = ~pv1213_0_ & ~new_n1960;
  assign new_n1962 = pv1213_0_ & new_n1960;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = new_n856 & ~new_n873;
  assign new_n1965 = ~new_n1935 & ~new_n1941;
  assign new_n1966 = ~new_n1942 & ~new_n1965;
  assign new_n1967 = ~new_n856 & ~new_n1966;
  assign new_n1968 = ~new_n1964 & ~new_n1967;
  assign new_n1969 = ~pv1213_2_ & ~new_n1968;
  assign new_n1970 = pv1213_2_ & new_n1968;
  assign new_n1971 = ~new_n1969 & ~new_n1970;
  assign new_n1972 = new_n856 & ~new_n859;
  assign new_n1973 = ~new_n856 & new_n1935;
  assign new_n1974 = ~new_n1972 & ~new_n1973;
  assign new_n1975 = ~pv1213_3_ & ~new_n1974;
  assign new_n1976 = pv1213_3_ & new_n1974;
  assign new_n1977 = ~new_n1975 & ~new_n1976;
  assign new_n1978 = new_n856 & ~new_n892;
  assign new_n1979 = ~new_n1942 & ~new_n1948;
  assign new_n1980 = ~new_n1949 & ~new_n1979;
  assign new_n1981 = ~new_n856 & ~new_n1980;
  assign new_n1982 = ~new_n1978 & ~new_n1981;
  assign new_n1983 = ~pv1213_1_ & ~new_n1982;
  assign new_n1984 = pv1213_1_ & new_n1982;
  assign new_n1985 = ~new_n1983 & ~new_n1984;
  assign new_n1986 = ~pv288_4_ & ~pv288_5_;
  assign new_n1987 = new_n1963 & new_n1971;
  assign new_n1988 = new_n1977 & new_n1987;
  assign new_n1989 = new_n1985 & new_n1988;
  assign new_n1990 = ~new_n842 & new_n1989;
  assign new_n1991 = ~new_n1986 & new_n1990;
  assign new_n1992 = ~pv1213_0_ & ~new_n1955;
  assign new_n1993 = pv1213_0_ & new_n1955;
  assign new_n1994 = ~new_n1992 & ~new_n1993;
  assign new_n1995 = ~pv1213_2_ & ~new_n1941;
  assign new_n1996 = pv1213_2_ & new_n1941;
  assign new_n1997 = ~new_n1995 & ~new_n1996;
  assign new_n1998 = ~pv1213_3_ & ~new_n1935;
  assign new_n1999 = pv1213_3_ & new_n1935;
  assign new_n2000 = ~new_n1998 & ~new_n1999;
  assign new_n2001 = ~pv1213_1_ & ~new_n1948;
  assign new_n2002 = pv1213_1_ & new_n1948;
  assign new_n2003 = ~new_n2001 & ~new_n2002;
  assign new_n2004 = new_n1994 & new_n1997;
  assign new_n2005 = new_n2000 & new_n2004;
  assign new_n2006 = new_n2003 & new_n2005;
  assign new_n2007 = ~new_n842 & new_n2006;
  assign new_n2008 = pv288_4_ & new_n2007;
  assign new_n2009 = ~new_n1991 & ~new_n2008;
  assign new_n2010 = new_n616 & new_n2009;
  assign new_n2011 = ~new_n956 & ~new_n1057;
  assign new_n2012 = new_n616 & new_n2011;
  assign new_n2013 = new_n2010 & new_n2012;
  assign new_n2014 = new_n881 & ~new_n2013;
  assign new_n2015 = ~new_n1765 & ~new_n1848;
  assign new_n2016 = ~new_n1931 & ~new_n2014;
  assign new_n2017 = new_n2015 & new_n2016;
  assign new_n2018 = ~pv172_0_ & pv240_0_;
  assign pv1719 = ~new_n699 & new_n2018;
  assign new_n2020 = pv1243_7_ & pv1243_9_;
  assign new_n2021 = ~new_n2017 & new_n2020;
  assign new_n2022 = pv1243_8_ & new_n2021;
  assign new_n2023 = ~pv248_0_ & new_n2022;
  assign new_n2024 = pv1719 & new_n2023;
  assign new_n2025 = pv243_0_ & pv244_0_;
  assign new_n2026 = pv245_0_ & new_n2025;
  assign new_n2027 = pv246_0_ & new_n2026;
  assign new_n2028 = pv247_0_ & new_n2027;
  assign new_n2029 = pv1719 & new_n2028;
  assign new_n2030 = ~pv248_0_ & new_n2029;
  assign new_n2031 = new_n1380 & pv1719;
  assign new_n2032 = ~pv248_0_ & new_n2031;
  assign new_n2033 = ~new_n2024 & ~new_n2030;
  assign pv393_0_ = new_n2032 | ~new_n2033;
  assign pv500_0_ = pv271_0_ | ~pv14_0_;
  assign pv544 = new_n491 & pv1213_7_;
  assign new_n2037 = pv257_2_ & pv257_1_;
  assign new_n2038 = pv257_5_ & new_n2037;
  assign new_n2039 = pv257_3_ & new_n2038;
  assign new_n2040 = pv257_7_ & new_n2039;
  assign new_n2041 = pv257_4_ & new_n2040;
  assign new_n2042 = pv257_6_ & new_n2041;
  assign new_n2043 = pv257_0_ & ~new_n2042;
  assign new_n2044 = ~pv257_0_ & new_n2042;
  assign pv650 = new_n2043 | new_n2044;
  assign new_n2046 = pv213_3_ & new_n1704;
  assign new_n2047 = ~new_n1589 & new_n2046;
  assign new_n2048 = pv165_5_ & new_n1586;
  assign pv1297_2_ = new_n2047 | new_n2048;
  assign new_n2050 = ~pv88_3_ & new_n572;
  assign new_n2051 = ~pv134_1_ & ~new_n572;
  assign pv1771_1_ = new_n2050 | new_n2051;
  assign new_n2053 = pv100_0_ & new_n1721;
  assign new_n2054 = pv124_0_ & new_n1725;
  assign new_n2055 = pv213_0_ & new_n1728;
  assign new_n2056 = pv108_0_ & new_n1732;
  assign new_n2057 = ~new_n2053 & ~new_n2054;
  assign new_n2058 = ~new_n2055 & ~new_n2056;
  assign pv1921_0_ = ~new_n2057 | ~new_n2058;
  assign new_n2060 = pv802_0_ & ~new_n639;
  assign new_n2061 = ~new_n1388 & ~new_n2060;
  assign new_n2062 = pv134_1_ & ~pv134_0_;
  assign new_n2063 = ~pv134_1_ & pv134_0_;
  assign new_n2064 = ~new_n2062 & ~new_n2063;
  assign new_n2065 = ~new_n2060 & ~new_n2061;
  assign new_n2066 = new_n1388 & new_n2065;
  assign new_n2067 = ~new_n2064 & new_n2066;
  assign new_n2068 = new_n1388 & ~new_n2060;
  assign new_n2069 = ~new_n1388 & ~new_n2068;
  assign new_n2070 = ~new_n2060 & new_n2069;
  assign new_n2071 = pv134_0_ & new_n2070;
  assign pv1992_0_ = new_n2067 | new_n2071;
  assign pv541 = new_n491 & pv1213_4_;
  assign new_n2074 = ~pv214_0_ & ~new_n699;
  assign new_n2075 = new_n1285 & new_n2074;
  assign new_n2076 = ~new_n704 & new_n2075;
  assign new_n2077 = ~new_n557 & ~new_n1279;
  assign new_n2078 = pv59_0_ & ~new_n699;
  assign new_n2079 = ~new_n2077 & new_n2078;
  assign new_n2080 = ~pv214_0_ & new_n2079;
  assign new_n2081 = pv62_0_ & ~new_n699;
  assign new_n2082 = new_n1132 & new_n2081;
  assign new_n2083 = ~pv214_0_ & new_n2082;
  assign new_n2084 = ~new_n2076 & ~new_n2080;
  assign pv620 = ~new_n2083 & new_n2084;
  assign new_n2086 = pv62_0_ & new_n758;
  assign new_n2087 = new_n557 & new_n2086;
  assign new_n2088 = pv14_0_ & new_n2087;
  assign new_n2089 = ~new_n491 & ~new_n1280;
  assign new_n2090 = ~new_n573 & ~new_n773;
  assign new_n2091 = new_n2089 & new_n2090;
  assign new_n2092 = ~new_n494 & ~new_n575;
  assign new_n2093 = ~new_n766 & new_n2092;
  assign new_n2094 = new_n2091 & new_n2093;
  assign new_n2095 = ~pv174_0_ & new_n585;
  assign new_n2096 = new_n2094 & ~new_n2095;
  assign new_n2097 = pv59_0_ & new_n2096;
  assign new_n2098 = ~new_n713 & new_n2097;
  assign new_n2099 = ~pv1719 & new_n2098;
  assign new_n2100 = pv14_0_ & new_n2099;
  assign new_n2101 = ~new_n841 & new_n2100;
  assign new_n2102 = new_n758 & new_n2101;
  assign pv1274_0_ = new_n2088 | new_n2102;
  assign new_n2104 = pv213_4_ & new_n1704;
  assign new_n2105 = ~new_n1589 & new_n2104;
  assign new_n2106 = pv165_6_ & new_n1586;
  assign pv1297_3_ = new_n2105 | new_n2106;
  assign pv1432 = pv66_0_ & new_n1628;
  assign new_n2109 = pv242_0_ & new_n639;
  assign new_n2110 = pv14_0_ & new_n2109;
  assign new_n2111 = ~pv1536_0_ & new_n1381;
  assign new_n2112 = ~new_n640 & new_n2111;
  assign pv1726_0_ = new_n2110 | new_n2112;
  assign new_n2114 = pv100_3_ & new_n1721;
  assign new_n2115 = pv124_3_ & new_n1725;
  assign new_n2116 = pv213_3_ & new_n1728;
  assign new_n2117 = pv108_3_ & new_n1732;
  assign new_n2118 = ~new_n2114 & ~new_n2115;
  assign new_n2119 = ~new_n2116 & ~new_n2117;
  assign pv1921_3_ = ~new_n2118 | ~new_n2119;
  assign new_n2121 = pv101_0_ & new_n1152;
  assign new_n2122 = ~pv108_4_ & new_n2121;
  assign new_n2123 = pv56_0_ & new_n1096;
  assign new_n2124 = pv14_0_ & ~new_n2122;
  assign new_n2125 = ~new_n2123 & new_n2124;
  assign new_n2126 = pv110_0_ & new_n2125;
  assign new_n2127 = ~pv102_0_ & ~pv1758_0_;
  assign new_n2128 = new_n510 & ~new_n2127;
  assign new_n2129 = ~pv110_0_ & new_n2128;
  assign pv1968_0_ = new_n2126 | new_n2129;
  assign new_n2131 = ~pv134_1_ & new_n2066;
  assign new_n2132 = pv134_1_ & new_n2070;
  assign pv1992_1_ = new_n2131 | new_n2132;
  assign new_n2134 = ~new_n1759 & ~new_n2008;
  assign new_n2135 = ~new_n1842 & new_n2134;
  assign new_n2136 = ~new_n1925 & new_n2135;
  assign new_n2137 = new_n616 & new_n2136;
  assign new_n2138 = ~new_n939 & new_n2137;
  assign new_n2139 = ~new_n1005 & new_n2138;
  assign new_n2140 = ~new_n848 & new_n2139;
  assign pv357 = ~new_n956 & new_n2140;
  assign new_n2142 = new_n505 & new_n616;
  assign new_n2143 = new_n545 & new_n2142;
  assign new_n2144 = new_n549 & new_n2143;
  assign new_n2145 = pv802_0_ & ~new_n2144;
  assign new_n2146 = ~new_n557 & new_n774;
  assign new_n2147 = ~pv174_0_ & ~new_n555;
  assign new_n2148 = new_n2146 & new_n2147;
  assign new_n2149 = pv56_0_ & ~new_n2148;
  assign new_n2150 = new_n616 & new_n1215;
  assign new_n2151 = pv59_0_ & ~new_n2150;
  assign new_n2152 = pv70_0_ & ~new_n616;
  assign new_n2153 = pv802_0_ & new_n1502;
  assign new_n2154 = ~pv215_0_ & pv66_0_;
  assign new_n2155 = pv763 & new_n2154;
  assign new_n2156 = ~new_n699 & new_n2155;
  assign new_n2157 = ~new_n2145 & ~new_n2149;
  assign new_n2158 = ~new_n1212 & ~new_n2151;
  assign new_n2159 = new_n2157 & new_n2158;
  assign new_n2160 = ~new_n2152 & ~new_n2153;
  assign new_n2161 = ~pv1719 & ~new_n2156;
  assign new_n2162 = new_n2160 & new_n2161;
  assign pv423_0_ = ~new_n2159 | ~new_n2162;
  assign pv542 = new_n491 & pv1213_5_;
  assign new_n2165 = pv41_0_ & ~pv45_0_;
  assign new_n2166 = ~pv41_0_ & pv45_0_;
  assign new_n2167 = ~new_n2165 & ~new_n2166;
  assign pv621 = pv293_0_ & new_n2167;
  assign new_n2169 = pv62_0_ & new_n572;
  assign new_n2170 = pv56_0_ & new_n572;
  assign new_n2171 = ~new_n491 & ~new_n573;
  assign new_n2172 = ~new_n575 & new_n2171;
  assign new_n2173 = pv802_0_ & ~new_n2172;
  assign new_n2174 = new_n507 & new_n2173;
  assign new_n2175 = new_n507 & ~new_n732;
  assign new_n2176 = pv59_0_ & new_n2175;
  assign new_n2177 = ~new_n2170 & ~new_n2174;
  assign new_n2178 = ~pv270_0_ & ~new_n2176;
  assign new_n2179 = new_n2177 & new_n2178;
  assign new_n2180 = ~pv302_0_ & ~new_n2169;
  assign pv630 = ~new_n2179 & new_n2180;
  assign new_n2182 = pv213_5_ & new_n1704;
  assign new_n2183 = ~new_n1589 & new_n2182;
  assign new_n2184 = pv165_7_ & new_n1586;
  assign pv1297_4_ = new_n2183 | new_n2184;
  assign new_n2186 = pv100_2_ & new_n1721;
  assign new_n2187 = pv124_2_ & new_n1725;
  assign new_n2188 = pv213_2_ & new_n1728;
  assign new_n2189 = pv108_2_ & new_n1732;
  assign new_n2190 = ~new_n2186 & ~new_n2187;
  assign new_n2191 = ~new_n2188 & ~new_n2189;
  assign pv1921_2_ = ~new_n2190 | ~new_n2191;
  assign pv547 = new_n491 & pv1213_10_;
  assign new_n2194 = pv257_6_ & pv257_7_;
  assign new_n2195 = pv257_5_ & ~new_n2194;
  assign new_n2196 = ~pv257_5_ & new_n2194;
  assign pv655 = new_n2195 | new_n2196;
  assign new_n2198 = ~pv259_0_ & new_n1661;
  assign new_n2199 = pv259_0_ & new_n1663;
  assign new_n2200 = ~new_n2198 & ~new_n2199;
  assign new_n2201 = pv14_0_ & new_n2200;
  assign new_n2202 = pv260_0_ & new_n2201;
  assign new_n2203 = pv14_0_ & ~new_n2200;
  assign new_n2204 = ~pv260_0_ & new_n2203;
  assign pv1467_0_ = new_n2202 | new_n2204;
  assign new_n2206 = pv62_0_ & pv91_1_;
  assign new_n2207 = pv59_0_ & pv91_0_;
  assign new_n2208 = ~new_n2206 & ~new_n2207;
  assign new_n2209 = new_n1223 & ~new_n2208;
  assign new_n2210 = ~pv294_0_ & ~new_n1279;
  assign new_n2211 = ~new_n1132 & new_n2210;
  assign new_n2212 = new_n2167 & ~new_n2209;
  assign pv1629_0_ = new_n2211 | ~new_n2212;
  assign new_n2214 = pv108_0_ & ~new_n1714;
  assign new_n2215 = ~new_n1278 & ~new_n2214;
  assign pv1896_0_ = new_n1153 | ~new_n2215;
  assign new_n2217 = pv213_5_ & new_n1728;
  assign new_n2218 = pv100_5_ & new_n1721;
  assign new_n2219 = pv124_5_ & new_n1725;
  assign new_n2220 = ~new_n2217 & ~new_n2218;
  assign pv1921_5_ = new_n2219 | ~new_n2220;
  assign new_n2222 = ~pv35_0_ & ~new_n1496;
  assign pv377 = pv203_0_ & ~new_n2222;
  assign pv548 = new_n491 & pv1213_11_;
  assign new_n2225 = pv257_6_ & pv257_5_;
  assign new_n2226 = pv257_7_ & new_n2225;
  assign new_n2227 = pv257_4_ & ~new_n2226;
  assign new_n2228 = ~pv257_4_ & new_n2226;
  assign pv654 = new_n2227 | new_n2228;
  assign new_n2230 = new_n494 & pv802_0_;
  assign new_n2231 = ~pv279_0_ & ~new_n2230;
  assign new_n2232 = pv149_5_ & new_n2230;
  assign pv821_0_ = new_n2231 | new_n2232;
  assign new_n2234 = new_n491 & new_n1278;
  assign new_n2235 = pv108_1_ & ~new_n1714;
  assign pv1897_0_ = new_n2234 | new_n2235;
  assign new_n2237 = pv100_4_ & new_n1721;
  assign new_n2238 = pv124_4_ & new_n1725;
  assign new_n2239 = pv213_4_ & new_n1728;
  assign new_n2240 = pv108_4_ & new_n1732;
  assign new_n2241 = ~new_n2237 & ~new_n2238;
  assign new_n2242 = ~new_n2239 & ~new_n2240;
  assign pv1921_4_ = ~new_n2241 | ~new_n2242;
  assign new_n2244 = pv56_0_ & new_n773;
  assign new_n2245 = pv59_0_ & ~new_n545;
  assign new_n2246 = ~new_n554 & new_n2245;
  assign new_n2247 = pv56_0_ & new_n766;
  assign new_n2248 = pv59_0_ & ~new_n505;
  assign new_n2249 = ~new_n786 & ~new_n2244;
  assign new_n2250 = ~new_n2246 & new_n2249;
  assign new_n2251 = ~new_n2247 & new_n2250;
  assign new_n2252 = ~new_n1212 & new_n2251;
  assign new_n2253 = ~new_n2248 & new_n2252;
  assign new_n2254 = ~pv43_0_ & ~new_n699;
  assign new_n2255 = ~pv214_0_ & new_n2254;
  assign new_n2256 = ~new_n2253 & new_n2255;
  assign pv527 = ~new_n704 & new_n2256;
  assign pv538 = new_n491 & pv1213_1_;
  assign pv545 = new_n491 & pv1213_8_;
  assign new_n2260 = pv257_4_ & new_n2225;
  assign new_n2261 = pv257_7_ & new_n2260;
  assign new_n2262 = pv257_3_ & ~new_n2261;
  assign new_n2263 = ~pv257_3_ & new_n2261;
  assign pv653 = new_n2262 | new_n2263;
  assign new_n2265 = pv37_0_ & ~pv1213_2_;
  assign new_n2266 = ~pv37_0_ & pv321_2_;
  assign pv1829_0_ = new_n2265 | new_n2266;
  assign new_n2268 = new_n490 & new_n719;
  assign new_n2269 = pv108_2_ & ~new_n1714;
  assign pv1898_0_ = new_n2268 | new_n2269;
  assign pv537 = new_n491 & pv1213_0_;
  assign pv546 = new_n491 & pv1213_9_;
  assign new_n2273 = ~new_n1689 & ~new_n2025;
  assign new_n2274 = pv245_0_ & new_n2273;
  assign new_n2275 = ~new_n1689 & new_n2025;
  assign new_n2276 = ~pv245_0_ & new_n2275;
  assign pv597_0_ = new_n2274 | new_n2276;
  assign new_n2278 = pv257_4_ & pv257_6_;
  assign new_n2279 = pv257_5_ & new_n2278;
  assign new_n2280 = pv257_3_ & new_n2279;
  assign new_n2281 = pv257_7_ & new_n2280;
  assign new_n2282 = pv257_2_ & ~new_n2281;
  assign new_n2283 = ~pv257_2_ & new_n2281;
  assign pv652 = new_n2282 | new_n2283;
  assign pv801 = new_n579 & new_n586;
  assign new_n2286 = new_n510 & new_n719;
  assign new_n2287 = pv108_3_ & ~new_n1714;
  assign pv1899_0_ = new_n2286 | new_n2287;
  assign new_n2289 = ~pv802_0_ & new_n1502;
  assign new_n2290 = ~new_n1392 & ~new_n2289;
  assign new_n2291 = new_n575 & pv802_0_;
  assign new_n2292 = new_n2290 & ~new_n2291;
  assign new_n2293 = pv802_0_ & new_n2292;
  assign new_n2294 = new_n491 & new_n2293;
  assign new_n2295 = pv1243_8_ & new_n2294;
  assign new_n2296 = new_n491 & pv802_0_;
  assign new_n2297 = ~pv199_4_ & pv199_3_;
  assign new_n2298 = pv199_4_ & ~pv199_3_;
  assign new_n2299 = ~new_n2297 & ~new_n2298;
  assign new_n2300 = ~new_n2291 & ~new_n2296;
  assign new_n2301 = ~new_n2290 & new_n2300;
  assign new_n2302 = ~new_n2299 & new_n2301;
  assign pv572_8_ = new_n2295 | new_n2302;
  assign new_n2304 = ~new_n510 & ~new_n567;
  assign new_n2305 = pv290_0_ & ~new_n2304;
  assign new_n2306 = new_n699 & new_n2305;
  assign new_n2307 = pv56_0_ & new_n1718;
  assign new_n2308 = pv14_0_ & ~new_n2306;
  assign new_n2309 = pv100_2_ & new_n2308;
  assign new_n2310 = ~new_n2307 & new_n2309;
  assign new_n2311 = pv165_4_ & new_n2306;
  assign pv1709_1_ = new_n2310 | new_n2311;
  assign pv373 = pv10_0_ & pv13_0_;
  assign new_n2314 = pv1243_7_ & new_n2294;
  assign new_n2315 = pv199_4_ & pv199_3_;
  assign new_n2316 = pv199_2_ & ~new_n2315;
  assign new_n2317 = ~pv199_2_ & new_n2315;
  assign new_n2318 = ~new_n2316 & ~new_n2317;
  assign new_n2319 = new_n2301 & ~new_n2318;
  assign pv572_7_ = new_n2314 | new_n2319;
  assign new_n2321 = ~pv149_6_ & new_n582;
  assign new_n2322 = pv14_0_ & ~new_n491;
  assign new_n2323 = pv277_0_ & new_n2322;
  assign pv1439_0_ = new_n2321 | new_n2323;
  assign new_n2325 = pv100_1_ & new_n2308;
  assign new_n2326 = ~new_n2307 & new_n2325;
  assign new_n2327 = pv165_3_ & new_n2306;
  assign pv1709_0_ = new_n2326 | new_n2327;
  assign new_n2329 = pv1243_6_ & new_n2294;
  assign new_n2330 = pv199_3_ & pv199_2_;
  assign new_n2331 = pv199_4_ & new_n2330;
  assign new_n2332 = pv199_1_ & ~new_n2331;
  assign new_n2333 = ~pv199_1_ & new_n2331;
  assign new_n2334 = ~new_n2332 & ~new_n2333;
  assign new_n2335 = new_n2301 & ~new_n2334;
  assign pv572_6_ = new_n2329 | new_n2335;
  assign new_n2337 = ~pv69_0_ & ~pv50_0_;
  assign pv1539 = new_n1628 & ~new_n2337;
  assign new_n2339 = pv1243_5_ & new_n2294;
  assign new_n2340 = pv199_1_ & new_n2330;
  assign new_n2341 = pv199_4_ & new_n2340;
  assign new_n2342 = pv199_0_ & ~new_n2341;
  assign new_n2343 = ~pv199_0_ & new_n2341;
  assign new_n2344 = ~new_n2342 & ~new_n2343;
  assign new_n2345 = new_n2301 & ~new_n2344;
  assign pv572_5_ = new_n2339 | new_n2345;
  assign new_n2347 = pv165_3_ & ~pv165_5_;
  assign new_n2348 = new_n758 & new_n2347;
  assign new_n2349 = pv763 & new_n2348;
  assign new_n2350 = pv14_0_ & new_n2349;
  assign new_n2351 = pv70_0_ & new_n2350;
  assign new_n2352 = ~pv165_4_ & new_n2351;
  assign new_n2353 = pv165_6_ & new_n2352;
  assign new_n2354 = pv65_0_ & ~new_n555;
  assign new_n2355 = new_n758 & new_n2354;
  assign new_n2356 = ~new_n1132 & new_n2355;
  assign new_n2357 = pv14_0_ & new_n2356;
  assign pv1392_0_ = new_n2353 | new_n2357;
  assign new_n2359 = pv258_0_ & ~pv259_0_;
  assign new_n2360 = ~pv260_0_ & new_n2359;
  assign new_n2361 = ~pv59_0_ & new_n2360;
  assign new_n2362 = pv262_0_ & ~new_n2361;
  assign new_n2363 = pv14_0_ & new_n2362;
  assign pv1679_0_ = ~new_n615 | new_n2363;
  assign new_n2365 = new_n616 & ~new_n842;
  assign new_n2366 = ~new_n1755 & ~new_n1991;
  assign new_n2367 = ~new_n1825 & new_n2366;
  assign new_n2368 = ~new_n1908 & new_n2367;
  assign new_n2369 = new_n2365 & new_n2368;
  assign new_n2370 = ~new_n1083 & new_n2369;
  assign new_n2371 = ~new_n1031 & new_n2370;
  assign new_n2372 = ~new_n854 & new_n2371;
  assign pv356 = ~new_n1057 & new_n2372;
  assign new_n2374 = pv215_0_ & pv66_0_;
  assign new_n2375 = pv66_0_ & new_n762;
  assign new_n2376 = pv66_0_ & pv763;
  assign new_n2377 = new_n493 & pv802_0_;
  assign new_n2378 = ~new_n491 & ~new_n511;
  assign new_n2379 = ~pv763 & ~new_n2378;
  assign new_n2380 = pv802_0_ & new_n2379;
  assign new_n2381 = ~new_n713 & ~new_n1132;
  assign new_n2382 = ~new_n1133 & ~new_n1223;
  assign new_n2383 = new_n2381 & new_n2382;
  assign new_n2384 = pv56_0_ & ~new_n2383;
  assign new_n2385 = ~new_n2375 & ~new_n2376;
  assign new_n2386 = ~new_n2377 & new_n2385;
  assign new_n2387 = ~new_n2380 & ~new_n2384;
  assign new_n2388 = new_n2386 & new_n2387;
  assign new_n2389 = ~pv32_1_ & ~new_n997;
  assign new_n2390 = pv32_1_ & new_n997;
  assign new_n2391 = ~new_n2389 & ~new_n2390;
  assign new_n2392 = ~pv32_0_ & ~new_n973;
  assign new_n2393 = pv32_0_ & new_n973;
  assign new_n2394 = ~new_n2392 & ~new_n2393;
  assign new_n2395 = ~pv32_2_ & ~new_n982;
  assign new_n2396 = pv32_2_ & new_n982;
  assign new_n2397 = ~new_n2395 & ~new_n2396;
  assign new_n2398 = new_n988 & new_n2391;
  assign new_n2399 = new_n2394 & new_n2398;
  assign new_n2400 = pv32_3_ & new_n2399;
  assign new_n2401 = new_n2397 & new_n2400;
  assign new_n2402 = new_n2390 & new_n2394;
  assign new_n2403 = new_n982 & new_n2394;
  assign new_n2404 = pv32_2_ & new_n2403;
  assign new_n2405 = new_n2391 & new_n2404;
  assign new_n2406 = ~new_n2393 & ~new_n2401;
  assign new_n2407 = ~new_n2402 & ~new_n2405;
  assign new_n2408 = new_n2406 & new_n2407;
  assign new_n2409 = ~new_n2388 & ~new_n2408;
  assign new_n2410 = new_n1496 & pv1719;
  assign new_n2411 = new_n702 & pv1719;
  assign new_n2412 = pv302_0_ & pv1719;
  assign new_n2413 = ~new_n554 & ~pv763;
  assign new_n2414 = pv802_0_ & ~new_n2413;
  assign new_n2415 = ~new_n2374 & ~new_n2409;
  assign new_n2416 = ~pv43_0_ & new_n2415;
  assign new_n2417 = new_n616 & new_n2416;
  assign new_n2418 = ~pv214_0_ & new_n2417;
  assign new_n2419 = ~new_n2032 & new_n2418;
  assign new_n2420 = ~new_n2024 & new_n2419;
  assign new_n2421 = ~new_n2410 & new_n2420;
  assign new_n2422 = ~new_n2030 & new_n2421;
  assign new_n2423 = ~new_n2411 & new_n2422;
  assign new_n2424 = ~new_n2412 & new_n2423;
  assign new_n2425 = pv423_0_ & new_n2424;
  assign new_n2426 = ~new_n1278 & new_n2425;
  assign new_n2427 = ~new_n704 & new_n2426;
  assign new_n2428 = ~pv1757_0_ & new_n2427;
  assign pv432 = ~new_n2414 & new_n2428;
  assign pv435_0_ = pv630 | pv432;
  assign new_n2431 = pv216_0_ & ~pv214_0_;
  assign new_n2432 = ~pv68_0_ & ~pv69_0_;
  assign new_n2433 = ~pv66_0_ & new_n2432;
  assign new_n2434 = ~pv70_0_ & new_n2433;
  assign new_n2435 = pv14_0_ & new_n730;
  assign new_n2436 = ~new_n2434 & new_n2435;
  assign new_n2437 = pv215_0_ & new_n2436;
  assign pv1492_0_ = new_n2431 | new_n2437;
  assign pv1537 = pv68_0_ & new_n1628;
  assign new_n2440 = ~pv43_0_ & pv45_0_;
  assign pv511_0_ = pv40_0_ | new_n2440;
  assign pv540 = new_n491 & pv1213_3_;
  assign new_n2443 = ~new_n1689 & ~new_n2027;
  assign new_n2444 = pv247_0_ & new_n2443;
  assign new_n2445 = ~new_n1689 & new_n2027;
  assign new_n2446 = ~pv247_0_ & new_n2445;
  assign pv609_0_ = new_n2444 | new_n2446;
  assign pv1426 = pv1_0_ & new_n692;
  assign new_n2449 = ~pv302_0_ & pv292_0_;
  assign new_n2450 = pv174_0_ & new_n699;
  assign new_n2451 = pv174_0_ & ~new_n755;
  assign new_n2452 = ~new_n579 & ~new_n2449;
  assign new_n2453 = ~new_n2450 & ~new_n2451;
  assign pv1620_0_ = ~new_n2452 | ~new_n2453;
  assign new_n2455 = ~pv290_0_ & ~pv802_0_;
  assign new_n2456 = new_n702 & new_n2455;
  assign new_n2457 = new_n732 & new_n2456;
  assign pv1736 = ~pv289_0_ & new_n2457;
  assign pv1429 = pv1_0_ & pv12_0_;
  assign new_n2460 = ~new_n1490 & ~new_n2363;
  assign new_n2461 = pv262_0_ & new_n2460;
  assign new_n2462 = pv261_0_ & ~new_n2461;
  assign new_n2463 = ~new_n1662 & ~new_n2462;
  assign pv1832 = pv14_0_ & ~new_n2463;
  assign new_n2465 = pv1243_9_ & new_n2294;
  assign new_n2466 = ~pv199_4_ & new_n2301;
  assign pv572_9_ = new_n2465 | new_n2466;
  assign new_n2468 = pv213_1_ & new_n1704;
  assign new_n2469 = ~new_n1589 & new_n2468;
  assign new_n2470 = pv165_3_ & new_n1586;
  assign pv1297_0_ = new_n2469 | new_n2470;
  assign pv1428 = pv1_0_ & pv11_0_;
  assign new_n2473 = new_n1583 & ~new_n2304;
  assign new_n2474 = ~new_n2306 & ~new_n2473;
  assign new_n2475 = pv14_0_ & new_n2474;
  assign new_n2476 = pv100_0_ & new_n2475;
  assign new_n2477 = ~new_n2307 & new_n2476;
  assign new_n2478 = ~new_n1595 & ~new_n2474;
  assign pv1693_0_ = new_n2477 | new_n2478;
  assign new_n2480 = pv108_5_ & ~new_n1404;
  assign pv1901_0_ = new_n1308 | new_n2480;
  assign new_n2482 = pv194_0_ & ~new_n1380;
  assign new_n2483 = ~pv194_0_ & new_n1380;
  assign new_n2484 = ~new_n2482 & ~new_n2483;
  assign new_n2485 = new_n2301 & ~new_n2484;
  assign new_n2486 = new_n2290 & ~new_n2296;
  assign new_n2487 = pv802_0_ & new_n2486;
  assign new_n2488 = new_n575 & new_n2487;
  assign new_n2489 = pv149_4_ & new_n2488;
  assign new_n2490 = ~pv321_2_ & new_n2294;
  assign new_n2491 = ~new_n2485 & ~new_n2489;
  assign pv572_0_ = new_n2490 | ~new_n2491;
  assign new_n2493 = pv239_4_ & ~pv239_3_;
  assign new_n2494 = ~pv239_4_ & pv239_3_;
  assign new_n2495 = ~new_n2493 & ~new_n2494;
  assign new_n2496 = ~pv802_0_ & ~new_n694;
  assign new_n2497 = new_n494 & new_n2496;
  assign new_n2498 = ~new_n2495 & new_n2497;
  assign new_n2499 = new_n494 & ~pv802_0_;
  assign new_n2500 = new_n694 & ~new_n2499;
  assign new_n2501 = pv1243_8_ & new_n2500;
  assign pv1552_0_ = new_n2498 | new_n2501;
  assign new_n2503 = pv33_0_ & ~new_n490;
  assign new_n2504 = pv289_0_ & new_n2503;
  assign pv1745_0_ = new_n585 | ~new_n2504;
  assign new_n2506 = pv37_0_ & ~pv1243_9_;
  assign pv1829_9_ = new_n2266 | new_n2506;
  assign new_n2508 = pv149_3_ & ~new_n1093;
  assign new_n2509 = ~new_n1713 & new_n2508;
  assign new_n2510 = new_n567 & new_n2509;
  assign new_n2511 = ~new_n841 & new_n2510;
  assign new_n2512 = pv149_5_ & new_n567;
  assign new_n2513 = ~pv149_3_ & new_n2512;
  assign new_n2514 = pv149_4_ & new_n2513;
  assign new_n2515 = ~pv149_7_ & new_n2514;
  assign new_n2516 = ~pv149_6_ & new_n2515;
  assign new_n2517 = ~pv149_6_ & new_n1717;
  assign new_n2518 = ~new_n2511 & ~new_n2516;
  assign new_n2519 = ~new_n2517 & new_n2518;
  assign new_n2520 = ~pv302_0_ & ~new_n2519;
  assign new_n2521 = pv149_0_ & pv149_1_;
  assign new_n2522 = ~pv149_2_ & new_n2521;
  assign new_n2523 = pv149_0_ & pv149_2_;
  assign new_n2524 = ~pv149_1_ & new_n2523;
  assign new_n2525 = pv149_2_ & new_n2521;
  assign new_n2526 = ~new_n2522 & ~new_n2524;
  assign new_n2527 = new_n2519 & new_n2526;
  assign new_n2528 = ~new_n2525 & new_n2527;
  assign new_n2529 = ~new_n2520 & ~new_n2528;
  assign new_n2530 = new_n616 & new_n2529;
  assign new_n2531 = pv65_0_ & new_n1132;
  assign new_n2532 = pv258_0_ & ~pv260_0_;
  assign new_n2533 = ~new_n616 & new_n2532;
  assign new_n2534 = ~pv259_0_ & new_n2533;
  assign new_n2535 = ~pv59_0_ & new_n2534;
  assign new_n2536 = ~new_n1718 & ~new_n2535;
  assign new_n2537 = ~new_n1224 & new_n2536;
  assign new_n2538 = ~new_n1095 & new_n2537;
  assign new_n2539 = ~new_n2321 & new_n2538;
  assign new_n2540 = ~new_n1096 & new_n2539;
  assign new_n2541 = ~new_n1588 & new_n2540;
  assign new_n2542 = pv56_0_ & ~new_n2541;
  assign new_n2543 = pv62_0_ & ~new_n2382;
  assign new_n2544 = ~new_n2531 & ~new_n2542;
  assign new_n2545 = ~new_n2543 & new_n2544;
  assign new_n2546 = ~pv1741_0_ & ~new_n2545;
  assign new_n2547 = ~new_n702 & new_n2546;
  assign new_n2548 = new_n758 & ~new_n1496;
  assign new_n2549 = ~new_n732 & ~new_n2548;
  assign new_n2550 = pv290_0_ & ~new_n699;
  assign new_n2551 = ~pv289_0_ & ~new_n2547;
  assign new_n2552 = ~pv214_0_ & ~new_n2549;
  assign new_n2553 = new_n2551 & new_n2552;
  assign new_n2554 = ~pv302_0_ & ~new_n701;
  assign new_n2555 = ~new_n2550 & new_n2554;
  assign new_n2556 = new_n2553 & new_n2555;
  assign new_n2557 = ~new_n2530 & new_n2556;
  assign pv798_0_ = ~pv14_0_ | ~new_n2557;
  assign new_n2559 = ~pv239_4_ & new_n2497;
  assign new_n2560 = pv1243_9_ & new_n2500;
  assign pv1552_1_ = new_n2559 | new_n2560;
  assign new_n2562 = pv802_0_ & new_n791;
  assign new_n2563 = ~new_n1580 & ~new_n2562;
  assign pv1645_0_ = new_n2409 | ~new_n2563;
  assign new_n2565 = new_n507 & ~new_n2172;
  assign new_n2566 = pv295_0_ & ~new_n2565;
  assign new_n2567 = new_n616 & new_n2566;
  assign new_n2568 = ~pv249_0_ & new_n2567;
  assign new_n2569 = ~pv289_0_ & new_n2568;
  assign pv1652_0_ = pv290_0_ | ~new_n2569;
  assign new_n2571 = ~new_n1689 & ~new_n2026;
  assign new_n2572 = pv246_0_ & new_n2571;
  assign new_n2573 = ~new_n1689 & new_n2026;
  assign new_n2574 = ~pv246_0_ & new_n2573;
  assign pv603_0_ = new_n2572 | new_n2574;
  assign new_n2576 = pv7_0_ & new_n2060;
  assign pv1378 = new_n692 & new_n2576;
  assign new_n2578 = pv1243_4_ & new_n2294;
  assign new_n2579 = pv199_1_ & pv199_3_;
  assign new_n2580 = pv199_2_ & new_n2579;
  assign new_n2581 = pv199_0_ & new_n2580;
  assign new_n2582 = pv199_4_ & new_n2581;
  assign new_n2583 = pv194_4_ & ~new_n2582;
  assign new_n2584 = ~pv194_4_ & new_n2582;
  assign new_n2585 = ~new_n2583 & ~new_n2584;
  assign new_n2586 = new_n2301 & ~new_n2585;
  assign pv572_4_ = new_n2578 | new_n2586;
  assign new_n2588 = pv149_4_ & new_n2230;
  assign new_n2589 = pv279_0_ & ~new_n2230;
  assign new_n2590 = pv280_0_ & new_n2589;
  assign new_n2591 = ~pv280_0_ & new_n2231;
  assign new_n2592 = ~new_n2588 & ~new_n2590;
  assign pv826_0_ = new_n2591 | ~new_n2592;
  assign new_n2594 = ~pv802_0_ & new_n702;
  assign new_n2595 = ~pv289_0_ & new_n2594;
  assign new_n2596 = pv262_0_ & new_n2363;
  assign new_n2597 = new_n615 & ~new_n2596;
  assign new_n2598 = ~new_n1095 & ~new_n1588;
  assign new_n2599 = ~new_n1096 & ~new_n1718;
  assign new_n2600 = new_n2598 & new_n2599;
  assign new_n2601 = ~new_n1224 & ~new_n2321;
  assign new_n2602 = new_n2597 & new_n2601;
  assign new_n2603 = new_n2600 & new_n2602;
  assign new_n2604 = pv1741_0_ & new_n2603;
  assign new_n2605 = ~pv289_0_ & new_n2604;
  assign new_n2606 = ~new_n1132 & new_n2597;
  assign new_n2607 = ~new_n1133 & new_n2606;
  assign new_n2608 = new_n2603 & new_n2607;
  assign new_n2609 = ~new_n1223 & new_n2608;
  assign new_n2610 = ~new_n701 & ~new_n2609;
  assign new_n2611 = new_n2545 & new_n2610;
  assign new_n2612 = new_n755 & new_n2611;
  assign new_n2613 = ~pv289_0_ & new_n2612;
  assign new_n2614 = ~new_n2595 & ~new_n2605;
  assign new_n2615 = ~new_n2613 & new_n2614;
  assign pv1669 = ~new_n2375 & new_n2615;
  assign new_n2617 = pv199_1_ & pv194_4_;
  assign new_n2618 = pv199_2_ & new_n2617;
  assign new_n2619 = pv199_0_ & new_n2618;
  assign new_n2620 = pv199_4_ & new_n2619;
  assign new_n2621 = pv199_3_ & new_n2620;
  assign new_n2622 = pv194_3_ & ~new_n2621;
  assign new_n2623 = ~pv194_3_ & new_n2621;
  assign new_n2624 = ~new_n2622 & ~new_n2623;
  assign new_n2625 = new_n2301 & ~new_n2624;
  assign new_n2626 = pv149_7_ & new_n2488;
  assign new_n2627 = pv1243_3_ & new_n2294;
  assign new_n2628 = ~new_n2625 & ~new_n2626;
  assign pv572_3_ = new_n2627 | ~new_n2628;
  assign new_n2630 = pv244_0_ & pv587;
  assign new_n2631 = pv243_0_ & ~new_n1689;
  assign new_n2632 = ~pv244_0_ & new_n2631;
  assign pv591_0_ = new_n2630 | new_n2632;
  assign new_n2634 = new_n579 & ~new_n586;
  assign new_n2635 = pv802_0_ & ~new_n2530;
  assign new_n2636 = pv763 & ~new_n1701;
  assign new_n2637 = ~new_n586 & new_n2636;
  assign new_n2638 = pv56_0_ & new_n2637;
  assign new_n2639 = pv56_0_ & ~new_n2519;
  assign new_n2640 = ~new_n2634 & ~new_n2635;
  assign new_n2641 = ~new_n2638 & ~new_n2639;
  assign new_n2642 = new_n2640 & new_n2641;
  assign pv966 = new_n1628 & ~new_n2642;
  assign new_n2644 = pv100_5_ & new_n2308;
  assign new_n2645 = ~new_n2307 & new_n2644;
  assign new_n2646 = pv165_7_ & new_n2306;
  assign pv1709_4_ = new_n2645 | new_n2646;
  assign new_n2648 = pv248_0_ & pv1719;
  assign new_n2649 = ~pv423_0_ & ~new_n2648;
  assign new_n2650 = ~pv43_0_ & ~new_n2411;
  assign new_n2651 = ~new_n2414 & new_n2650;
  assign new_n2652 = ~new_n2649 & new_n2651;
  assign new_n2653 = ~pv214_0_ & new_n2652;
  assign new_n2654 = ~new_n2030 & new_n2653;
  assign new_n2655 = ~new_n2024 & new_n2654;
  assign new_n2656 = ~new_n2410 & new_n2655;
  assign new_n2657 = ~new_n2412 & new_n2656;
  assign pv398_0_ = new_n2032 | ~new_n2657;
  assign new_n2659 = pv194_4_ & pv194_3_;
  assign new_n2660 = pv199_2_ & new_n2659;
  assign new_n2661 = pv199_0_ & new_n2660;
  assign new_n2662 = pv199_4_ & new_n2661;
  assign new_n2663 = pv199_1_ & new_n2662;
  assign new_n2664 = pv199_3_ & new_n2663;
  assign new_n2665 = pv194_2_ & ~new_n2664;
  assign new_n2666 = ~pv194_2_ & new_n2664;
  assign new_n2667 = ~new_n2665 & ~new_n2666;
  assign new_n2668 = new_n2301 & ~new_n2667;
  assign new_n2669 = pv149_6_ & new_n2488;
  assign new_n2670 = pv1243_2_ & new_n2294;
  assign new_n2671 = ~new_n2668 & ~new_n2669;
  assign pv572_2_ = new_n2670 | ~new_n2671;
  assign pv640_0_ = pv271_0_ | new_n1525;
  assign new_n2674 = new_n755 & new_n1699;
  assign new_n2675 = pv1536_0_ & ~new_n2674;
  assign new_n2676 = ~new_n1842 & new_n1926;
  assign new_n2677 = ~new_n939 & new_n2676;
  assign new_n2678 = ~new_n1005 & new_n2677;
  assign new_n2679 = ~new_n1031 & new_n2678;
  assign new_n2680 = ~new_n1083 & new_n2679;
  assign new_n2681 = ~new_n1825 & new_n2680;
  assign new_n2682 = ~pv1536_0_ & ~new_n2681;
  assign pv1512_1_ = new_n2675 | new_n2682;
  assign new_n2684 = pv100_4_ & new_n2308;
  assign new_n2685 = ~new_n2307 & new_n2684;
  assign new_n2686 = pv165_6_ & new_n2306;
  assign pv1709_3_ = new_n2685 | new_n2686;
  assign new_n2688 = pv194_3_ & pv194_2_;
  assign new_n2689 = pv199_2_ & new_n2688;
  assign new_n2690 = pv199_0_ & new_n2689;
  assign new_n2691 = pv199_4_ & new_n2690;
  assign new_n2692 = pv199_3_ & new_n2691;
  assign new_n2693 = pv194_4_ & new_n2692;
  assign new_n2694 = pv199_1_ & new_n2693;
  assign new_n2695 = pv194_1_ & ~new_n2694;
  assign new_n2696 = ~pv194_1_ & new_n2694;
  assign new_n2697 = ~new_n2695 & ~new_n2696;
  assign new_n2698 = new_n2301 & ~new_n2697;
  assign new_n2699 = pv149_5_ & new_n2488;
  assign new_n2700 = pv1243_1_ & new_n2294;
  assign new_n2701 = ~new_n2698 & ~new_n2699;
  assign pv572_1_ = new_n2700 | ~new_n2701;
  assign new_n2703 = new_n2519 & ~new_n2638;
  assign new_n2704 = new_n2541 & new_n2703;
  assign new_n2705 = pv56_0_ & new_n2704;
  assign new_n2706 = pv62_0_ & ~new_n616;
  assign new_n2707 = ~new_n494 & new_n640;
  assign new_n2708 = ~new_n1280 & new_n2707;
  assign new_n2709 = pv59_0_ & ~new_n2708;
  assign new_n2710 = ~new_n2705 & ~new_n2706;
  assign new_n2711 = ~new_n2709 & new_n2710;
  assign pv986 = new_n1628 & ~new_n2711;
  assign new_n2713 = ~new_n1491 & ~new_n1662;
  assign new_n2714 = pv258_0_ & pv14_0_;
  assign new_n2715 = new_n2713 & new_n2714;
  assign new_n2716 = ~pv258_0_ & pv14_0_;
  assign new_n2717 = ~new_n2713 & new_n2716;
  assign pv1451_0_ = new_n2715 | new_n2717;
  assign new_n2719 = new_n755 & ~new_n793;
  assign new_n2720 = ~new_n1699 & new_n2719;
  assign new_n2721 = pv1536_0_ & ~new_n2720;
  assign new_n2722 = ~new_n1842 & new_n2009;
  assign new_n2723 = ~new_n956 & new_n2722;
  assign new_n2724 = ~new_n1005 & new_n2723;
  assign new_n2725 = ~new_n1031 & new_n2724;
  assign new_n2726 = ~new_n1057 & new_n2725;
  assign new_n2727 = ~new_n1825 & new_n2726;
  assign new_n2728 = ~pv1536_0_ & ~new_n2727;
  assign pv1512_2_ = new_n2721 | new_n2728;
  assign new_n2730 = pv1921_1_ & ~pv1921_0_;
  assign new_n2731 = ~pv1921_1_ & pv1921_0_;
  assign new_n2732 = ~new_n2730 & ~new_n2731;
  assign new_n2733 = pv1921_3_ & ~pv1921_2_;
  assign new_n2734 = ~pv1921_3_ & pv1921_2_;
  assign new_n2735 = ~new_n2733 & ~new_n2734;
  assign new_n2736 = new_n2732 & ~new_n2735;
  assign new_n2737 = ~new_n2732 & new_n2735;
  assign new_n2738 = ~new_n2736 & ~new_n2737;
  assign new_n2739 = pv1921_5_ & ~pv1921_4_;
  assign new_n2740 = ~pv1921_5_ & pv1921_4_;
  assign new_n2741 = ~new_n2739 & ~new_n2740;
  assign new_n2742 = ~pv1953_0_ & pv1953_1_;
  assign new_n2743 = pv1953_0_ & ~pv1953_1_;
  assign new_n2744 = ~new_n2742 & ~new_n2743;
  assign new_n2745 = new_n2741 & ~new_n2744;
  assign new_n2746 = ~new_n2741 & new_n2744;
  assign new_n2747 = ~new_n2745 & ~new_n2746;
  assign new_n2748 = new_n2738 & ~new_n2747;
  assign new_n2749 = ~new_n2738 & new_n2747;
  assign pv1613_0_ = ~new_n2748 & ~new_n2749;
  assign new_n2751 = pv100_3_ & new_n2308;
  assign new_n2752 = ~new_n2307 & new_n2751;
  assign new_n2753 = pv165_5_ & new_n2306;
  assign pv1709_2_ = new_n2752 | new_n2753;
  assign pv1243_0_ = ~pv321_2_;
  assign pv657 = ~pv257_7_;
  assign pv1375 = ~pv268_5_;
  assign pv1481_0_ = ~pv214_0_;
  assign pv1671_0_ = ~pv205_0_;
  assign pv1863_0_ = ~pv301_0_;
  assign pv1864_0_ = ~pv302_0_;
  assign pv585_0_ = ~pv34_0_;
  assign pv1760_0_ = ~pv101_0_;
  assign pv1833_0_ = ~pv261_0_;
  assign pv1495_0_ = ~pv175_0_;
endmodule


