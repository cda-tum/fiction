// Benchmark "top" written by ABC on Mon Feb 19 11:52:43 2024

module top ( 
    pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_, pv128_6_,
    pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_,
    pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_  );
  input  pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_,
    pv128_6_, pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_;
  output pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_;
  wire new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n326, new_n327, new_n328, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n374, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n426, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n477, new_n478, new_n479, new_n480, new_n481, new_n482, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779;
  assign new_n267 = ~pv199_1_ & pv199_0_;
  assign new_n268 = pv32_10_ & new_n267;
  assign new_n269 = pv199_1_ & pv199_0_;
  assign new_n270 = pv64_10_ & new_n269;
  assign new_n271 = ~pv199_1_ & ~pv199_0_;
  assign new_n272 = pv96_10_ & new_n271;
  assign new_n273 = pv199_1_ & ~pv199_0_;
  assign new_n274 = ~pv96_10_ & new_n273;
  assign new_n275 = ~new_n272 & ~new_n274;
  assign new_n276 = ~new_n268 & ~new_n270;
  assign pv227_10_ = ~new_n275 | ~new_n276;
  assign new_n278 = pv32_23_ & new_n267;
  assign new_n279 = pv64_23_ & new_n269;
  assign new_n280 = pv96_23_ & new_n271;
  assign new_n281 = ~pv96_23_ & new_n273;
  assign new_n282 = ~new_n280 & ~new_n281;
  assign new_n283 = ~new_n278 & ~new_n279;
  assign pv227_23_ = ~new_n282 | ~new_n283;
  assign new_n285 = ~pv199_0_ & pv199_3_;
  assign new_n286 = pv199_1_ & new_n285;
  assign new_n287 = pv195_0_ & new_n286;
  assign new_n288 = ~pv199_1_ & new_n285;
  assign new_n289 = pv195_0_ & new_n288;
  assign pv266_6_ = new_n287 | new_n289;
  assign new_n291 = pv32_0_ & new_n267;
  assign new_n292 = pv64_0_ & new_n269;
  assign new_n293 = pv96_0_ & new_n271;
  assign new_n294 = ~pv96_0_ & new_n273;
  assign new_n295 = ~new_n293 & ~new_n294;
  assign new_n296 = ~new_n291 & ~new_n292;
  assign pv227_0_ = ~new_n295 | ~new_n296;
  assign new_n298 = pv32_24_ & new_n267;
  assign new_n299 = pv64_24_ & new_n269;
  assign new_n300 = pv96_24_ & new_n271;
  assign new_n301 = ~pv96_24_ & new_n273;
  assign new_n302 = ~new_n300 & ~new_n301;
  assign new_n303 = ~new_n298 & ~new_n299;
  assign pv227_24_ = ~new_n302 | ~new_n303;
  assign new_n305 = pv32_21_ & new_n267;
  assign new_n306 = pv64_21_ & new_n269;
  assign new_n307 = pv96_21_ & new_n271;
  assign new_n308 = ~pv96_21_ & new_n273;
  assign new_n309 = ~new_n307 & ~new_n308;
  assign new_n310 = ~new_n305 & ~new_n306;
  assign pv227_21_ = ~new_n309 | ~new_n310;
  assign new_n312 = pv199_1_ & ~pv199_3_;
  assign new_n313 = pv199_3_ & new_n269;
  assign new_n314 = pv194_0_ & new_n288;
  assign new_n315 = ~pv194_0_ & new_n286;
  assign new_n316 = ~new_n314 & ~new_n315;
  assign new_n317 = ~new_n312 & ~new_n313;
  assign pv266_4_ = ~new_n316 | ~new_n317;
  assign new_n319 = pv32_22_ & new_n267;
  assign new_n320 = pv64_22_ & new_n269;
  assign new_n321 = pv96_22_ & new_n271;
  assign new_n322 = ~pv96_22_ & new_n273;
  assign new_n323 = ~new_n321 & ~new_n322;
  assign new_n324 = ~new_n319 & ~new_n320;
  assign pv227_22_ = ~new_n323 | ~new_n324;
  assign new_n326 = pv194_1_ & new_n288;
  assign new_n327 = ~pv194_1_ & new_n286;
  assign new_n328 = ~new_n326 & ~new_n327;
  assign pv266_5_ = ~new_n317 | ~new_n328;
  assign new_n330 = pv32_27_ & new_n267;
  assign new_n331 = pv64_27_ & new_n269;
  assign new_n332 = pv96_27_ & new_n271;
  assign new_n333 = ~pv96_27_ & new_n273;
  assign new_n334 = ~new_n332 & ~new_n333;
  assign new_n335 = ~new_n330 & ~new_n331;
  assign pv227_27_ = ~new_n334 | ~new_n335;
  assign new_n337 = pv199_4_ & ~pv199_0_;
  assign new_n338 = ~pv199_1_ & new_n337;
  assign new_n339 = pv96_28_ & new_n338;
  assign new_n340 = pv199_4_ & pv199_0_;
  assign new_n341 = ~pv199_1_ & new_n340;
  assign new_n342 = pv32_28_ & new_n341;
  assign new_n343 = pv199_1_ & new_n337;
  assign new_n344 = ~pv96_28_ & new_n343;
  assign new_n345 = pv199_1_ & new_n340;
  assign new_n346 = pv64_28_ & new_n345;
  assign new_n347 = ~pv199_4_ & pv199_1_;
  assign new_n348 = ~new_n346 & ~new_n347;
  assign new_n349 = ~new_n339 & ~new_n342;
  assign new_n350 = ~new_n344 & new_n349;
  assign pv259_0_ = ~new_n348 | ~new_n350;
  assign new_n352 = pv32_25_ & new_n267;
  assign new_n353 = pv64_25_ & new_n269;
  assign new_n354 = pv96_25_ & new_n271;
  assign new_n355 = ~pv96_25_ & new_n273;
  assign new_n356 = ~new_n354 & ~new_n355;
  assign new_n357 = ~new_n352 & ~new_n353;
  assign pv227_25_ = ~new_n356 | ~new_n357;
  assign new_n359 = pv96_30_ & new_n338;
  assign new_n360 = pv32_30_ & new_n341;
  assign new_n361 = ~pv96_30_ & new_n343;
  assign new_n362 = pv64_30_ & new_n345;
  assign new_n363 = ~new_n347 & ~new_n362;
  assign new_n364 = ~new_n359 & ~new_n360;
  assign new_n365 = ~new_n361 & new_n364;
  assign pv259_2_ = ~new_n363 | ~new_n365;
  assign new_n367 = pv32_26_ & new_n267;
  assign new_n368 = pv64_26_ & new_n269;
  assign new_n369 = pv96_26_ & new_n271;
  assign new_n370 = ~pv96_26_ & new_n273;
  assign new_n371 = ~new_n369 & ~new_n370;
  assign new_n372 = ~new_n367 & ~new_n368;
  assign pv227_26_ = ~new_n371 | ~new_n372;
  assign new_n374 = pv96_29_ & new_n338;
  assign new_n375 = pv32_29_ & new_n341;
  assign new_n376 = ~pv96_29_ & new_n343;
  assign new_n377 = pv64_29_ & new_n345;
  assign new_n378 = ~new_n347 & ~new_n377;
  assign new_n379 = ~new_n374 & ~new_n375;
  assign new_n380 = ~new_n376 & new_n379;
  assign pv259_1_ = ~new_n378 | ~new_n380;
  assign new_n382 = pv32_7_ & new_n267;
  assign new_n383 = pv64_7_ & new_n269;
  assign new_n384 = pv96_7_ & new_n271;
  assign new_n385 = ~pv96_7_ & new_n273;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = ~new_n382 & ~new_n383;
  assign pv227_7_ = ~new_n386 | ~new_n387;
  assign new_n389 = pv32_18_ & new_n267;
  assign new_n390 = pv64_18_ & new_n269;
  assign new_n391 = pv96_18_ & new_n271;
  assign new_n392 = ~pv96_18_ & new_n273;
  assign new_n393 = ~new_n391 & ~new_n392;
  assign new_n394 = ~new_n389 & ~new_n390;
  assign pv227_18_ = ~new_n393 | ~new_n394;
  assign new_n396 = pv192_13_ & new_n338;
  assign new_n397 = pv128_13_ & new_n341;
  assign new_n398 = ~pv192_13_ & new_n343;
  assign new_n399 = pv160_13_ & new_n345;
  assign new_n400 = ~new_n347 & ~new_n399;
  assign new_n401 = ~new_n396 & ~new_n397;
  assign new_n402 = ~new_n398 & new_n401;
  assign pv259_17_ = ~new_n400 | ~new_n402;
  assign new_n404 = pv32_8_ & new_n267;
  assign new_n405 = pv64_8_ & new_n269;
  assign new_n406 = pv96_8_ & new_n271;
  assign new_n407 = ~pv96_8_ & new_n273;
  assign new_n408 = ~new_n406 & ~new_n407;
  assign new_n409 = ~new_n404 & ~new_n405;
  assign pv227_8_ = ~new_n408 | ~new_n409;
  assign new_n411 = pv32_17_ & new_n267;
  assign new_n412 = pv64_17_ & new_n269;
  assign new_n413 = pv96_17_ & new_n271;
  assign new_n414 = ~pv96_17_ & new_n273;
  assign new_n415 = ~new_n413 & ~new_n414;
  assign new_n416 = ~new_n411 & ~new_n412;
  assign pv227_17_ = ~new_n415 | ~new_n416;
  assign new_n418 = pv192_12_ & new_n338;
  assign new_n419 = pv128_12_ & new_n341;
  assign new_n420 = ~pv192_12_ & new_n343;
  assign new_n421 = pv160_12_ & new_n345;
  assign new_n422 = ~new_n347 & ~new_n421;
  assign new_n423 = ~new_n418 & ~new_n419;
  assign new_n424 = ~new_n420 & new_n423;
  assign pv259_16_ = ~new_n422 | ~new_n424;
  assign new_n426 = pv32_5_ & new_n267;
  assign new_n427 = pv64_5_ & new_n269;
  assign new_n428 = pv96_5_ & new_n271;
  assign new_n429 = ~pv96_5_ & new_n273;
  assign new_n430 = ~new_n428 & ~new_n429;
  assign new_n431 = ~new_n426 & ~new_n427;
  assign pv227_5_ = ~new_n430 | ~new_n431;
  assign new_n433 = pv32_16_ & new_n267;
  assign new_n434 = pv64_16_ & new_n269;
  assign new_n435 = pv96_16_ & new_n271;
  assign new_n436 = ~pv96_16_ & new_n273;
  assign new_n437 = ~new_n435 & ~new_n436;
  assign new_n438 = ~new_n433 & ~new_n434;
  assign pv227_16_ = ~new_n437 | ~new_n438;
  assign new_n440 = pv192_15_ & new_n338;
  assign new_n441 = pv128_15_ & new_n341;
  assign new_n442 = ~pv192_15_ & new_n343;
  assign new_n443 = pv160_15_ & new_n345;
  assign new_n444 = ~new_n347 & ~new_n443;
  assign new_n445 = ~new_n440 & ~new_n441;
  assign new_n446 = ~new_n442 & new_n445;
  assign pv259_19_ = ~new_n444 | ~new_n446;
  assign new_n448 = pv32_6_ & new_n267;
  assign new_n449 = pv64_6_ & new_n269;
  assign new_n450 = pv96_6_ & new_n271;
  assign new_n451 = ~pv96_6_ & new_n273;
  assign new_n452 = ~new_n450 & ~new_n451;
  assign new_n453 = ~new_n448 & ~new_n449;
  assign pv227_6_ = ~new_n452 | ~new_n453;
  assign new_n455 = pv32_15_ & new_n267;
  assign new_n456 = pv64_15_ & new_n269;
  assign new_n457 = pv96_15_ & new_n271;
  assign new_n458 = ~pv96_15_ & new_n273;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = ~new_n455 & ~new_n456;
  assign pv227_15_ = ~new_n459 | ~new_n460;
  assign new_n462 = pv192_14_ & new_n338;
  assign new_n463 = pv128_14_ & new_n341;
  assign new_n464 = ~pv192_14_ & new_n343;
  assign new_n465 = pv160_14_ & new_n345;
  assign new_n466 = ~new_n347 & ~new_n465;
  assign new_n467 = ~new_n462 & ~new_n463;
  assign new_n468 = ~new_n464 & new_n467;
  assign pv259_18_ = ~new_n466 | ~new_n468;
  assign new_n470 = pv32_3_ & new_n267;
  assign new_n471 = pv64_3_ & new_n269;
  assign new_n472 = pv96_3_ & new_n271;
  assign new_n473 = ~pv96_3_ & new_n273;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign new_n475 = ~new_n470 & ~new_n471;
  assign pv227_3_ = ~new_n474 | ~new_n475;
  assign new_n477 = pv32_14_ & new_n267;
  assign new_n478 = pv64_14_ & new_n269;
  assign new_n479 = pv96_14_ & new_n271;
  assign new_n480 = ~pv96_14_ & new_n273;
  assign new_n481 = ~new_n479 & ~new_n480;
  assign new_n482 = ~new_n477 & ~new_n478;
  assign pv227_14_ = ~new_n481 | ~new_n482;
  assign new_n484 = pv192_22_ & new_n338;
  assign new_n485 = pv128_22_ & new_n341;
  assign new_n486 = ~pv192_22_ & new_n343;
  assign new_n487 = pv160_22_ & new_n345;
  assign new_n488 = ~new_n347 & ~new_n487;
  assign new_n489 = ~new_n484 & ~new_n485;
  assign new_n490 = ~new_n486 & new_n489;
  assign pv259_26_ = ~new_n488 | ~new_n490;
  assign new_n492 = pv192_30_ & new_n288;
  assign new_n493 = pv199_0_ & pv199_3_;
  assign new_n494 = ~pv199_1_ & new_n493;
  assign new_n495 = pv128_30_ & new_n494;
  assign new_n496 = ~pv192_30_ & new_n286;
  assign new_n497 = pv160_30_ & new_n313;
  assign new_n498 = ~new_n312 & ~new_n497;
  assign new_n499 = ~new_n492 & ~new_n495;
  assign new_n500 = ~new_n496 & new_n499;
  assign pv266_2_ = ~new_n498 | ~new_n500;
  assign new_n502 = pv32_4_ & new_n267;
  assign new_n503 = pv64_4_ & new_n269;
  assign new_n504 = pv96_4_ & new_n271;
  assign new_n505 = ~pv96_4_ & new_n273;
  assign new_n506 = ~new_n504 & ~new_n505;
  assign new_n507 = ~new_n502 & ~new_n503;
  assign pv227_4_ = ~new_n506 | ~new_n507;
  assign new_n509 = pv32_13_ & new_n267;
  assign new_n510 = pv64_13_ & new_n269;
  assign new_n511 = pv96_13_ & new_n271;
  assign new_n512 = ~pv96_13_ & new_n273;
  assign new_n513 = ~new_n511 & ~new_n512;
  assign new_n514 = ~new_n509 & ~new_n510;
  assign pv227_13_ = ~new_n513 | ~new_n514;
  assign new_n516 = pv32_20_ & new_n267;
  assign new_n517 = pv64_20_ & new_n269;
  assign new_n518 = pv96_20_ & new_n271;
  assign new_n519 = ~pv96_20_ & new_n273;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = ~new_n516 & ~new_n517;
  assign pv227_20_ = ~new_n520 | ~new_n521;
  assign new_n523 = pv192_23_ & new_n338;
  assign new_n524 = pv128_23_ & new_n341;
  assign new_n525 = ~pv192_23_ & new_n343;
  assign new_n526 = pv160_23_ & new_n345;
  assign new_n527 = ~new_n347 & ~new_n526;
  assign new_n528 = ~new_n523 & ~new_n524;
  assign new_n529 = ~new_n525 & new_n528;
  assign pv259_27_ = ~new_n527 | ~new_n529;
  assign new_n531 = pv192_31_ & new_n288;
  assign new_n532 = pv128_31_ & new_n494;
  assign new_n533 = ~pv192_31_ & new_n286;
  assign new_n534 = pv160_31_ & new_n313;
  assign new_n535 = ~new_n312 & ~new_n534;
  assign new_n536 = ~new_n531 & ~new_n532;
  assign new_n537 = ~new_n533 & new_n536;
  assign pv266_3_ = ~new_n535 | ~new_n537;
  assign new_n539 = pv32_1_ & new_n267;
  assign new_n540 = pv64_1_ & new_n269;
  assign new_n541 = pv96_1_ & new_n271;
  assign new_n542 = ~pv96_1_ & new_n273;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign new_n544 = ~new_n539 & ~new_n540;
  assign pv227_1_ = ~new_n543 | ~new_n544;
  assign new_n546 = pv32_12_ & new_n267;
  assign new_n547 = pv64_12_ & new_n269;
  assign new_n548 = pv96_12_ & new_n271;
  assign new_n549 = ~pv96_12_ & new_n273;
  assign new_n550 = ~new_n548 & ~new_n549;
  assign new_n551 = ~new_n546 & ~new_n547;
  assign pv227_12_ = ~new_n550 | ~new_n551;
  assign new_n553 = pv192_24_ & new_n338;
  assign new_n554 = pv128_24_ & new_n341;
  assign new_n555 = ~pv192_24_ & new_n343;
  assign new_n556 = pv160_24_ & new_n345;
  assign new_n557 = ~new_n347 & ~new_n556;
  assign new_n558 = ~new_n553 & ~new_n554;
  assign new_n559 = ~new_n555 & new_n558;
  assign pv259_28_ = ~new_n557 | ~new_n559;
  assign new_n561 = pv192_28_ & new_n288;
  assign new_n562 = pv128_28_ & new_n494;
  assign new_n563 = ~pv192_28_ & new_n286;
  assign new_n564 = pv160_28_ & new_n313;
  assign new_n565 = ~new_n312 & ~new_n564;
  assign new_n566 = ~new_n561 & ~new_n562;
  assign new_n567 = ~new_n563 & new_n566;
  assign pv266_0_ = ~new_n565 | ~new_n567;
  assign new_n569 = pv32_2_ & new_n267;
  assign new_n570 = pv64_2_ & new_n269;
  assign new_n571 = pv96_2_ & new_n271;
  assign new_n572 = ~pv96_2_ & new_n273;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = ~new_n569 & ~new_n570;
  assign pv227_2_ = ~new_n573 | ~new_n574;
  assign new_n576 = pv32_11_ & new_n267;
  assign new_n577 = pv64_11_ & new_n269;
  assign new_n578 = pv96_11_ & new_n271;
  assign new_n579 = ~pv96_11_ & new_n273;
  assign new_n580 = ~new_n578 & ~new_n579;
  assign new_n581 = ~new_n576 & ~new_n577;
  assign pv227_11_ = ~new_n580 | ~new_n581;
  assign new_n583 = pv192_25_ & new_n338;
  assign new_n584 = pv128_25_ & new_n341;
  assign new_n585 = ~pv192_25_ & new_n343;
  assign new_n586 = pv160_25_ & new_n345;
  assign new_n587 = ~new_n347 & ~new_n586;
  assign new_n588 = ~new_n583 & ~new_n584;
  assign new_n589 = ~new_n585 & new_n588;
  assign pv259_29_ = ~new_n587 | ~new_n589;
  assign new_n591 = pv192_29_ & new_n288;
  assign new_n592 = pv128_29_ & new_n494;
  assign new_n593 = ~pv192_29_ & new_n286;
  assign new_n594 = pv160_29_ & new_n313;
  assign new_n595 = ~new_n312 & ~new_n594;
  assign new_n596 = ~new_n591 & ~new_n592;
  assign new_n597 = ~new_n593 & new_n596;
  assign pv266_1_ = ~new_n595 | ~new_n597;
  assign new_n599 = pv192_18_ & new_n338;
  assign new_n600 = pv128_18_ & new_n341;
  assign new_n601 = ~pv192_18_ & new_n343;
  assign new_n602 = pv160_18_ & new_n345;
  assign new_n603 = ~new_n347 & ~new_n602;
  assign new_n604 = ~new_n599 & ~new_n600;
  assign new_n605 = ~new_n601 & new_n604;
  assign pv259_22_ = ~new_n603 | ~new_n605;
  assign new_n607 = pv192_19_ & new_n338;
  assign new_n608 = pv128_19_ & new_n341;
  assign new_n609 = ~pv192_19_ & new_n343;
  assign new_n610 = pv160_19_ & new_n345;
  assign new_n611 = ~new_n347 & ~new_n610;
  assign new_n612 = ~new_n607 & ~new_n608;
  assign new_n613 = ~new_n609 & new_n612;
  assign pv259_23_ = ~new_n611 | ~new_n613;
  assign new_n615 = pv192_7_ & new_n338;
  assign new_n616 = pv128_7_ & new_n341;
  assign new_n617 = ~pv192_7_ & new_n343;
  assign new_n618 = pv160_7_ & new_n345;
  assign new_n619 = ~new_n347 & ~new_n618;
  assign new_n620 = ~new_n615 & ~new_n616;
  assign new_n621 = ~new_n617 & new_n620;
  assign pv259_11_ = ~new_n619 | ~new_n621;
  assign new_n623 = pv192_20_ & new_n338;
  assign new_n624 = pv128_20_ & new_n341;
  assign new_n625 = ~pv192_20_ & new_n343;
  assign new_n626 = pv160_20_ & new_n345;
  assign new_n627 = ~new_n347 & ~new_n626;
  assign new_n628 = ~new_n623 & ~new_n624;
  assign new_n629 = ~new_n625 & new_n628;
  assign pv259_24_ = ~new_n627 | ~new_n629;
  assign new_n631 = pv192_6_ & new_n338;
  assign new_n632 = pv128_6_ & new_n341;
  assign new_n633 = ~pv192_6_ & new_n343;
  assign new_n634 = pv160_6_ & new_n345;
  assign new_n635 = ~new_n347 & ~new_n634;
  assign new_n636 = ~new_n631 & ~new_n632;
  assign new_n637 = ~new_n633 & new_n636;
  assign pv259_10_ = ~new_n635 | ~new_n637;
  assign new_n639 = pv192_21_ & new_n338;
  assign new_n640 = pv128_21_ & new_n341;
  assign new_n641 = ~pv192_21_ & new_n343;
  assign new_n642 = pv160_21_ & new_n345;
  assign new_n643 = ~new_n347 & ~new_n642;
  assign new_n644 = ~new_n639 & ~new_n640;
  assign new_n645 = ~new_n641 & new_n644;
  assign pv259_25_ = ~new_n643 | ~new_n645;
  assign new_n647 = pv192_9_ & new_n338;
  assign new_n648 = pv128_9_ & new_n341;
  assign new_n649 = ~pv192_9_ & new_n343;
  assign new_n650 = pv160_9_ & new_n345;
  assign new_n651 = ~new_n347 & ~new_n650;
  assign new_n652 = ~new_n647 & ~new_n648;
  assign new_n653 = ~new_n649 & new_n652;
  assign pv259_13_ = ~new_n651 | ~new_n653;
  assign new_n655 = pv192_27_ & new_n338;
  assign new_n656 = pv128_27_ & new_n341;
  assign new_n657 = ~pv192_27_ & new_n343;
  assign new_n658 = pv160_27_ & new_n345;
  assign new_n659 = ~new_n347 & ~new_n658;
  assign new_n660 = ~new_n655 & ~new_n656;
  assign new_n661 = ~new_n657 & new_n660;
  assign pv259_31_ = ~new_n659 | ~new_n661;
  assign new_n663 = pv192_8_ & new_n338;
  assign new_n664 = pv128_8_ & new_n341;
  assign new_n665 = ~pv192_8_ & new_n343;
  assign new_n666 = pv160_8_ & new_n345;
  assign new_n667 = ~new_n347 & ~new_n666;
  assign new_n668 = ~new_n663 & ~new_n664;
  assign new_n669 = ~new_n665 & new_n668;
  assign pv259_12_ = ~new_n667 | ~new_n669;
  assign new_n671 = pv192_26_ & new_n338;
  assign new_n672 = pv128_26_ & new_n341;
  assign new_n673 = ~pv192_26_ & new_n343;
  assign new_n674 = pv160_26_ & new_n345;
  assign new_n675 = ~new_n347 & ~new_n674;
  assign new_n676 = ~new_n671 & ~new_n672;
  assign new_n677 = ~new_n673 & new_n676;
  assign pv259_30_ = ~new_n675 | ~new_n677;
  assign new_n679 = pv32_9_ & new_n267;
  assign new_n680 = pv64_9_ & new_n269;
  assign new_n681 = pv96_9_ & new_n271;
  assign new_n682 = ~pv96_9_ & new_n273;
  assign new_n683 = ~new_n681 & ~new_n682;
  assign new_n684 = ~new_n679 & ~new_n680;
  assign pv227_9_ = ~new_n683 | ~new_n684;
  assign new_n686 = pv192_11_ & new_n338;
  assign new_n687 = pv128_11_ & new_n341;
  assign new_n688 = ~pv192_11_ & new_n343;
  assign new_n689 = pv160_11_ & new_n345;
  assign new_n690 = ~new_n347 & ~new_n689;
  assign new_n691 = ~new_n686 & ~new_n687;
  assign new_n692 = ~new_n688 & new_n691;
  assign pv259_15_ = ~new_n690 | ~new_n692;
  assign new_n694 = pv192_16_ & new_n338;
  assign new_n695 = pv128_16_ & new_n341;
  assign new_n696 = ~pv192_16_ & new_n343;
  assign new_n697 = pv160_16_ & new_n345;
  assign new_n698 = ~new_n347 & ~new_n697;
  assign new_n699 = ~new_n694 & ~new_n695;
  assign new_n700 = ~new_n696 & new_n699;
  assign pv259_20_ = ~new_n698 | ~new_n700;
  assign new_n702 = pv32_19_ & new_n267;
  assign new_n703 = pv64_19_ & new_n269;
  assign new_n704 = pv96_19_ & new_n271;
  assign new_n705 = ~pv96_19_ & new_n273;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = ~new_n702 & ~new_n703;
  assign pv227_19_ = ~new_n706 | ~new_n707;
  assign new_n709 = pv192_10_ & new_n338;
  assign new_n710 = pv128_10_ & new_n341;
  assign new_n711 = ~pv192_10_ & new_n343;
  assign new_n712 = pv160_10_ & new_n345;
  assign new_n713 = ~new_n347 & ~new_n712;
  assign new_n714 = ~new_n709 & ~new_n710;
  assign new_n715 = ~new_n711 & new_n714;
  assign pv259_14_ = ~new_n713 | ~new_n715;
  assign new_n717 = pv192_17_ & new_n338;
  assign new_n718 = pv128_17_ & new_n341;
  assign new_n719 = ~pv192_17_ & new_n343;
  assign new_n720 = pv160_17_ & new_n345;
  assign new_n721 = ~new_n347 & ~new_n720;
  assign new_n722 = ~new_n717 & ~new_n718;
  assign new_n723 = ~new_n719 & new_n722;
  assign pv259_21_ = ~new_n721 | ~new_n723;
  assign new_n725 = pv192_0_ & new_n338;
  assign new_n726 = pv128_0_ & new_n341;
  assign new_n727 = ~pv192_0_ & new_n343;
  assign new_n728 = pv160_0_ & new_n345;
  assign new_n729 = ~new_n347 & ~new_n728;
  assign new_n730 = ~new_n725 & ~new_n726;
  assign new_n731 = ~new_n727 & new_n730;
  assign pv259_4_ = ~new_n729 | ~new_n731;
  assign new_n733 = pv96_31_ & new_n338;
  assign new_n734 = pv32_31_ & new_n341;
  assign new_n735 = ~pv96_31_ & new_n343;
  assign new_n736 = pv64_31_ & new_n345;
  assign new_n737 = ~new_n347 & ~new_n736;
  assign new_n738 = ~new_n733 & ~new_n734;
  assign new_n739 = ~new_n735 & new_n738;
  assign pv259_3_ = ~new_n737 | ~new_n739;
  assign new_n741 = pv192_2_ & new_n338;
  assign new_n742 = pv128_2_ & new_n341;
  assign new_n743 = ~pv192_2_ & new_n343;
  assign new_n744 = pv160_2_ & new_n345;
  assign new_n745 = ~new_n347 & ~new_n744;
  assign new_n746 = ~new_n741 & ~new_n742;
  assign new_n747 = ~new_n743 & new_n746;
  assign pv259_6_ = ~new_n745 | ~new_n747;
  assign new_n749 = pv192_1_ & new_n338;
  assign new_n750 = pv128_1_ & new_n341;
  assign new_n751 = ~pv192_1_ & new_n343;
  assign new_n752 = pv160_1_ & new_n345;
  assign new_n753 = ~new_n347 & ~new_n752;
  assign new_n754 = ~new_n749 & ~new_n750;
  assign new_n755 = ~new_n751 & new_n754;
  assign pv259_5_ = ~new_n753 | ~new_n755;
  assign new_n757 = pv192_4_ & new_n338;
  assign new_n758 = pv128_4_ & new_n341;
  assign new_n759 = ~pv192_4_ & new_n343;
  assign new_n760 = pv160_4_ & new_n345;
  assign new_n761 = ~new_n347 & ~new_n760;
  assign new_n762 = ~new_n757 & ~new_n758;
  assign new_n763 = ~new_n759 & new_n762;
  assign pv259_8_ = ~new_n761 | ~new_n763;
  assign new_n765 = pv192_3_ & new_n338;
  assign new_n766 = pv128_3_ & new_n341;
  assign new_n767 = ~pv192_3_ & new_n343;
  assign new_n768 = pv160_3_ & new_n345;
  assign new_n769 = ~new_n347 & ~new_n768;
  assign new_n770 = ~new_n765 & ~new_n766;
  assign new_n771 = ~new_n767 & new_n770;
  assign pv259_7_ = ~new_n769 | ~new_n771;
  assign new_n773 = pv192_5_ & new_n338;
  assign new_n774 = pv128_5_ & new_n341;
  assign new_n775 = ~pv192_5_ & new_n343;
  assign new_n776 = pv160_5_ & new_n345;
  assign new_n777 = ~new_n347 & ~new_n776;
  assign new_n778 = ~new_n773 & ~new_n774;
  assign new_n779 = ~new_n775 & new_n778;
  assign pv259_9_ = ~new_n777 | ~new_n779;
endmodule


