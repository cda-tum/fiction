// Benchmark "top" written by ABC on Mon Feb 19 11:52:45 2024

module top ( 
    pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, ph0, px,
    pi0, py, pj0, pz, pk0, pl0, pm0, pa, pb, pc, pd, pe, pf, pg, ph, pi,
    pj, pk, pl, pm, pn, po,
    pn0, po0, pp0  );
  input  pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw,
    ph0, px, pi0, py, pj0, pz, pk0, pl0, pm0, pa, pb, pc, pd, pe, pf, pg,
    ph, pi, pj, pk, pl, pm, pn, po;
  output pn0, po0, pp0;
  wire new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48,
    new_n49, new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56,
    new_n57, new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64,
    new_n65, new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72,
    new_n73, new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1454, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2715,
    new_n2716, new_n2717, new_n2718, new_n2719, new_n2720, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2830, new_n2831, new_n2832, new_n2833, new_n2834, new_n2835,
    new_n2836, new_n2837, new_n2838, new_n2839, new_n2840, new_n2841,
    new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847,
    new_n2848, new_n2849, new_n2850, new_n2851, new_n2852, new_n2853,
    new_n2854, new_n2855, new_n2856, new_n2857, new_n2858, new_n2859,
    new_n2860, new_n2861, new_n2862, new_n2863, new_n2864, new_n2865,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040,
    new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046,
    new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052,
    new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058,
    new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064,
    new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070,
    new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076,
    new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082,
    new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088,
    new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112,
    new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118,
    new_n3119, new_n3120, new_n3121, new_n3122, new_n3123, new_n3124,
    new_n3125, new_n3126, new_n3127, new_n3128, new_n3129, new_n3130,
    new_n3131, new_n3132, new_n3133, new_n3134, new_n3135, new_n3136,
    new_n3137, new_n3138, new_n3139, new_n3140, new_n3141, new_n3142,
    new_n3143, new_n3144, new_n3145, new_n3146, new_n3147, new_n3148,
    new_n3149, new_n3150, new_n3151, new_n3152, new_n3153, new_n3154,
    new_n3155, new_n3156, new_n3157, new_n3158, new_n3159, new_n3160,
    new_n3161, new_n3162, new_n3163, new_n3164, new_n3165, new_n3166,
    new_n3167, new_n3168, new_n3169, new_n3170, new_n3171, new_n3172,
    new_n3173, new_n3174, new_n3175, new_n3176, new_n3177, new_n3178,
    new_n3179, new_n3180, new_n3181, new_n3182, new_n3183, new_n3184,
    new_n3185, new_n3186, new_n3187, new_n3188, new_n3189, new_n3190,
    new_n3191, new_n3192, new_n3193, new_n3194, new_n3195, new_n3196,
    new_n3197, new_n3198, new_n3199, new_n3200, new_n3201, new_n3202,
    new_n3203, new_n3204, new_n3205, new_n3206, new_n3207, new_n3208,
    new_n3209, new_n3210, new_n3211, new_n3212, new_n3213, new_n3214,
    new_n3215, new_n3216, new_n3217, new_n3218, new_n3219, new_n3220,
    new_n3221, new_n3222, new_n3223, new_n3224, new_n3225, new_n3226,
    new_n3227, new_n3228, new_n3229, new_n3230, new_n3231, new_n3232,
    new_n3233, new_n3234, new_n3235, new_n3236, new_n3237, new_n3238,
    new_n3239, new_n3240, new_n3241, new_n3242, new_n3243, new_n3244,
    new_n3245, new_n3246, new_n3247, new_n3248, new_n3249, new_n3250,
    new_n3251, new_n3252, new_n3253, new_n3254, new_n3255, new_n3256,
    new_n3257, new_n3258, new_n3259, new_n3260, new_n3261, new_n3262,
    new_n3263, new_n3264, new_n3265, new_n3266, new_n3267, new_n3268,
    new_n3269, new_n3270, new_n3271, new_n3272, new_n3273, new_n3274,
    new_n3275, new_n3276, new_n3277, new_n3278, new_n3279, new_n3280,
    new_n3281, new_n3282, new_n3283, new_n3284, new_n3285, new_n3286,
    new_n3287, new_n3288, new_n3289, new_n3290, new_n3291, new_n3292,
    new_n3293, new_n3294, new_n3295, new_n3296, new_n3297, new_n3298,
    new_n3299, new_n3300, new_n3301, new_n3302, new_n3303, new_n3304,
    new_n3305, new_n3306, new_n3307, new_n3308, new_n3309, new_n3310,
    new_n3311, new_n3312, new_n3313, new_n3314, new_n3315, new_n3316,
    new_n3317, new_n3318, new_n3319, new_n3320, new_n3321, new_n3322,
    new_n3323, new_n3324, new_n3325, new_n3326, new_n3327, new_n3328,
    new_n3329, new_n3330, new_n3331, new_n3332, new_n3333, new_n3334,
    new_n3335, new_n3336, new_n3337, new_n3338, new_n3339, new_n3340,
    new_n3341, new_n3342, new_n3343, new_n3344, new_n3345, new_n3346,
    new_n3347, new_n3348, new_n3349, new_n3350, new_n3351, new_n3352,
    new_n3353, new_n3354, new_n3355, new_n3356, new_n3357, new_n3358,
    new_n3359, new_n3360, new_n3361, new_n3362, new_n3363, new_n3364,
    new_n3365, new_n3366, new_n3367, new_n3368, new_n3369, new_n3370,
    new_n3371, new_n3372, new_n3373, new_n3374, new_n3375, new_n3376,
    new_n3377, new_n3378, new_n3379, new_n3380, new_n3381, new_n3382,
    new_n3383, new_n3384, new_n3385, new_n3386, new_n3387, new_n3388,
    new_n3389, new_n3390, new_n3391, new_n3392, new_n3393, new_n3394,
    new_n3395, new_n3396, new_n3397, new_n3398, new_n3399, new_n3400,
    new_n3401, new_n3402, new_n3403, new_n3404, new_n3405, new_n3406,
    new_n3407, new_n3408, new_n3409, new_n3410, new_n3411, new_n3412,
    new_n3413, new_n3414, new_n3415, new_n3416, new_n3417, new_n3418,
    new_n3419, new_n3420, new_n3421, new_n3422, new_n3423, new_n3424,
    new_n3425, new_n3426, new_n3427, new_n3428, new_n3429, new_n3430,
    new_n3431, new_n3432, new_n3433, new_n3434, new_n3435, new_n3436,
    new_n3437, new_n3438, new_n3439, new_n3440, new_n3441, new_n3442,
    new_n3443, new_n3444, new_n3445, new_n3446, new_n3447, new_n3448,
    new_n3449, new_n3450, new_n3451, new_n3452, new_n3453, new_n3454,
    new_n3455, new_n3456, new_n3457, new_n3458, new_n3459, new_n3460,
    new_n3461, new_n3462, new_n3463, new_n3464, new_n3465, new_n3466,
    new_n3467, new_n3468, new_n3469, new_n3470, new_n3471, new_n3472,
    new_n3473, new_n3474, new_n3475, new_n3476, new_n3477, new_n3478,
    new_n3479, new_n3480, new_n3481, new_n3482, new_n3483, new_n3484,
    new_n3485, new_n3486, new_n3487, new_n3488, new_n3489, new_n3490,
    new_n3491, new_n3492, new_n3493, new_n3494, new_n3495, new_n3496,
    new_n3497, new_n3498, new_n3499, new_n3500, new_n3501, new_n3502,
    new_n3503, new_n3504, new_n3505, new_n3506, new_n3507, new_n3508,
    new_n3509, new_n3510, new_n3511, new_n3512, new_n3513, new_n3514,
    new_n3515, new_n3516, new_n3517, new_n3518, new_n3519, new_n3520,
    new_n3521, new_n3522, new_n3523, new_n3524, new_n3525, new_n3526,
    new_n3527, new_n3528, new_n3529, new_n3530, new_n3531, new_n3532,
    new_n3533, new_n3534, new_n3535, new_n3536, new_n3537, new_n3538,
    new_n3539, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544,
    new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550,
    new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556,
    new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562,
    new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568,
    new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574,
    new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580,
    new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586,
    new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592,
    new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598,
    new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604,
    new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610,
    new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616,
    new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300,
    new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306,
    new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312,
    new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318,
    new_n4319, new_n4320, new_n4321, new_n4322, new_n4323, new_n4324,
    new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330,
    new_n4331, new_n4332, new_n4333, new_n4334, new_n4335, new_n4336,
    new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342,
    new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414,
    new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420,
    new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426,
    new_n4427, new_n4428, new_n4429, new_n4430, new_n4431, new_n4432,
    new_n4433, new_n4434, new_n4435, new_n4436, new_n4437, new_n4438,
    new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444,
    new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450,
    new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456,
    new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462,
    new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468,
    new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474,
    new_n4475, new_n4476, new_n4477, new_n4478, new_n4479, new_n4480,
    new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486,
    new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492,
    new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498,
    new_n4499, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504,
    new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510,
    new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516,
    new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522,
    new_n4523, new_n4524, new_n4525, new_n4526, new_n4527, new_n4528,
    new_n4529, new_n4530, new_n4531, new_n4532, new_n4533, new_n4534,
    new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540,
    new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546,
    new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4552,
    new_n4553, new_n4554, new_n4555, new_n4556, new_n4557, new_n4558,
    new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564,
    new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570,
    new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576,
    new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582,
    new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588,
    new_n4589, new_n4590, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4634, new_n4635, new_n4636,
    new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642,
    new_n4643, new_n4644, new_n4645, new_n4646, new_n4647, new_n4648,
    new_n4649, new_n4650, new_n4651, new_n4652, new_n4653, new_n4654,
    new_n4655, new_n4656, new_n4657, new_n4658, new_n4659, new_n4660,
    new_n4661, new_n4662, new_n4663, new_n4664, new_n4665, new_n4666,
    new_n4667, new_n4668, new_n4669, new_n4670, new_n4671, new_n4672,
    new_n4673, new_n4674, new_n4675, new_n4676, new_n4677, new_n4678,
    new_n4679, new_n4680, new_n4681, new_n4682, new_n4683, new_n4684,
    new_n4685, new_n4686, new_n4687, new_n4688, new_n4689, new_n4690,
    new_n4691, new_n4692, new_n4693, new_n4694, new_n4695, new_n4696,
    new_n4697, new_n4698, new_n4699, new_n4700, new_n4701, new_n4702,
    new_n4703, new_n4704, new_n4705, new_n4706, new_n4707, new_n4708,
    new_n4709, new_n4710, new_n4711, new_n4712, new_n4713, new_n4714,
    new_n4715, new_n4716, new_n4717, new_n4718, new_n4719, new_n4720,
    new_n4721, new_n4722, new_n4723, new_n4724, new_n4725, new_n4726,
    new_n4727, new_n4728, new_n4729, new_n4730, new_n4731, new_n4732,
    new_n4733, new_n4734, new_n4735, new_n4736, new_n4737, new_n4738,
    new_n4739, new_n4740, new_n4741, new_n4742, new_n4743, new_n4744,
    new_n4745, new_n4746, new_n4747, new_n4748, new_n4749, new_n4750,
    new_n4751, new_n4752, new_n4753, new_n4754, new_n4755, new_n4756,
    new_n4757, new_n4758, new_n4759, new_n4760, new_n4761, new_n4762,
    new_n4763, new_n4764, new_n4765, new_n4766, new_n4767, new_n4768,
    new_n4769, new_n4770, new_n4771, new_n4772, new_n4773, new_n4774,
    new_n4775, new_n4776, new_n4777, new_n4778, new_n4779, new_n4780,
    new_n4781, new_n4782, new_n4783, new_n4784, new_n4785, new_n4786,
    new_n4787, new_n4788, new_n4789, new_n4790, new_n4791, new_n4792,
    new_n4793, new_n4794, new_n4795, new_n4796, new_n4797, new_n4798,
    new_n4799, new_n4800, new_n4801, new_n4802, new_n4803, new_n4804,
    new_n4805, new_n4806, new_n4807, new_n4808, new_n4809, new_n4810,
    new_n4811, new_n4812, new_n4813, new_n4814, new_n4815, new_n4816,
    new_n4817, new_n4818, new_n4819, new_n4820, new_n4821, new_n4822,
    new_n4823, new_n4824, new_n4825, new_n4826, new_n4827, new_n4828,
    new_n4829, new_n4830, new_n4831, new_n4832, new_n4833, new_n4834,
    new_n4835, new_n4836, new_n4837, new_n4838, new_n4839, new_n4840,
    new_n4841, new_n4842, new_n4843, new_n4844, new_n4845, new_n4846,
    new_n4847, new_n4848, new_n4849, new_n4850, new_n4851, new_n4852,
    new_n4853, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858,
    new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723,
    new_n5724, new_n5725, new_n5726, new_n5727, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822, new_n5823, new_n5824, new_n5825,
    new_n5826, new_n5827, new_n5828, new_n5829, new_n5830, new_n5831,
    new_n5832, new_n5833, new_n5834, new_n5835, new_n5836, new_n5837,
    new_n5838, new_n5839, new_n5840, new_n5841, new_n5842, new_n5843,
    new_n5844, new_n5845, new_n5846, new_n5847, new_n5848, new_n5849,
    new_n5850, new_n5851, new_n5852, new_n5853, new_n5854, new_n5855,
    new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861,
    new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867,
    new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5881, new_n5882, new_n5883, new_n5884, new_n5885,
    new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903,
    new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273, new_n6274, new_n6275,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6293,
    new_n6294, new_n6295, new_n6296, new_n6297, new_n6298, new_n6299,
    new_n6300, new_n6301, new_n6302, new_n6303, new_n6304, new_n6305,
    new_n6306, new_n6307, new_n6308, new_n6309, new_n6310, new_n6311,
    new_n6312, new_n6313, new_n6314, new_n6315, new_n6316, new_n6317,
    new_n6318, new_n6319, new_n6320, new_n6321, new_n6322, new_n6323,
    new_n6324, new_n6325, new_n6326, new_n6327, new_n6328, new_n6329,
    new_n6330, new_n6331, new_n6332, new_n6333, new_n6334, new_n6335,
    new_n6336, new_n6337, new_n6338, new_n6339, new_n6340, new_n6341,
    new_n6342, new_n6343, new_n6344, new_n6345, new_n6346, new_n6347,
    new_n6348, new_n6349, new_n6350, new_n6351, new_n6352, new_n6353,
    new_n6354, new_n6355, new_n6356, new_n6357, new_n6358, new_n6359,
    new_n6360, new_n6361, new_n6362, new_n6363, new_n6364, new_n6365,
    new_n6366, new_n6367, new_n6368, new_n6369, new_n6370, new_n6371,
    new_n6372, new_n6373, new_n6374, new_n6375, new_n6376, new_n6377,
    new_n6378, new_n6379, new_n6380, new_n6381, new_n6382, new_n6383,
    new_n6384, new_n6385, new_n6386, new_n6387, new_n6388, new_n6389,
    new_n6390, new_n6391, new_n6392, new_n6393, new_n6394, new_n6395,
    new_n6396, new_n6397, new_n6398, new_n6399, new_n6400, new_n6401,
    new_n6402, new_n6403, new_n6404, new_n6405, new_n6406, new_n6407,
    new_n6408, new_n6409, new_n6410, new_n6411, new_n6412, new_n6413,
    new_n6414, new_n6415, new_n6416, new_n6417, new_n6418, new_n6419,
    new_n6420, new_n6421, new_n6422, new_n6423, new_n6424, new_n6425,
    new_n6426, new_n6427, new_n6428, new_n6429, new_n6430, new_n6431,
    new_n6432, new_n6433, new_n6434, new_n6435, new_n6436, new_n6437,
    new_n6438, new_n6439, new_n6440, new_n6441, new_n6442, new_n6443,
    new_n6444, new_n6445, new_n6446, new_n6447, new_n6448, new_n6449,
    new_n6450, new_n6451, new_n6452, new_n6453, new_n6454, new_n6455,
    new_n6456, new_n6457, new_n6458, new_n6459, new_n6460, new_n6461,
    new_n6462, new_n6463, new_n6464, new_n6465, new_n6466, new_n6467,
    new_n6468, new_n6469, new_n6470, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502, new_n6503,
    new_n6504, new_n6505, new_n6506, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513, new_n6514, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556, new_n6557,
    new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587,
    new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611,
    new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653,
    new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860, new_n6861, new_n6862, new_n6863,
    new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875,
    new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730, new_n7731, new_n7732, new_n7733,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965, new_n7966, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285,
    new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303,
    new_n8304, new_n8305, new_n8306, new_n8307, new_n8308, new_n8309,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927,
    new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933,
    new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939,
    new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945,
    new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951,
    new_n8952, new_n8953, new_n8954, new_n8955, new_n8956, new_n8957,
    new_n8958, new_n8959, new_n8960, new_n8961, new_n8962, new_n8963,
    new_n8964, new_n8965, new_n8966, new_n8967, new_n8968, new_n8969,
    new_n8970, new_n8971, new_n8972, new_n8973, new_n8974, new_n8975,
    new_n8976, new_n8977, new_n8978, new_n8979, new_n8980, new_n8981,
    new_n8982, new_n8983, new_n8984, new_n8985, new_n8986, new_n8987,
    new_n8988, new_n8989, new_n8990, new_n8991, new_n8992, new_n8993,
    new_n8994, new_n8995, new_n8996, new_n8997, new_n8998, new_n8999,
    new_n9000, new_n9001, new_n9002, new_n9003, new_n9004, new_n9005,
    new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011,
    new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017,
    new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023,
    new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077,
    new_n9078, new_n9079, new_n9080, new_n9081, new_n9082, new_n9083,
    new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089,
    new_n9090, new_n9091, new_n9092, new_n9093, new_n9094, new_n9095,
    new_n9096, new_n9097, new_n9098, new_n9099, new_n9100, new_n9101,
    new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107,
    new_n9108, new_n9109, new_n9110, new_n9111, new_n9112, new_n9113,
    new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119,
    new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125,
    new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131,
    new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137,
    new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143,
    new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149,
    new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155,
    new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161,
    new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167,
    new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173,
    new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179,
    new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185,
    new_n9186, new_n9187, new_n9188, new_n9189, new_n9190, new_n9191,
    new_n9192, new_n9193, new_n9194, new_n9195, new_n9196, new_n9197,
    new_n9198, new_n9199, new_n9200, new_n9201, new_n9202, new_n9203,
    new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209,
    new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215,
    new_n9216, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221,
    new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022, new_n10023, new_n10024, new_n10025,
    new_n10026, new_n10027, new_n10028, new_n10029, new_n10030, new_n10031,
    new_n10032, new_n10033, new_n10034, new_n10035, new_n10036, new_n10037,
    new_n10038, new_n10039, new_n10040, new_n10041, new_n10042, new_n10043,
    new_n10044, new_n10045, new_n10046, new_n10047, new_n10048, new_n10049,
    new_n10050, new_n10051, new_n10052, new_n10053, new_n10054, new_n10055,
    new_n10056, new_n10057, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127,
    new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133,
    new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139,
    new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145,
    new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151,
    new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163,
    new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236, new_n10237, new_n10238, new_n10239, new_n10240, new_n10241,
    new_n10242, new_n10243, new_n10244, new_n10245, new_n10246, new_n10247,
    new_n10248, new_n10249, new_n10250, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261, new_n10262, new_n10263, new_n10264, new_n10265,
    new_n10266, new_n10267, new_n10268, new_n10269, new_n10270, new_n10271,
    new_n10272, new_n10273, new_n10274, new_n10275, new_n10276, new_n10277,
    new_n10278, new_n10279, new_n10280, new_n10281, new_n10282, new_n10283,
    new_n10284, new_n10285, new_n10286, new_n10287, new_n10288, new_n10289,
    new_n10290, new_n10291, new_n10292, new_n10293, new_n10294, new_n10295,
    new_n10296, new_n10297, new_n10298, new_n10299, new_n10300, new_n10301,
    new_n10302, new_n10303, new_n10304, new_n10305, new_n10306, new_n10307,
    new_n10308, new_n10309, new_n10310, new_n10311, new_n10312, new_n10313,
    new_n10314, new_n10315, new_n10316, new_n10317, new_n10318, new_n10319,
    new_n10320, new_n10321, new_n10322, new_n10323, new_n10324, new_n10325,
    new_n10326, new_n10327, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376;
  assign new_n42 = ~pj & pn;
  assign new_n43 = ~pf & new_n42;
  assign new_n44 = ~pg & new_n43;
  assign new_n45 = ~pe & new_n44;
  assign new_n46 = ~pa0 & new_n45;
  assign new_n47 = ~po & new_n46;
  assign new_n48 = pk0 & new_n47;
  assign new_n49 = ~pg0 & new_n48;
  assign new_n50 = ~pv & new_n49;
  assign new_n51 = ~py & new_n50;
  assign new_n52 = pd0 & new_n51;
  assign new_n53 = ~pj0 & new_n52;
  assign new_n54 = ~pc0 & new_n53;
  assign new_n55 = ~px & new_n54;
  assign new_n56 = ~pb0 & new_n55;
  assign new_n57 = ~pq & new_n56;
  assign new_n58 = ~pr & new_n57;
  assign new_n59 = ~pg & ~ph;
  assign new_n60 = ~pe & new_n59;
  assign new_n61 = ~pf & new_n60;
  assign new_n62 = ~pc & new_n61;
  assign new_n63 = pk0 & new_n62;
  assign new_n64 = ~po & new_n63;
  assign new_n65 = ~pc0 & new_n64;
  assign new_n66 = ~pd0 & new_n65;
  assign new_n67 = ~pi0 & new_n66;
  assign new_n68 = pj0 & new_n67;
  assign new_n69 = ~px & new_n68;
  assign new_n70 = ~pb0 & new_n69;
  assign new_n71 = ~pr & new_n70;
  assign new_n72 = pn & new_n71;
  assign new_n73 = ~pq & new_n72;
  assign new_n74 = ~pi & new_n73;
  assign new_n75 = ~pj & new_n74;
  assign new_n76 = ~pg & ~pn;
  assign new_n77 = ~pe & new_n76;
  assign new_n78 = ~pf & new_n77;
  assign new_n79 = ~pc & new_n78;
  assign new_n80 = ~pm & new_n79;
  assign new_n81 = pk0 & new_n80;
  assign new_n82 = ~pg0 & new_n81;
  assign new_n83 = ~py & new_n82;
  assign new_n84 = ~pf0 & new_n83;
  assign new_n85 = pi0 & new_n84;
  assign new_n86 = ~pj0 & new_n85;
  assign new_n87 = ~pd0 & new_n86;
  assign new_n88 = ~pb0 & new_n87;
  assign new_n89 = ~pc0 & new_n88;
  assign new_n90 = ~pq & new_n89;
  assign new_n91 = ~px & new_n90;
  assign new_n92 = ~px & pz;
  assign new_n93 = ~pq & new_n92;
  assign new_n94 = ~pr & new_n93;
  assign new_n95 = ~po & new_n94;
  assign new_n96 = pj0 & new_n95;
  assign new_n97 = ~pi0 & new_n96;
  assign new_n98 = ~pd0 & new_n97;
  assign new_n99 = ph0 & new_n98;
  assign new_n100 = ~pb0 & new_n99;
  assign new_n101 = ~pc0 & new_n100;
  assign new_n102 = ~pi & ~pj;
  assign new_n103 = ~pf & new_n102;
  assign new_n104 = ~pg & new_n103;
  assign new_n105 = ~pe & new_n104;
  assign new_n106 = ~pa0 & new_n105;
  assign new_n107 = ~pk & new_n106;
  assign new_n108 = ~pj0 & new_n107;
  assign new_n109 = pk0 & new_n108;
  assign new_n110 = ~pv & new_n109;
  assign new_n111 = ~py & new_n110;
  assign new_n112 = ~pc0 & new_n111;
  assign new_n113 = pd0 & new_n112;
  assign new_n114 = ~pb0 & new_n113;
  assign new_n115 = ~pr & new_n114;
  assign new_n116 = ~px & new_n115;
  assign new_n117 = ~pn & new_n116;
  assign new_n118 = ~pq & new_n117;
  assign new_n119 = ~pq & ~px;
  assign new_n120 = ~pf & new_n119;
  assign new_n121 = ~pg & new_n120;
  assign new_n122 = ~pe & new_n121;
  assign new_n123 = ~pm & new_n122;
  assign new_n124 = ~py & new_n123;
  assign new_n125 = ~pa0 & new_n124;
  assign new_n126 = ~po & new_n125;
  assign new_n127 = ~pf0 & new_n126;
  assign new_n128 = ~pg0 & new_n127;
  assign new_n129 = ~pv & new_n128;
  assign new_n130 = pk0 & new_n129;
  assign new_n131 = pd0 & new_n130;
  assign new_n132 = ~pj0 & new_n131;
  assign new_n133 = ~pb0 & new_n132;
  assign new_n134 = ~pc0 & new_n133;
  assign new_n135 = ~pg & ~pi;
  assign new_n136 = ~pe & new_n135;
  assign new_n137 = ~pf & new_n136;
  assign new_n138 = ~pc & new_n137;
  assign new_n139 = ~pm & new_n138;
  assign new_n140 = pk0 & new_n139;
  assign new_n141 = ~py & new_n140;
  assign new_n142 = ~pa0 & new_n141;
  assign new_n143 = ~pf0 & new_n142;
  assign new_n144 = ~pd0 & new_n143;
  assign new_n145 = ~pj0 & new_n144;
  assign new_n146 = ~pc0 & new_n145;
  assign new_n147 = ~px & new_n146;
  assign new_n148 = ~pb0 & new_n147;
  assign new_n149 = ~pn & new_n148;
  assign new_n150 = ~pq & new_n149;
  assign new_n151 = pu & ~pv;
  assign new_n152 = ~po & new_n151;
  assign new_n153 = ~pq & new_n152;
  assign new_n154 = ~pm & new_n153;
  assign new_n155 = ~pc0 & new_n154;
  assign new_n156 = pd0 & new_n155;
  assign new_n157 = ~pb0 & new_n156;
  assign new_n158 = ~py & new_n157;
  assign new_n159 = ~pa0 & new_n158;
  assign new_n160 = ~pw & new_n159;
  assign new_n161 = ~px & new_n160;
  assign new_n162 = ~pq & ~pg;
  assign new_n163 = ~pe & new_n162;
  assign new_n164 = ~pf & new_n163;
  assign new_n165 = ~pc & new_n164;
  assign new_n166 = ~pb & new_n165;
  assign new_n167 = ~pf0 & new_n166;
  assign new_n168 = pk0 & new_n167;
  assign new_n169 = ~pg0 & new_n168;
  assign new_n170 = ~py & new_n169;
  assign new_n171 = ~po & new_n170;
  assign new_n172 = pi0 & new_n171;
  assign new_n173 = ~pj0 & new_n172;
  assign new_n174 = ~pd0 & new_n173;
  assign new_n175 = ~pb0 & new_n174;
  assign new_n176 = ~pc0 & new_n175;
  assign new_n177 = ~pr & new_n176;
  assign new_n178 = ~px & new_n177;
  assign new_n179 = ~pq & ~pi;
  assign new_n180 = ~pf & new_n179;
  assign new_n181 = ~pg & new_n180;
  assign new_n182 = ~pe & new_n181;
  assign new_n183 = ~pm & new_n182;
  assign new_n184 = ~py & new_n183;
  assign new_n185 = ~pa0 & new_n184;
  assign new_n186 = ~po & new_n185;
  assign new_n187 = ~pf0 & new_n186;
  assign new_n188 = pk0 & new_n187;
  assign new_n189 = ~pv & new_n188;
  assign new_n190 = ~pj0 & new_n189;
  assign new_n191 = ~pc0 & new_n190;
  assign new_n192 = pd0 & new_n191;
  assign new_n193 = ~px & new_n192;
  assign new_n194 = ~pb0 & new_n193;
  assign new_n195 = ~pb & new_n62;
  assign new_n196 = ~pv & new_n195;
  assign new_n197 = ~py & new_n196;
  assign new_n198 = ~pa0 & new_n197;
  assign new_n199 = ~po & new_n198;
  assign new_n200 = pk0 & new_n199;
  assign new_n201 = ~pg0 & new_n200;
  assign new_n202 = ~pc0 & new_n201;
  assign new_n203 = ~px & new_n202;
  assign new_n204 = ~pb0 & new_n203;
  assign new_n205 = ~pq & new_n204;
  assign new_n206 = ~pr & new_n205;
  assign new_n207 = ~pb0 & ~px;
  assign new_n208 = ~pq & new_n207;
  assign new_n209 = ~pr & new_n208;
  assign new_n210 = ~ph & new_n209;
  assign new_n211 = ~pe0 & new_n210;
  assign new_n212 = ~pa0 & new_n211;
  assign new_n213 = ~po & new_n212;
  assign new_n214 = ~py & new_n213;
  assign new_n215 = pk0 & new_n214;
  assign new_n216 = ~pg0 & new_n215;
  assign new_n217 = ~pc0 & new_n216;
  assign new_n218 = ~pd0 & new_n217;
  assign new_n219 = ~pq & ~pr;
  assign new_n220 = ~pi & new_n219;
  assign new_n221 = ~pn & new_n220;
  assign new_n222 = ~ph & new_n221;
  assign new_n223 = ~pe0 & new_n222;
  assign new_n224 = pj0 & new_n223;
  assign new_n225 = pk0 & new_n224;
  assign new_n226 = ~pi0 & new_n225;
  assign new_n227 = ~pc0 & new_n226;
  assign new_n228 = ~pd0 & new_n227;
  assign new_n229 = ~px & new_n228;
  assign new_n230 = ~pb0 & new_n229;
  assign new_n231 = ~pq & ~pu;
  assign new_n232 = ~pm & new_n231;
  assign new_n233 = ~pn & new_n232;
  assign new_n234 = pc & new_n233;
  assign new_n235 = ~pc0 & new_n234;
  assign new_n236 = pd0 & new_n235;
  assign new_n237 = ~pb0 & new_n236;
  assign new_n238 = ~py & new_n237;
  assign new_n239 = ~pa0 & new_n238;
  assign new_n240 = ~pv & new_n239;
  assign new_n241 = ~px & new_n240;
  assign new_n242 = ~pj0 & new_n138;
  assign new_n243 = pk0 & new_n242;
  assign new_n244 = ~py & new_n243;
  assign new_n245 = ~pb0 & new_n244;
  assign new_n246 = ~pc0 & new_n245;
  assign new_n247 = ~pd0 & new_n246;
  assign new_n248 = pi0 & new_n247;
  assign new_n249 = ~pt & new_n248;
  assign new_n250 = ~px & new_n249;
  assign new_n251 = ~pr & new_n250;
  assign new_n252 = ~pn & new_n251;
  assign new_n253 = ~pq & new_n252;
  assign new_n254 = ~pj & new_n253;
  assign new_n255 = ~pl & new_n254;
  assign new_n256 = ~pm & new_n165;
  assign new_n257 = ~py & new_n256;
  assign new_n258 = ~pa0 & new_n257;
  assign new_n259 = ~po & new_n258;
  assign new_n260 = ~pf0 & new_n259;
  assign new_n261 = pk0 & new_n260;
  assign new_n262 = ~pg0 & new_n261;
  assign new_n263 = ~pj0 & new_n262;
  assign new_n264 = ~pc0 & new_n263;
  assign new_n265 = ~pd0 & new_n264;
  assign new_n266 = ~px & new_n265;
  assign new_n267 = ~pb0 & new_n266;
  assign new_n268 = ~pj0 & new_n139;
  assign new_n269 = pk0 & new_n268;
  assign new_n270 = ~py & new_n269;
  assign new_n271 = ~pf0 & new_n270;
  assign new_n272 = ~pd0 & new_n271;
  assign new_n273 = pi0 & new_n272;
  assign new_n274 = ~pc0 & new_n273;
  assign new_n275 = ~px & new_n274;
  assign new_n276 = ~pb0 & new_n275;
  assign new_n277 = ~pn & new_n276;
  assign new_n278 = ~pq & new_n277;
  assign new_n279 = ~pr & ~px;
  assign new_n280 = ~pi & new_n279;
  assign new_n281 = ~pq & new_n280;
  assign new_n282 = ~ph & new_n281;
  assign new_n283 = ~pe0 & new_n282;
  assign new_n284 = ~pa0 & new_n283;
  assign new_n285 = ~po & new_n284;
  assign new_n286 = ~py & new_n285;
  assign new_n287 = ~pd0 & new_n286;
  assign new_n288 = pk0 & new_n287;
  assign new_n289 = ~pb0 & new_n288;
  assign new_n290 = ~pc0 & new_n289;
  assign new_n291 = ~pn & new_n279;
  assign new_n292 = ~pq & new_n291;
  assign new_n293 = ~ph & new_n292;
  assign new_n294 = ~pe0 & new_n293;
  assign new_n295 = pk0 & new_n294;
  assign new_n296 = ~pg0 & new_n295;
  assign new_n297 = pj0 & new_n296;
  assign new_n298 = ~pd0 & new_n297;
  assign new_n299 = ~pi0 & new_n298;
  assign new_n300 = ~pb0 & new_n299;
  assign new_n301 = ~pc0 & new_n300;
  assign new_n302 = ~po & new_n92;
  assign new_n303 = ~pq & new_n302;
  assign new_n304 = ~pm & new_n303;
  assign new_n305 = pj0 & new_n304;
  assign new_n306 = ~pi0 & new_n305;
  assign new_n307 = ~pd0 & new_n306;
  assign new_n308 = ph0 & new_n307;
  assign new_n309 = ~pb0 & new_n308;
  assign new_n310 = ~pc0 & new_n309;
  assign new_n311 = ~pg & ~pj;
  assign new_n312 = ~pe & new_n311;
  assign new_n313 = ~pf & new_n312;
  assign new_n314 = ~pc & new_n313;
  assign new_n315 = ~pg0 & new_n314;
  assign new_n316 = ~py & new_n315;
  assign new_n317 = ~pa0 & new_n316;
  assign new_n318 = ~pj0 & new_n317;
  assign new_n319 = pk0 & new_n318;
  assign new_n320 = pd & new_n319;
  assign new_n321 = ~ps & new_n320;
  assign new_n322 = ~pc0 & new_n321;
  assign new_n323 = ~pd0 & new_n322;
  assign new_n324 = ~pb0 & new_n323;
  assign new_n325 = ~pr & new_n324;
  assign new_n326 = ~px & new_n325;
  assign new_n327 = ~pn & new_n326;
  assign new_n328 = ~pq & new_n327;
  assign new_n329 = ~py & new_n139;
  assign new_n330 = ~pa0 & new_n329;
  assign new_n331 = ~po & new_n330;
  assign new_n332 = ~pf0 & new_n331;
  assign new_n333 = ~pj0 & new_n332;
  assign new_n334 = pk0 & new_n333;
  assign new_n335 = ~pd0 & new_n334;
  assign new_n336 = ~pb0 & new_n335;
  assign new_n337 = ~pc0 & new_n336;
  assign new_n338 = ~pq & new_n337;
  assign new_n339 = ~px & new_n338;
  assign new_n340 = ~pg0 & new_n195;
  assign new_n341 = ~py & new_n340;
  assign new_n342 = ~pa0 & new_n341;
  assign new_n343 = ~po & new_n342;
  assign new_n344 = ~pd0 & new_n343;
  assign new_n345 = pk0 & new_n344;
  assign new_n346 = ~pc0 & new_n345;
  assign new_n347 = ~px & new_n346;
  assign new_n348 = ~pb0 & new_n347;
  assign new_n349 = ~pq & new_n348;
  assign new_n350 = ~pr & new_n349;
  assign new_n351 = ~py & new_n211;
  assign new_n352 = ~po & new_n351;
  assign new_n353 = ~pg0 & new_n352;
  assign new_n354 = pi0 & new_n353;
  assign new_n355 = pk0 & new_n354;
  assign new_n356 = ~pc0 & new_n355;
  assign new_n357 = ~pd0 & new_n356;
  assign new_n358 = pn & new_n207;
  assign new_n359 = ~pq & new_n358;
  assign new_n360 = ph & new_n359;
  assign new_n361 = ~pm & new_n360;
  assign new_n362 = pk & new_n361;
  assign new_n363 = pf0 & new_n362;
  assign new_n364 = ~po & new_n363;
  assign new_n365 = pi0 & new_n364;
  assign new_n366 = ~py & new_n365;
  assign new_n367 = ~pc0 & new_n366;
  assign new_n368 = ~pd0 & new_n367;
  assign new_n369 = ~pg0 & new_n256;
  assign new_n370 = ~py & new_n369;
  assign new_n371 = ~po & new_n370;
  assign new_n372 = ~pf0 & new_n371;
  assign new_n373 = ~pj0 & new_n372;
  assign new_n374 = pk0 & new_n373;
  assign new_n375 = pi0 & new_n374;
  assign new_n376 = ~pc0 & new_n375;
  assign new_n377 = ~pd0 & new_n376;
  assign new_n378 = ~px & new_n377;
  assign new_n379 = ~pb0 & new_n378;
  assign new_n380 = ~pc0 & new_n199;
  assign new_n381 = pk0 & new_n380;
  assign new_n382 = ~pb0 & new_n381;
  assign new_n383 = ~pr & new_n382;
  assign new_n384 = ~px & new_n383;
  assign new_n385 = ~pi & new_n384;
  assign new_n386 = ~pq & new_n385;
  assign new_n387 = ~py & new_n283;
  assign new_n388 = ~po & new_n387;
  assign new_n389 = pk0 & new_n388;
  assign new_n390 = ~pd0 & new_n389;
  assign new_n391 = pi0 & new_n390;
  assign new_n392 = ~pb0 & new_n391;
  assign new_n393 = ~pc0 & new_n392;
  assign new_n394 = pv & new_n364;
  assign new_n395 = ~py & new_n394;
  assign new_n396 = ~pc0 & new_n395;
  assign new_n397 = pi0 & new_n396;
  assign new_n398 = ~po & new_n232;
  assign new_n399 = pc & new_n398;
  assign new_n400 = ~pc0 & new_n399;
  assign new_n401 = pd0 & new_n400;
  assign new_n402 = ~pb0 & new_n401;
  assign new_n403 = ~py & new_n402;
  assign new_n404 = ~pa0 & new_n403;
  assign new_n405 = ~pv & new_n404;
  assign new_n406 = ~px & new_n405;
  assign new_n407 = ~po & new_n141;
  assign new_n408 = ~pf0 & new_n407;
  assign new_n409 = pi0 & new_n408;
  assign new_n410 = ~pj0 & new_n409;
  assign new_n411 = ~pd0 & new_n410;
  assign new_n412 = ~pb0 & new_n411;
  assign new_n413 = ~pc0 & new_n412;
  assign new_n414 = ~pq & new_n413;
  assign new_n415 = ~px & new_n414;
  assign new_n416 = pk0 & new_n195;
  assign new_n417 = ~pg0 & new_n416;
  assign new_n418 = ~py & new_n417;
  assign new_n419 = ~po & new_n418;
  assign new_n420 = ~pd0 & new_n419;
  assign new_n421 = pi0 & new_n420;
  assign new_n422 = ~pc0 & new_n421;
  assign new_n423 = ~px & new_n422;
  assign new_n424 = ~pb0 & new_n423;
  assign new_n425 = ~pq & new_n424;
  assign new_n426 = ~pr & new_n425;
  assign new_n427 = ~pg0 & new_n211;
  assign new_n428 = ~po & new_n427;
  assign new_n429 = pk0 & new_n428;
  assign new_n430 = ~pi0 & new_n429;
  assign new_n431 = pj0 & new_n430;
  assign new_n432 = ~pc0 & new_n431;
  assign new_n433 = ~pd0 & new_n432;
  assign new_n434 = ~pi0 & new_n364;
  assign new_n435 = pj0 & new_n434;
  assign new_n436 = ~pc0 & new_n435;
  assign new_n437 = ~pd0 & new_n436;
  assign new_n438 = ~pq & ~pn;
  assign new_n439 = ~pf & new_n438;
  assign new_n440 = ~pg & new_n439;
  assign new_n441 = ~pe & new_n440;
  assign new_n442 = ~pm & new_n441;
  assign new_n443 = ~pv & new_n442;
  assign new_n444 = ~py & new_n443;
  assign new_n445 = ~pa0 & new_n444;
  assign new_n446 = ~pf0 & new_n445;
  assign new_n447 = pk0 & new_n446;
  assign new_n448 = ~pg0 & new_n447;
  assign new_n449 = ~pj0 & new_n448;
  assign new_n450 = ~pc0 & new_n449;
  assign new_n451 = pd0 & new_n450;
  assign new_n452 = ~px & new_n451;
  assign new_n453 = ~pb0 & new_n452;
  assign new_n454 = ~py & new_n416;
  assign new_n455 = ~pa0 & new_n454;
  assign new_n456 = ~po & new_n455;
  assign new_n457 = ~pc0 & new_n456;
  assign new_n458 = ~pd0 & new_n457;
  assign new_n459 = ~pb0 & new_n458;
  assign new_n460 = ~pr & new_n459;
  assign new_n461 = ~px & new_n460;
  assign new_n462 = ~pi & new_n461;
  assign new_n463 = ~pq & new_n462;
  assign new_n464 = pk0 & new_n283;
  assign new_n465 = ~po & new_n464;
  assign new_n466 = pj0 & new_n465;
  assign new_n467 = ~pd0 & new_n466;
  assign new_n468 = ~pi0 & new_n467;
  assign new_n469 = ~pb0 & new_n468;
  assign new_n470 = ~pc0 & new_n469;
  assign new_n471 = pj0 & new_n364;
  assign new_n472 = pv & new_n471;
  assign new_n473 = ~pc0 & new_n472;
  assign new_n474 = ~pi0 & new_n473;
  assign new_n475 = ~pi & ~pn;
  assign new_n476 = ~pf & new_n475;
  assign new_n477 = ~pg & new_n476;
  assign new_n478 = ~pe & new_n477;
  assign new_n479 = ~pm & new_n478;
  assign new_n480 = ~pv & new_n479;
  assign new_n481 = ~py & new_n480;
  assign new_n482 = ~pa0 & new_n481;
  assign new_n483 = ~pf0 & new_n482;
  assign new_n484 = ~pj0 & new_n483;
  assign new_n485 = pk0 & new_n484;
  assign new_n486 = pd0 & new_n485;
  assign new_n487 = ~pb0 & new_n486;
  assign new_n488 = ~pc0 & new_n487;
  assign new_n489 = ~pq & new_n488;
  assign new_n490 = ~px & new_n489;
  assign new_n491 = ~py & new_n294;
  assign new_n492 = ~pa0 & new_n491;
  assign new_n493 = ~pg0 & new_n492;
  assign new_n494 = ~pd0 & new_n493;
  assign new_n495 = pk0 & new_n494;
  assign new_n496 = ~pb0 & new_n495;
  assign new_n497 = ~pc0 & new_n496;
  assign new_n498 = ~pq & ~pt;
  assign new_n499 = ~pl & new_n498;
  assign new_n500 = ~pn & new_n499;
  assign new_n501 = ph & new_n500;
  assign new_n502 = ~pm & new_n501;
  assign new_n503 = pk & new_n502;
  assign new_n504 = pf0 & new_n503;
  assign new_n505 = ~pa0 & new_n504;
  assign new_n506 = ~pc0 & new_n505;
  assign new_n507 = ~py & new_n506;
  assign new_n508 = ~px & new_n507;
  assign new_n509 = ~pb0 & new_n508;
  assign new_n510 = pv & ~py;
  assign new_n511 = ~pi0 & new_n510;
  assign new_n512 = ~pg0 & new_n511;
  assign new_n513 = ~pc0 & new_n512;
  assign new_n514 = ph0 & new_n513;
  assign new_n515 = ~pf0 & new_n514;
  assign new_n516 = ~pe0 & new_n515;
  assign new_n517 = ~pa0 & new_n516;
  assign new_n518 = po & new_n517;
  assign new_n519 = pv & ~pg0;
  assign new_n520 = ~pi0 & new_n519;
  assign new_n521 = pj0 & new_n520;
  assign new_n522 = ~pc0 & new_n521;
  assign new_n523 = ~pe0 & new_n522;
  assign new_n524 = ph0 & new_n523;
  assign new_n525 = po & new_n524;
  assign new_n526 = ~pf0 & new_n525;
  assign new_n527 = ~pe0 & ~pf0;
  assign new_n528 = ~pc0 & new_n527;
  assign new_n529 = pd0 & new_n528;
  assign new_n530 = pw & new_n529;
  assign new_n531 = pj0 & new_n530;
  assign new_n532 = ~pg0 & new_n531;
  assign new_n533 = ~pi0 & new_n532;
  assign new_n534 = ~pd0 & new_n528;
  assign new_n535 = pz & new_n534;
  assign new_n536 = ~pi0 & new_n535;
  assign new_n537 = pj0 & new_n536;
  assign new_n538 = ~pg0 & new_n537;
  assign new_n539 = ph0 & new_n538;
  assign new_n540 = pi0 & new_n195;
  assign new_n541 = pk0 & new_n540;
  assign new_n542 = ~py & new_n541;
  assign new_n543 = ~po & new_n542;
  assign new_n544 = ~pc0 & new_n543;
  assign new_n545 = ~pd0 & new_n544;
  assign new_n546 = ~pb0 & new_n545;
  assign new_n547 = ~pr & new_n546;
  assign new_n548 = ~px & new_n547;
  assign new_n549 = ~pi & new_n548;
  assign new_n550 = ~pq & new_n549;
  assign new_n551 = ~py & new_n223;
  assign new_n552 = ~pa0 & new_n551;
  assign new_n553 = pk0 & new_n552;
  assign new_n554 = ~pc0 & new_n553;
  assign new_n555 = ~pd0 & new_n554;
  assign new_n556 = ~px & new_n555;
  assign new_n557 = ~pb0 & new_n556;
  assign new_n558 = ~pn & new_n207;
  assign new_n559 = ~pq & new_n558;
  assign new_n560 = ph & new_n559;
  assign new_n561 = ~pm & new_n560;
  assign new_n562 = pk & new_n561;
  assign new_n563 = pf0 & new_n562;
  assign new_n564 = ~pa0 & new_n563;
  assign new_n565 = ~ps & new_n564;
  assign new_n566 = ~py & new_n565;
  assign new_n567 = ~pc0 & new_n566;
  assign new_n568 = pd & new_n567;
  assign new_n569 = ~pg0 & ~py;
  assign new_n570 = ~pd0 & new_n569;
  assign new_n571 = ~pi0 & new_n570;
  assign new_n572 = ~pc0 & new_n571;
  assign new_n573 = ph0 & new_n572;
  assign new_n574 = ~pf0 & new_n573;
  assign new_n575 = ~pe0 & new_n574;
  assign new_n576 = ~pa0 & new_n575;
  assign new_n577 = po & new_n576;
  assign new_n578 = ph0 & new_n522;
  assign new_n579 = pz & new_n578;
  assign new_n580 = ~pf0 & new_n579;
  assign new_n581 = ~pe0 & new_n580;
  assign new_n582 = ~px & ~py;
  assign new_n583 = ~pq & new_n582;
  assign new_n584 = ~pr & new_n583;
  assign new_n585 = ~po & new_n584;
  assign new_n586 = ph0 & new_n585;
  assign new_n587 = ~pb0 & new_n586;
  assign new_n588 = ~pc0 & new_n587;
  assign new_n589 = pz & new_n588;
  assign new_n590 = ~pa0 & new_n589;
  assign new_n591 = ~pc0 & ~pd0;
  assign new_n592 = pz & new_n591;
  assign new_n593 = ~pa0 & new_n592;
  assign new_n594 = ~py & new_n593;
  assign new_n595 = ~pi0 & new_n594;
  assign new_n596 = ~pg0 & new_n595;
  assign new_n597 = ph0 & new_n596;
  assign new_n598 = ~pe0 & new_n597;
  assign new_n599 = ~pf0 & new_n598;
  assign new_n600 = ~pg0 & new_n294;
  assign new_n601 = ~py & new_n600;
  assign new_n602 = pk0 & new_n601;
  assign new_n603 = ~pd0 & new_n602;
  assign new_n604 = pi0 & new_n603;
  assign new_n605 = ~pb0 & new_n604;
  assign new_n606 = ~pc0 & new_n605;
  assign new_n607 = pn & new_n279;
  assign new_n608 = ~pq & new_n607;
  assign new_n609 = ph & new_n608;
  assign new_n610 = pf0 & new_n609;
  assign new_n611 = ~po & new_n610;
  assign new_n612 = pk & new_n611;
  assign new_n613 = ~py & new_n612;
  assign new_n614 = ~pd0 & new_n613;
  assign new_n615 = pi0 & new_n614;
  assign new_n616 = ~pb0 & new_n615;
  assign new_n617 = ~pc0 & new_n616;
  assign new_n618 = ~pj & new_n207;
  assign new_n619 = ~pq & new_n618;
  assign new_n620 = ph & new_n619;
  assign new_n621 = pf0 & new_n620;
  assign new_n622 = ~pm & new_n621;
  assign new_n623 = ~po & new_n622;
  assign new_n624 = pj0 & new_n623;
  assign new_n625 = pv & new_n624;
  assign new_n626 = ~pc0 & new_n625;
  assign new_n627 = ~pi0 & new_n626;
  assign new_n628 = ~pc0 & new_n519;
  assign new_n629 = pi0 & new_n628;
  assign new_n630 = ~px & new_n629;
  assign new_n631 = ph0 & new_n630;
  assign new_n632 = ~pf0 & new_n631;
  assign new_n633 = ~pe0 & new_n632;
  assign new_n634 = ~py & new_n633;
  assign new_n635 = po & new_n634;
  assign new_n636 = ~pi0 & pj0;
  assign new_n637 = ~pc0 & new_n636;
  assign new_n638 = ~pd0 & new_n637;
  assign new_n639 = ~ph & new_n638;
  assign new_n640 = ~pf0 & new_n639;
  assign new_n641 = ~pe0 & new_n640;
  assign new_n642 = pk0 & new_n641;
  assign new_n643 = ~pg0 & new_n642;
  assign new_n644 = pw & ~px;
  assign new_n645 = ~po & new_n644;
  assign new_n646 = ~pq & new_n645;
  assign new_n647 = ~pm & new_n646;
  assign new_n648 = pd0 & new_n647;
  assign new_n649 = ~pb0 & new_n648;
  assign new_n650 = ~pc0 & new_n649;
  assign new_n651 = ~py & new_n650;
  assign new_n652 = ~pa0 & new_n651;
  assign new_n653 = ~py & new_n591;
  assign new_n654 = pz & new_n653;
  assign new_n655 = ~px & new_n654;
  assign new_n656 = pi0 & new_n655;
  assign new_n657 = ~pg0 & new_n656;
  assign new_n658 = ph0 & new_n657;
  assign new_n659 = ~pe0 & new_n658;
  assign new_n660 = ~pf0 & new_n659;
  assign new_n661 = pk0 & new_n223;
  assign new_n662 = ~py & new_n661;
  assign new_n663 = pi0 & new_n662;
  assign new_n664 = ~pc0 & new_n663;
  assign new_n665 = ~pd0 & new_n664;
  assign new_n666 = ~px & new_n665;
  assign new_n667 = ~pb0 & new_n666;
  assign new_n668 = pi0 & new_n613;
  assign new_n669 = pv & new_n668;
  assign new_n670 = ~pb0 & new_n669;
  assign new_n671 = ~pc0 & new_n670;
  assign new_n672 = pi0 & new_n623;
  assign new_n673 = ~py & new_n672;
  assign new_n674 = ~pc0 & new_n673;
  assign new_n675 = ~pd0 & new_n674;
  assign new_n676 = ~pb0 & ~pc0;
  assign new_n677 = ~pq & new_n676;
  assign new_n678 = ~px & new_n677;
  assign new_n679 = ~pn & new_n678;
  assign new_n680 = ph0 & new_n679;
  assign new_n681 = po & new_n680;
  assign new_n682 = ~pm & new_n681;
  assign new_n683 = ~py & new_n682;
  assign new_n684 = ~pa0 & new_n683;
  assign new_n685 = ~pg0 & pj0;
  assign new_n686 = pd0 & new_n685;
  assign new_n687 = ~pi0 & new_n686;
  assign new_n688 = ~pc0 & new_n687;
  assign new_n689 = ~pe0 & new_n688;
  assign new_n690 = pu & new_n689;
  assign new_n691 = ~pv & new_n690;
  assign new_n692 = ~pf0 & new_n691;
  assign new_n693 = ~pn & new_n644;
  assign new_n694 = ~pq & new_n693;
  assign new_n695 = ~pm & new_n694;
  assign new_n696 = pi0 & new_n695;
  assign new_n697 = ~pc0 & new_n696;
  assign new_n698 = pd0 & new_n697;
  assign new_n699 = ~py & new_n698;
  assign new_n700 = ~pb0 & new_n699;
  assign new_n701 = po & new_n534;
  assign new_n702 = ~pi0 & new_n701;
  assign new_n703 = pj0 & new_n702;
  assign new_n704 = ~pg0 & new_n703;
  assign new_n705 = ph0 & new_n704;
  assign new_n706 = ~pj & new_n279;
  assign new_n707 = ~pq & new_n706;
  assign new_n708 = ph & new_n707;
  assign new_n709 = ~po & new_n708;
  assign new_n710 = pf0 & new_n709;
  assign new_n711 = pv & new_n710;
  assign new_n712 = ~pi0 & new_n711;
  assign new_n713 = pj0 & new_n712;
  assign new_n714 = ~pb0 & new_n713;
  assign new_n715 = ~pc0 & new_n714;
  assign new_n716 = ~pc0 & ~pi0;
  assign new_n717 = ~px & new_n716;
  assign new_n718 = ~pb0 & new_n717;
  assign new_n719 = ~pq & new_n718;
  assign new_n720 = pz & new_n719;
  assign new_n721 = ph0 & new_n720;
  assign new_n722 = ~po & new_n721;
  assign new_n723 = ~pm & new_n722;
  assign new_n724 = pj0 & new_n723;
  assign new_n725 = pv & new_n724;
  assign new_n726 = ~pn & new_n209;
  assign new_n727 = ph0 & new_n726;
  assign new_n728 = ~pa0 & new_n727;
  assign new_n729 = po & new_n728;
  assign new_n730 = ~pc0 & new_n729;
  assign new_n731 = ~py & new_n730;
  assign new_n732 = ~pc0 & pd0;
  assign new_n733 = ~px & new_n732;
  assign new_n734 = ~py & new_n733;
  assign new_n735 = pw & new_n734;
  assign new_n736 = ~pg0 & new_n735;
  assign new_n737 = pi0 & new_n736;
  assign new_n738 = ~pe0 & new_n737;
  assign new_n739 = ~pf0 & new_n738;
  assign new_n740 = ~pq & new_n644;
  assign new_n741 = ~pr & new_n740;
  assign new_n742 = ~po & new_n741;
  assign new_n743 = pi0 & new_n742;
  assign new_n744 = ~pc0 & new_n743;
  assign new_n745 = pd0 & new_n744;
  assign new_n746 = ~py & new_n745;
  assign new_n747 = ~pb0 & new_n746;
  assign new_n748 = pj0 & new_n695;
  assign new_n749 = pd0 & new_n748;
  assign new_n750 = ~pi0 & new_n749;
  assign new_n751 = ~pb0 & new_n750;
  assign new_n752 = ~pc0 & new_n751;
  assign new_n753 = pj0 & new_n710;
  assign new_n754 = ~pd0 & new_n753;
  assign new_n755 = ~pi0 & new_n754;
  assign new_n756 = ~pb0 & new_n755;
  assign new_n757 = ~pc0 & new_n756;
  assign new_n758 = ~pc0 & pi0;
  assign new_n759 = ~px & new_n758;
  assign new_n760 = ~pb0 & new_n759;
  assign new_n761 = ~pq & new_n760;
  assign new_n762 = pz & new_n761;
  assign new_n763 = ph0 & new_n762;
  assign new_n764 = ~po & new_n763;
  assign new_n765 = ~pm & new_n764;
  assign new_n766 = pv & new_n765;
  assign new_n767 = ~py & new_n766;
  assign new_n768 = ~pv & ~pg0;
  assign new_n769 = pd0 & new_n768;
  assign new_n770 = ~pi0 & new_n769;
  assign new_n771 = ~pc0 & new_n770;
  assign new_n772 = pu & new_n771;
  assign new_n773 = ~pf0 & new_n772;
  assign new_n774 = ~pe0 & new_n773;
  assign new_n775 = ~py & new_n774;
  assign new_n776 = ~pa0 & new_n775;
  assign new_n777 = ~pn & new_n741;
  assign new_n778 = pd0 & new_n777;
  assign new_n779 = ~pb0 & new_n778;
  assign new_n780 = ~pc0 & new_n779;
  assign new_n781 = ~py & new_n780;
  assign new_n782 = ~pa0 & new_n781;
  assign new_n783 = pi0 & new_n647;
  assign new_n784 = ~pc0 & new_n783;
  assign new_n785 = pd0 & new_n784;
  assign new_n786 = ~py & new_n785;
  assign new_n787 = ~pb0 & new_n786;
  assign new_n788 = ~po & new_n582;
  assign new_n789 = ~pq & new_n788;
  assign new_n790 = ~pm & new_n789;
  assign new_n791 = pi0 & new_n790;
  assign new_n792 = ph0 & new_n791;
  assign new_n793 = ~pc0 & new_n792;
  assign new_n794 = ~pd0 & new_n793;
  assign new_n795 = pz & new_n794;
  assign new_n796 = ~pb0 & new_n795;
  assign new_n797 = pu & new_n679;
  assign new_n798 = ~pm & new_n797;
  assign new_n799 = ~pv & new_n798;
  assign new_n800 = ~py & new_n799;
  assign new_n801 = pd0 & new_n800;
  assign new_n802 = pi0 & new_n801;
  assign new_n803 = pz & new_n630;
  assign new_n804 = ~pe0 & new_n803;
  assign new_n805 = ph0 & new_n804;
  assign new_n806 = ~py & new_n805;
  assign new_n807 = ~pf0 & new_n806;
  assign new_n808 = ~pg0 & pi0;
  assign new_n809 = ~pc0 & new_n808;
  assign new_n810 = pd0 & new_n809;
  assign new_n811 = ~px & new_n810;
  assign new_n812 = pu & new_n811;
  assign new_n813 = ~pf0 & new_n812;
  assign new_n814 = ~pe0 & new_n813;
  assign new_n815 = ~pv & new_n814;
  assign new_n816 = ~py & new_n815;
  assign new_n817 = ~py & new_n732;
  assign new_n818 = ~pa0 & new_n817;
  assign new_n819 = pw & new_n818;
  assign new_n820 = ~pg0 & new_n819;
  assign new_n821 = ~pi0 & new_n820;
  assign new_n822 = ~pe0 & new_n821;
  assign new_n823 = ~pf0 & new_n822;
  assign new_n824 = ~px & new_n591;
  assign new_n825 = ~py & new_n824;
  assign new_n826 = po & new_n825;
  assign new_n827 = pi0 & new_n826;
  assign new_n828 = ~pg0 & new_n827;
  assign new_n829 = ph0 & new_n828;
  assign new_n830 = ~pe0 & new_n829;
  assign new_n831 = ~pf0 & new_n830;
  assign new_n832 = pj0 & new_n777;
  assign new_n833 = pd0 & new_n832;
  assign new_n834 = ~pi0 & new_n833;
  assign new_n835 = ~pb0 & new_n834;
  assign new_n836 = ~pc0 & new_n835;
  assign new_n837 = pj0 & new_n798;
  assign new_n838 = ~pv & new_n837;
  assign new_n839 = pd0 & new_n838;
  assign new_n840 = ~pi0 & new_n839;
  assign new_n841 = pz & new_n513;
  assign new_n842 = ~pe0 & new_n841;
  assign new_n843 = ph0 & new_n842;
  assign new_n844 = ~pa0 & new_n843;
  assign new_n845 = ~pf0 & new_n844;
  assign new_n846 = ~pj0 & pk0;
  assign new_n847 = ~pd0 & new_n846;
  assign new_n848 = ~pi0 & new_n847;
  assign new_n849 = ~pc0 & new_n848;
  assign new_n850 = ~pe0 & new_n849;
  assign new_n851 = ~pa0 & new_n850;
  assign new_n852 = ~pf0 & new_n851;
  assign new_n853 = ~pg0 & new_n852;
  assign new_n854 = ~py & new_n853;
  assign new_n855 = pd0 & new_n695;
  assign new_n856 = ~pb0 & new_n855;
  assign new_n857 = ~pc0 & new_n856;
  assign new_n858 = ~py & new_n857;
  assign new_n859 = ~pa0 & new_n858;
  assign new_n860 = ph0 & new_n790;
  assign new_n861 = ~pb0 & new_n860;
  assign new_n862 = ~pc0 & new_n861;
  assign new_n863 = pz & new_n862;
  assign new_n864 = ~pa0 & new_n863;
  assign new_n865 = pi0 & new_n585;
  assign new_n866 = ph0 & new_n865;
  assign new_n867 = ~pc0 & new_n866;
  assign new_n868 = ~pd0 & new_n867;
  assign new_n869 = pz & new_n868;
  assign new_n870 = ~pb0 & new_n869;
  assign new_n871 = ~pg0 & new_n541;
  assign new_n872 = ~py & new_n871;
  assign new_n873 = ~pc0 & new_n872;
  assign new_n874 = ~pd0 & new_n873;
  assign new_n875 = ~pb0 & new_n874;
  assign new_n876 = ~pr & new_n875;
  assign new_n877 = ~px & new_n876;
  assign new_n878 = ~pn & new_n877;
  assign new_n879 = ~pq & new_n878;
  assign new_n880 = pj0 & new_n62;
  assign new_n881 = pk0 & new_n880;
  assign new_n882 = ~po & new_n881;
  assign new_n883 = ~pm & new_n882;
  assign new_n884 = ~pd0 & new_n883;
  assign new_n885 = ~pi0 & new_n884;
  assign new_n886 = ~pc0 & new_n885;
  assign new_n887 = ~px & new_n886;
  assign new_n888 = ~pb0 & new_n887;
  assign new_n889 = ~pi & new_n888;
  assign new_n890 = ~pq & new_n889;
  assign new_n891 = ~pc & new_n292;
  assign new_n892 = ~pa0 & new_n891;
  assign new_n893 = ~pf0 & new_n892;
  assign new_n894 = ~pe0 & new_n893;
  assign new_n895 = ~pv & new_n894;
  assign new_n896 = ~py & new_n895;
  assign new_n897 = ~pg0 & new_n896;
  assign new_n898 = ~pj0 & new_n897;
  assign new_n899 = pk0 & new_n898;
  assign new_n900 = ~pb0 & new_n899;
  assign new_n901 = ~pc0 & new_n900;
  assign new_n902 = ~pi & new_n209;
  assign new_n903 = ~pf0 & new_n902;
  assign new_n904 = ~pe0 & new_n903;
  assign new_n905 = ~py & new_n904;
  assign new_n906 = ~po & new_n905;
  assign new_n907 = pk0 & new_n906;
  assign new_n908 = pi0 & new_n907;
  assign new_n909 = ~pj0 & new_n908;
  assign new_n910 = ~pc0 & new_n909;
  assign new_n911 = ~pd0 & new_n910;
  assign new_n912 = ~pl & new_n219;
  assign new_n913 = ~pn & new_n912;
  assign new_n914 = ph & new_n913;
  assign new_n915 = pf0 & new_n914;
  assign new_n916 = ~pa0 & new_n915;
  assign new_n917 = pk & new_n916;
  assign new_n918 = ~py & new_n917;
  assign new_n919 = ~pb0 & new_n918;
  assign new_n920 = ~pc0 & new_n919;
  assign new_n921 = ~pt & new_n920;
  assign new_n922 = ~px & new_n921;
  assign new_n923 = ~pj & new_n119;
  assign new_n924 = ~pn & new_n923;
  assign new_n925 = ph & new_n924;
  assign new_n926 = pf0 & new_n925;
  assign new_n927 = ~pm & new_n926;
  assign new_n928 = pj0 & new_n927;
  assign new_n929 = ~pd0 & new_n928;
  assign new_n930 = ~pi0 & new_n929;
  assign new_n931 = ~pb0 & new_n930;
  assign new_n932 = ~pc0 & new_n931;
  assign new_n933 = pa & new_n679;
  assign new_n934 = ~pm & new_n933;
  assign new_n935 = ~py & new_n934;
  assign new_n936 = ~pa0 & new_n935;
  assign new_n937 = pd0 & new_n936;
  assign new_n938 = ~pv & new_n937;
  assign new_n939 = ~pb0 & new_n733;
  assign new_n940 = ~pq & new_n939;
  assign new_n941 = pu & new_n940;
  assign new_n942 = ~pm & new_n941;
  assign new_n943 = ~py & new_n942;
  assign new_n944 = ~po & new_n943;
  assign new_n945 = pi0 & new_n944;
  assign new_n946 = ~pv & new_n945;
  assign new_n947 = ~pj & new_n219;
  assign new_n948 = ~pn & new_n947;
  assign new_n949 = ph & new_n948;
  assign new_n950 = pf0 & new_n949;
  assign new_n951 = ~pa0 & new_n950;
  assign new_n952 = ~pc0 & new_n951;
  assign new_n953 = ~py & new_n952;
  assign new_n954 = ~px & new_n953;
  assign new_n955 = ~pb0 & new_n954;
  assign new_n956 = pi0 & ~pj0;
  assign new_n957 = ~pc0 & new_n956;
  assign new_n958 = ~pd0 & new_n957;
  assign new_n959 = ~px & new_n958;
  assign new_n960 = ~pe0 & new_n959;
  assign new_n961 = ~py & new_n960;
  assign new_n962 = ~pf0 & new_n961;
  assign new_n963 = pk0 & new_n962;
  assign new_n964 = ~pg0 & new_n963;
  assign new_n965 = pi0 & new_n777;
  assign new_n966 = ~pc0 & new_n965;
  assign new_n967 = pd0 & new_n966;
  assign new_n968 = ~py & new_n967;
  assign new_n969 = ~pb0 & new_n968;
  assign new_n970 = ~pd0 & new_n195;
  assign new_n971 = pi0 & new_n970;
  assign new_n972 = pk0 & new_n971;
  assign new_n973 = ~py & new_n972;
  assign new_n974 = ~pb0 & new_n973;
  assign new_n975 = ~pc0 & new_n974;
  assign new_n976 = ~px & new_n975;
  assign new_n977 = ~pq & new_n976;
  assign new_n978 = ~pr & new_n977;
  assign new_n979 = ~pi & new_n978;
  assign new_n980 = ~pn & new_n979;
  assign new_n981 = ~pg0 & new_n63;
  assign new_n982 = ~po & new_n981;
  assign new_n983 = ~pm & new_n982;
  assign new_n984 = ~pi0 & new_n983;
  assign new_n985 = pj0 & new_n984;
  assign new_n986 = ~pd0 & new_n985;
  assign new_n987 = ~pb0 & new_n986;
  assign new_n988 = ~pc0 & new_n987;
  assign new_n989 = ~pq & new_n988;
  assign new_n990 = ~px & new_n989;
  assign new_n991 = ~pc & new_n221;
  assign new_n992 = ~pa0 & new_n991;
  assign new_n993 = ~pf0 & new_n992;
  assign new_n994 = ~pe0 & new_n993;
  assign new_n995 = ~pv & new_n994;
  assign new_n996 = ~py & new_n995;
  assign new_n997 = pk0 & new_n996;
  assign new_n998 = ~pc0 & new_n997;
  assign new_n999 = ~pj0 & new_n998;
  assign new_n1000 = ~px & new_n999;
  assign new_n1001 = ~pb0 & new_n1000;
  assign new_n1002 = ~pa0 & new_n904;
  assign new_n1003 = ~po & new_n1002;
  assign new_n1004 = ~py & new_n1003;
  assign new_n1005 = ~pj0 & new_n1004;
  assign new_n1006 = pk0 & new_n1005;
  assign new_n1007 = ~pc0 & new_n1006;
  assign new_n1008 = ~pd0 & new_n1007;
  assign new_n1009 = ph & new_n292;
  assign new_n1010 = pf0 & new_n1009;
  assign new_n1011 = ~pa0 & new_n1010;
  assign new_n1012 = pk & new_n1011;
  assign new_n1013 = ~py & new_n1012;
  assign new_n1014 = pd & new_n1013;
  assign new_n1015 = ~ps & new_n1014;
  assign new_n1016 = ~pb0 & new_n1015;
  assign new_n1017 = ~pc0 & new_n1016;
  assign new_n1018 = pk & new_n609;
  assign new_n1019 = pf0 & new_n1018;
  assign new_n1020 = ~po & new_n1019;
  assign new_n1021 = ~py & new_n1020;
  assign new_n1022 = ~pa0 & new_n1021;
  assign new_n1023 = ~pb0 & new_n1022;
  assign new_n1024 = ~pc0 & new_n1023;
  assign new_n1025 = pa & new_n940;
  assign new_n1026 = ~pm & new_n1025;
  assign new_n1027 = ~pa0 & new_n1026;
  assign new_n1028 = ~po & new_n1027;
  assign new_n1029 = ~pv & new_n1028;
  assign new_n1030 = ~py & new_n1029;
  assign new_n1031 = ~pv & new_n942;
  assign new_n1032 = ~po & new_n1031;
  assign new_n1033 = ~pi0 & new_n1032;
  assign new_n1034 = pj0 & new_n1033;
  assign new_n1035 = pf0 & new_n708;
  assign new_n1036 = ~po & new_n1035;
  assign new_n1037 = ~py & new_n1036;
  assign new_n1038 = ~pa0 & new_n1037;
  assign new_n1039 = ~pb0 & new_n1038;
  assign new_n1040 = ~pc0 & new_n1039;
  assign new_n1041 = ~pd0 & pi0;
  assign new_n1042 = ~px & new_n1041;
  assign new_n1043 = ~pc0 & new_n1042;
  assign new_n1044 = ~ph & new_n1043;
  assign new_n1045 = ~pe0 & new_n1044;
  assign new_n1046 = ~py & new_n1045;
  assign new_n1047 = ~pf0 & new_n1046;
  assign new_n1048 = pk0 & new_n1047;
  assign new_n1049 = ~pg0 & new_n1048;
  assign new_n1050 = pd0 & new_n742;
  assign new_n1051 = ~pb0 & new_n1050;
  assign new_n1052 = ~pc0 & new_n1051;
  assign new_n1053 = ~py & new_n1052;
  assign new_n1054 = ~pa0 & new_n1053;
  assign new_n1055 = ~ph & ~pi;
  assign new_n1056 = ~pf & new_n1055;
  assign new_n1057 = ~pg & new_n1056;
  assign new_n1058 = ~pe & new_n1057;
  assign new_n1059 = ~pv & new_n1058;
  assign new_n1060 = ~py & new_n1059;
  assign new_n1061 = ~pa0 & new_n1060;
  assign new_n1062 = ~pb0 & new_n1061;
  assign new_n1063 = ~pc0 & new_n1062;
  assign new_n1064 = pd0 & new_n1063;
  assign new_n1065 = pk0 & new_n1064;
  assign new_n1066 = ~pt & new_n1065;
  assign new_n1067 = ~px & new_n1066;
  assign new_n1068 = ~pr & new_n1067;
  assign new_n1069 = ~pn & new_n1068;
  assign new_n1070 = ~pq & new_n1069;
  assign new_n1071 = ~pj & new_n1070;
  assign new_n1072 = ~pl & new_n1071;
  assign new_n1073 = ~pi0 & new_n195;
  assign new_n1074 = pj0 & new_n1073;
  assign new_n1075 = pk0 & new_n1074;
  assign new_n1076 = ~pg0 & new_n1075;
  assign new_n1077 = ~pc0 & new_n1076;
  assign new_n1078 = ~pd0 & new_n1077;
  assign new_n1079 = ~pb0 & new_n1078;
  assign new_n1080 = ~pr & new_n1079;
  assign new_n1081 = ~px & new_n1080;
  assign new_n1082 = ~pn & new_n1081;
  assign new_n1083 = ~pq & new_n1082;
  assign new_n1084 = ~pm & new_n1061;
  assign new_n1085 = pd0 & new_n1084;
  assign new_n1086 = pk0 & new_n1085;
  assign new_n1087 = ~pc0 & new_n1086;
  assign new_n1088 = ~px & new_n1087;
  assign new_n1089 = ~pb0 & new_n1088;
  assign new_n1090 = ~pn & new_n1089;
  assign new_n1091 = ~pq & new_n1090;
  assign new_n1092 = ~pc & new_n209;
  assign new_n1093 = ~po & new_n1092;
  assign new_n1094 = ~pf0 & new_n1093;
  assign new_n1095 = ~pe0 & new_n1094;
  assign new_n1096 = ~py & new_n1095;
  assign new_n1097 = ~pa0 & new_n1096;
  assign new_n1098 = ~pv & new_n1097;
  assign new_n1099 = pk0 & new_n1098;
  assign new_n1100 = ~pg0 & new_n1099;
  assign new_n1101 = ~pc0 & new_n1100;
  assign new_n1102 = ~pj0 & new_n1101;
  assign new_n1103 = ~pi & new_n559;
  assign new_n1104 = ~pm & new_n1103;
  assign new_n1105 = ~pe0 & new_n1104;
  assign new_n1106 = ~py & new_n1105;
  assign new_n1107 = ~pf0 & new_n1106;
  assign new_n1108 = pk0 & new_n1107;
  assign new_n1109 = pi0 & new_n1108;
  assign new_n1110 = ~pj0 & new_n1109;
  assign new_n1111 = ~pc0 & new_n1110;
  assign new_n1112 = ~pd0 & new_n1111;
  assign new_n1113 = pj0 & new_n612;
  assign new_n1114 = ~pd0 & new_n1113;
  assign new_n1115 = ~pi0 & new_n1114;
  assign new_n1116 = ~pb0 & new_n1115;
  assign new_n1117 = ~pc0 & new_n1116;
  assign new_n1118 = ~py & new_n710;
  assign new_n1119 = pi0 & new_n1118;
  assign new_n1120 = pv & new_n1119;
  assign new_n1121 = ~pb0 & new_n1120;
  assign new_n1122 = ~pc0 & new_n1121;
  assign new_n1123 = pa & new_n726;
  assign new_n1124 = ~pa0 & new_n1123;
  assign new_n1125 = ~pv & new_n1124;
  assign new_n1126 = ~py & new_n1125;
  assign new_n1127 = ~pc0 & new_n1126;
  assign new_n1128 = pd0 & new_n1127;
  assign new_n1129 = po & new_n727;
  assign new_n1130 = pv & new_n1129;
  assign new_n1131 = ~py & new_n1130;
  assign new_n1132 = ~pc0 & new_n1131;
  assign new_n1133 = pi0 & new_n1132;
  assign new_n1134 = ~pm & new_n925;
  assign new_n1135 = pf0 & new_n1134;
  assign new_n1136 = ~py & new_n1135;
  assign new_n1137 = ~pa0 & new_n1136;
  assign new_n1138 = ~pb0 & new_n1137;
  assign new_n1139 = ~pc0 & new_n1138;
  assign new_n1140 = po & new_n279;
  assign new_n1141 = ~pq & new_n1140;
  assign new_n1142 = ~pn & new_n1141;
  assign new_n1143 = pi0 & new_n1142;
  assign new_n1144 = ph0 & new_n1143;
  assign new_n1145 = ~pc0 & new_n1144;
  assign new_n1146 = ~pd0 & new_n1145;
  assign new_n1147 = ~py & new_n1146;
  assign new_n1148 = ~pb0 & new_n1147;
  assign new_n1149 = pj0 & new_n647;
  assign new_n1150 = pd0 & new_n1149;
  assign new_n1151 = ~pi0 & new_n1150;
  assign new_n1152 = ~pb0 & new_n1151;
  assign new_n1153 = ~pc0 & new_n1152;
  assign new_n1154 = pd & new_n62;
  assign new_n1155 = ~ps & new_n1154;
  assign new_n1156 = ~py & new_n1155;
  assign new_n1157 = ~pc0 & new_n1156;
  assign new_n1158 = ~pd0 & new_n1157;
  assign new_n1159 = pi0 & new_n1158;
  assign new_n1160 = pk0 & new_n1159;
  assign new_n1161 = ~px & new_n1160;
  assign new_n1162 = ~pb0 & new_n1161;
  assign new_n1163 = ~pr & new_n1162;
  assign new_n1164 = ~pn & new_n1163;
  assign new_n1165 = ~pq & new_n1164;
  assign new_n1166 = ~pi & new_n1165;
  assign new_n1167 = ~pj & new_n1166;
  assign new_n1168 = ~pi0 & new_n970;
  assign new_n1169 = pj0 & new_n1168;
  assign new_n1170 = pk0 & new_n1169;
  assign new_n1171 = ~pb0 & new_n1170;
  assign new_n1172 = ~pc0 & new_n1171;
  assign new_n1173 = ~px & new_n1172;
  assign new_n1174 = ~pq & new_n1173;
  assign new_n1175 = ~pr & new_n1174;
  assign new_n1176 = ~pi & new_n1175;
  assign new_n1177 = ~pn & new_n1176;
  assign new_n1178 = ~ph & ~pn;
  assign new_n1179 = ~pf & new_n1178;
  assign new_n1180 = ~pg & new_n1179;
  assign new_n1181 = ~pe & new_n1180;
  assign new_n1182 = ~pv & new_n1181;
  assign new_n1183 = ~py & new_n1182;
  assign new_n1184 = ~pa0 & new_n1183;
  assign new_n1185 = ~pm & new_n1184;
  assign new_n1186 = pk0 & new_n1185;
  assign new_n1187 = ~pg0 & new_n1186;
  assign new_n1188 = pd0 & new_n1187;
  assign new_n1189 = ~pb0 & new_n1188;
  assign new_n1190 = ~pc0 & new_n1189;
  assign new_n1191 = ~pq & new_n1190;
  assign new_n1192 = ~px & new_n1191;
  assign new_n1193 = ~pc & new_n281;
  assign new_n1194 = ~po & new_n1193;
  assign new_n1195 = ~pf0 & new_n1194;
  assign new_n1196 = ~pe0 & new_n1195;
  assign new_n1197 = ~py & new_n1196;
  assign new_n1198 = ~pa0 & new_n1197;
  assign new_n1199 = ~pv & new_n1198;
  assign new_n1200 = ~pj0 & new_n1199;
  assign new_n1201 = pk0 & new_n1200;
  assign new_n1202 = ~pb0 & new_n1201;
  assign new_n1203 = ~pc0 & new_n1202;
  assign new_n1204 = ~pa0 & new_n1105;
  assign new_n1205 = ~pf0 & new_n1204;
  assign new_n1206 = ~py & new_n1205;
  assign new_n1207 = ~pj0 & new_n1206;
  assign new_n1208 = pk0 & new_n1207;
  assign new_n1209 = ~pc0 & new_n1208;
  assign new_n1210 = ~pd0 & new_n1209;
  assign new_n1211 = pv & new_n612;
  assign new_n1212 = ~pi0 & new_n1211;
  assign new_n1213 = pj0 & new_n1212;
  assign new_n1214 = ~pb0 & new_n1213;
  assign new_n1215 = ~pc0 & new_n1214;
  assign new_n1216 = ~pd0 & new_n1118;
  assign new_n1217 = pi0 & new_n1216;
  assign new_n1218 = ~pb0 & new_n1217;
  assign new_n1219 = ~pc0 & new_n1218;
  assign new_n1220 = ~pr & new_n676;
  assign new_n1221 = ~px & new_n1220;
  assign new_n1222 = ~pq & new_n1221;
  assign new_n1223 = pa & new_n1222;
  assign new_n1224 = ~po & new_n1223;
  assign new_n1225 = ~py & new_n1224;
  assign new_n1226 = ~pa0 & new_n1225;
  assign new_n1227 = pd0 & new_n1226;
  assign new_n1228 = ~pv & new_n1227;
  assign new_n1229 = pj0 & new_n1129;
  assign new_n1230 = pv & new_n1229;
  assign new_n1231 = ~pc0 & new_n1230;
  assign new_n1232 = ~pi0 & new_n1231;
  assign new_n1233 = ~pm & new_n620;
  assign new_n1234 = pf0 & new_n1233;
  assign new_n1235 = ~pa0 & new_n1234;
  assign new_n1236 = ~po & new_n1235;
  assign new_n1237 = ~pc0 & new_n1236;
  assign new_n1238 = ~py & new_n1237;
  assign new_n1239 = ~pn & new_n119;
  assign new_n1240 = po & new_n1239;
  assign new_n1241 = ~pm & new_n1240;
  assign new_n1242 = pi0 & new_n1241;
  assign new_n1243 = ph0 & new_n1242;
  assign new_n1244 = ~pc0 & new_n1243;
  assign new_n1245 = ~pd0 & new_n1244;
  assign new_n1246 = ~py & new_n1245;
  assign new_n1247 = ~pb0 & new_n1246;
  assign new_n1248 = pj0 & new_n742;
  assign new_n1249 = pd0 & new_n1248;
  assign new_n1250 = ~pi0 & new_n1249;
  assign new_n1251 = ~pb0 & new_n1250;
  assign new_n1252 = ~pc0 & new_n1251;
  assign new_n1253 = ~pb & new_n138;
  assign new_n1254 = ~pf0 & new_n1253;
  assign new_n1255 = pk0 & new_n1254;
  assign new_n1256 = ~py & new_n1255;
  assign new_n1257 = ~pa0 & new_n1256;
  assign new_n1258 = ~po & new_n1257;
  assign new_n1259 = ~pd0 & new_n1258;
  assign new_n1260 = ~pj0 & new_n1259;
  assign new_n1261 = ~pc0 & new_n1260;
  assign new_n1262 = ~px & new_n1261;
  assign new_n1263 = ~pb0 & new_n1262;
  assign new_n1264 = ~pq & new_n1263;
  assign new_n1265 = ~pr & new_n1264;
  assign new_n1266 = pf0 & new_n560;
  assign new_n1267 = ~pm & new_n1266;
  assign new_n1268 = ~py & new_n1267;
  assign new_n1269 = pk & new_n1268;
  assign new_n1270 = pv & new_n1269;
  assign new_n1271 = pd & new_n1270;
  assign new_n1272 = ~ps & new_n1271;
  assign new_n1273 = ~pc0 & new_n1272;
  assign new_n1274 = pi0 & new_n1273;
  assign new_n1275 = pk & new_n914;
  assign new_n1276 = pf0 & new_n1275;
  assign new_n1277 = pi0 & new_n1276;
  assign new_n1278 = ~py & new_n1277;
  assign new_n1279 = ~pd0 & new_n1278;
  assign new_n1280 = ~pb0 & new_n1279;
  assign new_n1281 = ~pc0 & new_n1280;
  assign new_n1282 = ~pt & new_n1281;
  assign new_n1283 = ~px & new_n1282;
  assign new_n1284 = ~ph & new_n678;
  assign new_n1285 = ~pe0 & new_n1284;
  assign new_n1286 = ~po & new_n1285;
  assign new_n1287 = ~pm & new_n1286;
  assign new_n1288 = ~py & new_n1287;
  assign new_n1289 = pk0 & new_n1288;
  assign new_n1290 = ~pg0 & new_n1289;
  assign new_n1291 = ~pd0 & new_n1290;
  assign new_n1292 = pi0 & new_n1291;
  assign new_n1293 = ~pi & new_n119;
  assign new_n1294 = ~pn & new_n1293;
  assign new_n1295 = ~ph & new_n1294;
  assign new_n1296 = ~pe0 & new_n1295;
  assign new_n1297 = pk0 & new_n1296;
  assign new_n1298 = ~pm & new_n1297;
  assign new_n1299 = pj0 & new_n1298;
  assign new_n1300 = ~pd0 & new_n1299;
  assign new_n1301 = ~pi0 & new_n1300;
  assign new_n1302 = ~pb0 & new_n1301;
  assign new_n1303 = ~pc0 & new_n1302;
  assign new_n1304 = pv & new_n623;
  assign new_n1305 = ~py & new_n1304;
  assign new_n1306 = ~pc0 & new_n1305;
  assign new_n1307 = pi0 & new_n1306;
  assign new_n1308 = ~pi0 & new_n623;
  assign new_n1309 = pj0 & new_n1308;
  assign new_n1310 = ~pc0 & new_n1309;
  assign new_n1311 = ~pd0 & new_n1310;
  assign new_n1312 = ~py & new_n949;
  assign new_n1313 = pf0 & new_n1312;
  assign new_n1314 = pi0 & new_n1313;
  assign new_n1315 = ~pc0 & new_n1314;
  assign new_n1316 = ~pd0 & new_n1315;
  assign new_n1317 = ~px & new_n1316;
  assign new_n1318 = ~pb0 & new_n1317;
  assign new_n1319 = ~pm & new_n680;
  assign new_n1320 = ~py & new_n1319;
  assign new_n1321 = po & new_n1320;
  assign new_n1322 = pi0 & new_n1321;
  assign new_n1323 = pv & new_n1322;
  assign new_n1324 = pu & new_n726;
  assign new_n1325 = ~pv & new_n1324;
  assign new_n1326 = ~pi0 & new_n1325;
  assign new_n1327 = pj0 & new_n1326;
  assign new_n1328 = ~pc0 & new_n1327;
  assign new_n1329 = pd0 & new_n1328;
  assign new_n1330 = ~ph & ~pj;
  assign new_n1331 = ~pf & new_n1330;
  assign new_n1332 = ~pg & new_n1331;
  assign new_n1333 = ~pe & new_n1332;
  assign new_n1334 = ~pa0 & new_n1333;
  assign new_n1335 = ~pk & new_n1334;
  assign new_n1336 = pk0 & new_n1335;
  assign new_n1337 = ~pg0 & new_n1336;
  assign new_n1338 = ~pv & new_n1337;
  assign new_n1339 = ~py & new_n1338;
  assign new_n1340 = ~pc0 & new_n1339;
  assign new_n1341 = pd0 & new_n1340;
  assign new_n1342 = ~pb0 & new_n1341;
  assign new_n1343 = ~pr & new_n1342;
  assign new_n1344 = ~px & new_n1343;
  assign new_n1345 = ~pn & new_n1344;
  assign new_n1346 = ~pq & new_n1345;
  assign new_n1347 = pf0 & new_n501;
  assign new_n1348 = ~pm & new_n1347;
  assign new_n1349 = ~py & new_n1348;
  assign new_n1350 = pk & new_n1349;
  assign new_n1351 = pv & new_n1350;
  assign new_n1352 = ~pc0 & new_n1351;
  assign new_n1353 = pi0 & new_n1352;
  assign new_n1354 = ~px & new_n1353;
  assign new_n1355 = ~pb0 & new_n1354;
  assign new_n1356 = pk & new_n1009;
  assign new_n1357 = pf0 & new_n1356;
  assign new_n1358 = ~ps & new_n1357;
  assign new_n1359 = ~py & new_n1358;
  assign new_n1360 = pd & new_n1359;
  assign new_n1361 = ~pd0 & new_n1360;
  assign new_n1362 = pi0 & new_n1361;
  assign new_n1363 = ~pb0 & new_n1362;
  assign new_n1364 = ~pc0 & new_n1363;
  assign new_n1365 = ~pi & new_n207;
  assign new_n1366 = ~pq & new_n1365;
  assign new_n1367 = ~ph & new_n1366;
  assign new_n1368 = ~pe0 & new_n1367;
  assign new_n1369 = ~po & new_n1368;
  assign new_n1370 = ~pm & new_n1369;
  assign new_n1371 = ~py & new_n1370;
  assign new_n1372 = pi0 & new_n1371;
  assign new_n1373 = pk0 & new_n1372;
  assign new_n1374 = ~pc0 & new_n1373;
  assign new_n1375 = ~pd0 & new_n1374;
  assign new_n1376 = ~ph & new_n559;
  assign new_n1377 = ~pe0 & new_n1376;
  assign new_n1378 = ~pg0 & new_n1377;
  assign new_n1379 = ~pm & new_n1378;
  assign new_n1380 = pk0 & new_n1379;
  assign new_n1381 = ~pi0 & new_n1380;
  assign new_n1382 = pj0 & new_n1381;
  assign new_n1383 = ~pc0 & new_n1382;
  assign new_n1384 = ~pd0 & new_n1383;
  assign new_n1385 = pf0 & new_n360;
  assign new_n1386 = ~pm & new_n1385;
  assign new_n1387 = pk & new_n1386;
  assign new_n1388 = ~pa0 & new_n1387;
  assign new_n1389 = ~po & new_n1388;
  assign new_n1390 = ~pc0 & new_n1389;
  assign new_n1391 = ~py & new_n1390;
  assign new_n1392 = ~py & new_n927;
  assign new_n1393 = pi0 & new_n1392;
  assign new_n1394 = pv & new_n1393;
  assign new_n1395 = ~pb0 & new_n1394;
  assign new_n1396 = ~pc0 & new_n1395;
  assign new_n1397 = pv & new_n1313;
  assign new_n1398 = ~pc0 & new_n1397;
  assign new_n1399 = pi0 & new_n1398;
  assign new_n1400 = ~px & new_n1399;
  assign new_n1401 = ~pb0 & new_n1400;
  assign new_n1402 = pv & new_n1319;
  assign new_n1403 = po & new_n1402;
  assign new_n1404 = ~pi0 & new_n1403;
  assign new_n1405 = pj0 & new_n1404;
  assign new_n1406 = ~py & new_n1324;
  assign new_n1407 = pi0 & new_n1406;
  assign new_n1408 = ~pv & new_n1407;
  assign new_n1409 = ~pc0 & new_n1408;
  assign new_n1410 = pd0 & new_n1409;
  assign new_n1411 = ~pk & new_n63;
  assign new_n1412 = ~pc0 & new_n1411;
  assign new_n1413 = ~pd0 & new_n1412;
  assign new_n1414 = ~pi0 & new_n1413;
  assign new_n1415 = pj0 & new_n1414;
  assign new_n1416 = ~px & new_n1415;
  assign new_n1417 = ~pb0 & new_n1416;
  assign new_n1418 = ~pr & new_n1417;
  assign new_n1419 = ~pn & new_n1418;
  assign new_n1420 = ~pq & new_n1419;
  assign new_n1421 = ~pi & new_n1420;
  assign new_n1422 = ~pj & new_n1421;
  assign new_n1423 = ~ps & new_n1269;
  assign new_n1424 = pi0 & new_n1423;
  assign new_n1425 = pd & new_n1424;
  assign new_n1426 = ~pc0 & new_n1425;
  assign new_n1427 = ~pd0 & new_n1426;
  assign new_n1428 = pj0 & new_n1276;
  assign new_n1429 = pv & new_n1428;
  assign new_n1430 = ~pi0 & new_n1429;
  assign new_n1431 = ~pb0 & new_n1430;
  assign new_n1432 = ~pc0 & new_n1431;
  assign new_n1433 = ~pt & new_n1432;
  assign new_n1434 = ~px & new_n1433;
  assign new_n1435 = ~pa0 & new_n1287;
  assign new_n1436 = ~pg0 & new_n1435;
  assign new_n1437 = ~py & new_n1436;
  assign new_n1438 = ~pd0 & new_n1437;
  assign new_n1439 = pk0 & new_n1438;
  assign new_n1440 = ~py & new_n1296;
  assign new_n1441 = ~pm & new_n1440;
  assign new_n1442 = pk0 & new_n1441;
  assign new_n1443 = ~pd0 & new_n1442;
  assign new_n1444 = pi0 & new_n1443;
  assign new_n1445 = ~pb0 & new_n1444;
  assign new_n1446 = ~pc0 & new_n1445;
  assign new_n1447 = pn & new_n947;
  assign new_n1448 = pc & new_n1447;
  assign new_n1449 = ~po & new_n1448;
  assign new_n1450 = ~py & new_n1449;
  assign new_n1451 = ~pa0 & new_n1450;
  assign new_n1452 = ~pv & new_n1451;
  assign new_n1453 = ~pc0 & new_n1452;
  assign new_n1454 = pd0 & new_n1453;
  assign new_n1455 = ~px & new_n1454;
  assign new_n1456 = ~pb0 & new_n1455;
  assign new_n1457 = ~pd0 & new_n1392;
  assign new_n1458 = pi0 & new_n1457;
  assign new_n1459 = ~pb0 & new_n1458;
  assign new_n1460 = ~pc0 & new_n1459;
  assign new_n1461 = pj0 & new_n949;
  assign new_n1462 = pf0 & new_n1461;
  assign new_n1463 = ~pi0 & new_n1462;
  assign new_n1464 = ~pc0 & new_n1463;
  assign new_n1465 = ~pd0 & new_n1464;
  assign new_n1466 = ~px & new_n1465;
  assign new_n1467 = ~pb0 & new_n1466;
  assign new_n1468 = pz & new_n1222;
  assign new_n1469 = ph0 & new_n1468;
  assign new_n1470 = ~py & new_n1469;
  assign new_n1471 = ~po & new_n1470;
  assign new_n1472 = pi0 & new_n1471;
  assign new_n1473 = pv & new_n1472;
  assign new_n1474 = pu & new_n1222;
  assign new_n1475 = ~po & new_n1474;
  assign new_n1476 = pj0 & new_n1475;
  assign new_n1477 = ~pv & new_n1476;
  assign new_n1478 = pd0 & new_n1477;
  assign new_n1479 = ~pi0 & new_n1478;
  assign new_n1480 = ~py & new_n62;
  assign new_n1481 = ~po & new_n1480;
  assign new_n1482 = ~pc0 & new_n1481;
  assign new_n1483 = ~pd0 & new_n1482;
  assign new_n1484 = pi0 & new_n1483;
  assign new_n1485 = pk0 & new_n1484;
  assign new_n1486 = ~px & new_n1485;
  assign new_n1487 = ~pb0 & new_n1486;
  assign new_n1488 = ~pr & new_n1487;
  assign new_n1489 = pn & new_n1488;
  assign new_n1490 = ~pq & new_n1489;
  assign new_n1491 = ~pi & new_n1490;
  assign new_n1492 = ~pj & new_n1491;
  assign new_n1493 = pi0 & new_n1350;
  assign new_n1494 = ~pc0 & new_n1493;
  assign new_n1495 = ~pd0 & new_n1494;
  assign new_n1496 = ~px & new_n1495;
  assign new_n1497 = ~pb0 & new_n1496;
  assign new_n1498 = pv & new_n1358;
  assign new_n1499 = pd & new_n1498;
  assign new_n1500 = ~pi0 & new_n1499;
  assign new_n1501 = pj0 & new_n1500;
  assign new_n1502 = ~pb0 & new_n1501;
  assign new_n1503 = ~pc0 & new_n1502;
  assign new_n1504 = ~pa0 & new_n1370;
  assign new_n1505 = pk0 & new_n1504;
  assign new_n1506 = ~py & new_n1505;
  assign new_n1507 = ~pc0 & new_n1506;
  assign new_n1508 = ~pd0 & new_n1507;
  assign new_n1509 = ~py & new_n1377;
  assign new_n1510 = ~pm & new_n1509;
  assign new_n1511 = ~pg0 & new_n1510;
  assign new_n1512 = pi0 & new_n1511;
  assign new_n1513 = pk0 & new_n1512;
  assign new_n1514 = ~pc0 & new_n1513;
  assign new_n1515 = ~pd0 & new_n1514;
  assign new_n1516 = pc & new_n948;
  assign new_n1517 = ~pk & new_n1516;
  assign new_n1518 = ~py & new_n1517;
  assign new_n1519 = ~pa0 & new_n1518;
  assign new_n1520 = ~pv & new_n1519;
  assign new_n1521 = ~pc0 & new_n1520;
  assign new_n1522 = pd0 & new_n1521;
  assign new_n1523 = ~px & new_n1522;
  assign new_n1524 = ~pb0 & new_n1523;
  assign new_n1525 = pv & new_n927;
  assign new_n1526 = ~pi0 & new_n1525;
  assign new_n1527 = pj0 & new_n1526;
  assign new_n1528 = ~pb0 & new_n1527;
  assign new_n1529 = ~pc0 & new_n1528;
  assign new_n1530 = pv & new_n949;
  assign new_n1531 = pf0 & new_n1530;
  assign new_n1532 = pj0 & new_n1531;
  assign new_n1533 = ~pc0 & new_n1532;
  assign new_n1534 = ~pi0 & new_n1533;
  assign new_n1535 = ~px & new_n1534;
  assign new_n1536 = ~pb0 & new_n1535;
  assign new_n1537 = pv & new_n1469;
  assign new_n1538 = ~po & new_n1537;
  assign new_n1539 = ~pi0 & new_n1538;
  assign new_n1540 = pj0 & new_n1539;
  assign new_n1541 = ~pv & new_n1475;
  assign new_n1542 = ~py & new_n1541;
  assign new_n1543 = pd0 & new_n1542;
  assign new_n1544 = pi0 & new_n1543;
  assign new_n1545 = ~pv & new_n1333;
  assign new_n1546 = ~py & new_n1545;
  assign new_n1547 = ~pa0 & new_n1546;
  assign new_n1548 = pk0 & new_n1547;
  assign new_n1549 = pd & new_n1548;
  assign new_n1550 = ~ps & new_n1549;
  assign new_n1551 = ~pg0 & new_n1550;
  assign new_n1552 = ~pc0 & new_n1551;
  assign new_n1553 = pd0 & new_n1552;
  assign new_n1554 = ~pb0 & new_n1553;
  assign new_n1555 = ~pr & new_n1554;
  assign new_n1556 = ~px & new_n1555;
  assign new_n1557 = ~pn & new_n1556;
  assign new_n1558 = ~pq & new_n1557;
  assign new_n1559 = ~ps & new_n314;
  assign new_n1560 = ~pg0 & new_n1559;
  assign new_n1561 = ~py & new_n1560;
  assign new_n1562 = pi0 & new_n1561;
  assign new_n1563 = ~pj0 & new_n1562;
  assign new_n1564 = pk0 & new_n1563;
  assign new_n1565 = pd & new_n1564;
  assign new_n1566 = ~pc0 & new_n1565;
  assign new_n1567 = ~pd0 & new_n1566;
  assign new_n1568 = ~pb0 & new_n1567;
  assign new_n1569 = ~pr & new_n1568;
  assign new_n1570 = ~px & new_n1569;
  assign new_n1571 = ~pn & new_n1570;
  assign new_n1572 = ~pq & new_n1571;
  assign new_n1573 = ~pi0 & new_n62;
  assign new_n1574 = pj0 & new_n1573;
  assign new_n1575 = pk0 & new_n1574;
  assign new_n1576 = ~px & new_n1575;
  assign new_n1577 = ~pb0 & new_n1576;
  assign new_n1578 = ~pc0 & new_n1577;
  assign new_n1579 = ~pd0 & new_n1578;
  assign new_n1580 = ~pr & new_n1579;
  assign new_n1581 = ~pt & new_n1580;
  assign new_n1582 = ~pq & new_n1581;
  assign new_n1583 = ~pl & new_n1582;
  assign new_n1584 = ~pn & new_n1583;
  assign new_n1585 = ~pi & new_n1584;
  assign new_n1586 = ~pj & new_n1585;
  assign new_n1587 = ~pb & new_n79;
  assign new_n1588 = ~pf0 & new_n1587;
  assign new_n1589 = ~pj0 & new_n1588;
  assign new_n1590 = pk0 & new_n1589;
  assign new_n1591 = ~pg0 & new_n1590;
  assign new_n1592 = ~py & new_n1591;
  assign new_n1593 = ~pd0 & new_n1592;
  assign new_n1594 = pi0 & new_n1593;
  assign new_n1595 = ~pc0 & new_n1594;
  assign new_n1596 = ~px & new_n1595;
  assign new_n1597 = ~pb0 & new_n1596;
  assign new_n1598 = ~pq & new_n1597;
  assign new_n1599 = ~pr & new_n1598;
  assign new_n1600 = ~pk & new_n1480;
  assign new_n1601 = ~pc0 & new_n1600;
  assign new_n1602 = ~pd0 & new_n1601;
  assign new_n1603 = pi0 & new_n1602;
  assign new_n1604 = pk0 & new_n1603;
  assign new_n1605 = ~px & new_n1604;
  assign new_n1606 = ~pb0 & new_n1605;
  assign new_n1607 = ~pr & new_n1606;
  assign new_n1608 = ~pn & new_n1607;
  assign new_n1609 = ~pq & new_n1608;
  assign new_n1610 = ~pi & new_n1609;
  assign new_n1611 = ~pj & new_n1610;
  assign new_n1612 = ~py & new_n138;
  assign new_n1613 = ~po & new_n1612;
  assign new_n1614 = ~pd0 & new_n1613;
  assign new_n1615 = pi0 & new_n1614;
  assign new_n1616 = ~pj0 & new_n1615;
  assign new_n1617 = pk0 & new_n1616;
  assign new_n1618 = ~pb0 & new_n1617;
  assign new_n1619 = ~pc0 & new_n1618;
  assign new_n1620 = ~px & new_n1619;
  assign new_n1621 = ~pq & new_n1620;
  assign new_n1622 = ~pr & new_n1621;
  assign new_n1623 = ~pj & new_n1622;
  assign new_n1624 = pn & new_n1623;
  assign new_n1625 = ~pg0 & new_n62;
  assign new_n1626 = ~py & new_n1625;
  assign new_n1627 = ~pa0 & new_n1626;
  assign new_n1628 = ~pm & new_n1627;
  assign new_n1629 = ~pd0 & new_n1628;
  assign new_n1630 = pk0 & new_n1629;
  assign new_n1631 = ~pc0 & new_n1630;
  assign new_n1632 = ~px & new_n1631;
  assign new_n1633 = ~pb0 & new_n1632;
  assign new_n1634 = ~pn & new_n1633;
  assign new_n1635 = ~pq & new_n1634;
  assign new_n1636 = ~pi & new_n678;
  assign new_n1637 = ~pm & new_n1636;
  assign new_n1638 = ~pe0 & new_n1637;
  assign new_n1639 = ~po & new_n1638;
  assign new_n1640 = ~pf0 & new_n1639;
  assign new_n1641 = ~pa0 & new_n1640;
  assign new_n1642 = ~pv & new_n1641;
  assign new_n1643 = ~py & new_n1642;
  assign new_n1644 = ~pj0 & new_n1643;
  assign new_n1645 = pk0 & new_n1644;
  assign new_n1646 = ~ph & new_n279;
  assign new_n1647 = ~pq & new_n1646;
  assign new_n1648 = ~pc & new_n1647;
  assign new_n1649 = ~po & new_n1648;
  assign new_n1650 = ~pe0 & new_n1649;
  assign new_n1651 = ~py & new_n1650;
  assign new_n1652 = ~pa0 & new_n1651;
  assign new_n1653 = ~pv & new_n1652;
  assign new_n1654 = pk0 & new_n1653;
  assign new_n1655 = ~pg0 & new_n1654;
  assign new_n1656 = ~pb0 & new_n1655;
  assign new_n1657 = ~pc0 & new_n1656;
  assign new_n1658 = pj0 & new_n1348;
  assign new_n1659 = pk & new_n1658;
  assign new_n1660 = ~pi0 & new_n1659;
  assign new_n1661 = ~pc0 & new_n1660;
  assign new_n1662 = ~pd0 & new_n1661;
  assign new_n1663 = ~px & new_n1662;
  assign new_n1664 = ~pb0 & new_n1663;
  assign new_n1665 = ~pv & new_n1435;
  assign new_n1666 = ~py & new_n1665;
  assign new_n1667 = pk0 & new_n1666;
  assign new_n1668 = ~pg0 & new_n1667;
  assign new_n1669 = ~pa0 & new_n1296;
  assign new_n1670 = ~pm & new_n1669;
  assign new_n1671 = ~py & new_n1670;
  assign new_n1672 = ~pd0 & new_n1671;
  assign new_n1673 = pk0 & new_n1672;
  assign new_n1674 = ~pb0 & new_n1673;
  assign new_n1675 = ~pc0 & new_n1674;
  assign new_n1676 = ~pj & ~pl;
  assign new_n1677 = ~pf & new_n1676;
  assign new_n1678 = ~pg & new_n1677;
  assign new_n1679 = ~pe & new_n1678;
  assign new_n1680 = ~pv & new_n1679;
  assign new_n1681 = ~py & new_n1680;
  assign new_n1682 = ~pa0 & new_n1681;
  assign new_n1683 = pd0 & new_n1682;
  assign new_n1684 = ~pj0 & new_n1683;
  assign new_n1685 = pk0 & new_n1684;
  assign new_n1686 = ~pg0 & new_n1685;
  assign new_n1687 = ~pb0 & new_n1686;
  assign new_n1688 = ~pc0 & new_n1687;
  assign new_n1689 = ~px & new_n1688;
  assign new_n1690 = ~pr & new_n1689;
  assign new_n1691 = ~pt & new_n1690;
  assign new_n1692 = ~pn & new_n1691;
  assign new_n1693 = ~pq & new_n1692;
  assign new_n1694 = pk0 & new_n138;
  assign new_n1695 = ~py & new_n1694;
  assign new_n1696 = ~pa0 & new_n1695;
  assign new_n1697 = ~pb0 & new_n1696;
  assign new_n1698 = ~pc0 & new_n1697;
  assign new_n1699 = ~pd0 & new_n1698;
  assign new_n1700 = ~pj0 & new_n1699;
  assign new_n1701 = ~pt & new_n1700;
  assign new_n1702 = ~px & new_n1701;
  assign new_n1703 = ~pr & new_n1702;
  assign new_n1704 = ~pn & new_n1703;
  assign new_n1705 = ~pq & new_n1704;
  assign new_n1706 = ~pj & new_n1705;
  assign new_n1707 = ~pl & new_n1706;
  assign new_n1708 = ~pv & new_n167;
  assign new_n1709 = ~py & new_n1708;
  assign new_n1710 = ~pa0 & new_n1709;
  assign new_n1711 = ~po & new_n1710;
  assign new_n1712 = pk0 & new_n1711;
  assign new_n1713 = ~pg0 & new_n1712;
  assign new_n1714 = ~pj0 & new_n1713;
  assign new_n1715 = ~pb0 & new_n1714;
  assign new_n1716 = ~pc0 & new_n1715;
  assign new_n1717 = ~pr & new_n1716;
  assign new_n1718 = ~px & new_n1717;
  assign new_n1719 = ~pj0 & new_n1254;
  assign new_n1720 = pk0 & new_n1719;
  assign new_n1721 = ~py & new_n1720;
  assign new_n1722 = ~pa0 & new_n1721;
  assign new_n1723 = ~pc0 & new_n1722;
  assign new_n1724 = ~pd0 & new_n1723;
  assign new_n1725 = ~pb0 & new_n1724;
  assign new_n1726 = ~pr & new_n1725;
  assign new_n1727 = ~px & new_n1726;
  assign new_n1728 = ~pn & new_n1727;
  assign new_n1729 = ~pq & new_n1728;
  assign new_n1730 = ~pk & new_n1625;
  assign new_n1731 = ~pd0 & new_n1730;
  assign new_n1732 = ~pi0 & new_n1731;
  assign new_n1733 = pj0 & new_n1732;
  assign new_n1734 = pk0 & new_n1733;
  assign new_n1735 = ~pb0 & new_n1734;
  assign new_n1736 = ~pc0 & new_n1735;
  assign new_n1737 = ~px & new_n1736;
  assign new_n1738 = ~pq & new_n1737;
  assign new_n1739 = ~pr & new_n1738;
  assign new_n1740 = ~pj & new_n1739;
  assign new_n1741 = ~pn & new_n1740;
  assign new_n1742 = ~pd0 & new_n1481;
  assign new_n1743 = pi0 & new_n1742;
  assign new_n1744 = pk0 & new_n1743;
  assign new_n1745 = ~pg0 & new_n1744;
  assign new_n1746 = ~pb0 & new_n1745;
  assign new_n1747 = ~pc0 & new_n1746;
  assign new_n1748 = ~px & new_n1747;
  assign new_n1749 = ~pq & new_n1748;
  assign new_n1750 = ~pr & new_n1749;
  assign new_n1751 = ~pj & new_n1750;
  assign new_n1752 = pn & new_n1751;
  assign new_n1753 = ~py & new_n63;
  assign new_n1754 = ~pa0 & new_n1753;
  assign new_n1755 = ~pm & new_n1754;
  assign new_n1756 = ~pc0 & new_n1755;
  assign new_n1757 = ~pd0 & new_n1756;
  assign new_n1758 = ~pb0 & new_n1757;
  assign new_n1759 = ~pq & new_n1758;
  assign new_n1760 = ~px & new_n1759;
  assign new_n1761 = ~pi & new_n1760;
  assign new_n1762 = ~pn & new_n1761;
  assign new_n1763 = ~pc0 & ~pj0;
  assign new_n1764 = ~px & new_n1763;
  assign new_n1765 = ~pb0 & new_n1764;
  assign new_n1766 = ~pq & new_n1765;
  assign new_n1767 = ~pm & new_n1766;
  assign new_n1768 = ~pe0 & new_n1767;
  assign new_n1769 = ~po & new_n1768;
  assign new_n1770 = ~pf0 & new_n1769;
  assign new_n1771 = ~pa0 & new_n1770;
  assign new_n1772 = ~pv & new_n1771;
  assign new_n1773 = ~py & new_n1772;
  assign new_n1774 = pk0 & new_n1773;
  assign new_n1775 = ~pg0 & new_n1774;
  assign new_n1776 = ~ph & new_n219;
  assign new_n1777 = ~pi & new_n1776;
  assign new_n1778 = ~pc & new_n1777;
  assign new_n1779 = ~po & new_n1778;
  assign new_n1780 = ~pe0 & new_n1779;
  assign new_n1781 = ~py & new_n1780;
  assign new_n1782 = ~pa0 & new_n1781;
  assign new_n1783 = ~pv & new_n1782;
  assign new_n1784 = ~pc0 & new_n1783;
  assign new_n1785 = pk0 & new_n1784;
  assign new_n1786 = ~px & new_n1785;
  assign new_n1787 = ~pb0 & new_n1786;
  assign new_n1788 = ~ps & new_n1267;
  assign new_n1789 = pk & new_n1788;
  assign new_n1790 = pd & new_n1789;
  assign new_n1791 = ~pi0 & new_n1790;
  assign new_n1792 = pj0 & new_n1791;
  assign new_n1793 = ~pc0 & new_n1792;
  assign new_n1794 = ~pd0 & new_n1793;
  assign new_n1795 = ~pv & new_n1504;
  assign new_n1796 = ~py & new_n1795;
  assign new_n1797 = ~pc0 & new_n1796;
  assign new_n1798 = pk0 & new_n1797;
  assign new_n1799 = ~pa0 & new_n1377;
  assign new_n1800 = ~pm & new_n1799;
  assign new_n1801 = ~py & new_n1800;
  assign new_n1802 = pk0 & new_n1801;
  assign new_n1803 = ~pg0 & new_n1802;
  assign new_n1804 = ~pc0 & new_n1803;
  assign new_n1805 = ~pd0 & new_n1804;
  assign new_n1806 = ~ps & new_n138;
  assign new_n1807 = ~py & new_n1806;
  assign new_n1808 = ~pa0 & new_n1807;
  assign new_n1809 = ~pd0 & new_n1808;
  assign new_n1810 = ~pj0 & new_n1809;
  assign new_n1811 = pk0 & new_n1810;
  assign new_n1812 = pd & new_n1811;
  assign new_n1813 = ~pb0 & new_n1812;
  assign new_n1814 = ~pc0 & new_n1813;
  assign new_n1815 = ~px & new_n1814;
  assign new_n1816 = ~pq & new_n1815;
  assign new_n1817 = ~pr & new_n1816;
  assign new_n1818 = ~pj & new_n1817;
  assign new_n1819 = ~pn & new_n1818;
  assign new_n1820 = ~pv & new_n1254;
  assign new_n1821 = ~py & new_n1820;
  assign new_n1822 = ~pa0 & new_n1821;
  assign new_n1823 = ~po & new_n1822;
  assign new_n1824 = ~pj0 & new_n1823;
  assign new_n1825 = pk0 & new_n1824;
  assign new_n1826 = ~pc0 & new_n1825;
  assign new_n1827 = ~px & new_n1826;
  assign new_n1828 = ~pb0 & new_n1827;
  assign new_n1829 = ~pq & new_n1828;
  assign new_n1830 = ~pr & new_n1829;
  assign new_n1831 = ~pj & ~pn;
  assign new_n1832 = ~pf & new_n1831;
  assign new_n1833 = ~pg & new_n1832;
  assign new_n1834 = ~pe & new_n1833;
  assign new_n1835 = ~pa0 & new_n1834;
  assign new_n1836 = ~pk & new_n1835;
  assign new_n1837 = pk0 & new_n1836;
  assign new_n1838 = ~pg0 & new_n1837;
  assign new_n1839 = ~pv & new_n1838;
  assign new_n1840 = ~py & new_n1839;
  assign new_n1841 = pd0 & new_n1840;
  assign new_n1842 = ~pj0 & new_n1841;
  assign new_n1843 = ~pc0 & new_n1842;
  assign new_n1844 = ~px & new_n1843;
  assign new_n1845 = ~pb0 & new_n1844;
  assign new_n1846 = ~pq & new_n1845;
  assign new_n1847 = ~pr & new_n1846;
  assign new_n1848 = ~pd0 & new_n1600;
  assign new_n1849 = pi0 & new_n1848;
  assign new_n1850 = pk0 & new_n1849;
  assign new_n1851 = ~pg0 & new_n1850;
  assign new_n1852 = ~pb0 & new_n1851;
  assign new_n1853 = ~pc0 & new_n1852;
  assign new_n1854 = ~px & new_n1853;
  assign new_n1855 = ~pq & new_n1854;
  assign new_n1856 = ~pr & new_n1855;
  assign new_n1857 = ~pj & new_n1856;
  assign new_n1858 = ~pn & new_n1857;
  assign new_n1859 = ~py & new_n314;
  assign new_n1860 = ~po & new_n1859;
  assign new_n1861 = pi0 & new_n1860;
  assign new_n1862 = ~pj0 & new_n1861;
  assign new_n1863 = pk0 & new_n1862;
  assign new_n1864 = ~pg0 & new_n1863;
  assign new_n1865 = ~pc0 & new_n1864;
  assign new_n1866 = ~pd0 & new_n1865;
  assign new_n1867 = ~pb0 & new_n1866;
  assign new_n1868 = ~pr & new_n1867;
  assign new_n1869 = ~px & new_n1868;
  assign new_n1870 = pn & new_n1869;
  assign new_n1871 = ~pq & new_n1870;
  assign new_n1872 = pj0 & new_n195;
  assign new_n1873 = pk0 & new_n1872;
  assign new_n1874 = ~pg0 & new_n1873;
  assign new_n1875 = ~po & new_n1874;
  assign new_n1876 = ~pd0 & new_n1875;
  assign new_n1877 = ~pi0 & new_n1876;
  assign new_n1878 = ~pc0 & new_n1877;
  assign new_n1879 = ~px & new_n1878;
  assign new_n1880 = ~pb0 & new_n1879;
  assign new_n1881 = ~pq & new_n1880;
  assign new_n1882 = ~pr & new_n1881;
  assign new_n1883 = ~py & new_n1058;
  assign new_n1884 = ~pa0 & new_n1883;
  assign new_n1885 = ~po & new_n1884;
  assign new_n1886 = ~pm & new_n1885;
  assign new_n1887 = pk0 & new_n1886;
  assign new_n1888 = ~pv & new_n1887;
  assign new_n1889 = pd0 & new_n1888;
  assign new_n1890 = ~pb0 & new_n1889;
  assign new_n1891 = ~pc0 & new_n1890;
  assign new_n1892 = ~pq & new_n1891;
  assign new_n1893 = ~px & new_n1892;
  assign new_n1894 = ~pn & new_n1776;
  assign new_n1895 = ~pc & new_n1894;
  assign new_n1896 = ~pa0 & new_n1895;
  assign new_n1897 = ~pe0 & new_n1896;
  assign new_n1898 = ~pv & new_n1897;
  assign new_n1899 = ~py & new_n1898;
  assign new_n1900 = ~pg0 & new_n1899;
  assign new_n1901 = ~pc0 & new_n1900;
  assign new_n1902 = pk0 & new_n1901;
  assign new_n1903 = ~px & new_n1902;
  assign new_n1904 = ~pb0 & new_n1903;
  assign new_n1905 = pv & new_n1276;
  assign new_n1906 = ~py & new_n1905;
  assign new_n1907 = pi0 & new_n1906;
  assign new_n1908 = ~pb0 & new_n1907;
  assign new_n1909 = ~pc0 & new_n1908;
  assign new_n1910 = ~pt & new_n1909;
  assign new_n1911 = ~px & new_n1910;
  assign new_n1912 = ~py & new_n1516;
  assign new_n1913 = ~pa0 & new_n1912;
  assign new_n1914 = ~ps & new_n1913;
  assign new_n1915 = ~pv & new_n1914;
  assign new_n1916 = pd & new_n1915;
  assign new_n1917 = ~pc0 & new_n1916;
  assign new_n1918 = pd0 & new_n1917;
  assign new_n1919 = ~px & new_n1918;
  assign new_n1920 = ~pb0 & new_n1919;
  assign new_n1921 = pk0 & new_n1671;
  assign new_n1922 = ~pv & new_n1921;
  assign new_n1923 = ~pb0 & new_n1922;
  assign new_n1924 = ~pc0 & new_n1923;
  assign new_n1925 = pj0 & new_n1142;
  assign new_n1926 = ~pi0 & new_n1925;
  assign new_n1927 = ~pd0 & new_n1926;
  assign new_n1928 = ph0 & new_n1927;
  assign new_n1929 = ~pb0 & new_n1928;
  assign new_n1930 = ~pc0 & new_n1929;
  assign new_n1931 = ~pv & new_n1834;
  assign new_n1932 = ~py & new_n1931;
  assign new_n1933 = ~pa0 & new_n1932;
  assign new_n1934 = pk0 & new_n1933;
  assign new_n1935 = pd & new_n1934;
  assign new_n1936 = ~ps & new_n1935;
  assign new_n1937 = ~pg0 & new_n1936;
  assign new_n1938 = pd0 & new_n1937;
  assign new_n1939 = ~pj0 & new_n1938;
  assign new_n1940 = ~pc0 & new_n1939;
  assign new_n1941 = ~px & new_n1940;
  assign new_n1942 = ~pb0 & new_n1941;
  assign new_n1943 = ~pq & new_n1942;
  assign new_n1944 = ~pr & new_n1943;
  assign new_n1945 = ~pc0 & new_n317;
  assign new_n1946 = ~pd0 & new_n1945;
  assign new_n1947 = ~pj0 & new_n1946;
  assign new_n1948 = pk0 & new_n1947;
  assign new_n1949 = ~px & new_n1948;
  assign new_n1950 = ~pb0 & new_n1949;
  assign new_n1951 = ~pt & new_n1950;
  assign new_n1952 = ~pq & new_n1951;
  assign new_n1953 = ~pr & new_n1952;
  assign new_n1954 = ~pl & new_n1953;
  assign new_n1955 = ~pn & new_n1954;
  assign new_n1956 = ~pg0 & new_n167;
  assign new_n1957 = ~py & new_n1956;
  assign new_n1958 = ~pa0 & new_n1957;
  assign new_n1959 = ~po & new_n1958;
  assign new_n1960 = ~pj0 & new_n1959;
  assign new_n1961 = pk0 & new_n1960;
  assign new_n1962 = ~pd0 & new_n1961;
  assign new_n1963 = ~pb0 & new_n1962;
  assign new_n1964 = ~pc0 & new_n1963;
  assign new_n1965 = ~pr & new_n1964;
  assign new_n1966 = ~px & new_n1965;
  assign new_n1967 = pi0 & new_n1254;
  assign new_n1968 = ~pj0 & new_n1967;
  assign new_n1969 = pk0 & new_n1968;
  assign new_n1970 = ~py & new_n1969;
  assign new_n1971 = ~pc0 & new_n1970;
  assign new_n1972 = ~pd0 & new_n1971;
  assign new_n1973 = ~pb0 & new_n1972;
  assign new_n1974 = ~pr & new_n1973;
  assign new_n1975 = ~px & new_n1974;
  assign new_n1976 = ~pn & new_n1975;
  assign new_n1977 = ~pq & new_n1976;
  assign new_n1978 = ~pk & new_n1612;
  assign new_n1979 = ~pd0 & new_n1978;
  assign new_n1980 = pi0 & new_n1979;
  assign new_n1981 = ~pj0 & new_n1980;
  assign new_n1982 = pk0 & new_n1981;
  assign new_n1983 = ~pb0 & new_n1982;
  assign new_n1984 = ~pc0 & new_n1983;
  assign new_n1985 = ~px & new_n1984;
  assign new_n1986 = ~pq & new_n1985;
  assign new_n1987 = ~pr & new_n1986;
  assign new_n1988 = ~pj & new_n1987;
  assign new_n1989 = ~pn & new_n1988;
  assign new_n1990 = ~pa0 & new_n138;
  assign new_n1991 = ~po & new_n1990;
  assign new_n1992 = ~pd0 & new_n1991;
  assign new_n1993 = ~pj0 & new_n1992;
  assign new_n1994 = pk0 & new_n1993;
  assign new_n1995 = ~py & new_n1994;
  assign new_n1996 = ~pb0 & new_n1995;
  assign new_n1997 = ~pc0 & new_n1996;
  assign new_n1998 = ~px & new_n1997;
  assign new_n1999 = ~pq & new_n1998;
  assign new_n2000 = ~pr & new_n1999;
  assign new_n2001 = ~pj & new_n2000;
  assign new_n2002 = pn & new_n2001;
  assign new_n2003 = ~po & new_n1075;
  assign new_n2004 = ~pc0 & new_n2003;
  assign new_n2005 = ~pd0 & new_n2004;
  assign new_n2006 = ~pb0 & new_n2005;
  assign new_n2007 = ~pr & new_n2006;
  assign new_n2008 = ~px & new_n2007;
  assign new_n2009 = ~pi & new_n2008;
  assign new_n2010 = ~pq & new_n2009;
  assign new_n2011 = ~pq & ~ph;
  assign new_n2012 = ~pf & new_n2011;
  assign new_n2013 = ~pg & new_n2012;
  assign new_n2014 = ~pe & new_n2013;
  assign new_n2015 = ~py & new_n2014;
  assign new_n2016 = ~pa0 & new_n2015;
  assign new_n2017 = ~po & new_n2016;
  assign new_n2018 = ~pm & new_n2017;
  assign new_n2019 = ~pg0 & new_n2018;
  assign new_n2020 = ~pv & new_n2019;
  assign new_n2021 = pk0 & new_n2020;
  assign new_n2022 = ~pc0 & new_n2021;
  assign new_n2023 = pd0 & new_n2022;
  assign new_n2024 = ~px & new_n2023;
  assign new_n2025 = ~pb0 & new_n2024;
  assign new_n2026 = ~ph & new_n438;
  assign new_n2027 = ~pi & new_n2026;
  assign new_n2028 = ~pc & new_n2027;
  assign new_n2029 = ~pa0 & new_n2028;
  assign new_n2030 = ~pe0 & new_n2029;
  assign new_n2031 = ~pv & new_n2030;
  assign new_n2032 = ~py & new_n2031;
  assign new_n2033 = pk0 & new_n2032;
  assign new_n2034 = ~pb0 & new_n2033;
  assign new_n2035 = ~pc0 & new_n2034;
  assign new_n2036 = ~pr & new_n2035;
  assign new_n2037 = ~px & new_n2036;
  assign new_n2038 = pv & new_n1357;
  assign new_n2039 = ~py & new_n2038;
  assign new_n2040 = ~ps & new_n2039;
  assign new_n2041 = pi0 & new_n2040;
  assign new_n2042 = pd & new_n2041;
  assign new_n2043 = ~pb0 & new_n2042;
  assign new_n2044 = ~pc0 & new_n2043;
  assign new_n2045 = ~pj & new_n438;
  assign new_n2046 = ~pl & new_n2045;
  assign new_n2047 = pc & new_n2046;
  assign new_n2048 = ~py & new_n2047;
  assign new_n2049 = ~pa0 & new_n2048;
  assign new_n2050 = pd0 & new_n2049;
  assign new_n2051 = ~pv & new_n2050;
  assign new_n2052 = ~pc0 & new_n2051;
  assign new_n2053 = ~px & new_n2052;
  assign new_n2054 = ~pb0 & new_n2053;
  assign new_n2055 = ~pr & new_n2054;
  assign new_n2056 = ~pt & new_n2055;
  assign new_n2057 = ~pg0 & new_n1801;
  assign new_n2058 = ~pv & new_n2057;
  assign new_n2059 = ~pc0 & new_n2058;
  assign new_n2060 = pk0 & new_n2059;
  assign new_n2061 = pd0 & new_n1061;
  assign new_n2062 = pk0 & new_n2061;
  assign new_n2063 = pd & new_n2062;
  assign new_n2064 = ~ps & new_n2063;
  assign new_n2065 = ~pb0 & new_n2064;
  assign new_n2066 = ~pc0 & new_n2065;
  assign new_n2067 = ~px & new_n2066;
  assign new_n2068 = ~pq & new_n2067;
  assign new_n2069 = ~pr & new_n2068;
  assign new_n2070 = ~pj & new_n2069;
  assign new_n2071 = ~pn & new_n2070;
  assign new_n2072 = pd & new_n138;
  assign new_n2073 = ~ps & new_n2072;
  assign new_n2074 = ~py & new_n2073;
  assign new_n2075 = ~pd0 & new_n2074;
  assign new_n2076 = pi0 & new_n2075;
  assign new_n2077 = ~pj0 & new_n2076;
  assign new_n2078 = pk0 & new_n2077;
  assign new_n2079 = ~pb0 & new_n2078;
  assign new_n2080 = ~pc0 & new_n2079;
  assign new_n2081 = ~px & new_n2080;
  assign new_n2082 = ~pq & new_n2081;
  assign new_n2083 = ~pr & new_n2082;
  assign new_n2084 = ~pj & new_n2083;
  assign new_n2085 = ~pn & new_n2084;
  assign new_n2086 = pi0 & new_n62;
  assign new_n2087 = pk0 & new_n2086;
  assign new_n2088 = ~py & new_n2087;
  assign new_n2089 = ~px & new_n2088;
  assign new_n2090 = ~pb0 & new_n2089;
  assign new_n2091 = ~pc0 & new_n2090;
  assign new_n2092 = ~pd0 & new_n2091;
  assign new_n2093 = ~pr & new_n2092;
  assign new_n2094 = ~pt & new_n2093;
  assign new_n2095 = ~pq & new_n2094;
  assign new_n2096 = ~pl & new_n2095;
  assign new_n2097 = ~pn & new_n2096;
  assign new_n2098 = ~pi & new_n2097;
  assign new_n2099 = ~pj & new_n2098;
  assign new_n2100 = ~pg0 & new_n1588;
  assign new_n2101 = ~pv & new_n2100;
  assign new_n2102 = ~py & new_n2101;
  assign new_n2103 = ~pa0 & new_n2102;
  assign new_n2104 = ~pj0 & new_n2103;
  assign new_n2105 = pk0 & new_n2104;
  assign new_n2106 = ~pc0 & new_n2105;
  assign new_n2107 = ~px & new_n2106;
  assign new_n2108 = ~pb0 & new_n2107;
  assign new_n2109 = ~pq & new_n2108;
  assign new_n2110 = ~pr & new_n2109;
  assign new_n2111 = ~pk & new_n1990;
  assign new_n2112 = ~pd0 & new_n2111;
  assign new_n2113 = ~pj0 & new_n2112;
  assign new_n2114 = pk0 & new_n2113;
  assign new_n2115 = ~py & new_n2114;
  assign new_n2116 = ~pb0 & new_n2115;
  assign new_n2117 = ~pc0 & new_n2116;
  assign new_n2118 = ~px & new_n2117;
  assign new_n2119 = ~pq & new_n2118;
  assign new_n2120 = ~pr & new_n2119;
  assign new_n2121 = ~pj & new_n2120;
  assign new_n2122 = ~pn & new_n2121;
  assign new_n2123 = ~pa0 & new_n314;
  assign new_n2124 = ~po & new_n2123;
  assign new_n2125 = ~pj0 & new_n2124;
  assign new_n2126 = pk0 & new_n2125;
  assign new_n2127 = ~pg0 & new_n2126;
  assign new_n2128 = ~py & new_n2127;
  assign new_n2129 = ~pc0 & new_n2128;
  assign new_n2130 = ~pd0 & new_n2129;
  assign new_n2131 = ~pb0 & new_n2130;
  assign new_n2132 = ~pr & new_n2131;
  assign new_n2133 = ~px & new_n2132;
  assign new_n2134 = pn & new_n2133;
  assign new_n2135 = ~pq & new_n2134;
  assign new_n2136 = ~pv & new_n340;
  assign new_n2137 = ~py & new_n2136;
  assign new_n2138 = ~pa0 & new_n2137;
  assign new_n2139 = ~pc0 & new_n2138;
  assign new_n2140 = pk0 & new_n2139;
  assign new_n2141 = ~pb0 & new_n2140;
  assign new_n2142 = ~pr & new_n2141;
  assign new_n2143 = ~px & new_n2142;
  assign new_n2144 = ~pn & new_n2143;
  assign new_n2145 = ~pq & new_n2144;
  assign new_n2146 = ~pa0 & new_n1480;
  assign new_n2147 = ~po & new_n2146;
  assign new_n2148 = ~pm & new_n2147;
  assign new_n2149 = ~pd0 & new_n2148;
  assign new_n2150 = pk0 & new_n2149;
  assign new_n2151 = ~pc0 & new_n2150;
  assign new_n2152 = ~px & new_n2151;
  assign new_n2153 = ~pb0 & new_n2152;
  assign new_n2154 = ~pi & new_n2153;
  assign new_n2155 = ~pq & new_n2154;
  assign new_n2156 = ~pg0 & new_n881;
  assign new_n2157 = ~pm & new_n2156;
  assign new_n2158 = ~pd0 & new_n2157;
  assign new_n2159 = ~pi0 & new_n2158;
  assign new_n2160 = ~pc0 & new_n2159;
  assign new_n2161 = ~px & new_n2160;
  assign new_n2162 = ~pb0 & new_n2161;
  assign new_n2163 = ~pn & new_n2162;
  assign new_n2164 = ~pq & new_n2163;
  assign new_n2165 = pk0 & new_n1206;
  assign new_n2166 = ~pv & new_n2165;
  assign new_n2167 = ~pc0 & new_n2166;
  assign new_n2168 = ~pj0 & new_n2167;
  assign new_n2169 = pd & new_n1357;
  assign new_n2170 = ~ps & new_n2169;
  assign new_n2171 = pj0 & new_n2170;
  assign new_n2172 = ~pd0 & new_n2171;
  assign new_n2173 = ~pi0 & new_n2172;
  assign new_n2174 = ~pb0 & new_n2173;
  assign new_n2175 = ~pc0 & new_n2174;
  assign new_n2176 = pk0 & new_n1370;
  assign new_n2177 = ~pi0 & new_n2176;
  assign new_n2178 = pj0 & new_n2177;
  assign new_n2179 = ~pc0 & new_n2178;
  assign new_n2180 = ~pd0 & new_n2179;
  assign new_n2181 = ~pq & new_n151;
  assign new_n2182 = ~pr & new_n2181;
  assign new_n2183 = ~pn & new_n2182;
  assign new_n2184 = ~pc0 & new_n2183;
  assign new_n2185 = pd0 & new_n2184;
  assign new_n2186 = ~pb0 & new_n2185;
  assign new_n2187 = ~py & new_n2186;
  assign new_n2188 = ~pa0 & new_n2187;
  assign new_n2189 = ~pw & new_n2188;
  assign new_n2190 = ~px & new_n2189;
  assign new_n2191 = ~pv & new_n105;
  assign new_n2192 = ~py & new_n2191;
  assign new_n2193 = ~pa0 & new_n2192;
  assign new_n2194 = ~pc0 & new_n2193;
  assign new_n2195 = pd0 & new_n2194;
  assign new_n2196 = ~pj0 & new_n2195;
  assign new_n2197 = pk0 & new_n2196;
  assign new_n2198 = ~px & new_n2197;
  assign new_n2199 = ~pb0 & new_n2198;
  assign new_n2200 = ~pt & new_n2199;
  assign new_n2201 = ~pq & new_n2200;
  assign new_n2202 = ~pr & new_n2201;
  assign new_n2203 = ~pl & new_n2202;
  assign new_n2204 = ~pn & new_n2203;
  assign new_n2205 = ~py & new_n981;
  assign new_n2206 = ~pb0 & new_n2205;
  assign new_n2207 = ~pc0 & new_n2206;
  assign new_n2208 = ~pd0 & new_n2207;
  assign new_n2209 = pi0 & new_n2208;
  assign new_n2210 = ~pt & new_n2209;
  assign new_n2211 = ~px & new_n2210;
  assign new_n2212 = ~pr & new_n2211;
  assign new_n2213 = ~pn & new_n2212;
  assign new_n2214 = ~pq & new_n2213;
  assign new_n2215 = ~pj & new_n2214;
  assign new_n2216 = ~pl & new_n2215;
  assign new_n2217 = ~pg0 & new_n1155;
  assign new_n2218 = ~pd0 & new_n2217;
  assign new_n2219 = ~pi0 & new_n2218;
  assign new_n2220 = pj0 & new_n2219;
  assign new_n2221 = pk0 & new_n2220;
  assign new_n2222 = ~pb0 & new_n2221;
  assign new_n2223 = ~pc0 & new_n2222;
  assign new_n2224 = ~px & new_n2223;
  assign new_n2225 = ~pq & new_n2224;
  assign new_n2226 = ~pr & new_n2225;
  assign new_n2227 = ~pj & new_n2226;
  assign new_n2228 = ~pn & new_n2227;
  assign new_n2229 = ~po & new_n1721;
  assign new_n2230 = ~pd0 & new_n2229;
  assign new_n2231 = pi0 & new_n2230;
  assign new_n2232 = ~pc0 & new_n2231;
  assign new_n2233 = ~px & new_n2232;
  assign new_n2234 = ~pb0 & new_n2233;
  assign new_n2235 = ~pq & new_n2234;
  assign new_n2236 = ~pr & new_n2235;
  assign new_n2237 = ~pk & new_n1859;
  assign new_n2238 = pi0 & new_n2237;
  assign new_n2239 = ~pj0 & new_n2238;
  assign new_n2240 = pk0 & new_n2239;
  assign new_n2241 = ~pg0 & new_n2240;
  assign new_n2242 = ~pc0 & new_n2241;
  assign new_n2243 = ~pd0 & new_n2242;
  assign new_n2244 = ~pb0 & new_n2243;
  assign new_n2245 = ~pr & new_n2244;
  assign new_n2246 = ~px & new_n2245;
  assign new_n2247 = ~pn & new_n2246;
  assign new_n2248 = ~pq & new_n2247;
  assign new_n2249 = ~pa0 & new_n1058;
  assign new_n2250 = ~po & new_n2249;
  assign new_n2251 = pd0 & new_n2250;
  assign new_n2252 = pk0 & new_n2251;
  assign new_n2253 = ~pv & new_n2252;
  assign new_n2254 = ~py & new_n2253;
  assign new_n2255 = ~pb0 & new_n2254;
  assign new_n2256 = ~pc0 & new_n2255;
  assign new_n2257 = ~px & new_n2256;
  assign new_n2258 = ~pq & new_n2257;
  assign new_n2259 = ~pr & new_n2258;
  assign new_n2260 = ~pj & new_n2259;
  assign new_n2261 = pn & new_n2260;
  assign new_n2262 = ~pv & new_n416;
  assign new_n2263 = ~py & new_n2262;
  assign new_n2264 = ~pa0 & new_n2263;
  assign new_n2265 = ~pb0 & new_n2264;
  assign new_n2266 = ~pc0 & new_n2265;
  assign new_n2267 = ~px & new_n2266;
  assign new_n2268 = ~pq & new_n2267;
  assign new_n2269 = ~pr & new_n2268;
  assign new_n2270 = ~pi & new_n2269;
  assign new_n2271 = ~pn & new_n2270;
  assign new_n2272 = pk0 & new_n2148;
  assign new_n2273 = ~pg0 & new_n2272;
  assign new_n2274 = ~pd0 & new_n2273;
  assign new_n2275 = ~pb0 & new_n2274;
  assign new_n2276 = ~pc0 & new_n2275;
  assign new_n2277 = ~pq & new_n2276;
  assign new_n2278 = ~px & new_n2277;
  assign new_n2279 = ~pm & new_n1575;
  assign new_n2280 = ~pc0 & new_n2279;
  assign new_n2281 = ~pd0 & new_n2280;
  assign new_n2282 = ~pb0 & new_n2281;
  assign new_n2283 = ~pq & new_n2282;
  assign new_n2284 = ~px & new_n2283;
  assign new_n2285 = ~pi & new_n2284;
  assign new_n2286 = ~pn & new_n2285;
  assign new_n2287 = ~pm & new_n679;
  assign new_n2288 = ~pe0 & new_n2287;
  assign new_n2289 = ~pa0 & new_n2288;
  assign new_n2290 = ~pf0 & new_n2289;
  assign new_n2291 = ~py & new_n2290;
  assign new_n2292 = ~pg0 & new_n2291;
  assign new_n2293 = ~pv & new_n2292;
  assign new_n2294 = ~pj0 & new_n2293;
  assign new_n2295 = pk0 & new_n2294;
  assign new_n2296 = ~pi0 & new_n1276;
  assign new_n2297 = pj0 & new_n2296;
  assign new_n2298 = ~pd0 & new_n2297;
  assign new_n2299 = ~pb0 & new_n2298;
  assign new_n2300 = ~pc0 & new_n2299;
  assign new_n2301 = ~pt & new_n2300;
  assign new_n2302 = ~px & new_n2301;
  assign new_n2303 = ~pg0 & new_n1287;
  assign new_n2304 = pj0 & new_n2303;
  assign new_n2305 = pk0 & new_n2304;
  assign new_n2306 = ~pd0 & new_n2305;
  assign new_n2307 = ~pi0 & new_n2306;
  assign new_n2308 = pj0 & new_n1241;
  assign new_n2309 = ~pi0 & new_n2308;
  assign new_n2310 = ~pd0 & new_n2309;
  assign new_n2311 = ph0 & new_n2310;
  assign new_n2312 = ~pb0 & new_n2311;
  assign new_n2313 = ~pc0 & new_n2312;
  assign new_n2314 = ~pc0 & new_n1547;
  assign new_n2315 = pd0 & new_n2314;
  assign new_n2316 = pk0 & new_n2315;
  assign new_n2317 = ~pg0 & new_n2316;
  assign new_n2318 = ~px & new_n2317;
  assign new_n2319 = ~pb0 & new_n2318;
  assign new_n2320 = ~pt & new_n2319;
  assign new_n2321 = ~pq & new_n2320;
  assign new_n2322 = ~pr & new_n2321;
  assign new_n2323 = ~pl & new_n2322;
  assign new_n2324 = ~pn & new_n2323;
  assign new_n2325 = pk0 & new_n314;
  assign new_n2326 = ~pg0 & new_n2325;
  assign new_n2327 = ~py & new_n2326;
  assign new_n2328 = ~pc0 & new_n2327;
  assign new_n2329 = ~pd0 & new_n2328;
  assign new_n2330 = pi0 & new_n2329;
  assign new_n2331 = ~pj0 & new_n2330;
  assign new_n2332 = ~px & new_n2331;
  assign new_n2333 = ~pb0 & new_n2332;
  assign new_n2334 = ~pt & new_n2333;
  assign new_n2335 = ~pq & new_n2334;
  assign new_n2336 = ~pr & new_n2335;
  assign new_n2337 = ~pl & new_n2336;
  assign new_n2338 = ~pn & new_n2337;
  assign new_n2339 = ~pb0 & new_n2156;
  assign new_n2340 = ~pc0 & new_n2339;
  assign new_n2341 = ~pd0 & new_n2340;
  assign new_n2342 = ~pi0 & new_n2341;
  assign new_n2343 = ~pt & new_n2342;
  assign new_n2344 = ~px & new_n2343;
  assign new_n2345 = ~pr & new_n2344;
  assign new_n2346 = ~pn & new_n2345;
  assign new_n2347 = ~pq & new_n2346;
  assign new_n2348 = ~pj & new_n2347;
  assign new_n2349 = ~pl & new_n2348;
  assign new_n2350 = pk0 & new_n1588;
  assign new_n2351 = ~pg0 & new_n2350;
  assign new_n2352 = ~py & new_n2351;
  assign new_n2353 = ~pa0 & new_n2352;
  assign new_n2354 = ~pd0 & new_n2353;
  assign new_n2355 = ~pj0 & new_n2354;
  assign new_n2356 = ~pc0 & new_n2355;
  assign new_n2357 = ~px & new_n2356;
  assign new_n2358 = ~pb0 & new_n2357;
  assign new_n2359 = ~pq & new_n2358;
  assign new_n2360 = ~pr & new_n2359;
  assign new_n2361 = ~pk & new_n2249;
  assign new_n2362 = pd0 & new_n2361;
  assign new_n2363 = pk0 & new_n2362;
  assign new_n2364 = ~pv & new_n2363;
  assign new_n2365 = ~py & new_n2364;
  assign new_n2366 = ~pb0 & new_n2365;
  assign new_n2367 = ~pc0 & new_n2366;
  assign new_n2368 = ~px & new_n2367;
  assign new_n2369 = ~pq & new_n2368;
  assign new_n2370 = ~pr & new_n2369;
  assign new_n2371 = ~pj & new_n2370;
  assign new_n2372 = ~pn & new_n2371;
  assign new_n2373 = ~po & new_n106;
  assign new_n2374 = ~pj0 & new_n2373;
  assign new_n2375 = pk0 & new_n2374;
  assign new_n2376 = ~pv & new_n2375;
  assign new_n2377 = ~py & new_n2376;
  assign new_n2378 = ~pc0 & new_n2377;
  assign new_n2379 = pd0 & new_n2378;
  assign new_n2380 = ~pb0 & new_n2379;
  assign new_n2381 = ~pr & new_n2380;
  assign new_n2382 = ~px & new_n2381;
  assign new_n2383 = pn & new_n2382;
  assign new_n2384 = ~pq & new_n2383;
  assign new_n2385 = ~pg0 & new_n80;
  assign new_n2386 = ~py & new_n2385;
  assign new_n2387 = ~pa0 & new_n2386;
  assign new_n2388 = ~pf0 & new_n2387;
  assign new_n2389 = ~pj0 & new_n2388;
  assign new_n2390 = pk0 & new_n2389;
  assign new_n2391 = ~pd0 & new_n2390;
  assign new_n2392 = ~pb0 & new_n2391;
  assign new_n2393 = ~pc0 & new_n2392;
  assign new_n2394 = ~pq & new_n2393;
  assign new_n2395 = ~px & new_n2394;
  assign new_n2396 = ~pa0 & new_n418;
  assign new_n2397 = ~pc0 & new_n2396;
  assign new_n2398 = ~pd0 & new_n2397;
  assign new_n2399 = ~pb0 & new_n2398;
  assign new_n2400 = ~pr & new_n2399;
  assign new_n2401 = ~px & new_n2400;
  assign new_n2402 = ~pn & new_n2401;
  assign new_n2403 = ~pq & new_n2402;
  assign new_n2404 = ~po & new_n1753;
  assign new_n2405 = ~pm & new_n2404;
  assign new_n2406 = ~pd0 & new_n2405;
  assign new_n2407 = pi0 & new_n2406;
  assign new_n2408 = ~pc0 & new_n2407;
  assign new_n2409 = ~px & new_n2408;
  assign new_n2410 = ~pb0 & new_n2409;
  assign new_n2411 = ~pi & new_n2410;
  assign new_n2412 = ~pq & new_n2411;
  assign new_n2413 = ~pm & new_n2205;
  assign new_n2414 = ~pd0 & new_n2413;
  assign new_n2415 = pi0 & new_n2414;
  assign new_n2416 = ~pc0 & new_n2415;
  assign new_n2417 = ~px & new_n2416;
  assign new_n2418 = ~pb0 & new_n2417;
  assign new_n2419 = ~pn & new_n2418;
  assign new_n2420 = ~pq & new_n2419;
  assign new_n2421 = ~py & new_n1640;
  assign new_n2422 = ~pj0 & new_n2421;
  assign new_n2423 = pk0 & new_n2422;
  assign new_n2424 = ~pd0 & new_n2423;
  assign new_n2425 = pi0 & new_n2424;
  assign new_n2426 = ~pi & new_n292;
  assign new_n2427 = ~pf0 & new_n2426;
  assign new_n2428 = ~pe0 & new_n2427;
  assign new_n2429 = ~py & new_n2428;
  assign new_n2430 = ~pa0 & new_n2429;
  assign new_n2431 = pk0 & new_n2430;
  assign new_n2432 = ~pd0 & new_n2431;
  assign new_n2433 = ~pj0 & new_n2432;
  assign new_n2434 = ~pb0 & new_n2433;
  assign new_n2435 = ~pc0 & new_n2434;
  assign new_n2436 = pv & new_n1348;
  assign new_n2437 = pk & new_n2436;
  assign new_n2438 = pj0 & new_n2437;
  assign new_n2439 = ~pc0 & new_n2438;
  assign new_n2440 = ~pi0 & new_n2439;
  assign new_n2441 = ~px & new_n2440;
  assign new_n2442 = ~pb0 & new_n2441;
  assign new_n2443 = ~po & new_n2182;
  assign new_n2444 = ~pc0 & new_n2443;
  assign new_n2445 = pd0 & new_n2444;
  assign new_n2446 = ~pb0 & new_n2445;
  assign new_n2447 = ~py & new_n2446;
  assign new_n2448 = ~pa0 & new_n2447;
  assign new_n2449 = ~pw & new_n2448;
  assign new_n2450 = ~px & new_n2449;
  assign new_n2451 = ~pj0 & new_n2193;
  assign new_n2452 = pk0 & new_n2451;
  assign new_n2453 = pd & new_n2452;
  assign new_n2454 = ~ps & new_n2453;
  assign new_n2455 = ~pc0 & new_n2454;
  assign new_n2456 = pd0 & new_n2455;
  assign new_n2457 = ~pb0 & new_n2456;
  assign new_n2458 = ~pr & new_n2457;
  assign new_n2459 = ~px & new_n2458;
  assign new_n2460 = ~pn & new_n2459;
  assign new_n2461 = ~pq & new_n2460;
  assign new_n2462 = ~ps & new_n62;
  assign new_n2463 = ~pg0 & new_n2462;
  assign new_n2464 = ~py & new_n2463;
  assign new_n2465 = ~pd0 & new_n2464;
  assign new_n2466 = pi0 & new_n2465;
  assign new_n2467 = pk0 & new_n2466;
  assign new_n2468 = pd & new_n2467;
  assign new_n2469 = ~pb0 & new_n2468;
  assign new_n2470 = ~pc0 & new_n2469;
  assign new_n2471 = ~px & new_n2470;
  assign new_n2472 = ~pq & new_n2471;
  assign new_n2473 = ~pr & new_n2472;
  assign new_n2474 = ~pj & new_n2473;
  assign new_n2475 = ~pn & new_n2474;
  assign new_n2476 = pd & new_n63;
  assign new_n2477 = ~ps & new_n2476;
  assign new_n2478 = ~pc0 & new_n2477;
  assign new_n2479 = ~pd0 & new_n2478;
  assign new_n2480 = ~pi0 & new_n2479;
  assign new_n2481 = pj0 & new_n2480;
  assign new_n2482 = ~px & new_n2481;
  assign new_n2483 = ~pb0 & new_n2482;
  assign new_n2484 = ~pr & new_n2483;
  assign new_n2485 = ~pn & new_n2484;
  assign new_n2486 = ~pq & new_n2485;
  assign new_n2487 = ~pi & new_n2486;
  assign new_n2488 = ~pj & new_n2487;
  assign new_n2489 = ~pv & new_n1255;
  assign new_n2490 = ~py & new_n2489;
  assign new_n2491 = ~pa0 & new_n2490;
  assign new_n2492 = ~pc0 & new_n2491;
  assign new_n2493 = ~pj0 & new_n2492;
  assign new_n2494 = ~pb0 & new_n2493;
  assign new_n2495 = ~pr & new_n2494;
  assign new_n2496 = ~px & new_n2495;
  assign new_n2497 = ~pn & new_n2496;
  assign new_n2498 = ~pq & new_n2497;
  assign new_n2499 = ~pk & new_n2123;
  assign new_n2500 = ~pj0 & new_n2499;
  assign new_n2501 = pk0 & new_n2500;
  assign new_n2502 = ~pg0 & new_n2501;
  assign new_n2503 = ~py & new_n2502;
  assign new_n2504 = ~pc0 & new_n2503;
  assign new_n2505 = ~pd0 & new_n2504;
  assign new_n2506 = ~pb0 & new_n2505;
  assign new_n2507 = ~pr & new_n2506;
  assign new_n2508 = ~px & new_n2507;
  assign new_n2509 = ~pn & new_n2508;
  assign new_n2510 = ~pq & new_n2509;
  assign new_n2511 = ~po & new_n1334;
  assign new_n2512 = pk0 & new_n2511;
  assign new_n2513 = ~pg0 & new_n2512;
  assign new_n2514 = ~pv & new_n2513;
  assign new_n2515 = ~py & new_n2514;
  assign new_n2516 = ~pc0 & new_n2515;
  assign new_n2517 = pd0 & new_n2516;
  assign new_n2518 = ~pb0 & new_n2517;
  assign new_n2519 = ~pr & new_n2518;
  assign new_n2520 = ~px & new_n2519;
  assign new_n2521 = pn & new_n2520;
  assign new_n2522 = ~pq & new_n2521;
  assign new_n2523 = ~po & new_n1625;
  assign new_n2524 = ~pd0 & new_n2523;
  assign new_n2525 = ~pi0 & new_n2524;
  assign new_n2526 = pj0 & new_n2525;
  assign new_n2527 = pk0 & new_n2526;
  assign new_n2528 = ~pb0 & new_n2527;
  assign new_n2529 = ~pc0 & new_n2528;
  assign new_n2530 = ~px & new_n2529;
  assign new_n2531 = ~pq & new_n2530;
  assign new_n2532 = ~pr & new_n2531;
  assign new_n2533 = ~pj & new_n2532;
  assign new_n2534 = pn & new_n2533;
  assign new_n2535 = pk0 & new_n970;
  assign new_n2536 = ~py & new_n2535;
  assign new_n2537 = ~pa0 & new_n2536;
  assign new_n2538 = ~pb0 & new_n2537;
  assign new_n2539 = ~pc0 & new_n2538;
  assign new_n2540 = ~px & new_n2539;
  assign new_n2541 = ~pq & new_n2540;
  assign new_n2542 = ~pr & new_n2541;
  assign new_n2543 = ~pi & new_n2542;
  assign new_n2544 = ~pn & new_n2543;
  assign new_n2545 = ~po & new_n1626;
  assign new_n2546 = ~pm & new_n2545;
  assign new_n2547 = pi0 & new_n2546;
  assign new_n2548 = pk0 & new_n2547;
  assign new_n2549 = ~pd0 & new_n2548;
  assign new_n2550 = ~pb0 & new_n2549;
  assign new_n2551 = ~pc0 & new_n2550;
  assign new_n2552 = ~pq & new_n2551;
  assign new_n2553 = ~px & new_n2552;
  assign new_n2554 = ~pm & new_n2088;
  assign new_n2555 = ~pc0 & new_n2554;
  assign new_n2556 = ~pd0 & new_n2555;
  assign new_n2557 = ~pb0 & new_n2556;
  assign new_n2558 = ~pq & new_n2557;
  assign new_n2559 = ~px & new_n2558;
  assign new_n2560 = ~pi & new_n2559;
  assign new_n2561 = ~pn & new_n2560;
  assign new_n2562 = pk0 & new_n1641;
  assign new_n2563 = ~py & new_n2562;
  assign new_n2564 = ~pd0 & new_n2563;
  assign new_n2565 = ~pj0 & new_n2564;
  assign new_n2566 = pk0 & new_n2428;
  assign new_n2567 = ~py & new_n2566;
  assign new_n2568 = ~pj0 & new_n2567;
  assign new_n2569 = ~pd0 & new_n2568;
  assign new_n2570 = pi0 & new_n2569;
  assign new_n2571 = ~pb0 & new_n2570;
  assign new_n2572 = ~pc0 & new_n2571;
  assign new_n2573 = pv & new_n1267;
  assign new_n2574 = pk & new_n2573;
  assign new_n2575 = ~ps & new_n2574;
  assign new_n2576 = pj0 & new_n2575;
  assign new_n2577 = pd & new_n2576;
  assign new_n2578 = ~pc0 & new_n2577;
  assign new_n2579 = ~pi0 & new_n2578;
  assign new_n2580 = ~pn & new_n151;
  assign new_n2581 = ~pq & new_n2580;
  assign new_n2582 = ~pm & new_n2581;
  assign new_n2583 = ~pc0 & new_n2582;
  assign new_n2584 = pd0 & new_n2583;
  assign new_n2585 = ~pb0 & new_n2584;
  assign new_n2586 = ~py & new_n2585;
  assign new_n2587 = ~pa0 & new_n2586;
  assign new_n2588 = ~pw & new_n2587;
  assign new_n2589 = ~px & new_n2588;
  assign new_n2590 = ~new_n2579 & ~new_n2589;
  assign new_n2591 = ~new_n2565 & ~new_n2572;
  assign new_n2592 = new_n2590 & new_n2591;
  assign new_n2593 = ~new_n2553 & ~new_n2561;
  assign new_n2594 = ~new_n2534 & ~new_n2544;
  assign new_n2595 = new_n2593 & new_n2594;
  assign new_n2596 = new_n2592 & new_n2595;
  assign new_n2597 = ~new_n2510 & ~new_n2522;
  assign new_n2598 = ~new_n2488 & ~new_n2498;
  assign new_n2599 = new_n2597 & new_n2598;
  assign new_n2600 = ~new_n2461 & ~new_n2475;
  assign new_n2601 = ~new_n2435 & ~new_n2442;
  assign new_n2602 = ~new_n2450 & new_n2601;
  assign new_n2603 = new_n2600 & new_n2602;
  assign new_n2604 = new_n2599 & new_n2603;
  assign new_n2605 = new_n2596 & new_n2604;
  assign new_n2606 = ~new_n2420 & ~new_n2425;
  assign new_n2607 = ~new_n2403 & ~new_n2412;
  assign new_n2608 = new_n2606 & new_n2607;
  assign new_n2609 = ~new_n2384 & ~new_n2395;
  assign new_n2610 = ~new_n2360 & ~new_n2372;
  assign new_n2611 = new_n2609 & new_n2610;
  assign new_n2612 = new_n2608 & new_n2611;
  assign new_n2613 = ~new_n2338 & ~new_n2349;
  assign new_n2614 = ~new_n2313 & ~new_n2324;
  assign new_n2615 = new_n2613 & new_n2614;
  assign new_n2616 = ~new_n2302 & ~new_n2307;
  assign new_n2617 = ~new_n2278 & ~new_n2286;
  assign new_n2618 = ~new_n2295 & new_n2617;
  assign new_n2619 = new_n2616 & new_n2618;
  assign new_n2620 = new_n2615 & new_n2619;
  assign new_n2621 = new_n2612 & new_n2620;
  assign new_n2622 = new_n2605 & new_n2621;
  assign new_n2623 = ~new_n2261 & ~new_n2271;
  assign new_n2624 = ~new_n2236 & ~new_n2248;
  assign new_n2625 = new_n2623 & new_n2624;
  assign new_n2626 = ~new_n2216 & ~new_n2228;
  assign new_n2627 = ~new_n2190 & ~new_n2204;
  assign new_n2628 = new_n2626 & new_n2627;
  assign new_n2629 = new_n2625 & new_n2628;
  assign new_n2630 = ~new_n2175 & ~new_n2180;
  assign new_n2631 = ~new_n2164 & ~new_n2168;
  assign new_n2632 = new_n2630 & new_n2631;
  assign new_n2633 = ~new_n2145 & ~new_n2155;
  assign new_n2634 = ~new_n2110 & ~new_n2122;
  assign new_n2635 = ~new_n2135 & new_n2634;
  assign new_n2636 = new_n2633 & new_n2635;
  assign new_n2637 = new_n2632 & new_n2636;
  assign new_n2638 = new_n2629 & new_n2637;
  assign new_n2639 = ~new_n2085 & ~new_n2099;
  assign new_n2640 = ~new_n2060 & ~new_n2071;
  assign new_n2641 = new_n2639 & new_n2640;
  assign new_n2642 = ~new_n2044 & ~new_n2056;
  assign new_n2643 = ~new_n2010 & ~new_n2025;
  assign new_n2644 = ~new_n2037 & new_n2643;
  assign new_n2645 = new_n2642 & new_n2644;
  assign new_n2646 = new_n2641 & new_n2645;
  assign new_n2647 = ~new_n1989 & ~new_n2002;
  assign new_n2648 = ~new_n1966 & ~new_n1977;
  assign new_n2649 = new_n2647 & new_n2648;
  assign new_n2650 = ~new_n1944 & ~new_n1955;
  assign new_n2651 = ~new_n1920 & ~new_n1924;
  assign new_n2652 = ~new_n1930 & new_n2651;
  assign new_n2653 = new_n2650 & new_n2652;
  assign new_n2654 = new_n2649 & new_n2653;
  assign new_n2655 = new_n2646 & new_n2654;
  assign new_n2656 = new_n2638 & new_n2655;
  assign new_n2657 = new_n2622 & new_n2656;
  assign new_n2658 = ~new_n1904 & ~new_n1911;
  assign new_n2659 = ~new_n1882 & ~new_n1893;
  assign new_n2660 = new_n2658 & new_n2659;
  assign new_n2661 = ~new_n1830 & ~new_n1847;
  assign new_n2662 = ~new_n1858 & ~new_n1871;
  assign new_n2663 = new_n2661 & new_n2662;
  assign new_n2664 = new_n2660 & new_n2663;
  assign new_n2665 = ~new_n1805 & ~new_n1819;
  assign new_n2666 = ~new_n1794 & ~new_n1798;
  assign new_n2667 = new_n2665 & new_n2666;
  assign new_n2668 = ~new_n1775 & ~new_n1787;
  assign new_n2669 = ~new_n1741 & ~new_n1752;
  assign new_n2670 = ~new_n1762 & new_n2669;
  assign new_n2671 = new_n2668 & new_n2670;
  assign new_n2672 = new_n2667 & new_n2671;
  assign new_n2673 = new_n2664 & new_n2672;
  assign new_n2674 = ~new_n1718 & ~new_n1729;
  assign new_n2675 = ~new_n1693 & ~new_n1707;
  assign new_n2676 = new_n2674 & new_n2675;
  assign new_n2677 = ~new_n1668 & ~new_n1675;
  assign new_n2678 = ~new_n1645 & ~new_n1657;
  assign new_n2679 = ~new_n1664 & new_n2678;
  assign new_n2680 = new_n2677 & new_n2679;
  assign new_n2681 = new_n2676 & new_n2680;
  assign new_n2682 = ~new_n1624 & ~new_n1635;
  assign new_n2683 = ~new_n1599 & ~new_n1611;
  assign new_n2684 = new_n2682 & new_n2683;
  assign new_n2685 = ~new_n1572 & ~new_n1586;
  assign new_n2686 = ~new_n1540 & ~new_n1544;
  assign new_n2687 = ~new_n1558 & new_n2686;
  assign new_n2688 = new_n2685 & new_n2687;
  assign new_n2689 = new_n2684 & new_n2688;
  assign new_n2690 = new_n2681 & new_n2689;
  assign new_n2691 = new_n2673 & new_n2690;
  assign new_n2692 = ~new_n1529 & ~new_n1536;
  assign new_n2693 = ~new_n1515 & ~new_n1524;
  assign new_n2694 = new_n2692 & new_n2693;
  assign new_n2695 = ~new_n1503 & ~new_n1508;
  assign new_n2696 = ~new_n1492 & ~new_n1497;
  assign new_n2697 = new_n2695 & new_n2696;
  assign new_n2698 = new_n2694 & new_n2697;
  assign new_n2699 = ~new_n1473 & ~new_n1479;
  assign new_n2700 = ~new_n1460 & ~new_n1467;
  assign new_n2701 = new_n2699 & new_n2700;
  assign new_n2702 = ~new_n1446 & ~new_n1456;
  assign new_n2703 = ~new_n1427 & ~new_n1434;
  assign new_n2704 = ~new_n1439 & new_n2703;
  assign new_n2705 = new_n2702 & new_n2704;
  assign new_n2706 = new_n2701 & new_n2705;
  assign new_n2707 = new_n2698 & new_n2706;
  assign new_n2708 = ~new_n1410 & ~new_n1422;
  assign new_n2709 = ~new_n1401 & ~new_n1405;
  assign new_n2710 = new_n2708 & new_n2709;
  assign new_n2711 = ~new_n1391 & ~new_n1396;
  assign new_n2712 = ~new_n1364 & ~new_n1375;
  assign new_n2713 = ~new_n1384 & new_n2712;
  assign new_n2714 = new_n2711 & new_n2713;
  assign new_n2715 = new_n2710 & new_n2714;
  assign new_n2716 = ~new_n1346 & ~new_n1355;
  assign new_n2717 = ~new_n1323 & ~new_n1329;
  assign new_n2718 = new_n2716 & new_n2717;
  assign new_n2719 = ~new_n1311 & ~new_n1318;
  assign new_n2720 = ~new_n1292 & ~new_n1303;
  assign new_n2721 = ~new_n1307 & new_n2720;
  assign new_n2722 = new_n2719 & new_n2721;
  assign new_n2723 = new_n2718 & new_n2722;
  assign new_n2724 = new_n2715 & new_n2723;
  assign new_n2725 = new_n2707 & new_n2724;
  assign new_n2726 = new_n2691 & new_n2725;
  assign new_n2727 = new_n2657 & new_n2726;
  assign new_n2728 = ~new_n1274 & ~new_n1283;
  assign new_n2729 = ~new_n1252 & ~new_n1265;
  assign new_n2730 = new_n2728 & new_n2729;
  assign new_n2731 = ~new_n1238 & ~new_n1247;
  assign new_n2732 = ~new_n1228 & ~new_n1232;
  assign new_n2733 = new_n2731 & new_n2732;
  assign new_n2734 = new_n2730 & new_n2733;
  assign new_n2735 = ~new_n1215 & ~new_n1219;
  assign new_n2736 = ~new_n1203 & ~new_n1210;
  assign new_n2737 = new_n2735 & new_n2736;
  assign new_n2738 = ~new_n1177 & ~new_n1192;
  assign new_n2739 = ~new_n1148 & ~new_n1153;
  assign new_n2740 = ~new_n1167 & new_n2739;
  assign new_n2741 = new_n2738 & new_n2740;
  assign new_n2742 = new_n2737 & new_n2741;
  assign new_n2743 = new_n2734 & new_n2742;
  assign new_n2744 = ~new_n1133 & ~new_n1139;
  assign new_n2745 = ~new_n1122 & ~new_n1128;
  assign new_n2746 = new_n2744 & new_n2745;
  assign new_n2747 = ~new_n1112 & ~new_n1117;
  assign new_n2748 = ~new_n1091 & ~new_n1102;
  assign new_n2749 = new_n2747 & new_n2748;
  assign new_n2750 = new_n2746 & new_n2749;
  assign new_n2751 = ~new_n1072 & ~new_n1083;
  assign new_n2752 = ~new_n1049 & ~new_n1054;
  assign new_n2753 = new_n2751 & new_n2752;
  assign new_n2754 = ~new_n1034 & ~new_n1040;
  assign new_n2755 = ~new_n1017 & ~new_n1024;
  assign new_n2756 = ~new_n1030 & new_n2755;
  assign new_n2757 = new_n2754 & new_n2756;
  assign new_n2758 = new_n2753 & new_n2757;
  assign new_n2759 = new_n2750 & new_n2758;
  assign new_n2760 = new_n2743 & new_n2759;
  assign new_n2761 = ~new_n964 & ~new_n969;
  assign new_n2762 = ~new_n946 & ~new_n955;
  assign new_n2763 = new_n2761 & new_n2762;
  assign new_n2764 = ~new_n980 & ~new_n990;
  assign new_n2765 = ~new_n1001 & ~new_n1008;
  assign new_n2766 = new_n2764 & new_n2765;
  assign new_n2767 = new_n2763 & new_n2766;
  assign new_n2768 = ~new_n932 & ~new_n938;
  assign new_n2769 = ~new_n911 & ~new_n922;
  assign new_n2770 = new_n2768 & new_n2769;
  assign new_n2771 = ~new_n890 & ~new_n901;
  assign new_n2772 = ~new_n864 & ~new_n870;
  assign new_n2773 = ~new_n879 & new_n2772;
  assign new_n2774 = new_n2771 & new_n2773;
  assign new_n2775 = new_n2770 & new_n2774;
  assign new_n2776 = new_n2767 & new_n2775;
  assign new_n2777 = ~new_n840 & ~new_n845;
  assign new_n2778 = ~new_n854 & ~new_n859;
  assign new_n2779 = new_n2777 & new_n2778;
  assign new_n2780 = ~new_n831 & ~new_n836;
  assign new_n2781 = ~new_n807 & ~new_n816;
  assign new_n2782 = ~new_n823 & new_n2781;
  assign new_n2783 = new_n2780 & new_n2782;
  assign new_n2784 = new_n2779 & new_n2783;
  assign new_n2785 = ~new_n796 & ~new_n802;
  assign new_n2786 = ~new_n782 & ~new_n787;
  assign new_n2787 = new_n2785 & new_n2786;
  assign new_n2788 = ~new_n767 & ~new_n776;
  assign new_n2789 = ~new_n747 & ~new_n752;
  assign new_n2790 = ~new_n757 & new_n2789;
  assign new_n2791 = new_n2788 & new_n2790;
  assign new_n2792 = new_n2787 & new_n2791;
  assign new_n2793 = new_n2784 & new_n2792;
  assign new_n2794 = new_n2776 & new_n2793;
  assign new_n2795 = new_n2760 & new_n2794;
  assign new_n2796 = ~new_n700 & ~new_n705;
  assign new_n2797 = ~new_n684 & ~new_n692;
  assign new_n2798 = new_n2796 & new_n2797;
  assign new_n2799 = ~new_n715 & ~new_n725;
  assign new_n2800 = ~new_n731 & ~new_n739;
  assign new_n2801 = new_n2799 & new_n2800;
  assign new_n2802 = new_n2798 & new_n2801;
  assign new_n2803 = ~new_n671 & ~new_n675;
  assign new_n2804 = ~new_n660 & ~new_n667;
  assign new_n2805 = new_n2803 & new_n2804;
  assign new_n2806 = ~new_n643 & ~new_n652;
  assign new_n2807 = ~new_n617 & ~new_n627;
  assign new_n2808 = ~new_n635 & new_n2807;
  assign new_n2809 = new_n2806 & new_n2808;
  assign new_n2810 = new_n2805 & new_n2809;
  assign new_n2811 = new_n2802 & new_n2810;
  assign new_n2812 = ~new_n599 & ~new_n606;
  assign new_n2813 = ~new_n581 & ~new_n590;
  assign new_n2814 = new_n2812 & new_n2813;
  assign new_n2815 = ~new_n568 & ~new_n577;
  assign new_n2816 = ~new_n539 & ~new_n550;
  assign new_n2817 = ~new_n557 & new_n2816;
  assign new_n2818 = new_n2815 & new_n2817;
  assign new_n2819 = new_n2814 & new_n2818;
  assign new_n2820 = ~new_n526 & ~new_n533;
  assign new_n2821 = ~new_n509 & ~new_n518;
  assign new_n2822 = new_n2820 & new_n2821;
  assign new_n2823 = ~new_n490 & ~new_n497;
  assign new_n2824 = ~new_n463 & ~new_n470;
  assign new_n2825 = ~new_n474 & new_n2824;
  assign new_n2826 = new_n2823 & new_n2825;
  assign new_n2827 = new_n2822 & new_n2826;
  assign new_n2828 = new_n2819 & new_n2827;
  assign new_n2829 = new_n2811 & new_n2828;
  assign new_n2830 = ~new_n437 & ~new_n453;
  assign new_n2831 = ~new_n426 & ~new_n433;
  assign new_n2832 = new_n2830 & new_n2831;
  assign new_n2833 = ~new_n406 & ~new_n415;
  assign new_n2834 = ~new_n393 & ~new_n397;
  assign new_n2835 = new_n2833 & new_n2834;
  assign new_n2836 = new_n2832 & new_n2835;
  assign new_n2837 = ~new_n379 & ~new_n386;
  assign new_n2838 = ~new_n357 & ~new_n368;
  assign new_n2839 = new_n2837 & new_n2838;
  assign new_n2840 = ~new_n339 & ~new_n350;
  assign new_n2841 = ~new_n301 & ~new_n310;
  assign new_n2842 = ~new_n328 & new_n2841;
  assign new_n2843 = new_n2840 & new_n2842;
  assign new_n2844 = new_n2839 & new_n2843;
  assign new_n2845 = new_n2836 & new_n2844;
  assign new_n2846 = ~new_n161 & ~new_n178;
  assign new_n2847 = ~new_n134 & ~new_n150;
  assign new_n2848 = new_n2846 & new_n2847;
  assign new_n2849 = ~new_n101 & ~new_n118;
  assign new_n2850 = ~new_n58 & ~new_n75;
  assign new_n2851 = ~new_n91 & new_n2850;
  assign new_n2852 = new_n2849 & new_n2851;
  assign new_n2853 = new_n2848 & new_n2852;
  assign new_n2854 = ~new_n278 & ~new_n290;
  assign new_n2855 = ~new_n255 & ~new_n267;
  assign new_n2856 = new_n2854 & new_n2855;
  assign new_n2857 = ~new_n230 & ~new_n241;
  assign new_n2858 = ~new_n194 & ~new_n206;
  assign new_n2859 = ~new_n218 & new_n2858;
  assign new_n2860 = new_n2857 & new_n2859;
  assign new_n2861 = new_n2856 & new_n2860;
  assign new_n2862 = new_n2853 & new_n2861;
  assign new_n2863 = new_n2845 & new_n2862;
  assign new_n2864 = new_n2829 & new_n2863;
  assign new_n2865 = new_n2795 & new_n2864;
  assign pn0 = ~new_n2727 | ~new_n2865;
  assign new_n2867 = ~pa & new_n61;
  assign new_n2868 = pl0 & new_n2867;
  assign new_n2869 = pd & new_n2868;
  assign new_n2870 = ~ps & new_n2869;
  assign new_n2871 = ~po & new_n2870;
  assign new_n2872 = ~pa0 & new_n2871;
  assign new_n2873 = ~pb0 & new_n2872;
  assign new_n2874 = ~pc0 & new_n2873;
  assign new_n2875 = pd0 & new_n2874;
  assign new_n2876 = ~px & new_n2875;
  assign new_n2877 = ~py & new_n2876;
  assign new_n2878 = ~pu & new_n2877;
  assign new_n2879 = ~pq & new_n2878;
  assign new_n2880 = ~pr & new_n2879;
  assign new_n2881 = ~pi & new_n2880;
  assign new_n2882 = ~pj & new_n2881;
  assign new_n2883 = ~pc & new_n1058;
  assign new_n2884 = pi0 & new_n2883;
  assign new_n2885 = ~pk & new_n2884;
  assign new_n2886 = ~pc0 & new_n2885;
  assign new_n2887 = ~pd0 & new_n2886;
  assign new_n2888 = ~ph0 & new_n2887;
  assign new_n2889 = pl0 & new_n2888;
  assign new_n2890 = ~py & new_n2889;
  assign new_n2891 = ~pb0 & new_n2890;
  assign new_n2892 = ~px & new_n2891;
  assign new_n2893 = ~pq & new_n2892;
  assign new_n2894 = ~pr & new_n2893;
  assign new_n2895 = ~pj & new_n2894;
  assign new_n2896 = ~pn & new_n2895;
  assign new_n2897 = ~pq & ~pj;
  assign new_n2898 = ~pf & new_n2897;
  assign new_n2899 = ~pg & new_n2898;
  assign new_n2900 = ~pe & new_n2899;
  assign new_n2901 = ~po & new_n2900;
  assign new_n2902 = ~pc & new_n2901;
  assign new_n2903 = pi0 & new_n2902;
  assign new_n2904 = pd & new_n2903;
  assign new_n2905 = ~ps & new_n2904;
  assign new_n2906 = ~pg0 & new_n2905;
  assign new_n2907 = ~pj0 & new_n2906;
  assign new_n2908 = ~pd0 & new_n2907;
  assign new_n2909 = pl0 & new_n2908;
  assign new_n2910 = ~pc0 & new_n2909;
  assign new_n2911 = ~py & new_n2910;
  assign new_n2912 = ~pb0 & new_n2911;
  assign new_n2913 = ~pr & new_n2912;
  assign new_n2914 = ~px & new_n2913;
  assign new_n2915 = ~ps & new_n1834;
  assign new_n2916 = ~pg0 & new_n2915;
  assign new_n2917 = ~pj0 & new_n2916;
  assign new_n2918 = ~pc & new_n2917;
  assign new_n2919 = ~pd0 & new_n2918;
  assign new_n2920 = ~ph0 & new_n2919;
  assign new_n2921 = pl0 & new_n2920;
  assign new_n2922 = pd & new_n2921;
  assign new_n2923 = ~pb0 & new_n2922;
  assign new_n2924 = ~pc0 & new_n2923;
  assign new_n2925 = ~pa0 & new_n2924;
  assign new_n2926 = ~px & new_n2925;
  assign new_n2927 = ~py & new_n2926;
  assign new_n2928 = ~pq & new_n2927;
  assign new_n2929 = ~pr & new_n2928;
  assign new_n2930 = ~pj0 & new_n1834;
  assign new_n2931 = ~pc & new_n2930;
  assign new_n2932 = ~pk & new_n2931;
  assign new_n2933 = ~pd0 & new_n2932;
  assign new_n2934 = ~ph0 & new_n2933;
  assign new_n2935 = pl0 & new_n2934;
  assign new_n2936 = ~pg0 & new_n2935;
  assign new_n2937 = ~pb0 & new_n2936;
  assign new_n2938 = ~pc0 & new_n2937;
  assign new_n2939 = ~pa0 & new_n2938;
  assign new_n2940 = ~px & new_n2939;
  assign new_n2941 = ~py & new_n2940;
  assign new_n2942 = ~pq & new_n2941;
  assign new_n2943 = ~pr & new_n2942;
  assign new_n2944 = ~po & new_n1058;
  assign new_n2945 = ~pc & new_n2944;
  assign new_n2946 = ~pi0 & new_n2945;
  assign new_n2947 = ~pc0 & new_n2946;
  assign new_n2948 = ~pd0 & new_n2947;
  assign new_n2949 = pl0 & new_n2948;
  assign new_n2950 = pj0 & new_n2949;
  assign new_n2951 = ~px & new_n2950;
  assign new_n2952 = ~pb0 & new_n2951;
  assign new_n2953 = ~pt & new_n2952;
  assign new_n2954 = ~pq & new_n2953;
  assign new_n2955 = ~pr & new_n2954;
  assign new_n2956 = ~pj & new_n2955;
  assign new_n2957 = ~pl & new_n2956;
  assign new_n2958 = ~ps & new_n1058;
  assign new_n2959 = pj0 & new_n2958;
  assign new_n2960 = ~pc & new_n2959;
  assign new_n2961 = ~pi0 & new_n2960;
  assign new_n2962 = ~pd0 & new_n2961;
  assign new_n2963 = ~ph0 & new_n2962;
  assign new_n2964 = pl0 & new_n2963;
  assign new_n2965 = pd & new_n2964;
  assign new_n2966 = ~pb0 & new_n2965;
  assign new_n2967 = ~pc0 & new_n2966;
  assign new_n2968 = ~px & new_n2967;
  assign new_n2969 = ~pq & new_n2968;
  assign new_n2970 = ~pr & new_n2969;
  assign new_n2971 = ~pj & new_n2970;
  assign new_n2972 = ~pn & new_n2971;
  assign new_n2973 = ~pj0 & new_n105;
  assign new_n2974 = ~pc & new_n2973;
  assign new_n2975 = ~pk & new_n2974;
  assign new_n2976 = ~pc0 & new_n2975;
  assign new_n2977 = ~pd0 & new_n2976;
  assign new_n2978 = ~ph0 & new_n2977;
  assign new_n2979 = pl0 & new_n2978;
  assign new_n2980 = ~pa0 & new_n2979;
  assign new_n2981 = ~pb0 & new_n2980;
  assign new_n2982 = ~py & new_n2981;
  assign new_n2983 = ~pr & new_n2982;
  assign new_n2984 = ~px & new_n2983;
  assign new_n2985 = ~pn & new_n2984;
  assign new_n2986 = ~pq & new_n2985;
  assign new_n2987 = ~po & new_n105;
  assign new_n2988 = ~pc & new_n2987;
  assign new_n2989 = pi0 & new_n2988;
  assign new_n2990 = pl0 & new_n2989;
  assign new_n2991 = pd & new_n2990;
  assign new_n2992 = ~ps & new_n2991;
  assign new_n2993 = ~pj0 & new_n2992;
  assign new_n2994 = ~pc0 & new_n2993;
  assign new_n2995 = ~pd0 & new_n2994;
  assign new_n2996 = ~pb0 & new_n2995;
  assign new_n2997 = ~px & new_n2996;
  assign new_n2998 = ~py & new_n2997;
  assign new_n2999 = ~pq & new_n2998;
  assign new_n3000 = ~pr & new_n2999;
  assign new_n3001 = ~pn & new_n584;
  assign new_n3002 = ~pe0 & new_n3001;
  assign new_n3003 = pf0 & new_n3002;
  assign new_n3004 = ~pg0 & new_n3003;
  assign new_n3005 = pi0 & new_n3004;
  assign new_n3006 = pl0 & new_n3005;
  assign new_n3007 = ~pd0 & new_n3006;
  assign new_n3008 = ~ph0 & new_n3007;
  assign new_n3009 = ~pb0 & new_n3008;
  assign new_n3010 = ~pc0 & new_n3009;
  assign new_n3011 = pi0 & new_n2426;
  assign new_n3012 = ~pe0 & new_n3011;
  assign new_n3013 = pl0 & new_n3012;
  assign new_n3014 = ~pj0 & new_n3013;
  assign new_n3015 = ~ph0 & new_n3014;
  assign new_n3016 = ~pc0 & new_n3015;
  assign new_n3017 = ~pd0 & new_n3016;
  assign new_n3018 = ~py & new_n3017;
  assign new_n3019 = ~pb0 & new_n3018;
  assign new_n3020 = ~ph0 & new_n2867;
  assign new_n3021 = pl0 & new_n3020;
  assign new_n3022 = pd & new_n3021;
  assign new_n3023 = ~ps & new_n3022;
  assign new_n3024 = ~pa0 & new_n3023;
  assign new_n3025 = ~pb0 & new_n3024;
  assign new_n3026 = ~pc0 & new_n3025;
  assign new_n3027 = pd0 & new_n3026;
  assign new_n3028 = ~px & new_n3027;
  assign new_n3029 = ~pg0 & new_n3028;
  assign new_n3030 = ~py & new_n3029;
  assign new_n3031 = ~pu & new_n3030;
  assign new_n3032 = ~pq & new_n3031;
  assign new_n3033 = ~pr & new_n3032;
  assign new_n3034 = ~pj & new_n3033;
  assign new_n3035 = ~pn & new_n3034;
  assign new_n3036 = ~pa & new_n313;
  assign new_n3037 = ~pj0 & new_n3036;
  assign new_n3038 = ~po & new_n3037;
  assign new_n3039 = ~pk & new_n3038;
  assign new_n3040 = ~pc0 & new_n3039;
  assign new_n3041 = pd0 & new_n3040;
  assign new_n3042 = pl0 & new_n3041;
  assign new_n3043 = ~pg0 & new_n3042;
  assign new_n3044 = ~pa0 & new_n3043;
  assign new_n3045 = ~pb0 & new_n3044;
  assign new_n3046 = ~py & new_n3045;
  assign new_n3047 = ~pu & new_n3046;
  assign new_n3048 = ~px & new_n3047;
  assign new_n3049 = ~pq & new_n3048;
  assign new_n3050 = ~pr & new_n3049;
  assign new_n3051 = ~po & new_n1679;
  assign new_n3052 = ~pc & new_n3051;
  assign new_n3053 = pi0 & new_n3052;
  assign new_n3054 = ~pd0 & new_n3053;
  assign new_n3055 = pl0 & new_n3054;
  assign new_n3056 = ~pg0 & new_n3055;
  assign new_n3057 = ~pj0 & new_n3056;
  assign new_n3058 = ~pb0 & new_n3057;
  assign new_n3059 = ~pc0 & new_n3058;
  assign new_n3060 = ~py & new_n3059;
  assign new_n3061 = ~pt & new_n3060;
  assign new_n3062 = ~px & new_n3061;
  assign new_n3063 = ~pq & new_n3062;
  assign new_n3064 = ~pr & new_n3063;
  assign new_n3065 = pl0 & new_n3003;
  assign new_n3066 = ~pg0 & new_n3065;
  assign new_n3067 = ~ph0 & new_n3066;
  assign new_n3068 = ~pc0 & new_n3067;
  assign new_n3069 = ~pd0 & new_n3068;
  assign new_n3070 = ~pa0 & new_n3069;
  assign new_n3071 = ~pb0 & new_n3070;
  assign new_n3072 = ~pi0 & new_n222;
  assign new_n3073 = ~pe0 & new_n3072;
  assign new_n3074 = pl0 & new_n3073;
  assign new_n3075 = pj0 & new_n3074;
  assign new_n3076 = ~ph0 & new_n3075;
  assign new_n3077 = ~pc0 & new_n3076;
  assign new_n3078 = ~pd0 & new_n3077;
  assign new_n3079 = ~px & new_n3078;
  assign new_n3080 = ~pb0 & new_n3079;
  assign new_n3081 = ~pa & new_n137;
  assign new_n3082 = ~pj0 & new_n3081;
  assign new_n3083 = ~po & new_n3082;
  assign new_n3084 = ~pk & new_n3083;
  assign new_n3085 = ~pb0 & new_n3084;
  assign new_n3086 = ~pc0 & new_n3085;
  assign new_n3087 = pd0 & new_n3086;
  assign new_n3088 = pl0 & new_n3087;
  assign new_n3089 = ~py & new_n3088;
  assign new_n3090 = ~pa0 & new_n3089;
  assign new_n3091 = ~px & new_n3090;
  assign new_n3092 = ~pr & new_n3091;
  assign new_n3093 = ~pu & new_n3092;
  assign new_n3094 = ~pj & new_n3093;
  assign new_n3095 = ~pq & new_n3094;
  assign new_n3096 = ~po & new_n1333;
  assign new_n3097 = ~pc & new_n3096;
  assign new_n3098 = pi0 & new_n3097;
  assign new_n3099 = pl0 & new_n3098;
  assign new_n3100 = pd & new_n3099;
  assign new_n3101 = ~ps & new_n3100;
  assign new_n3102 = ~pg0 & new_n3101;
  assign new_n3103 = ~pc0 & new_n3102;
  assign new_n3104 = ~pd0 & new_n3103;
  assign new_n3105 = ~pb0 & new_n3104;
  assign new_n3106 = ~px & new_n3105;
  assign new_n3107 = ~py & new_n3106;
  assign new_n3108 = ~pq & new_n3107;
  assign new_n3109 = ~pr & new_n3108;
  assign new_n3110 = ~pm & new_n1295;
  assign new_n3111 = ~pe0 & new_n3110;
  assign new_n3112 = pj0 & new_n3111;
  assign new_n3113 = ~pi0 & new_n3112;
  assign new_n3114 = pl0 & new_n3113;
  assign new_n3115 = ~pd0 & new_n3114;
  assign new_n3116 = ~ph0 & new_n3115;
  assign new_n3117 = ~pb0 & new_n3116;
  assign new_n3118 = ~pc0 & new_n3117;
  assign new_n3119 = ~pu & ~px;
  assign new_n3120 = ~pq & new_n3119;
  assign new_n3121 = ~pr & new_n3120;
  assign new_n3122 = ~pa & new_n3121;
  assign new_n3123 = ~po & new_n3122;
  assign new_n3124 = ~pe0 & new_n3123;
  assign new_n3125 = ~pg0 & new_n3124;
  assign new_n3126 = ~pj0 & new_n3125;
  assign new_n3127 = pl0 & new_n3126;
  assign new_n3128 = ~pb0 & new_n3127;
  assign new_n3129 = ~pc0 & new_n3128;
  assign new_n3130 = ~py & new_n3129;
  assign new_n3131 = ~pa0 & new_n3130;
  assign new_n3132 = ~pg0 & new_n2867;
  assign new_n3133 = ~po & new_n3132;
  assign new_n3134 = ~pk & new_n3133;
  assign new_n3135 = ~pb0 & new_n3134;
  assign new_n3136 = ~pc0 & new_n3135;
  assign new_n3137 = pd0 & new_n3136;
  assign new_n3138 = pl0 & new_n3137;
  assign new_n3139 = ~py & new_n3138;
  assign new_n3140 = ~pa0 & new_n3139;
  assign new_n3141 = ~px & new_n3140;
  assign new_n3142 = ~pr & new_n3141;
  assign new_n3143 = ~pu & new_n3142;
  assign new_n3144 = ~pj & new_n3143;
  assign new_n3145 = ~pq & new_n3144;
  assign new_n3146 = ~pc0 & new_n2989;
  assign new_n3147 = ~pd0 & new_n3146;
  assign new_n3148 = pl0 & new_n3147;
  assign new_n3149 = ~pj0 & new_n3148;
  assign new_n3150 = ~py & new_n3149;
  assign new_n3151 = ~pb0 & new_n3150;
  assign new_n3152 = ~px & new_n3151;
  assign new_n3153 = ~pr & new_n3152;
  assign new_n3154 = ~pt & new_n3153;
  assign new_n3155 = ~pl & new_n3154;
  assign new_n3156 = ~pq & new_n3155;
  assign new_n3157 = ~pn & new_n582;
  assign new_n3158 = ~pq & new_n3157;
  assign new_n3159 = ~pi & new_n3158;
  assign new_n3160 = ~pm & new_n3159;
  assign new_n3161 = ~pe0 & new_n3160;
  assign new_n3162 = ~pj0 & new_n3161;
  assign new_n3163 = pi0 & new_n3162;
  assign new_n3164 = pl0 & new_n3163;
  assign new_n3165 = ~pd0 & new_n3164;
  assign new_n3166 = ~ph0 & new_n3165;
  assign new_n3167 = ~pb0 & new_n3166;
  assign new_n3168 = ~pc0 & new_n3167;
  assign new_n3169 = pi0 & new_n222;
  assign new_n3170 = ~pe0 & new_n3169;
  assign new_n3171 = ~ph0 & new_n3170;
  assign new_n3172 = pl0 & new_n3171;
  assign new_n3173 = ~pd0 & new_n3172;
  assign new_n3174 = ~pb0 & new_n3173;
  assign new_n3175 = ~pc0 & new_n3174;
  assign new_n3176 = ~px & new_n3175;
  assign new_n3177 = ~py & new_n3176;
  assign new_n3178 = ~po & new_n2868;
  assign new_n3179 = ~pk & new_n3178;
  assign new_n3180 = ~pa0 & new_n3179;
  assign new_n3181 = ~pb0 & new_n3180;
  assign new_n3182 = ~pc0 & new_n3181;
  assign new_n3183 = pd0 & new_n3182;
  assign new_n3184 = ~px & new_n3183;
  assign new_n3185 = ~py & new_n3184;
  assign new_n3186 = ~pu & new_n3185;
  assign new_n3187 = ~pq & new_n3186;
  assign new_n3188 = ~pr & new_n3187;
  assign new_n3189 = ~pi & new_n3188;
  assign new_n3190 = ~pj & new_n3189;
  assign new_n3191 = pi0 & new_n2945;
  assign new_n3192 = ~pd0 & new_n3191;
  assign new_n3193 = pl0 & new_n3192;
  assign new_n3194 = pd & new_n3193;
  assign new_n3195 = ~ps & new_n3194;
  assign new_n3196 = ~pb0 & new_n3195;
  assign new_n3197 = ~pc0 & new_n3196;
  assign new_n3198 = ~py & new_n3197;
  assign new_n3199 = ~pr & new_n3198;
  assign new_n3200 = ~px & new_n3199;
  assign new_n3201 = ~pj & new_n3200;
  assign new_n3202 = ~pq & new_n3201;
  assign new_n3203 = pl0 & new_n3111;
  assign new_n3204 = pi0 & new_n3203;
  assign new_n3205 = ~ph0 & new_n3204;
  assign new_n3206 = ~pc0 & new_n3205;
  assign new_n3207 = ~pd0 & new_n3206;
  assign new_n3208 = ~py & new_n3207;
  assign new_n3209 = ~pb0 & new_n3208;
  assign new_n3210 = ~pr & ~pu;
  assign new_n3211 = ~ph & new_n3210;
  assign new_n3212 = ~pq & new_n3211;
  assign new_n3213 = ~pa & new_n3212;
  assign new_n3214 = ~po & new_n3213;
  assign new_n3215 = ~pe0 & new_n3214;
  assign new_n3216 = pl0 & new_n3215;
  assign new_n3217 = ~pg0 & new_n3216;
  assign new_n3218 = ~pc0 & new_n3217;
  assign new_n3219 = ~pa0 & new_n3218;
  assign new_n3220 = ~pb0 & new_n3219;
  assign new_n3221 = ~px & new_n3220;
  assign new_n3222 = ~py & new_n3221;
  assign new_n3223 = ~pi0 & new_n3097;
  assign new_n3224 = pd & new_n3223;
  assign new_n3225 = ~ps & new_n3224;
  assign new_n3226 = ~pg0 & new_n3225;
  assign new_n3227 = pj0 & new_n3226;
  assign new_n3228 = ~pd0 & new_n3227;
  assign new_n3229 = pl0 & new_n3228;
  assign new_n3230 = ~pc0 & new_n3229;
  assign new_n3231 = ~px & new_n3230;
  assign new_n3232 = ~pb0 & new_n3231;
  assign new_n3233 = ~pq & new_n3232;
  assign new_n3234 = ~pr & new_n3233;
  assign new_n3235 = ~pc0 & new_n3098;
  assign new_n3236 = ~pd0 & new_n3235;
  assign new_n3237 = pl0 & new_n3236;
  assign new_n3238 = ~pg0 & new_n3237;
  assign new_n3239 = ~py & new_n3238;
  assign new_n3240 = ~pb0 & new_n3239;
  assign new_n3241 = ~px & new_n3240;
  assign new_n3242 = ~pr & new_n3241;
  assign new_n3243 = ~pt & new_n3242;
  assign new_n3244 = ~pl & new_n3243;
  assign new_n3245 = ~pq & new_n3244;
  assign new_n3246 = ~pu & new_n583;
  assign new_n3247 = ~pa & new_n3246;
  assign new_n3248 = ~pm & new_n3247;
  assign new_n3249 = ~pe0 & new_n3248;
  assign new_n3250 = ~pj0 & new_n3249;
  assign new_n3251 = ~po & new_n3250;
  assign new_n3252 = ~pg0 & new_n3251;
  assign new_n3253 = ~pc0 & new_n3252;
  assign new_n3254 = pl0 & new_n3253;
  assign new_n3255 = ~pa0 & new_n3254;
  assign new_n3256 = ~pb0 & new_n3255;
  assign new_n3257 = ~pi & new_n3210;
  assign new_n3258 = ~pq & new_n3257;
  assign new_n3259 = ~pa & new_n3258;
  assign new_n3260 = ~po & new_n3259;
  assign new_n3261 = ~pe0 & new_n3260;
  assign new_n3262 = pl0 & new_n3261;
  assign new_n3263 = ~pj0 & new_n3262;
  assign new_n3264 = ~pc0 & new_n3263;
  assign new_n3265 = ~pa0 & new_n3264;
  assign new_n3266 = ~pb0 & new_n3265;
  assign new_n3267 = ~px & new_n3266;
  assign new_n3268 = ~py & new_n3267;
  assign new_n3269 = ~pd0 & new_n3223;
  assign new_n3270 = pl0 & new_n3269;
  assign new_n3271 = ~pg0 & new_n3270;
  assign new_n3272 = pj0 & new_n3271;
  assign new_n3273 = ~pb0 & new_n3272;
  assign new_n3274 = ~pc0 & new_n3273;
  assign new_n3275 = ~px & new_n3274;
  assign new_n3276 = ~pr & new_n3275;
  assign new_n3277 = ~pt & new_n3276;
  assign new_n3278 = ~pl & new_n3277;
  assign new_n3279 = ~pq & new_n3278;
  assign new_n3280 = ~pi & new_n3119;
  assign new_n3281 = ~pq & new_n3280;
  assign new_n3282 = ~pa & new_n3281;
  assign new_n3283 = ~pm & new_n3282;
  assign new_n3284 = ~pe0 & new_n3283;
  assign new_n3285 = ~pj0 & new_n3284;
  assign new_n3286 = ~po & new_n3285;
  assign new_n3287 = pl0 & new_n3286;
  assign new_n3288 = ~pb0 & new_n3287;
  assign new_n3289 = ~pc0 & new_n3288;
  assign new_n3290 = ~py & new_n3289;
  assign new_n3291 = ~pa0 & new_n3290;
  assign new_n3292 = ~pj0 & new_n2426;
  assign new_n3293 = ~pe0 & new_n3292;
  assign new_n3294 = ~ph0 & new_n3293;
  assign new_n3295 = pl0 & new_n3294;
  assign new_n3296 = ~pd0 & new_n3295;
  assign new_n3297 = ~pb0 & new_n3296;
  assign new_n3298 = ~pc0 & new_n3297;
  assign new_n3299 = ~py & new_n3298;
  assign new_n3300 = ~pa0 & new_n3299;
  assign new_n3301 = ~px & new_n676;
  assign new_n3302 = ~py & new_n3301;
  assign new_n3303 = ~pq & new_n3302;
  assign new_n3304 = pv & new_n3303;
  assign new_n3305 = pi0 & new_n3304;
  assign new_n3306 = ~pm & new_n3305;
  assign new_n3307 = pd0 & new_n3306;
  assign new_n3308 = ~po & new_n3307;
  assign new_n3309 = ~ph0 & pl0;
  assign new_n3310 = ~pc0 & new_n3309;
  assign new_n3311 = ~pd0 & new_n3310;
  assign new_n3312 = ~ph & new_n3311;
  assign new_n3313 = ~pf0 & new_n3312;
  assign new_n3314 = ~pi0 & new_n3313;
  assign new_n3315 = ~pe0 & new_n3314;
  assign new_n3316 = ~pg0 & new_n3315;
  assign new_n3317 = pj0 & new_n3316;
  assign new_n3318 = pv & ~pw;
  assign new_n3319 = ~pq & new_n3318;
  assign new_n3320 = ~pr & new_n3319;
  assign new_n3321 = ~pn & new_n3320;
  assign new_n3322 = pd0 & new_n3321;
  assign new_n3323 = ~pc0 & new_n3322;
  assign new_n3324 = ~pa0 & new_n3323;
  assign new_n3325 = ~pb0 & new_n3324;
  assign new_n3326 = ~px & new_n3325;
  assign new_n3327 = ~py & new_n3326;
  assign new_n3328 = ~pb0 & new_n3191;
  assign new_n3329 = ~pc0 & new_n3328;
  assign new_n3330 = ~pd0 & new_n3329;
  assign new_n3331 = pl0 & new_n3330;
  assign new_n3332 = ~px & new_n3331;
  assign new_n3333 = ~py & new_n3332;
  assign new_n3334 = ~pt & new_n3333;
  assign new_n3335 = ~pq & new_n3334;
  assign new_n3336 = ~pr & new_n3335;
  assign new_n3337 = ~pj & new_n3336;
  assign new_n3338 = ~pl & new_n3337;
  assign new_n3339 = ~ph & new_n3119;
  assign new_n3340 = ~pq & new_n3339;
  assign new_n3341 = ~pa & new_n3340;
  assign new_n3342 = ~pm & new_n3341;
  assign new_n3343 = ~pe0 & new_n3342;
  assign new_n3344 = ~pg0 & new_n3343;
  assign new_n3345 = ~po & new_n3344;
  assign new_n3346 = pl0 & new_n3345;
  assign new_n3347 = ~pb0 & new_n3346;
  assign new_n3348 = ~pc0 & new_n3347;
  assign new_n3349 = ~py & new_n3348;
  assign new_n3350 = ~pa0 & new_n3349;
  assign new_n3351 = ~pa & new_n1777;
  assign new_n3352 = ~po & new_n3351;
  assign new_n3353 = ~pe0 & new_n3352;
  assign new_n3354 = ~pc0 & new_n3353;
  assign new_n3355 = pl0 & new_n3354;
  assign new_n3356 = ~pb0 & new_n3355;
  assign new_n3357 = ~py & new_n3356;
  assign new_n3358 = ~pa0 & new_n3357;
  assign new_n3359 = ~pu & new_n3358;
  assign new_n3360 = ~px & new_n3359;
  assign new_n3361 = ~pb0 & ~py;
  assign new_n3362 = ~pq & new_n3361;
  assign new_n3363 = ~px & new_n3362;
  assign new_n3364 = ~pn & new_n3363;
  assign new_n3365 = pv & new_n3364;
  assign new_n3366 = pi0 & new_n3365;
  assign new_n3367 = ~pm & new_n3366;
  assign new_n3368 = ~pc0 & new_n3367;
  assign new_n3369 = pd0 & new_n3368;
  assign new_n3370 = ~pg0 & pl0;
  assign new_n3371 = ~pc0 & new_n3370;
  assign new_n3372 = ~pd0 & new_n3371;
  assign new_n3373 = ~ph & new_n3372;
  assign new_n3374 = ~pf0 & new_n3373;
  assign new_n3375 = ~pi0 & new_n3374;
  assign new_n3376 = ~pe0 & new_n3375;
  assign new_n3377 = pj0 & new_n3376;
  assign new_n3378 = ~po & new_n3377;
  assign new_n3379 = ~ph & new_n231;
  assign new_n3380 = ~pi & new_n3379;
  assign new_n3381 = ~pa & new_n3380;
  assign new_n3382 = ~pm & new_n3381;
  assign new_n3383 = ~pe0 & new_n3382;
  assign new_n3384 = pl0 & new_n3383;
  assign new_n3385 = ~po & new_n3384;
  assign new_n3386 = ~pc0 & new_n3385;
  assign new_n3387 = ~pa0 & new_n3386;
  assign new_n3388 = ~pb0 & new_n3387;
  assign new_n3389 = ~px & new_n3388;
  assign new_n3390 = ~py & new_n3389;
  assign new_n3391 = pf0 & new_n3303;
  assign new_n3392 = ~pm & new_n3391;
  assign new_n3393 = ~pe0 & new_n3392;
  assign new_n3394 = pi0 & new_n3393;
  assign new_n3395 = ~pg0 & new_n3394;
  assign new_n3396 = ~po & new_n3395;
  assign new_n3397 = ~pd0 & new_n3396;
  assign new_n3398 = pl0 & new_n3397;
  assign new_n3399 = ~pi & new_n584;
  assign new_n3400 = ~pe0 & new_n3399;
  assign new_n3401 = ~po & new_n3400;
  assign new_n3402 = pi0 & new_n3401;
  assign new_n3403 = ~pj0 & new_n3402;
  assign new_n3404 = ~pd0 & new_n3403;
  assign new_n3405 = pl0 & new_n3404;
  assign new_n3406 = ~pb0 & new_n3405;
  assign new_n3407 = ~pc0 & new_n3406;
  assign new_n3408 = pv & new_n1222;
  assign new_n3409 = ~po & new_n3408;
  assign new_n3410 = ~pi0 & new_n3409;
  assign new_n3411 = pd0 & new_n3410;
  assign new_n3412 = pj0 & new_n3411;
  assign new_n3413 = ph & new_n3158;
  assign new_n3414 = pf0 & new_n3413;
  assign new_n3415 = ~pc0 & new_n3414;
  assign new_n3416 = ~pm & new_n3415;
  assign new_n3417 = ~pa0 & new_n3416;
  assign new_n3418 = ~pb0 & new_n3417;
  assign new_n3419 = pl0 & new_n3161;
  assign new_n3420 = ~pj0 & new_n3419;
  assign new_n3421 = ~ph0 & new_n3420;
  assign new_n3422 = ~pc0 & new_n3421;
  assign new_n3423 = ~pd0 & new_n3422;
  assign new_n3424 = ~pa0 & new_n3423;
  assign new_n3425 = ~pb0 & new_n3424;
  assign new_n3426 = ~pb0 & new_n824;
  assign new_n3427 = ~pq & new_n3426;
  assign new_n3428 = pf0 & new_n3427;
  assign new_n3429 = ~pm & new_n3428;
  assign new_n3430 = ~pe0 & new_n3429;
  assign new_n3431 = ~pi0 & new_n3430;
  assign new_n3432 = pj0 & new_n3431;
  assign new_n3433 = ~po & new_n3432;
  assign new_n3434 = pl0 & new_n3433;
  assign new_n3435 = ~pg0 & new_n3434;
  assign new_n3436 = ~po & new_n283;
  assign new_n3437 = ~pi0 & new_n3436;
  assign new_n3438 = pj0 & new_n3437;
  assign new_n3439 = ~pd0 & new_n3438;
  assign new_n3440 = pl0 & new_n3439;
  assign new_n3441 = ~pb0 & new_n3440;
  assign new_n3442 = ~pc0 & new_n3441;
  assign new_n3443 = pv & new_n726;
  assign new_n3444 = pj0 & new_n3443;
  assign new_n3445 = ~pi0 & new_n3444;
  assign new_n3446 = ~pc0 & new_n3445;
  assign new_n3447 = pd0 & new_n3446;
  assign new_n3448 = ~pa0 & ~py;
  assign new_n3449 = ~pq & new_n3448;
  assign new_n3450 = ~px & new_n3449;
  assign new_n3451 = ph & new_n3450;
  assign new_n3452 = pf0 & new_n3451;
  assign new_n3453 = ~po & new_n3452;
  assign new_n3454 = ~pm & new_n3453;
  assign new_n3455 = ~pb0 & new_n3454;
  assign new_n3456 = ~pc0 & new_n3455;
  assign new_n3457 = ~pr & new_n207;
  assign new_n3458 = pu & new_n3457;
  assign new_n3459 = ~pq & new_n3458;
  assign new_n3460 = pz & new_n3459;
  assign new_n3461 = ~pi0 & new_n3460;
  assign new_n3462 = pj0 & new_n3461;
  assign new_n3463 = ~po & new_n3462;
  assign new_n3464 = ~pc0 & new_n3463;
  assign new_n3465 = ph0 & new_n3464;
  assign new_n3466 = ~ph & new_n825;
  assign new_n3467 = ~pf0 & new_n3466;
  assign new_n3468 = ~pe0 & new_n3467;
  assign new_n3469 = ~pg0 & new_n3468;
  assign new_n3470 = pi0 & new_n3469;
  assign new_n3471 = ~ph0 & new_n3470;
  assign new_n3472 = pl0 & new_n3471;
  assign new_n3473 = ~pr & new_n3361;
  assign new_n3474 = ~px & new_n3473;
  assign new_n3475 = ~pq & new_n3474;
  assign new_n3476 = pv & new_n3475;
  assign new_n3477 = ~po & new_n3476;
  assign new_n3478 = pi0 & new_n3477;
  assign new_n3479 = ~pc0 & new_n3478;
  assign new_n3480 = pd0 & new_n3479;
  assign new_n3481 = ~pb0 & new_n1010;
  assign new_n3482 = ~pc0 & new_n3481;
  assign new_n3483 = ~py & new_n3482;
  assign new_n3484 = ~pa0 & new_n3483;
  assign new_n3485 = ~po & new_n3320;
  assign new_n3486 = pd0 & new_n3485;
  assign new_n3487 = ~pc0 & new_n3486;
  assign new_n3488 = ~pa0 & new_n3487;
  assign new_n3489 = ~pb0 & new_n3488;
  assign new_n3490 = ~px & new_n3489;
  assign new_n3491 = ~py & new_n3490;
  assign new_n3492 = pz & new_n726;
  assign new_n3493 = ~pi0 & new_n3492;
  assign new_n3494 = ph0 & new_n3493;
  assign new_n3495 = pj0 & new_n3494;
  assign new_n3496 = ~pc0 & new_n3495;
  assign new_n3497 = ~pd0 & new_n3496;
  assign new_n3498 = ~pd0 & ~ph0;
  assign new_n3499 = ~py & new_n3498;
  assign new_n3500 = ~pc0 & new_n3499;
  assign new_n3501 = ~px & new_n3500;
  assign new_n3502 = ~pf0 & new_n3501;
  assign new_n3503 = ~pe0 & new_n3502;
  assign new_n3504 = ~pj0 & new_n3503;
  assign new_n3505 = pi0 & new_n3504;
  assign new_n3506 = pl0 & new_n3505;
  assign new_n3507 = ~pg0 & new_n3506;
  assign new_n3508 = pv & new_n3001;
  assign new_n3509 = pd0 & new_n3508;
  assign new_n3510 = pi0 & new_n3509;
  assign new_n3511 = ~pb0 & new_n3510;
  assign new_n3512 = ~pc0 & new_n3511;
  assign new_n3513 = ph & new_n584;
  assign new_n3514 = pf0 & new_n3513;
  assign new_n3515 = ~pc0 & new_n3514;
  assign new_n3516 = ~po & new_n3515;
  assign new_n3517 = ~pa0 & new_n3516;
  assign new_n3518 = ~pb0 & new_n3517;
  assign new_n3519 = ph & new_n209;
  assign new_n3520 = pf0 & new_n3519;
  assign new_n3521 = ~pi0 & new_n3520;
  assign new_n3522 = pj0 & new_n3521;
  assign new_n3523 = ~po & new_n3522;
  assign new_n3524 = ~pc0 & new_n3523;
  assign new_n3525 = ~pd0 & new_n3524;
  assign new_n3526 = pv & new_n679;
  assign new_n3527 = ~pi0 & new_n3526;
  assign new_n3528 = ~pm & new_n3527;
  assign new_n3529 = pd0 & new_n3528;
  assign new_n3530 = pj0 & new_n3529;
  assign new_n3531 = ~pc0 & ph0;
  assign new_n3532 = ~py & new_n3531;
  assign new_n3533 = ~pa0 & new_n3532;
  assign new_n3534 = pu & new_n3533;
  assign new_n3535 = pz & new_n3534;
  assign new_n3536 = ~pe0 & new_n3535;
  assign new_n3537 = ~pf0 & new_n3536;
  assign new_n3538 = ~pg0 & new_n3537;
  assign new_n3539 = ~pi0 & new_n3538;
  assign new_n3540 = pd0 & ~pg0;
  assign new_n3541 = ~py & new_n3540;
  assign new_n3542 = ~pc0 & new_n3541;
  assign new_n3543 = ~px & new_n3542;
  assign new_n3544 = ~pf0 & new_n3543;
  assign new_n3545 = pv & new_n3544;
  assign new_n3546 = pi0 & new_n3545;
  assign new_n3547 = ~pe0 & new_n3546;
  assign new_n3548 = pu & ~px;
  assign new_n3549 = ~pq & new_n3548;
  assign new_n3550 = ~pr & new_n3549;
  assign new_n3551 = ph & new_n3550;
  assign new_n3552 = pf0 & new_n3551;
  assign new_n3553 = ~pi0 & new_n3552;
  assign new_n3554 = pj0 & new_n3553;
  assign new_n3555 = ~po & new_n3554;
  assign new_n3556 = ~pb0 & new_n3555;
  assign new_n3557 = ~pc0 & new_n3556;
  assign new_n3558 = pv & new_n940;
  assign new_n3559 = ~pi0 & new_n3558;
  assign new_n3560 = ~pm & new_n3559;
  assign new_n3561 = pj0 & new_n3560;
  assign new_n3562 = ~po & new_n3561;
  assign new_n3563 = ~px & new_n3531;
  assign new_n3564 = ~py & new_n3563;
  assign new_n3565 = pu & new_n3564;
  assign new_n3566 = pz & new_n3565;
  assign new_n3567 = ~pe0 & new_n3566;
  assign new_n3568 = ~pf0 & new_n3567;
  assign new_n3569 = ~pg0 & new_n3568;
  assign new_n3570 = pi0 & new_n3569;
  assign new_n3571 = ~pa0 & new_n3540;
  assign new_n3572 = ~pc0 & new_n3571;
  assign new_n3573 = ~py & new_n3572;
  assign new_n3574 = ~pf0 & new_n3573;
  assign new_n3575 = pv & new_n3574;
  assign new_n3576 = ~pi0 & new_n3575;
  assign new_n3577 = ~pe0 & new_n3576;
  assign new_n3578 = ~pn & new_n3318;
  assign new_n3579 = ~pq & new_n3578;
  assign new_n3580 = ~pm & new_n3579;
  assign new_n3581 = pd0 & new_n3580;
  assign new_n3582 = ~pc0 & new_n3581;
  assign new_n3583 = ~pa0 & new_n3582;
  assign new_n3584 = ~pb0 & new_n3583;
  assign new_n3585 = ~px & new_n3584;
  assign new_n3586 = ~py & new_n3585;
  assign new_n3587 = ~pg0 & new_n2868;
  assign new_n3588 = ~po & new_n3587;
  assign new_n3589 = ~pa0 & new_n3588;
  assign new_n3590 = ~pb0 & new_n3589;
  assign new_n3591 = ~pc0 & new_n3590;
  assign new_n3592 = pd0 & new_n3591;
  assign new_n3593 = ~px & new_n3592;
  assign new_n3594 = ~py & new_n3593;
  assign new_n3595 = ~pu & new_n3594;
  assign new_n3596 = ~pq & new_n3595;
  assign new_n3597 = ~pr & new_n3596;
  assign new_n3598 = ~pj & new_n3597;
  assign new_n3599 = pn & new_n3598;
  assign new_n3600 = pi0 & new_n1058;
  assign new_n3601 = ~pb & new_n3600;
  assign new_n3602 = ~pd0 & new_n3601;
  assign new_n3603 = ~ph0 & new_n3602;
  assign new_n3604 = pl0 & new_n3603;
  assign new_n3605 = ~pc & new_n3604;
  assign new_n3606 = ~pb0 & new_n3605;
  assign new_n3607 = ~pc0 & new_n3606;
  assign new_n3608 = ~py & new_n3607;
  assign new_n3609 = ~pr & new_n3608;
  assign new_n3610 = ~px & new_n3609;
  assign new_n3611 = ~pn & new_n3610;
  assign new_n3612 = ~pq & new_n3611;
  assign new_n3613 = pi0 & new_n1333;
  assign new_n3614 = ~pk & new_n3613;
  assign new_n3615 = pl0 & new_n3614;
  assign new_n3616 = ~pg0 & new_n3615;
  assign new_n3617 = ~po & new_n3616;
  assign new_n3618 = ~pc & new_n3617;
  assign new_n3619 = ~pc0 & new_n3618;
  assign new_n3620 = ~pd0 & new_n3619;
  assign new_n3621 = ~pb0 & new_n3620;
  assign new_n3622 = ~px & new_n3621;
  assign new_n3623 = ~py & new_n3622;
  assign new_n3624 = ~pq & new_n3623;
  assign new_n3625 = ~pr & new_n3624;
  assign new_n3626 = ~pc0 & new_n2988;
  assign new_n3627 = ~pd0 & new_n3626;
  assign new_n3628 = pl0 & new_n3627;
  assign new_n3629 = ~pj0 & new_n3628;
  assign new_n3630 = ~pa0 & new_n3629;
  assign new_n3631 = ~pb0 & new_n3630;
  assign new_n3632 = ~py & new_n3631;
  assign new_n3633 = ~pr & new_n3632;
  assign new_n3634 = ~px & new_n3633;
  assign new_n3635 = pn & new_n3634;
  assign new_n3636 = ~pq & new_n3635;
  assign new_n3637 = ~pr & new_n3448;
  assign new_n3638 = ~px & new_n3637;
  assign new_n3639 = ~pq & new_n3638;
  assign new_n3640 = pf0 & new_n3639;
  assign new_n3641 = ~po & new_n3640;
  assign new_n3642 = ~pe0 & new_n3641;
  assign new_n3643 = ~pg0 & new_n3642;
  assign new_n3644 = ~pd0 & new_n3643;
  assign new_n3645 = pl0 & new_n3644;
  assign new_n3646 = ~pb0 & new_n3645;
  assign new_n3647 = ~pc0 & new_n3646;
  assign new_n3648 = pu & new_n208;
  assign new_n3649 = ~pn & new_n3648;
  assign new_n3650 = pz & new_n3649;
  assign new_n3651 = ~pm & new_n3650;
  assign new_n3652 = pj0 & new_n3651;
  assign new_n3653 = ~pi0 & new_n3652;
  assign new_n3654 = ~pc0 & new_n3653;
  assign new_n3655 = ph0 & new_n3654;
  assign new_n3656 = ~pa0 & new_n3498;
  assign new_n3657 = ~pc0 & new_n3656;
  assign new_n3658 = ~py & new_n3657;
  assign new_n3659 = ~pf0 & new_n3658;
  assign new_n3660 = ~pe0 & new_n3659;
  assign new_n3661 = ~pj0 & new_n3660;
  assign new_n3662 = ~pi0 & new_n3661;
  assign new_n3663 = pl0 & new_n3662;
  assign new_n3664 = ~pg0 & new_n3663;
  assign new_n3665 = ~pm & new_n3414;
  assign new_n3666 = ~pd0 & new_n3665;
  assign new_n3667 = pi0 & new_n3666;
  assign new_n3668 = ~pb0 & new_n3667;
  assign new_n3669 = ~pc0 & new_n3668;
  assign new_n3670 = ~pn & new_n3121;
  assign new_n3671 = pc & new_n3670;
  assign new_n3672 = pd0 & new_n3671;
  assign new_n3673 = ~pb0 & new_n3672;
  assign new_n3674 = ~pc0 & new_n3673;
  assign new_n3675 = ~py & new_n3674;
  assign new_n3676 = ~pa0 & new_n3675;
  assign new_n3677 = ~pn & new_n3450;
  assign new_n3678 = pz & new_n3677;
  assign new_n3679 = ph0 & new_n3678;
  assign new_n3680 = ~pm & new_n3679;
  assign new_n3681 = ~pb0 & new_n3680;
  assign new_n3682 = ~pc0 & new_n3681;
  assign new_n3683 = pd0 & new_n636;
  assign new_n3684 = ~pg0 & new_n3683;
  assign new_n3685 = ~pc0 & new_n3684;
  assign new_n3686 = pv & new_n3685;
  assign new_n3687 = ~pe0 & new_n3686;
  assign new_n3688 = ~pf0 & new_n3687;
  assign new_n3689 = pd0 & new_n2867;
  assign new_n3690 = pl0 & new_n3689;
  assign new_n3691 = ~po & new_n3690;
  assign new_n3692 = ~py & new_n3691;
  assign new_n3693 = ~pa0 & new_n3692;
  assign new_n3694 = ~pb0 & new_n3693;
  assign new_n3695 = ~pc0 & new_n3694;
  assign new_n3696 = ~pu & new_n3695;
  assign new_n3697 = ~px & new_n3696;
  assign new_n3698 = ~pr & new_n3697;
  assign new_n3699 = pn & new_n3698;
  assign new_n3700 = ~pq & new_n3699;
  assign new_n3701 = ~pi & new_n3700;
  assign new_n3702 = ~pj & new_n3701;
  assign new_n3703 = pi0 & new_n1181;
  assign new_n3704 = ~pb & new_n3703;
  assign new_n3705 = ~ph0 & new_n3704;
  assign new_n3706 = pl0 & new_n3705;
  assign new_n3707 = ~pg0 & new_n3706;
  assign new_n3708 = ~pc & new_n3707;
  assign new_n3709 = ~pc0 & new_n3708;
  assign new_n3710 = ~pd0 & new_n3709;
  assign new_n3711 = ~pb0 & new_n3710;
  assign new_n3712 = ~px & new_n3711;
  assign new_n3713 = ~py & new_n3712;
  assign new_n3714 = ~pq & new_n3713;
  assign new_n3715 = ~pr & new_n3714;
  assign new_n3716 = ~pk & new_n3600;
  assign new_n3717 = ~pd0 & new_n3716;
  assign new_n3718 = pl0 & new_n3717;
  assign new_n3719 = ~po & new_n3718;
  assign new_n3720 = ~pc & new_n3719;
  assign new_n3721 = ~pb0 & new_n3720;
  assign new_n3722 = ~pc0 & new_n3721;
  assign new_n3723 = ~py & new_n3722;
  assign new_n3724 = ~pr & new_n3723;
  assign new_n3725 = ~px & new_n3724;
  assign new_n3726 = ~pj & new_n3725;
  assign new_n3727 = ~pq & new_n3726;
  assign new_n3728 = ~po & new_n45;
  assign new_n3729 = ~pc & new_n3728;
  assign new_n3730 = ~pd0 & new_n3729;
  assign new_n3731 = pl0 & new_n3730;
  assign new_n3732 = ~pg0 & new_n3731;
  assign new_n3733 = ~pj0 & new_n3732;
  assign new_n3734 = ~pb0 & new_n3733;
  assign new_n3735 = ~pc0 & new_n3734;
  assign new_n3736 = ~pa0 & new_n3735;
  assign new_n3737 = ~px & new_n3736;
  assign new_n3738 = ~py & new_n3737;
  assign new_n3739 = ~pq & new_n3738;
  assign new_n3740 = ~pr & new_n3739;
  assign new_n3741 = pf0 & new_n3475;
  assign new_n3742 = pi0 & new_n3741;
  assign new_n3743 = ~pe0 & new_n3742;
  assign new_n3744 = ~po & new_n3743;
  assign new_n3745 = pl0 & new_n3744;
  assign new_n3746 = ~pg0 & new_n3745;
  assign new_n3747 = ~pc0 & new_n3746;
  assign new_n3748 = ~pd0 & new_n3747;
  assign new_n3749 = pu & new_n3361;
  assign new_n3750 = ~px & new_n3749;
  assign new_n3751 = ~pq & new_n3750;
  assign new_n3752 = pz & new_n3751;
  assign new_n3753 = ~pm & new_n3752;
  assign new_n3754 = ~po & new_n3753;
  assign new_n3755 = pi0 & new_n3754;
  assign new_n3756 = ~pc0 & new_n3755;
  assign new_n3757 = ph0 & new_n3756;
  assign new_n3758 = ~pd0 & pl0;
  assign new_n3759 = ~pa0 & new_n3758;
  assign new_n3760 = ~pc0 & new_n3759;
  assign new_n3761 = ~py & new_n3760;
  assign new_n3762 = ~pf0 & new_n3761;
  assign new_n3763 = ~pe0 & new_n3762;
  assign new_n3764 = ~po & new_n3763;
  assign new_n3765 = ~pi0 & new_n3764;
  assign new_n3766 = ~pg0 & new_n3765;
  assign new_n3767 = ~pj0 & new_n3766;
  assign new_n3768 = ~pn & new_n3548;
  assign new_n3769 = ~pq & new_n3768;
  assign new_n3770 = ph & new_n3769;
  assign new_n3771 = pf0 & new_n3770;
  assign new_n3772 = ~pm & new_n3771;
  assign new_n3773 = ~pc0 & new_n3772;
  assign new_n3774 = pi0 & new_n3773;
  assign new_n3775 = ~py & new_n3774;
  assign new_n3776 = ~pb0 & new_n3775;
  assign new_n3777 = ~pr & new_n582;
  assign new_n3778 = ~pu & new_n3777;
  assign new_n3779 = ~pq & new_n3778;
  assign new_n3780 = pc & new_n3779;
  assign new_n3781 = ~po & new_n3780;
  assign new_n3782 = ~pc0 & new_n3781;
  assign new_n3783 = pd0 & new_n3782;
  assign new_n3784 = ~pa0 & new_n3783;
  assign new_n3785 = ~pb0 & new_n3784;
  assign new_n3786 = pz & new_n3001;
  assign new_n3787 = ~pc0 & new_n3786;
  assign new_n3788 = ph0 & new_n3787;
  assign new_n3789 = ~pa0 & new_n3788;
  assign new_n3790 = ~pb0 & new_n3789;
  assign new_n3791 = ~pc0 & new_n685;
  assign new_n3792 = ph0 & new_n3791;
  assign new_n3793 = pu & new_n3792;
  assign new_n3794 = ~pf0 & new_n3793;
  assign new_n3795 = pz & new_n3794;
  assign new_n3796 = ~pi0 & new_n3795;
  assign new_n3797 = ~pe0 & new_n3796;
  assign new_n3798 = ~pa & new_n78;
  assign new_n3799 = ~pj0 & new_n3798;
  assign new_n3800 = ~pm & new_n3799;
  assign new_n3801 = pd0 & new_n3800;
  assign new_n3802 = ~ph0 & new_n3801;
  assign new_n3803 = pl0 & new_n3802;
  assign new_n3804 = ~pg0 & new_n3803;
  assign new_n3805 = ~pb0 & new_n3804;
  assign new_n3806 = ~pc0 & new_n3805;
  assign new_n3807 = ~pa0 & new_n3806;
  assign new_n3808 = ~px & new_n3807;
  assign new_n3809 = ~py & new_n3808;
  assign new_n3810 = ~pq & new_n3809;
  assign new_n3811 = ~pu & new_n3810;
  assign new_n3812 = ~pc & new_n478;
  assign new_n3813 = ~pb & new_n3812;
  assign new_n3814 = ~pd0 & new_n3813;
  assign new_n3815 = ~ph0 & new_n3814;
  assign new_n3816 = pl0 & new_n3815;
  assign new_n3817 = ~pj0 & new_n3816;
  assign new_n3818 = ~pb0 & new_n3817;
  assign new_n3819 = ~pc0 & new_n3818;
  assign new_n3820 = ~pa0 & new_n3819;
  assign new_n3821 = ~px & new_n3820;
  assign new_n3822 = ~py & new_n3821;
  assign new_n3823 = ~pq & new_n3822;
  assign new_n3824 = ~pr & new_n3823;
  assign new_n3825 = pi0 & new_n2900;
  assign new_n3826 = ~pk & new_n3825;
  assign new_n3827 = ~pg0 & new_n3826;
  assign new_n3828 = ~pj0 & new_n3827;
  assign new_n3829 = ~po & new_n3828;
  assign new_n3830 = ~pc & new_n3829;
  assign new_n3831 = ~pd0 & new_n3830;
  assign new_n3832 = pl0 & new_n3831;
  assign new_n3833 = ~pc0 & new_n3832;
  assign new_n3834 = ~py & new_n3833;
  assign new_n3835 = ~pb0 & new_n3834;
  assign new_n3836 = ~pr & new_n3835;
  assign new_n3837 = ~px & new_n3836;
  assign new_n3838 = ~pc0 & new_n2884;
  assign new_n3839 = ~pd0 & new_n3838;
  assign new_n3840 = pl0 & new_n3839;
  assign new_n3841 = ~po & new_n3840;
  assign new_n3842 = ~py & new_n3841;
  assign new_n3843 = ~pb0 & new_n3842;
  assign new_n3844 = ~px & new_n3843;
  assign new_n3845 = ~pq & new_n3844;
  assign new_n3846 = ~pr & new_n3845;
  assign new_n3847 = ~pj & new_n3846;
  assign new_n3848 = pn & new_n3847;
  assign new_n3849 = pf0 & new_n1222;
  assign new_n3850 = ~pi0 & new_n3849;
  assign new_n3851 = ~pe0 & new_n3850;
  assign new_n3852 = ~po & new_n3851;
  assign new_n3853 = ~pg0 & new_n3852;
  assign new_n3854 = pj0 & new_n3853;
  assign new_n3855 = ~pd0 & new_n3854;
  assign new_n3856 = pl0 & new_n3855;
  assign new_n3857 = pz & new_n3364;
  assign new_n3858 = ~pm & new_n3857;
  assign new_n3859 = ph0 & new_n3858;
  assign new_n3860 = pi0 & new_n3859;
  assign new_n3861 = ~pc0 & new_n3860;
  assign new_n3862 = ~pd0 & new_n3861;
  assign new_n3863 = ~po & new_n3468;
  assign new_n3864 = pi0 & new_n3863;
  assign new_n3865 = pl0 & new_n3864;
  assign new_n3866 = ~pg0 & new_n3865;
  assign new_n3867 = ph & new_n3363;
  assign new_n3868 = pf0 & new_n3867;
  assign new_n3869 = ~pm & new_n3868;
  assign new_n3870 = ~po & new_n3869;
  assign new_n3871 = pi0 & new_n3870;
  assign new_n3872 = ~pc0 & new_n3871;
  assign new_n3873 = ~pd0 & new_n3872;
  assign new_n3874 = ~pr & pu;
  assign new_n3875 = ~pn & new_n3874;
  assign new_n3876 = ~pq & new_n3875;
  assign new_n3877 = ph & new_n3876;
  assign new_n3878 = pf0 & new_n3877;
  assign new_n3879 = pi0 & new_n3878;
  assign new_n3880 = ~pb0 & new_n3879;
  assign new_n3881 = ~pc0 & new_n3880;
  assign new_n3882 = ~px & new_n3881;
  assign new_n3883 = ~py & new_n3882;
  assign new_n3884 = ~pc0 & new_n3081;
  assign new_n3885 = pd0 & new_n3884;
  assign new_n3886 = ~ph0 & new_n3885;
  assign new_n3887 = pl0 & new_n3886;
  assign new_n3888 = ~px & new_n3887;
  assign new_n3889 = ~py & new_n3888;
  assign new_n3890 = ~pa0 & new_n3889;
  assign new_n3891 = ~pb0 & new_n3890;
  assign new_n3892 = ~pt & new_n3891;
  assign new_n3893 = ~pj0 & new_n3892;
  assign new_n3894 = ~pu & new_n3893;
  assign new_n3895 = ~pr & new_n3894;
  assign new_n3896 = ~pn & new_n3895;
  assign new_n3897 = ~pq & new_n3896;
  assign new_n3898 = ~pj & new_n3897;
  assign new_n3899 = ~pl & new_n3898;
  assign new_n3900 = ~pm & new_n3082;
  assign new_n3901 = ~pc0 & new_n3900;
  assign new_n3902 = pd0 & new_n3901;
  assign new_n3903 = ~ph0 & new_n3902;
  assign new_n3904 = pl0 & new_n3903;
  assign new_n3905 = ~pa0 & new_n3904;
  assign new_n3906 = ~pb0 & new_n3905;
  assign new_n3907 = ~py & new_n3906;
  assign new_n3908 = ~pu & new_n3907;
  assign new_n3909 = ~px & new_n3908;
  assign new_n3910 = ~pn & new_n3909;
  assign new_n3911 = ~pq & new_n3910;
  assign new_n3912 = ~pc & new_n441;
  assign new_n3913 = ~pb & new_n3912;
  assign new_n3914 = ~ph0 & new_n3913;
  assign new_n3915 = pl0 & new_n3914;
  assign new_n3916 = ~pg0 & new_n3915;
  assign new_n3917 = ~pj0 & new_n3916;
  assign new_n3918 = ~pc0 & new_n3917;
  assign new_n3919 = ~pd0 & new_n3918;
  assign new_n3920 = ~pb0 & new_n3919;
  assign new_n3921 = ~py & new_n3920;
  assign new_n3922 = ~pa0 & new_n3921;
  assign new_n3923 = ~pr & new_n3922;
  assign new_n3924 = ~px & new_n3923;
  assign new_n3925 = pi0 & new_n105;
  assign new_n3926 = ~pk & new_n3925;
  assign new_n3927 = pl0 & new_n3926;
  assign new_n3928 = ~pj0 & new_n3927;
  assign new_n3929 = ~po & new_n3928;
  assign new_n3930 = ~pc & new_n3929;
  assign new_n3931 = ~pc0 & new_n3930;
  assign new_n3932 = ~pd0 & new_n3931;
  assign new_n3933 = ~pb0 & new_n3932;
  assign new_n3934 = ~px & new_n3933;
  assign new_n3935 = ~py & new_n3934;
  assign new_n3936 = ~pq & new_n3935;
  assign new_n3937 = ~pr & new_n3936;
  assign new_n3938 = ~pc & new_n1333;
  assign new_n3939 = pi0 & new_n3938;
  assign new_n3940 = ~pd0 & new_n3939;
  assign new_n3941 = pl0 & new_n3940;
  assign new_n3942 = ~pg0 & new_n3941;
  assign new_n3943 = ~po & new_n3942;
  assign new_n3944 = ~pb0 & new_n3943;
  assign new_n3945 = ~pc0 & new_n3944;
  assign new_n3946 = ~py & new_n3945;
  assign new_n3947 = ~pr & new_n3946;
  assign new_n3948 = ~px & new_n3947;
  assign new_n3949 = pn & new_n3948;
  assign new_n3950 = ~pq & new_n3949;
  assign new_n3951 = ~pa0 & ~pb0;
  assign new_n3952 = ~px & new_n3951;
  assign new_n3953 = ~py & new_n3952;
  assign new_n3954 = ~pq & new_n3953;
  assign new_n3955 = pf0 & new_n3954;
  assign new_n3956 = ~pm & new_n3955;
  assign new_n3957 = ~pe0 & new_n3956;
  assign new_n3958 = ~po & new_n3957;
  assign new_n3959 = pl0 & new_n3958;
  assign new_n3960 = ~pg0 & new_n3959;
  assign new_n3961 = ~pc0 & new_n3960;
  assign new_n3962 = ~pd0 & new_n3961;
  assign new_n3963 = pu & new_n583;
  assign new_n3964 = ~pn & new_n3963;
  assign new_n3965 = pz & new_n3964;
  assign new_n3966 = ~pm & new_n3965;
  assign new_n3967 = ph0 & new_n3966;
  assign new_n3968 = pi0 & new_n3967;
  assign new_n3969 = ~pb0 & new_n3968;
  assign new_n3970 = ~pc0 & new_n3969;
  assign new_n3971 = ~py & new_n3758;
  assign new_n3972 = ~pc0 & new_n3971;
  assign new_n3973 = ~px & new_n3972;
  assign new_n3974 = ~pf0 & new_n3973;
  assign new_n3975 = ~pe0 & new_n3974;
  assign new_n3976 = ~po & new_n3975;
  assign new_n3977 = pi0 & new_n3976;
  assign new_n3978 = ~pg0 & new_n3977;
  assign new_n3979 = ~pj0 & new_n3978;
  assign new_n3980 = ph & new_n3963;
  assign new_n3981 = pf0 & new_n3980;
  assign new_n3982 = ~pm & new_n3981;
  assign new_n3983 = ~po & new_n3982;
  assign new_n3984 = pi0 & new_n3983;
  assign new_n3985 = ~pb0 & new_n3984;
  assign new_n3986 = ~pc0 & new_n3985;
  assign new_n3987 = pi0 & new_n1010;
  assign new_n3988 = ~pc0 & new_n3987;
  assign new_n3989 = ~pd0 & new_n3988;
  assign new_n3990 = ~py & new_n3989;
  assign new_n3991 = ~pb0 & new_n3990;
  assign new_n3992 = ~po & new_n3318;
  assign new_n3993 = ~pq & new_n3992;
  assign new_n3994 = ~pm & new_n3993;
  assign new_n3995 = pd0 & new_n3994;
  assign new_n3996 = ~pc0 & new_n3995;
  assign new_n3997 = ~pa0 & new_n3996;
  assign new_n3998 = ~pb0 & new_n3997;
  assign new_n3999 = ~px & new_n3998;
  assign new_n4000 = ~py & new_n3999;
  assign new_n4001 = ~pg0 & new_n1333;
  assign new_n4002 = pj0 & new_n4001;
  assign new_n4003 = ~pc & new_n4002;
  assign new_n4004 = ~pi0 & new_n4003;
  assign new_n4005 = ~pc0 & new_n4004;
  assign new_n4006 = ~pd0 & new_n4005;
  assign new_n4007 = ~ph0 & new_n4006;
  assign new_n4008 = pl0 & new_n4007;
  assign new_n4009 = ~px & new_n4008;
  assign new_n4010 = ~pb0 & new_n4009;
  assign new_n4011 = ~pt & new_n4010;
  assign new_n4012 = ~pq & new_n4011;
  assign new_n4013 = ~pr & new_n4012;
  assign new_n4014 = ~pl & new_n4013;
  assign new_n4015 = ~pn & new_n4014;
  assign new_n4016 = pl0 & new_n442;
  assign new_n4017 = ~pg0 & new_n4016;
  assign new_n4018 = ~pj0 & new_n4017;
  assign new_n4019 = ~pc & new_n4018;
  assign new_n4020 = ~pd0 & new_n4019;
  assign new_n4021 = ~ph0 & new_n4020;
  assign new_n4022 = ~pc0 & new_n4021;
  assign new_n4023 = ~pa0 & new_n4022;
  assign new_n4024 = ~pb0 & new_n4023;
  assign new_n4025 = ~px & new_n4024;
  assign new_n4026 = ~py & new_n4025;
  assign new_n4027 = ~pb & new_n1058;
  assign new_n4028 = pl0 & new_n4027;
  assign new_n4029 = ~po & new_n4028;
  assign new_n4030 = ~pc & new_n4029;
  assign new_n4031 = pi0 & new_n4030;
  assign new_n4032 = ~pc0 & new_n4031;
  assign new_n4033 = ~pd0 & new_n4032;
  assign new_n4034 = ~pb0 & new_n4033;
  assign new_n4035 = ~px & new_n4034;
  assign new_n4036 = ~py & new_n4035;
  assign new_n4037 = ~pq & new_n4036;
  assign new_n4038 = ~pr & new_n4037;
  assign new_n4039 = ~pn & new_n3119;
  assign new_n4040 = ~pq & new_n4039;
  assign new_n4041 = ~pa & new_n4040;
  assign new_n4042 = ~pj0 & new_n4041;
  assign new_n4043 = ~pm & new_n4042;
  assign new_n4044 = ~pe0 & new_n4043;
  assign new_n4045 = pl0 & new_n4044;
  assign new_n4046 = ~pg0 & new_n4045;
  assign new_n4047 = ~ph0 & new_n4046;
  assign new_n4048 = ~pb0 & new_n4047;
  assign new_n4049 = ~pc0 & new_n4048;
  assign new_n4050 = ~py & new_n4049;
  assign new_n4051 = ~pa0 & new_n4050;
  assign new_n4052 = ~pe0 & new_n726;
  assign new_n4053 = pf0 & new_n4052;
  assign new_n4054 = pj0 & new_n4053;
  assign new_n4055 = ~pi0 & new_n4054;
  assign new_n4056 = ~pg0 & new_n4055;
  assign new_n4057 = ~ph0 & new_n4056;
  assign new_n4058 = pl0 & new_n4057;
  assign new_n4059 = ~pc0 & new_n4058;
  assign new_n4060 = ~pd0 & new_n4059;
  assign new_n4061 = ~pi & new_n3450;
  assign new_n4062 = ~pe0 & new_n4061;
  assign new_n4063 = ~po & new_n4062;
  assign new_n4064 = ~pm & new_n4063;
  assign new_n4065 = ~pj0 & new_n4064;
  assign new_n4066 = ~pd0 & new_n4065;
  assign new_n4067 = pl0 & new_n4066;
  assign new_n4068 = ~pb0 & new_n4067;
  assign new_n4069 = ~pc0 & new_n4068;
  assign new_n4070 = pi0 & new_n3436;
  assign new_n4071 = pl0 & new_n4070;
  assign new_n4072 = ~pc0 & new_n4071;
  assign new_n4073 = ~pd0 & new_n4072;
  assign new_n4074 = ~py & new_n4073;
  assign new_n4075 = ~pb0 & new_n4074;
  assign new_n4076 = pu & new_n3777;
  assign new_n4077 = ~pq & new_n4076;
  assign new_n4078 = pz & new_n4077;
  assign new_n4079 = pi0 & new_n4078;
  assign new_n4080 = ph0 & new_n4079;
  assign new_n4081 = ~po & new_n4080;
  assign new_n4082 = ~pb0 & new_n4081;
  assign new_n4083 = ~pc0 & new_n4082;
  assign new_n4084 = pj0 & new_n1267;
  assign new_n4085 = ~pi0 & new_n4084;
  assign new_n4086 = ~pc0 & new_n4085;
  assign new_n4087 = ~pd0 & new_n4086;
  assign new_n4088 = pi0 & new_n3552;
  assign new_n4089 = ~pc0 & new_n4088;
  assign new_n4090 = ~po & new_n4089;
  assign new_n4091 = ~py & new_n4090;
  assign new_n4092 = ~pb0 & new_n4091;
  assign new_n4093 = ~ph0 & new_n1058;
  assign new_n4094 = pl0 & new_n4093;
  assign new_n4095 = ~pc & new_n4094;
  assign new_n4096 = pi0 & new_n4095;
  assign new_n4097 = ~py & new_n4096;
  assign new_n4098 = ~pb0 & new_n4097;
  assign new_n4099 = ~pc0 & new_n4098;
  assign new_n4100 = ~pd0 & new_n4099;
  assign new_n4101 = ~pt & new_n4100;
  assign new_n4102 = ~px & new_n4101;
  assign new_n4103 = ~pr & new_n4102;
  assign new_n4104 = ~pn & new_n4103;
  assign new_n4105 = ~pq & new_n4104;
  assign new_n4106 = ~pj & new_n4105;
  assign new_n4107 = ~pl & new_n4106;
  assign new_n4108 = ~ph0 & new_n479;
  assign new_n4109 = pl0 & new_n4108;
  assign new_n4110 = ~pj0 & new_n4109;
  assign new_n4111 = ~pc & new_n4110;
  assign new_n4112 = ~pc0 & new_n4111;
  assign new_n4113 = ~pd0 & new_n4112;
  assign new_n4114 = ~pb0 & new_n4113;
  assign new_n4115 = ~py & new_n4114;
  assign new_n4116 = ~pa0 & new_n4115;
  assign new_n4117 = ~pq & new_n4116;
  assign new_n4118 = ~px & new_n4117;
  assign new_n4119 = ~pb & new_n2014;
  assign new_n4120 = ~pg0 & new_n4119;
  assign new_n4121 = ~po & new_n4120;
  assign new_n4122 = ~pc & new_n4121;
  assign new_n4123 = pi0 & new_n4122;
  assign new_n4124 = ~pd0 & new_n4123;
  assign new_n4125 = pl0 & new_n4124;
  assign new_n4126 = ~pc0 & new_n4125;
  assign new_n4127 = ~py & new_n4126;
  assign new_n4128 = ~pb0 & new_n4127;
  assign new_n4129 = ~pr & new_n4128;
  assign new_n4130 = ~px & new_n4129;
  assign new_n4131 = ~pi & new_n231;
  assign new_n4132 = ~pn & new_n4131;
  assign new_n4133 = ~pa & new_n4132;
  assign new_n4134 = ~pj0 & new_n4133;
  assign new_n4135 = ~pm & new_n4134;
  assign new_n4136 = ~pe0 & new_n4135;
  assign new_n4137 = ~ph0 & new_n4136;
  assign new_n4138 = pl0 & new_n4137;
  assign new_n4139 = ~pc0 & new_n4138;
  assign new_n4140 = ~pa0 & new_n4139;
  assign new_n4141 = ~pb0 & new_n4140;
  assign new_n4142 = ~px & new_n4141;
  assign new_n4143 = ~py & new_n4142;
  assign new_n4144 = ~pe0 & new_n3677;
  assign new_n4145 = pf0 & new_n4144;
  assign new_n4146 = ~pg0 & new_n4145;
  assign new_n4147 = ~pm & new_n4146;
  assign new_n4148 = pl0 & new_n4147;
  assign new_n4149 = ~pd0 & new_n4148;
  assign new_n4150 = ~ph0 & new_n4149;
  assign new_n4151 = ~pb0 & new_n4150;
  assign new_n4152 = ~pc0 & new_n4151;
  assign new_n4153 = ~pi & new_n582;
  assign new_n4154 = ~pq & new_n4153;
  assign new_n4155 = ~ph & new_n4154;
  assign new_n4156 = ~pe0 & new_n4155;
  assign new_n4157 = pi0 & new_n4156;
  assign new_n4158 = ~pm & new_n4157;
  assign new_n4159 = ~po & new_n4158;
  assign new_n4160 = ~pd0 & new_n4159;
  assign new_n4161 = pl0 & new_n4160;
  assign new_n4162 = ~pb0 & new_n4161;
  assign new_n4163 = ~pc0 & new_n4162;
  assign new_n4164 = ~pj0 & new_n3400;
  assign new_n4165 = ~po & new_n4164;
  assign new_n4166 = pl0 & new_n4165;
  assign new_n4167 = ~pc0 & new_n4166;
  assign new_n4168 = ~pd0 & new_n4167;
  assign new_n4169 = ~pa0 & new_n4168;
  assign new_n4170 = ~pb0 & new_n4169;
  assign new_n4171 = ~pn & new_n3550;
  assign new_n4172 = pz & new_n4171;
  assign new_n4173 = ~pi0 & new_n4172;
  assign new_n4174 = ph0 & new_n4173;
  assign new_n4175 = pj0 & new_n4174;
  assign new_n4176 = ~pb0 & new_n4175;
  assign new_n4177 = ~pc0 & new_n4176;
  assign new_n4178 = pj0 & new_n3772;
  assign new_n4179 = ~pi0 & new_n4178;
  assign new_n4180 = ~pb0 & new_n4179;
  assign new_n4181 = ~pc0 & new_n4180;
  assign new_n4182 = pi0 & new_n3514;
  assign new_n4183 = ~pd0 & new_n4182;
  assign new_n4184 = ~po & new_n4183;
  assign new_n4185 = ~pb0 & new_n4184;
  assign new_n4186 = ~pc0 & new_n4185;
  assign new_n4187 = ~pg0 & new_n3690;
  assign new_n4188 = ~po & new_n4187;
  assign new_n4189 = ~py & new_n4188;
  assign new_n4190 = ~pa0 & new_n4189;
  assign new_n4191 = ~pb0 & new_n4190;
  assign new_n4192 = ~pc0 & new_n4191;
  assign new_n4193 = ~pu & new_n4192;
  assign new_n4194 = ~px & new_n4193;
  assign new_n4195 = ~pt & new_n4194;
  assign new_n4196 = ~pq & new_n4195;
  assign new_n4197 = ~pr & new_n4196;
  assign new_n4198 = ~pj & new_n4197;
  assign new_n4199 = ~pl & new_n4198;
  assign new_n4200 = ~pa & new_n164;
  assign new_n4201 = ~pm & new_n4200;
  assign new_n4202 = pl0 & new_n4201;
  assign new_n4203 = ~pg0 & new_n4202;
  assign new_n4204 = ~pj0 & new_n4203;
  assign new_n4205 = ~po & new_n4204;
  assign new_n4206 = ~pc0 & new_n4205;
  assign new_n4207 = pd0 & new_n4206;
  assign new_n4208 = ~pb0 & new_n4207;
  assign new_n4209 = ~py & new_n4208;
  assign new_n4210 = ~pa0 & new_n4209;
  assign new_n4211 = ~pu & new_n4210;
  assign new_n4212 = ~px & new_n4211;
  assign new_n4213 = ~pb & new_n182;
  assign new_n4214 = pl0 & new_n4213;
  assign new_n4215 = ~pj0 & new_n4214;
  assign new_n4216 = ~po & new_n4215;
  assign new_n4217 = ~pc & new_n4216;
  assign new_n4218 = ~pc0 & new_n4217;
  assign new_n4219 = ~pd0 & new_n4218;
  assign new_n4220 = ~pb0 & new_n4219;
  assign new_n4221 = ~py & new_n4220;
  assign new_n4222 = ~pa0 & new_n4221;
  assign new_n4223 = ~pr & new_n4222;
  assign new_n4224 = ~px & new_n4223;
  assign new_n4225 = ~pj0 & new_n122;
  assign new_n4226 = ~po & new_n4225;
  assign new_n4227 = ~pc & new_n4226;
  assign new_n4228 = ~pm & new_n4227;
  assign new_n4229 = pl0 & new_n4228;
  assign new_n4230 = ~pg0 & new_n4229;
  assign new_n4231 = ~pd0 & new_n4230;
  assign new_n4232 = ~pb0 & new_n4231;
  assign new_n4233 = ~pc0 & new_n4232;
  assign new_n4234 = ~py & new_n4233;
  assign new_n4235 = ~pa0 & new_n4234;
  assign new_n4236 = ~pe0 & new_n3364;
  assign new_n4237 = pf0 & new_n4236;
  assign new_n4238 = pi0 & new_n4237;
  assign new_n4239 = ~pm & new_n4238;
  assign new_n4240 = ~pg0 & new_n4239;
  assign new_n4241 = ~ph0 & new_n4240;
  assign new_n4242 = pl0 & new_n4241;
  assign new_n4243 = ~pc0 & new_n4242;
  assign new_n4244 = ~pd0 & new_n4243;
  assign new_n4245 = ~pi & new_n3363;
  assign new_n4246 = ~pe0 & new_n4245;
  assign new_n4247 = pi0 & new_n4246;
  assign new_n4248 = ~pm & new_n4247;
  assign new_n4249 = ~po & new_n4248;
  assign new_n4250 = pl0 & new_n4249;
  assign new_n4251 = ~pj0 & new_n4250;
  assign new_n4252 = ~pc0 & new_n4251;
  assign new_n4253 = ~pd0 & new_n4252;
  assign new_n4254 = pu & new_n676;
  assign new_n4255 = ~px & new_n4254;
  assign new_n4256 = ~pq & new_n4255;
  assign new_n4257 = pz & new_n4256;
  assign new_n4258 = ~pm & new_n4257;
  assign new_n4259 = ~po & new_n4258;
  assign new_n4260 = ~pi0 & new_n4259;
  assign new_n4261 = ph0 & new_n4260;
  assign new_n4262 = pj0 & new_n4261;
  assign new_n4263 = pi0 & new_n4172;
  assign new_n4264 = ~pc0 & new_n4263;
  assign new_n4265 = ph0 & new_n4264;
  assign new_n4266 = ~py & new_n4265;
  assign new_n4267 = ~pb0 & new_n4266;
  assign new_n4268 = ph & new_n678;
  assign new_n4269 = pf0 & new_n4268;
  assign new_n4270 = ~pm & new_n4269;
  assign new_n4271 = ~po & new_n4270;
  assign new_n4272 = ~pi0 & new_n4271;
  assign new_n4273 = ~pd0 & new_n4272;
  assign new_n4274 = pj0 & new_n4273;
  assign new_n4275 = ~pi0 & new_n3878;
  assign new_n4276 = ~pc0 & new_n4275;
  assign new_n4277 = pj0 & new_n4276;
  assign new_n4278 = ~px & new_n4277;
  assign new_n4279 = ~pb0 & new_n4278;
  assign new_n4280 = ~pc & new_n105;
  assign new_n4281 = pi0 & new_n4280;
  assign new_n4282 = ~pk & new_n4281;
  assign new_n4283 = ~pd0 & new_n4282;
  assign new_n4284 = ~ph0 & new_n4283;
  assign new_n4285 = pl0 & new_n4284;
  assign new_n4286 = ~pj0 & new_n4285;
  assign new_n4287 = ~pb0 & new_n4286;
  assign new_n4288 = ~pc0 & new_n4287;
  assign new_n4289 = ~py & new_n4288;
  assign new_n4290 = ~pr & new_n4289;
  assign new_n4291 = ~px & new_n4290;
  assign new_n4292 = ~pn & new_n4291;
  assign new_n4293 = ~pq & new_n4292;
  assign new_n4294 = ~pm & new_n3081;
  assign new_n4295 = pd0 & new_n4294;
  assign new_n4296 = pl0 & new_n4295;
  assign new_n4297 = ~pj0 & new_n4296;
  assign new_n4298 = ~po & new_n4297;
  assign new_n4299 = ~pb0 & new_n4298;
  assign new_n4300 = ~pc0 & new_n4299;
  assign new_n4301 = ~pa0 & new_n4300;
  assign new_n4302 = ~px & new_n4301;
  assign new_n4303 = ~py & new_n4302;
  assign new_n4304 = ~pq & new_n4303;
  assign new_n4305 = ~pu & new_n4304;
  assign new_n4306 = ~pf & new_n219;
  assign new_n4307 = ~pg & new_n4306;
  assign new_n4308 = ~pe & new_n4307;
  assign new_n4309 = ~pb & new_n4308;
  assign new_n4310 = ~pg0 & new_n4309;
  assign new_n4311 = ~pj0 & new_n4310;
  assign new_n4312 = ~po & new_n4311;
  assign new_n4313 = ~pc & new_n4312;
  assign new_n4314 = ~pd0 & new_n4313;
  assign new_n4315 = pl0 & new_n4314;
  assign new_n4316 = ~pc0 & new_n4315;
  assign new_n4317 = ~pa0 & new_n4316;
  assign new_n4318 = ~pb0 & new_n4317;
  assign new_n4319 = ~px & new_n4318;
  assign new_n4320 = ~py & new_n4319;
  assign new_n4321 = ~pj0 & new_n182;
  assign new_n4322 = ~po & new_n4321;
  assign new_n4323 = ~pc & new_n4322;
  assign new_n4324 = ~pm & new_n4323;
  assign new_n4325 = ~pd0 & new_n4324;
  assign new_n4326 = pl0 & new_n4325;
  assign new_n4327 = ~pc0 & new_n4326;
  assign new_n4328 = ~pa0 & new_n4327;
  assign new_n4329 = ~pb0 & new_n4328;
  assign new_n4330 = ~px & new_n4329;
  assign new_n4331 = ~py & new_n4330;
  assign new_n4332 = ~pe0 & new_n679;
  assign new_n4333 = pf0 & new_n4332;
  assign new_n4334 = ~pi0 & new_n4333;
  assign new_n4335 = ~pm & new_n4334;
  assign new_n4336 = pj0 & new_n4335;
  assign new_n4337 = pl0 & new_n4336;
  assign new_n4338 = ~pg0 & new_n4337;
  assign new_n4339 = ~pd0 & new_n4338;
  assign new_n4340 = ~ph0 & new_n4339;
  assign new_n4341 = ~pi0 & new_n1368;
  assign new_n4342 = ~pm & new_n4341;
  assign new_n4343 = ~po & new_n4342;
  assign new_n4344 = pl0 & new_n4343;
  assign new_n4345 = pj0 & new_n4344;
  assign new_n4346 = ~pc0 & new_n4345;
  assign new_n4347 = ~pd0 & new_n4346;
  assign new_n4348 = pz & new_n679;
  assign new_n4349 = ~pm & new_n4348;
  assign new_n4350 = pj0 & new_n4349;
  assign new_n4351 = ~pi0 & new_n4350;
  assign new_n4352 = ~pd0 & new_n4351;
  assign new_n4353 = ph0 & new_n4352;
  assign new_n4354 = pi0 & new_n3786;
  assign new_n4355 = ~pd0 & new_n4354;
  assign new_n4356 = ph0 & new_n4355;
  assign new_n4357 = ~pb0 & new_n4356;
  assign new_n4358 = ~pc0 & new_n4357;
  assign new_n4359 = ph & new_n3648;
  assign new_n4360 = pf0 & new_n4359;
  assign new_n4361 = ~pm & new_n4360;
  assign new_n4362 = ~po & new_n4361;
  assign new_n4363 = ~pi0 & new_n4362;
  assign new_n4364 = ~pc0 & new_n4363;
  assign new_n4365 = pj0 & new_n4364;
  assign new_n4366 = ~pi0 & new_n1010;
  assign new_n4367 = ~pd0 & new_n4366;
  assign new_n4368 = pj0 & new_n4367;
  assign new_n4369 = ~pb0 & new_n4368;
  assign new_n4370 = ~pc0 & new_n4369;
  assign new_n4371 = ~ph0 & new_n3081;
  assign new_n4372 = pl0 & new_n4371;
  assign new_n4373 = ~pj0 & new_n4372;
  assign new_n4374 = ~pk & new_n4373;
  assign new_n4375 = ~pa0 & new_n4374;
  assign new_n4376 = ~pb0 & new_n4375;
  assign new_n4377 = ~pc0 & new_n4376;
  assign new_n4378 = pd0 & new_n4377;
  assign new_n4379 = ~px & new_n4378;
  assign new_n4380 = ~py & new_n4379;
  assign new_n4381 = ~pu & new_n4380;
  assign new_n4382 = ~pq & new_n4381;
  assign new_n4383 = ~pr & new_n4382;
  assign new_n4384 = ~pj & new_n4383;
  assign new_n4385 = ~pn & new_n4384;
  assign new_n4386 = ~ps & new_n1333;
  assign new_n4387 = ~pg0 & new_n4386;
  assign new_n4388 = ~pc & new_n4387;
  assign new_n4389 = pi0 & new_n4388;
  assign new_n4390 = ~pd0 & new_n4389;
  assign new_n4391 = ~ph0 & new_n4390;
  assign new_n4392 = pl0 & new_n4391;
  assign new_n4393 = pd & new_n4392;
  assign new_n4394 = ~pb0 & new_n4393;
  assign new_n4395 = ~pc0 & new_n4394;
  assign new_n4396 = ~py & new_n4395;
  assign new_n4397 = ~pr & new_n4396;
  assign new_n4398 = ~px & new_n4397;
  assign new_n4399 = ~pn & new_n4398;
  assign new_n4400 = ~pq & new_n4399;
  assign new_n4401 = pd0 & new_n3081;
  assign new_n4402 = pl0 & new_n4401;
  assign new_n4403 = ~pj0 & new_n4402;
  assign new_n4404 = ~po & new_n4403;
  assign new_n4405 = ~py & new_n4404;
  assign new_n4406 = ~pa0 & new_n4405;
  assign new_n4407 = ~pb0 & new_n4406;
  assign new_n4408 = ~pc0 & new_n4407;
  assign new_n4409 = ~pu & new_n4408;
  assign new_n4410 = ~px & new_n4409;
  assign new_n4411 = ~pt & new_n4410;
  assign new_n4412 = ~pq & new_n4411;
  assign new_n4413 = ~pr & new_n4412;
  assign new_n4414 = ~pj & new_n4413;
  assign new_n4415 = ~pl & new_n4414;
  assign new_n4416 = ~pc & new_n1834;
  assign new_n4417 = pi0 & new_n4416;
  assign new_n4418 = ~pk & new_n4417;
  assign new_n4419 = ~ph0 & new_n4418;
  assign new_n4420 = pl0 & new_n4419;
  assign new_n4421 = ~pg0 & new_n4420;
  assign new_n4422 = ~pj0 & new_n4421;
  assign new_n4423 = ~pc0 & new_n4422;
  assign new_n4424 = ~pd0 & new_n4423;
  assign new_n4425 = ~pb0 & new_n4424;
  assign new_n4426 = ~px & new_n4425;
  assign new_n4427 = ~py & new_n4426;
  assign new_n4428 = ~pq & new_n4427;
  assign new_n4429 = ~pr & new_n4428;
  assign new_n4430 = ~po & new_n4200;
  assign new_n4431 = ~pb & new_n4430;
  assign new_n4432 = pd0 & new_n4431;
  assign new_n4433 = pl0 & new_n4432;
  assign new_n4434 = ~pg0 & new_n4433;
  assign new_n4435 = ~pj0 & new_n4434;
  assign new_n4436 = ~pb0 & new_n4435;
  assign new_n4437 = ~pc0 & new_n4436;
  assign new_n4438 = ~pa0 & new_n4437;
  assign new_n4439 = ~px & new_n4438;
  assign new_n4440 = ~py & new_n4439;
  assign new_n4441 = ~pr & new_n4440;
  assign new_n4442 = ~pu & new_n4441;
  assign new_n4443 = ~pk & new_n4280;
  assign new_n4444 = ~pd0 & new_n4443;
  assign new_n4445 = pl0 & new_n4444;
  assign new_n4446 = ~pj0 & new_n4445;
  assign new_n4447 = ~po & new_n4446;
  assign new_n4448 = ~pb0 & new_n4447;
  assign new_n4449 = ~pc0 & new_n4448;
  assign new_n4450 = ~pa0 & new_n4449;
  assign new_n4451 = ~px & new_n4450;
  assign new_n4452 = ~py & new_n4451;
  assign new_n4453 = ~pq & new_n4452;
  assign new_n4454 = ~pr & new_n4453;
  assign new_n4455 = ~pg0 & new_n442;
  assign new_n4456 = ~pj0 & new_n4455;
  assign new_n4457 = ~pc & new_n4456;
  assign new_n4458 = pi0 & new_n4457;
  assign new_n4459 = ~ph0 & new_n4458;
  assign new_n4460 = pl0 & new_n4459;
  assign new_n4461 = ~pd0 & new_n4460;
  assign new_n4462 = ~pb0 & new_n4461;
  assign new_n4463 = ~pc0 & new_n4462;
  assign new_n4464 = ~px & new_n4463;
  assign new_n4465 = ~py & new_n4464;
  assign new_n4466 = pj0 & new_n4027;
  assign new_n4467 = ~po & new_n4466;
  assign new_n4468 = ~pc & new_n4467;
  assign new_n4469 = ~pi0 & new_n4468;
  assign new_n4470 = ~pd0 & new_n4469;
  assign new_n4471 = pl0 & new_n4470;
  assign new_n4472 = ~pc0 & new_n4471;
  assign new_n4473 = ~px & new_n4472;
  assign new_n4474 = ~pb0 & new_n4473;
  assign new_n4475 = ~pq & new_n4474;
  assign new_n4476 = ~pr & new_n4475;
  assign new_n4477 = ~po & new_n2014;
  assign new_n4478 = ~pc & new_n4477;
  assign new_n4479 = pi0 & new_n4478;
  assign new_n4480 = ~pm & new_n4479;
  assign new_n4481 = pl0 & new_n4480;
  assign new_n4482 = ~pg0 & new_n4481;
  assign new_n4483 = ~pd0 & new_n4482;
  assign new_n4484 = ~pb0 & new_n4483;
  assign new_n4485 = ~pc0 & new_n4484;
  assign new_n4486 = ~px & new_n4485;
  assign new_n4487 = ~py & new_n4486;
  assign new_n4488 = ~pa & new_n2027;
  assign new_n4489 = ~ph0 & new_n4488;
  assign new_n4490 = pl0 & new_n4489;
  assign new_n4491 = ~pe0 & new_n4490;
  assign new_n4492 = ~pb0 & new_n4491;
  assign new_n4493 = ~pc0 & new_n4492;
  assign new_n4494 = ~pa0 & new_n4493;
  assign new_n4495 = ~px & new_n4494;
  assign new_n4496 = ~py & new_n4495;
  assign new_n4497 = ~pr & new_n4496;
  assign new_n4498 = ~pu & new_n4497;
  assign new_n4499 = ~pg0 & new_n3021;
  assign new_n4500 = ~pk & new_n4499;
  assign new_n4501 = ~pa0 & new_n4500;
  assign new_n4502 = ~pb0 & new_n4501;
  assign new_n4503 = ~pc0 & new_n4502;
  assign new_n4504 = pd0 & new_n4503;
  assign new_n4505 = ~px & new_n4504;
  assign new_n4506 = ~py & new_n4505;
  assign new_n4507 = ~pu & new_n4506;
  assign new_n4508 = ~pq & new_n4507;
  assign new_n4509 = ~pr & new_n4508;
  assign new_n4510 = ~pj & new_n4509;
  assign new_n4511 = ~pn & new_n4510;
  assign new_n4512 = pl0 & new_n105;
  assign new_n4513 = ~pj0 & new_n4512;
  assign new_n4514 = ~pc & new_n4513;
  assign new_n4515 = pi0 & new_n4514;
  assign new_n4516 = ~pb0 & new_n4515;
  assign new_n4517 = ~pc0 & new_n4516;
  assign new_n4518 = ~pd0 & new_n4517;
  assign new_n4519 = ~ph0 & new_n4518;
  assign new_n4520 = ~px & new_n4519;
  assign new_n4521 = ~py & new_n4520;
  assign new_n4522 = ~pt & new_n4521;
  assign new_n4523 = ~pq & new_n4522;
  assign new_n4524 = ~pr & new_n4523;
  assign new_n4525 = ~pl & new_n4524;
  assign new_n4526 = ~pn & new_n4525;
  assign new_n4527 = pd & new_n2867;
  assign new_n4528 = ~ps & new_n4527;
  assign new_n4529 = ~pg0 & new_n4528;
  assign new_n4530 = ~po & new_n4529;
  assign new_n4531 = ~pb0 & new_n4530;
  assign new_n4532 = ~pc0 & new_n4531;
  assign new_n4533 = pd0 & new_n4532;
  assign new_n4534 = pl0 & new_n4533;
  assign new_n4535 = ~py & new_n4534;
  assign new_n4536 = ~pa0 & new_n4535;
  assign new_n4537 = ~px & new_n4536;
  assign new_n4538 = ~pr & new_n4537;
  assign new_n4539 = ~pu & new_n4538;
  assign new_n4540 = ~pj & new_n4539;
  assign new_n4541 = ~pq & new_n4540;
  assign new_n4542 = ~pi0 & new_n2883;
  assign new_n4543 = ~pk & new_n4542;
  assign new_n4544 = ~pd0 & new_n4543;
  assign new_n4545 = ~ph0 & new_n4544;
  assign new_n4546 = pl0 & new_n4545;
  assign new_n4547 = pj0 & new_n4546;
  assign new_n4548 = ~pb0 & new_n4547;
  assign new_n4549 = ~pc0 & new_n4548;
  assign new_n4550 = ~px & new_n4549;
  assign new_n4551 = ~pq & new_n4550;
  assign new_n4552 = ~pr & new_n4551;
  assign new_n4553 = ~pj & new_n4552;
  assign new_n4554 = ~pn & new_n4553;
  assign new_n4555 = ~po & new_n3081;
  assign new_n4556 = ~pb & new_n4555;
  assign new_n4557 = ~pc0 & new_n4556;
  assign new_n4558 = pd0 & new_n4557;
  assign new_n4559 = pl0 & new_n4558;
  assign new_n4560 = ~pj0 & new_n4559;
  assign new_n4561 = ~pa0 & new_n4560;
  assign new_n4562 = ~pb0 & new_n4561;
  assign new_n4563 = ~py & new_n4562;
  assign new_n4564 = ~pu & new_n4563;
  assign new_n4565 = ~px & new_n4564;
  assign new_n4566 = ~pq & new_n4565;
  assign new_n4567 = ~pr & new_n4566;
  assign new_n4568 = ~pc & new_n2900;
  assign new_n4569 = ~pk & new_n4568;
  assign new_n4570 = pl0 & new_n4569;
  assign new_n4571 = ~pg0 & new_n4570;
  assign new_n4572 = ~pj0 & new_n4571;
  assign new_n4573 = ~po & new_n4572;
  assign new_n4574 = ~pc0 & new_n4573;
  assign new_n4575 = ~pd0 & new_n4574;
  assign new_n4576 = ~pb0 & new_n4575;
  assign new_n4577 = ~py & new_n4576;
  assign new_n4578 = ~pa0 & new_n4577;
  assign new_n4579 = ~pr & new_n4578;
  assign new_n4580 = ~px & new_n4579;
  assign new_n4581 = pl0 & new_n479;
  assign new_n4582 = ~pj0 & new_n4581;
  assign new_n4583 = ~pc & new_n4582;
  assign new_n4584 = pi0 & new_n4583;
  assign new_n4585 = ~pd0 & new_n4584;
  assign new_n4586 = ~ph0 & new_n4585;
  assign new_n4587 = ~pc0 & new_n4586;
  assign new_n4588 = ~py & new_n4587;
  assign new_n4589 = ~pb0 & new_n4588;
  assign new_n4590 = ~pq & new_n4589;
  assign new_n4591 = ~px & new_n4590;
  assign new_n4592 = pj0 & new_n4119;
  assign new_n4593 = ~po & new_n4592;
  assign new_n4594 = ~pc & new_n4593;
  assign new_n4595 = ~pi0 & new_n4594;
  assign new_n4596 = pl0 & new_n4595;
  assign new_n4597 = ~pg0 & new_n4596;
  assign new_n4598 = ~pd0 & new_n4597;
  assign new_n4599 = ~pb0 & new_n4598;
  assign new_n4600 = ~pc0 & new_n4599;
  assign new_n4601 = ~pr & new_n4600;
  assign new_n4602 = ~px & new_n4601;
  assign new_n4603 = ~pm & new_n3191;
  assign new_n4604 = ~pd0 & new_n4603;
  assign new_n4605 = pl0 & new_n4604;
  assign new_n4606 = ~pc0 & new_n4605;
  assign new_n4607 = ~py & new_n4606;
  assign new_n4608 = ~pb0 & new_n4607;
  assign new_n4609 = ~pq & new_n4608;
  assign new_n4610 = ~px & new_n4609;
  assign new_n4611 = ~pa & new_n1894;
  assign new_n4612 = pl0 & new_n4611;
  assign new_n4613 = ~pg0 & new_n4612;
  assign new_n4614 = ~pe0 & new_n4613;
  assign new_n4615 = ~pc0 & new_n4614;
  assign new_n4616 = ~ph0 & new_n4615;
  assign new_n4617 = ~pb0 & new_n4616;
  assign new_n4618 = ~py & new_n4617;
  assign new_n4619 = ~pa0 & new_n4618;
  assign new_n4620 = ~pu & new_n4619;
  assign new_n4621 = ~px & new_n4620;
  assign new_n4622 = ~ph0 & new_n3689;
  assign new_n4623 = pl0 & new_n4622;
  assign new_n4624 = ~pk & new_n4623;
  assign new_n4625 = ~py & new_n4624;
  assign new_n4626 = ~pa0 & new_n4625;
  assign new_n4627 = ~pb0 & new_n4626;
  assign new_n4628 = ~pc0 & new_n4627;
  assign new_n4629 = ~pu & new_n4628;
  assign new_n4630 = ~px & new_n4629;
  assign new_n4631 = ~pr & new_n4630;
  assign new_n4632 = ~pn & new_n4631;
  assign new_n4633 = ~pq & new_n4632;
  assign new_n4634 = ~pi & new_n4633;
  assign new_n4635 = ~pj & new_n4634;
  assign new_n4636 = pd & new_n1058;
  assign new_n4637 = ~ps & new_n4636;
  assign new_n4638 = ~pc & new_n4637;
  assign new_n4639 = pi0 & new_n4638;
  assign new_n4640 = ~pc0 & new_n4639;
  assign new_n4641 = ~pd0 & new_n4640;
  assign new_n4642 = ~ph0 & new_n4641;
  assign new_n4643 = pl0 & new_n4642;
  assign new_n4644 = ~py & new_n4643;
  assign new_n4645 = ~pb0 & new_n4644;
  assign new_n4646 = ~px & new_n4645;
  assign new_n4647 = ~pq & new_n4646;
  assign new_n4648 = ~pr & new_n4647;
  assign new_n4649 = ~pj & new_n4648;
  assign new_n4650 = ~pn & new_n4649;
  assign new_n4651 = pl0 & new_n3036;
  assign new_n4652 = ~pg0 & new_n4651;
  assign new_n4653 = ~pj0 & new_n4652;
  assign new_n4654 = ~po & new_n4653;
  assign new_n4655 = ~pa0 & new_n4654;
  assign new_n4656 = ~pb0 & new_n4655;
  assign new_n4657 = ~pc0 & new_n4656;
  assign new_n4658 = pd0 & new_n4657;
  assign new_n4659 = ~px & new_n4658;
  assign new_n4660 = ~py & new_n4659;
  assign new_n4661 = ~pu & new_n4660;
  assign new_n4662 = ~pr & new_n4661;
  assign new_n4663 = ~pt & new_n4662;
  assign new_n4664 = ~pl & new_n4663;
  assign new_n4665 = ~pq & new_n4664;
  assign new_n4666 = ~pi0 & new_n3938;
  assign new_n4667 = ~pk & new_n4666;
  assign new_n4668 = ~ph0 & new_n4667;
  assign new_n4669 = pl0 & new_n4668;
  assign new_n4670 = ~pg0 & new_n4669;
  assign new_n4671 = pj0 & new_n4670;
  assign new_n4672 = ~pc0 & new_n4671;
  assign new_n4673 = ~pd0 & new_n4672;
  assign new_n4674 = ~pb0 & new_n4673;
  assign new_n4675 = ~pr & new_n4674;
  assign new_n4676 = ~px & new_n4675;
  assign new_n4677 = ~pn & new_n4676;
  assign new_n4678 = ~pq & new_n4677;
  assign new_n4679 = ~pj0 & new_n2900;
  assign new_n4680 = ~po & new_n4679;
  assign new_n4681 = ~pc & new_n4680;
  assign new_n4682 = pl0 & new_n4681;
  assign new_n4683 = pd & new_n4682;
  assign new_n4684 = ~ps & new_n4683;
  assign new_n4685 = ~pg0 & new_n4684;
  assign new_n4686 = ~pc0 & new_n4685;
  assign new_n4687 = ~pd0 & new_n4686;
  assign new_n4688 = ~pb0 & new_n4687;
  assign new_n4689 = ~py & new_n4688;
  assign new_n4690 = ~pa0 & new_n4689;
  assign new_n4691 = ~pr & new_n4690;
  assign new_n4692 = ~px & new_n4691;
  assign new_n4693 = ~pm & new_n2868;
  assign new_n4694 = ~pb0 & new_n4693;
  assign new_n4695 = ~pc0 & new_n4694;
  assign new_n4696 = pd0 & new_n4695;
  assign new_n4697 = ~ph0 & new_n4696;
  assign new_n4698 = ~py & new_n4697;
  assign new_n4699 = ~pa0 & new_n4698;
  assign new_n4700 = ~px & new_n4699;
  assign new_n4701 = ~pq & new_n4700;
  assign new_n4702 = ~pu & new_n4701;
  assign new_n4703 = ~pi & new_n4702;
  assign new_n4704 = ~pn & new_n4703;
  assign new_n4705 = ~pm & new_n1181;
  assign new_n4706 = pl0 & new_n4705;
  assign new_n4707 = ~pg0 & new_n4706;
  assign new_n4708 = ~pc & new_n4707;
  assign new_n4709 = pi0 & new_n4708;
  assign new_n4710 = ~pd0 & new_n4709;
  assign new_n4711 = ~ph0 & new_n4710;
  assign new_n4712 = ~pc0 & new_n4711;
  assign new_n4713 = ~py & new_n4712;
  assign new_n4714 = ~pb0 & new_n4713;
  assign new_n4715 = ~pq & new_n4714;
  assign new_n4716 = ~px & new_n4715;
  assign new_n4717 = ~pj0 & new_n4213;
  assign new_n4718 = ~po & new_n4717;
  assign new_n4719 = ~pc & new_n4718;
  assign new_n4720 = pi0 & new_n4719;
  assign new_n4721 = ~pd0 & new_n4720;
  assign new_n4722 = pl0 & new_n4721;
  assign new_n4723 = ~pc0 & new_n4722;
  assign new_n4724 = ~py & new_n4723;
  assign new_n4725 = ~pb0 & new_n4724;
  assign new_n4726 = ~pr & new_n4725;
  assign new_n4727 = ~px & new_n4726;
  assign new_n4728 = ~po & new_n122;
  assign new_n4729 = ~pc & new_n4728;
  assign new_n4730 = pi0 & new_n4729;
  assign new_n4731 = ~pm & new_n4730;
  assign new_n4732 = ~pg0 & new_n4731;
  assign new_n4733 = ~pj0 & new_n4732;
  assign new_n4734 = pl0 & new_n4733;
  assign new_n4735 = ~pc0 & new_n4734;
  assign new_n4736 = ~pd0 & new_n4735;
  assign new_n4737 = ~py & new_n4736;
  assign new_n4738 = ~pb0 & new_n4737;
  assign new_n4739 = ~pa & new_n221;
  assign new_n4740 = pl0 & new_n4739;
  assign new_n4741 = ~pj0 & new_n4740;
  assign new_n4742 = ~pe0 & new_n4741;
  assign new_n4743 = ~pc0 & new_n4742;
  assign new_n4744 = ~ph0 & new_n4743;
  assign new_n4745 = ~pb0 & new_n4744;
  assign new_n4746 = ~py & new_n4745;
  assign new_n4747 = ~pa0 & new_n4746;
  assign new_n4748 = ~pu & new_n4747;
  assign new_n4749 = ~px & new_n4748;
  assign new_n4750 = ~ph0 & new_n4004;
  assign new_n4751 = pl0 & new_n4750;
  assign new_n4752 = pd & new_n4751;
  assign new_n4753 = ~ps & new_n4752;
  assign new_n4754 = ~pc0 & new_n4753;
  assign new_n4755 = ~pd0 & new_n4754;
  assign new_n4756 = ~pb0 & new_n4755;
  assign new_n4757 = ~pr & new_n4756;
  assign new_n4758 = ~px & new_n4757;
  assign new_n4759 = ~pn & new_n4758;
  assign new_n4760 = ~pq & new_n4759;
  assign new_n4761 = pl0 & new_n1333;
  assign new_n4762 = ~pg0 & new_n4761;
  assign new_n4763 = ~pc & new_n4762;
  assign new_n4764 = pi0 & new_n4763;
  assign new_n4765 = ~pb0 & new_n4764;
  assign new_n4766 = ~pc0 & new_n4765;
  assign new_n4767 = ~pd0 & new_n4766;
  assign new_n4768 = ~ph0 & new_n4767;
  assign new_n4769 = ~px & new_n4768;
  assign new_n4770 = ~py & new_n4769;
  assign new_n4771 = ~pt & new_n4770;
  assign new_n4772 = ~pq & new_n4771;
  assign new_n4773 = ~pr & new_n4772;
  assign new_n4774 = ~pl & new_n4773;
  assign new_n4775 = ~pn & new_n4774;
  assign new_n4776 = pd & new_n3081;
  assign new_n4777 = ~ps & new_n4776;
  assign new_n4778 = ~pj0 & new_n4777;
  assign new_n4779 = ~po & new_n4778;
  assign new_n4780 = ~pb0 & new_n4779;
  assign new_n4781 = ~pc0 & new_n4780;
  assign new_n4782 = pd0 & new_n4781;
  assign new_n4783 = pl0 & new_n4782;
  assign new_n4784 = ~py & new_n4783;
  assign new_n4785 = ~pa0 & new_n4784;
  assign new_n4786 = ~px & new_n4785;
  assign new_n4787 = ~pr & new_n4786;
  assign new_n4788 = ~pu & new_n4787;
  assign new_n4789 = ~pj & new_n4788;
  assign new_n4790 = ~pq & new_n4789;
  assign new_n4791 = ~pb & new_n3021;
  assign new_n4792 = ~pa0 & new_n4791;
  assign new_n4793 = ~pb0 & new_n4792;
  assign new_n4794 = ~pc0 & new_n4793;
  assign new_n4795 = pd0 & new_n4794;
  assign new_n4796 = ~px & new_n4795;
  assign new_n4797 = ~py & new_n4796;
  assign new_n4798 = ~pu & new_n4797;
  assign new_n4799 = ~pq & new_n4798;
  assign new_n4800 = ~pr & new_n4799;
  assign new_n4801 = ~pi & new_n4800;
  assign new_n4802 = ~pn & new_n4801;
  assign new_n4803 = ~pj0 & new_n1679;
  assign new_n4804 = ~po & new_n4803;
  assign new_n4805 = ~pc & new_n4804;
  assign new_n4806 = ~pc0 & new_n4805;
  assign new_n4807 = ~pd0 & new_n4806;
  assign new_n4808 = pl0 & new_n4807;
  assign new_n4809 = ~pg0 & new_n4808;
  assign new_n4810 = ~pa0 & new_n4809;
  assign new_n4811 = ~pb0 & new_n4810;
  assign new_n4812 = ~py & new_n4811;
  assign new_n4813 = ~pt & new_n4812;
  assign new_n4814 = ~px & new_n4813;
  assign new_n4815 = ~pq & new_n4814;
  assign new_n4816 = ~pr & new_n4815;
  assign new_n4817 = ~pm & new_n3132;
  assign new_n4818 = ~pc0 & new_n4817;
  assign new_n4819 = pd0 & new_n4818;
  assign new_n4820 = ~ph0 & new_n4819;
  assign new_n4821 = pl0 & new_n4820;
  assign new_n4822 = ~pa0 & new_n4821;
  assign new_n4823 = ~pb0 & new_n4822;
  assign new_n4824 = ~py & new_n4823;
  assign new_n4825 = ~pu & new_n4824;
  assign new_n4826 = ~px & new_n4825;
  assign new_n4827 = ~pn & new_n4826;
  assign new_n4828 = ~pq & new_n4827;
  assign new_n4829 = ~pm & new_n1058;
  assign new_n4830 = ~ph0 & new_n4829;
  assign new_n4831 = pl0 & new_n4830;
  assign new_n4832 = ~pc & new_n4831;
  assign new_n4833 = pi0 & new_n4832;
  assign new_n4834 = ~pc0 & new_n4833;
  assign new_n4835 = ~pd0 & new_n4834;
  assign new_n4836 = ~pb0 & new_n4835;
  assign new_n4837 = ~px & new_n4836;
  assign new_n4838 = ~py & new_n4837;
  assign new_n4839 = ~pn & new_n4838;
  assign new_n4840 = ~pq & new_n4839;
  assign new_n4841 = ~pj0 & new_n4309;
  assign new_n4842 = ~po & new_n4841;
  assign new_n4843 = ~pc & new_n4842;
  assign new_n4844 = pi0 & new_n4843;
  assign new_n4845 = pl0 & new_n4844;
  assign new_n4846 = ~pg0 & new_n4845;
  assign new_n4847 = ~pd0 & new_n4846;
  assign new_n4848 = ~pb0 & new_n4847;
  assign new_n4849 = ~pc0 & new_n4848;
  assign new_n4850 = ~px & new_n4849;
  assign new_n4851 = ~py & new_n4850;
  assign new_n4852 = ~po & new_n182;
  assign new_n4853 = ~pc & new_n4852;
  assign new_n4854 = pi0 & new_n4853;
  assign new_n4855 = ~pm & new_n4854;
  assign new_n4856 = pl0 & new_n4855;
  assign new_n4857 = ~pj0 & new_n4856;
  assign new_n4858 = ~pd0 & new_n4857;
  assign new_n4859 = ~pb0 & new_n4858;
  assign new_n4860 = ~pc0 & new_n4859;
  assign new_n4861 = ~px & new_n4860;
  assign new_n4862 = ~py & new_n4861;
  assign new_n4863 = ~pn & new_n3210;
  assign new_n4864 = ~pq & new_n4863;
  assign new_n4865 = ~pa & new_n4864;
  assign new_n4866 = ~pg0 & new_n4865;
  assign new_n4867 = ~pj0 & new_n4866;
  assign new_n4868 = ~pe0 & new_n4867;
  assign new_n4869 = ~ph0 & new_n4868;
  assign new_n4870 = pl0 & new_n4869;
  assign new_n4871 = ~pc0 & new_n4870;
  assign new_n4872 = ~pa0 & new_n4871;
  assign new_n4873 = ~pb0 & new_n4872;
  assign new_n4874 = ~px & new_n4873;
  assign new_n4875 = ~py & new_n4874;
  assign new_n4876 = pd & new_n4372;
  assign new_n4877 = ~ps & new_n4876;
  assign new_n4878 = ~pa0 & new_n4877;
  assign new_n4879 = ~pb0 & new_n4878;
  assign new_n4880 = ~pc0 & new_n4879;
  assign new_n4881 = pd0 & new_n4880;
  assign new_n4882 = ~px & new_n4881;
  assign new_n4883 = ~pj0 & new_n4882;
  assign new_n4884 = ~py & new_n4883;
  assign new_n4885 = ~pu & new_n4884;
  assign new_n4886 = ~pq & new_n4885;
  assign new_n4887 = ~pr & new_n4886;
  assign new_n4888 = ~pj & new_n4887;
  assign new_n4889 = ~pn & new_n4888;
  assign new_n4890 = ~pc0 & new_n2867;
  assign new_n4891 = pd0 & new_n4890;
  assign new_n4892 = ~ph0 & new_n4891;
  assign new_n4893 = pl0 & new_n4892;
  assign new_n4894 = ~px & new_n4893;
  assign new_n4895 = ~py & new_n4894;
  assign new_n4896 = ~pa0 & new_n4895;
  assign new_n4897 = ~pb0 & new_n4896;
  assign new_n4898 = ~pt & new_n4897;
  assign new_n4899 = ~pg0 & new_n4898;
  assign new_n4900 = ~pu & new_n4899;
  assign new_n4901 = ~pr & new_n4900;
  assign new_n4902 = ~pn & new_n4901;
  assign new_n4903 = ~pq & new_n4902;
  assign new_n4904 = ~pj & new_n4903;
  assign new_n4905 = ~pl & new_n4904;
  assign new_n4906 = ~pg0 & new_n1834;
  assign new_n4907 = ~pj0 & new_n4906;
  assign new_n4908 = ~pc & new_n4907;
  assign new_n4909 = pi0 & new_n4908;
  assign new_n4910 = ~ph0 & new_n4909;
  assign new_n4911 = pl0 & new_n4910;
  assign new_n4912 = pd & new_n4911;
  assign new_n4913 = ~ps & new_n4912;
  assign new_n4914 = ~pc0 & new_n4913;
  assign new_n4915 = ~pd0 & new_n4914;
  assign new_n4916 = ~pb0 & new_n4915;
  assign new_n4917 = ~px & new_n4916;
  assign new_n4918 = ~py & new_n4917;
  assign new_n4919 = ~pq & new_n4918;
  assign new_n4920 = ~pr & new_n4919;
  assign new_n4921 = ~ph0 & new_n105;
  assign new_n4922 = pl0 & new_n4921;
  assign new_n4923 = ~pj0 & new_n4922;
  assign new_n4924 = ~pc & new_n4923;
  assign new_n4925 = ~pa0 & new_n4924;
  assign new_n4926 = ~pb0 & new_n4925;
  assign new_n4927 = ~pc0 & new_n4926;
  assign new_n4928 = ~pd0 & new_n4927;
  assign new_n4929 = ~px & new_n4928;
  assign new_n4930 = ~py & new_n4929;
  assign new_n4931 = ~pt & new_n4930;
  assign new_n4932 = ~pq & new_n4931;
  assign new_n4933 = ~pr & new_n4932;
  assign new_n4934 = ~pl & new_n4933;
  assign new_n4935 = ~pn & new_n4934;
  assign new_n4936 = ~pb & new_n3587;
  assign new_n4937 = ~pb0 & new_n4936;
  assign new_n4938 = ~pc0 & new_n4937;
  assign new_n4939 = pd0 & new_n4938;
  assign new_n4940 = ~ph0 & new_n4939;
  assign new_n4941 = ~py & new_n4940;
  assign new_n4942 = ~pa0 & new_n4941;
  assign new_n4943 = ~px & new_n4942;
  assign new_n4944 = ~pr & new_n4943;
  assign new_n4945 = ~pu & new_n4944;
  assign new_n4946 = ~pn & new_n4945;
  assign new_n4947 = ~pq & new_n4946;
  assign new_n4948 = ~po & new_n2973;
  assign new_n4949 = ~pc & new_n4948;
  assign new_n4950 = ~pd0 & new_n4949;
  assign new_n4951 = pl0 & new_n4950;
  assign new_n4952 = pd & new_n4951;
  assign new_n4953 = ~ps & new_n4952;
  assign new_n4954 = ~pb0 & new_n4953;
  assign new_n4955 = ~pc0 & new_n4954;
  assign new_n4956 = ~pa0 & new_n4955;
  assign new_n4957 = ~px & new_n4956;
  assign new_n4958 = ~py & new_n4957;
  assign new_n4959 = ~pq & new_n4958;
  assign new_n4960 = ~pr & new_n4959;
  assign new_n4961 = ~pi0 & new_n1058;
  assign new_n4962 = ~pb & new_n4961;
  assign new_n4963 = ~ph0 & new_n4962;
  assign new_n4964 = pl0 & new_n4963;
  assign new_n4965 = pj0 & new_n4964;
  assign new_n4966 = ~pc & new_n4965;
  assign new_n4967 = ~pc0 & new_n4966;
  assign new_n4968 = ~pd0 & new_n4967;
  assign new_n4969 = ~pb0 & new_n4968;
  assign new_n4970 = ~pr & new_n4969;
  assign new_n4971 = ~px & new_n4970;
  assign new_n4972 = ~pn & new_n4971;
  assign new_n4973 = ~pq & new_n4972;
  assign new_n4974 = ~pi0 & new_n1333;
  assign new_n4975 = ~pk & new_n4974;
  assign new_n4976 = ~pg0 & new_n4975;
  assign new_n4977 = pj0 & new_n4976;
  assign new_n4978 = ~po & new_n4977;
  assign new_n4979 = ~pc & new_n4978;
  assign new_n4980 = ~pd0 & new_n4979;
  assign new_n4981 = pl0 & new_n4980;
  assign new_n4982 = ~pc0 & new_n4981;
  assign new_n4983 = ~px & new_n4982;
  assign new_n4984 = ~pb0 & new_n4983;
  assign new_n4985 = ~pq & new_n4984;
  assign new_n4986 = ~pr & new_n4985;
  assign new_n4987 = ~pd0 & new_n4281;
  assign new_n4988 = pl0 & new_n4987;
  assign new_n4989 = ~pj0 & new_n4988;
  assign new_n4990 = ~po & new_n4989;
  assign new_n4991 = ~pb0 & new_n4990;
  assign new_n4992 = ~pc0 & new_n4991;
  assign new_n4993 = ~py & new_n4992;
  assign new_n4994 = ~pr & new_n4993;
  assign new_n4995 = ~px & new_n4994;
  assign new_n4996 = pn & new_n4995;
  assign new_n4997 = ~pq & new_n4996;
  assign new_n4998 = ~pi0 & new_n4478;
  assign new_n4999 = ~pm & new_n4998;
  assign new_n5000 = ~pg0 & new_n4999;
  assign new_n5001 = pj0 & new_n5000;
  assign new_n5002 = pl0 & new_n5001;
  assign new_n5003 = ~pc0 & new_n5002;
  assign new_n5004 = ~pd0 & new_n5003;
  assign new_n5005 = ~px & new_n5004;
  assign new_n5006 = ~pb0 & new_n5005;
  assign new_n5007 = pl0 & new_n4488;
  assign new_n5008 = ~pm & new_n5007;
  assign new_n5009 = ~pe0 & new_n5008;
  assign new_n5010 = ~pc0 & new_n5009;
  assign new_n5011 = ~ph0 & new_n5010;
  assign new_n5012 = ~pb0 & new_n5011;
  assign new_n5013 = ~py & new_n5012;
  assign new_n5014 = ~pa0 & new_n5013;
  assign new_n5015 = ~pu & new_n5014;
  assign new_n5016 = ~px & new_n5015;
  assign new_n5017 = pd0 & new_n3036;
  assign new_n5018 = ~ph0 & new_n5017;
  assign new_n5019 = pl0 & new_n5018;
  assign new_n5020 = ~pg0 & new_n5019;
  assign new_n5021 = ~py & new_n5020;
  assign new_n5022 = ~pa0 & new_n5021;
  assign new_n5023 = ~pb0 & new_n5022;
  assign new_n5024 = ~pc0 & new_n5023;
  assign new_n5025 = ~pu & new_n5024;
  assign new_n5026 = ~pj0 & new_n5025;
  assign new_n5027 = ~px & new_n5026;
  assign new_n5028 = ~pt & new_n5027;
  assign new_n5029 = ~pq & new_n5028;
  assign new_n5030 = ~pr & new_n5029;
  assign new_n5031 = ~pl & new_n5030;
  assign new_n5032 = ~pn & new_n5031;
  assign new_n5033 = pd & new_n4623;
  assign new_n5034 = ~py & new_n5033;
  assign new_n5035 = ~pa0 & new_n5034;
  assign new_n5036 = ~pb0 & new_n5035;
  assign new_n5037 = ~pc0 & new_n5036;
  assign new_n5038 = ~pu & new_n5037;
  assign new_n5039 = ~ps & new_n5038;
  assign new_n5040 = ~px & new_n5039;
  assign new_n5041 = ~pr & new_n5040;
  assign new_n5042 = ~pn & new_n5041;
  assign new_n5043 = ~pq & new_n5042;
  assign new_n5044 = ~pi & new_n5043;
  assign new_n5045 = ~pj & new_n5044;
  assign new_n5046 = pl0 & new_n1058;
  assign new_n5047 = pj0 & new_n5046;
  assign new_n5048 = ~pc & new_n5047;
  assign new_n5049 = ~pi0 & new_n5048;
  assign new_n5050 = ~pb0 & new_n5049;
  assign new_n5051 = ~pc0 & new_n5050;
  assign new_n5052 = ~pd0 & new_n5051;
  assign new_n5053 = ~ph0 & new_n5052;
  assign new_n5054 = ~pt & new_n5053;
  assign new_n5055 = ~px & new_n5054;
  assign new_n5056 = ~pr & new_n5055;
  assign new_n5057 = ~pn & new_n5056;
  assign new_n5058 = ~pq & new_n5057;
  assign new_n5059 = ~pj & new_n5058;
  assign new_n5060 = ~pl & new_n5059;
  assign new_n5061 = ~ps & new_n3036;
  assign new_n5062 = ~pg0 & new_n5061;
  assign new_n5063 = ~pj0 & new_n5062;
  assign new_n5064 = ~po & new_n5063;
  assign new_n5065 = ~pc0 & new_n5064;
  assign new_n5066 = pd0 & new_n5065;
  assign new_n5067 = pl0 & new_n5066;
  assign new_n5068 = pd & new_n5067;
  assign new_n5069 = ~pa0 & new_n5068;
  assign new_n5070 = ~pb0 & new_n5069;
  assign new_n5071 = ~py & new_n5070;
  assign new_n5072 = ~pu & new_n5071;
  assign new_n5073 = ~px & new_n5072;
  assign new_n5074 = ~pq & new_n5073;
  assign new_n5075 = ~pr & new_n5074;
  assign new_n5076 = pl0 & new_n3081;
  assign new_n5077 = ~pj0 & new_n5076;
  assign new_n5078 = ~pb & new_n5077;
  assign new_n5079 = ~pb0 & new_n5078;
  assign new_n5080 = ~pc0 & new_n5079;
  assign new_n5081 = pd0 & new_n5080;
  assign new_n5082 = ~ph0 & new_n5081;
  assign new_n5083 = ~py & new_n5082;
  assign new_n5084 = ~pa0 & new_n5083;
  assign new_n5085 = ~px & new_n5084;
  assign new_n5086 = ~pr & new_n5085;
  assign new_n5087 = ~pu & new_n5086;
  assign new_n5088 = ~pn & new_n5087;
  assign new_n5089 = ~pq & new_n5088;
  assign new_n5090 = ~pb0 & new_n4949;
  assign new_n5091 = ~pc0 & new_n5090;
  assign new_n5092 = ~pd0 & new_n5091;
  assign new_n5093 = pl0 & new_n5092;
  assign new_n5094 = ~py & new_n5093;
  assign new_n5095 = ~pa0 & new_n5094;
  assign new_n5096 = ~px & new_n5095;
  assign new_n5097 = ~pr & new_n5096;
  assign new_n5098 = ~pt & new_n5097;
  assign new_n5099 = ~pl & new_n5098;
  assign new_n5100 = ~pq & new_n5099;
  assign new_n5101 = ~pi0 & new_n1181;
  assign new_n5102 = ~pb & new_n5101;
  assign new_n5103 = pl0 & new_n5102;
  assign new_n5104 = ~pg0 & new_n5103;
  assign new_n5105 = pj0 & new_n5104;
  assign new_n5106 = ~pc & new_n5105;
  assign new_n5107 = ~pd0 & new_n5106;
  assign new_n5108 = ~ph0 & new_n5107;
  assign new_n5109 = ~pc0 & new_n5108;
  assign new_n5110 = ~px & new_n5109;
  assign new_n5111 = ~pb0 & new_n5110;
  assign new_n5112 = ~pq & new_n5111;
  assign new_n5113 = ~pr & new_n5112;
  assign new_n5114 = ~pk & new_n4961;
  assign new_n5115 = pl0 & new_n5114;
  assign new_n5116 = pj0 & new_n5115;
  assign new_n5117 = ~po & new_n5116;
  assign new_n5118 = ~pc & new_n5117;
  assign new_n5119 = ~pc0 & new_n5118;
  assign new_n5120 = ~pd0 & new_n5119;
  assign new_n5121 = ~pb0 & new_n5120;
  assign new_n5122 = ~pr & new_n5121;
  assign new_n5123 = ~px & new_n5122;
  assign new_n5124 = ~pj & new_n5123;
  assign new_n5125 = ~pq & new_n5124;
  assign new_n5126 = ~pc & new_n45;
  assign new_n5127 = pi0 & new_n5126;
  assign new_n5128 = pl0 & new_n5127;
  assign new_n5129 = ~pg0 & new_n5128;
  assign new_n5130 = ~pj0 & new_n5129;
  assign new_n5131 = ~po & new_n5130;
  assign new_n5132 = ~pc0 & new_n5131;
  assign new_n5133 = ~pd0 & new_n5132;
  assign new_n5134 = ~pb0 & new_n5133;
  assign new_n5135 = ~px & new_n5134;
  assign new_n5136 = ~py & new_n5135;
  assign new_n5137 = ~pq & new_n5136;
  assign new_n5138 = ~pr & new_n5137;
  assign new_n5139 = ~pm & new_n2946;
  assign new_n5140 = pl0 & new_n5139;
  assign new_n5141 = pj0 & new_n5140;
  assign new_n5142 = ~pd0 & new_n5141;
  assign new_n5143 = ~pb0 & new_n5142;
  assign new_n5144 = ~pc0 & new_n5143;
  assign new_n5145 = ~pq & new_n5144;
  assign new_n5146 = ~px & new_n5145;
  assign new_n5147 = ~pn & new_n3379;
  assign new_n5148 = ~pa & new_n5147;
  assign new_n5149 = ~pg0 & new_n5148;
  assign new_n5150 = ~pm & new_n5149;
  assign new_n5151 = ~pe0 & new_n5150;
  assign new_n5152 = ~ph0 & new_n5151;
  assign new_n5153 = pl0 & new_n5152;
  assign new_n5154 = ~pc0 & new_n5153;
  assign new_n5155 = ~pa0 & new_n5154;
  assign new_n5156 = ~pb0 & new_n5155;
  assign new_n5157 = ~px & new_n5156;
  assign new_n5158 = ~py & new_n5157;
  assign new_n5159 = pd & new_n4651;
  assign new_n5160 = ~ps & new_n5159;
  assign new_n5161 = ~pg0 & new_n5160;
  assign new_n5162 = ~pb0 & new_n5161;
  assign new_n5163 = ~pc0 & new_n5162;
  assign new_n5164 = pd0 & new_n5163;
  assign new_n5165 = ~ph0 & new_n5164;
  assign new_n5166 = ~py & new_n5165;
  assign new_n5167 = ~pj0 & new_n5166;
  assign new_n5168 = ~pa0 & new_n5167;
  assign new_n5169 = ~px & new_n5168;
  assign new_n5170 = ~pr & new_n5169;
  assign new_n5171 = ~pu & new_n5170;
  assign new_n5172 = ~pn & new_n5171;
  assign new_n5173 = ~pq & new_n5172;
  assign new_n5174 = ~pb0 & new_n2867;
  assign new_n5175 = ~pc0 & new_n5174;
  assign new_n5176 = pd0 & new_n5175;
  assign new_n5177 = ~ph0 & new_n5176;
  assign new_n5178 = ~pu & new_n5177;
  assign new_n5179 = ~px & new_n5178;
  assign new_n5180 = ~py & new_n5179;
  assign new_n5181 = ~pa0 & new_n5180;
  assign new_n5182 = ~pr & new_n5181;
  assign new_n5183 = pl0 & new_n5182;
  assign new_n5184 = ~pt & new_n5183;
  assign new_n5185 = ~pq & new_n5184;
  assign new_n5186 = ~pl & new_n5185;
  assign new_n5187 = ~pn & new_n5186;
  assign new_n5188 = ~pi & new_n5187;
  assign new_n5189 = ~pj & new_n5188;
  assign new_n5190 = ~ps & new_n105;
  assign new_n5191 = ~pj0 & new_n5190;
  assign new_n5192 = ~pc & new_n5191;
  assign new_n5193 = pi0 & new_n5192;
  assign new_n5194 = ~pd0 & new_n5193;
  assign new_n5195 = ~ph0 & new_n5194;
  assign new_n5196 = pl0 & new_n5195;
  assign new_n5197 = pd & new_n5196;
  assign new_n5198 = ~pb0 & new_n5197;
  assign new_n5199 = ~pc0 & new_n5198;
  assign new_n5200 = ~py & new_n5199;
  assign new_n5201 = ~pr & new_n5200;
  assign new_n5202 = ~px & new_n5201;
  assign new_n5203 = ~pn & new_n5202;
  assign new_n5204 = ~pq & new_n5203;
  assign new_n5205 = pl0 & new_n1679;
  assign new_n5206 = ~pg0 & new_n5205;
  assign new_n5207 = ~pj0 & new_n5206;
  assign new_n5208 = ~pc & new_n5207;
  assign new_n5209 = ~pb0 & new_n5208;
  assign new_n5210 = ~pc0 & new_n5209;
  assign new_n5211 = ~pd0 & new_n5210;
  assign new_n5212 = ~ph0 & new_n5211;
  assign new_n5213 = ~py & new_n5212;
  assign new_n5214 = ~pa0 & new_n5213;
  assign new_n5215 = ~px & new_n5214;
  assign new_n5216 = ~pr & new_n5215;
  assign new_n5217 = ~pt & new_n5216;
  assign new_n5218 = ~pn & new_n5217;
  assign new_n5219 = ~pq & new_n5218;
  assign new_n5220 = ~pg0 & new_n3798;
  assign new_n5221 = ~pj0 & new_n5220;
  assign new_n5222 = ~pb & new_n5221;
  assign new_n5223 = ~pc0 & new_n5222;
  assign new_n5224 = pd0 & new_n5223;
  assign new_n5225 = ~ph0 & new_n5224;
  assign new_n5226 = pl0 & new_n5225;
  assign new_n5227 = ~pa0 & new_n5226;
  assign new_n5228 = ~pb0 & new_n5227;
  assign new_n5229 = ~py & new_n5228;
  assign new_n5230 = ~pu & new_n5229;
  assign new_n5231 = ~px & new_n5230;
  assign new_n5232 = ~pq & new_n5231;
  assign new_n5233 = ~pr & new_n5232;
  assign new_n5234 = pl0 & new_n2946;
  assign new_n5235 = pd & new_n5234;
  assign new_n5236 = ~ps & new_n5235;
  assign new_n5237 = pj0 & new_n5236;
  assign new_n5238 = ~pc0 & new_n5237;
  assign new_n5239 = ~pd0 & new_n5238;
  assign new_n5240 = ~pb0 & new_n5239;
  assign new_n5241 = ~pr & new_n5240;
  assign new_n5242 = ~px & new_n5241;
  assign new_n5243 = ~pj & new_n5242;
  assign new_n5244 = ~pq & new_n5243;
  assign new_n5245 = ~pg0 & new_n3036;
  assign new_n5246 = ~pj0 & new_n5245;
  assign new_n5247 = ~po & new_n5246;
  assign new_n5248 = ~pb0 & new_n5247;
  assign new_n5249 = ~pc0 & new_n5248;
  assign new_n5250 = pd0 & new_n5249;
  assign new_n5251 = pl0 & new_n5250;
  assign new_n5252 = ~py & new_n5251;
  assign new_n5253 = ~pa0 & new_n5252;
  assign new_n5254 = ~px & new_n5253;
  assign new_n5255 = ~pr & new_n5254;
  assign new_n5256 = ~pu & new_n5255;
  assign new_n5257 = pn & new_n5256;
  assign new_n5258 = ~pq & new_n5257;
  assign new_n5259 = pi0 & new_n478;
  assign new_n5260 = ~pb & new_n5259;
  assign new_n5261 = ~ph0 & new_n5260;
  assign new_n5262 = pl0 & new_n5261;
  assign new_n5263 = ~pj0 & new_n5262;
  assign new_n5264 = ~pc & new_n5263;
  assign new_n5265 = ~pc0 & new_n5264;
  assign new_n5266 = ~pd0 & new_n5265;
  assign new_n5267 = ~pb0 & new_n5266;
  assign new_n5268 = ~px & new_n5267;
  assign new_n5269 = ~py & new_n5268;
  assign new_n5270 = ~pq & new_n5269;
  assign new_n5271 = ~pr & new_n5270;
  assign new_n5272 = ~po & new_n2867;
  assign new_n5273 = ~pb & new_n5272;
  assign new_n5274 = ~pc0 & new_n5273;
  assign new_n5275 = pd0 & new_n5274;
  assign new_n5276 = pl0 & new_n5275;
  assign new_n5277 = ~pg0 & new_n5276;
  assign new_n5278 = ~pa0 & new_n5277;
  assign new_n5279 = ~pb0 & new_n5278;
  assign new_n5280 = ~py & new_n5279;
  assign new_n5281 = ~pu & new_n5280;
  assign new_n5282 = ~px & new_n5281;
  assign new_n5283 = ~pq & new_n5282;
  assign new_n5284 = ~pr & new_n5283;
  assign new_n5285 = ~pd0 & new_n4542;
  assign new_n5286 = pl0 & new_n5285;
  assign new_n5287 = pj0 & new_n5286;
  assign new_n5288 = ~po & new_n5287;
  assign new_n5289 = ~pb0 & new_n5288;
  assign new_n5290 = ~pc0 & new_n5289;
  assign new_n5291 = ~px & new_n5290;
  assign new_n5292 = ~pq & new_n5291;
  assign new_n5293 = ~pr & new_n5292;
  assign new_n5294 = ~pj & new_n5293;
  assign new_n5295 = pn & new_n5294;
  assign new_n5296 = ~pg0 & new_n4705;
  assign new_n5297 = pj0 & new_n5296;
  assign new_n5298 = ~pc & new_n5297;
  assign new_n5299 = ~pi0 & new_n5298;
  assign new_n5300 = ~ph0 & new_n5299;
  assign new_n5301 = pl0 & new_n5300;
  assign new_n5302 = ~pd0 & new_n5301;
  assign new_n5303 = ~pb0 & new_n5302;
  assign new_n5304 = ~pc0 & new_n5303;
  assign new_n5305 = ~pq & new_n5304;
  assign new_n5306 = ~px & new_n5305;
  assign new_n5307 = ~pm & new_n2867;
  assign new_n5308 = ~pc0 & new_n5307;
  assign new_n5309 = pd0 & new_n5308;
  assign new_n5310 = pl0 & new_n5309;
  assign new_n5311 = ~po & new_n5310;
  assign new_n5312 = ~pa0 & new_n5311;
  assign new_n5313 = ~pb0 & new_n5312;
  assign new_n5314 = ~py & new_n5313;
  assign new_n5315 = ~pu & new_n5314;
  assign new_n5316 = ~px & new_n5315;
  assign new_n5317 = ~pi & new_n5316;
  assign new_n5318 = ~pq & new_n5317;
  assign new_n5319 = ~pk & new_n4653;
  assign new_n5320 = ~pb0 & new_n5319;
  assign new_n5321 = ~pc0 & new_n5320;
  assign new_n5322 = pd0 & new_n5321;
  assign new_n5323 = ~ph0 & new_n5322;
  assign new_n5324 = ~py & new_n5323;
  assign new_n5325 = ~pa0 & new_n5324;
  assign new_n5326 = ~px & new_n5325;
  assign new_n5327 = ~pr & new_n5326;
  assign new_n5328 = ~pu & new_n5327;
  assign new_n5329 = ~pn & new_n5328;
  assign new_n5330 = ~pq & new_n5329;
  assign new_n5331 = ~pg0 & new_n1679;
  assign new_n5332 = ~pj0 & new_n5331;
  assign new_n5333 = ~pc & new_n5332;
  assign new_n5334 = pi0 & new_n5333;
  assign new_n5335 = ~pc0 & new_n5334;
  assign new_n5336 = ~pd0 & new_n5335;
  assign new_n5337 = ~ph0 & new_n5336;
  assign new_n5338 = pl0 & new_n5337;
  assign new_n5339 = ~py & new_n5338;
  assign new_n5340 = ~pb0 & new_n5339;
  assign new_n5341 = ~px & new_n5340;
  assign new_n5342 = ~pr & new_n5341;
  assign new_n5343 = ~pt & new_n5342;
  assign new_n5344 = ~pn & new_n5343;
  assign new_n5345 = ~pq & new_n5344;
  assign new_n5346 = pd & new_n105;
  assign new_n5347 = ~ps & new_n5346;
  assign new_n5348 = ~pj0 & new_n5347;
  assign new_n5349 = ~pc & new_n5348;
  assign new_n5350 = ~pc0 & new_n5349;
  assign new_n5351 = ~pd0 & new_n5350;
  assign new_n5352 = ~ph0 & new_n5351;
  assign new_n5353 = pl0 & new_n5352;
  assign new_n5354 = ~pa0 & new_n5353;
  assign new_n5355 = ~pb0 & new_n5354;
  assign new_n5356 = ~py & new_n5355;
  assign new_n5357 = ~pr & new_n5356;
  assign new_n5358 = ~px & new_n5357;
  assign new_n5359 = ~pn & new_n5358;
  assign new_n5360 = ~pq & new_n5359;
  assign new_n5361 = pl0 & new_n4891;
  assign new_n5362 = ~po & new_n5361;
  assign new_n5363 = ~px & new_n5362;
  assign new_n5364 = ~py & new_n5363;
  assign new_n5365 = ~pa0 & new_n5364;
  assign new_n5366 = ~pb0 & new_n5365;
  assign new_n5367 = ~pt & new_n5366;
  assign new_n5368 = ~pu & new_n5367;
  assign new_n5369 = ~pr & new_n5368;
  assign new_n5370 = ~pl & new_n5369;
  assign new_n5371 = ~pq & new_n5370;
  assign new_n5372 = ~pi & new_n5371;
  assign new_n5373 = ~pj & new_n5372;
  assign new_n5374 = ~pk & new_n3939;
  assign new_n5375 = ~pd0 & new_n5374;
  assign new_n5376 = ~ph0 & new_n5375;
  assign new_n5377 = pl0 & new_n5376;
  assign new_n5378 = ~pg0 & new_n5377;
  assign new_n5379 = ~pb0 & new_n5378;
  assign new_n5380 = ~pc0 & new_n5379;
  assign new_n5381 = ~py & new_n5380;
  assign new_n5382 = ~pr & new_n5381;
  assign new_n5383 = ~px & new_n5382;
  assign new_n5384 = ~pn & new_n5383;
  assign new_n5385 = ~pq & new_n5384;
  assign new_n5386 = ~po & new_n5077;
  assign new_n5387 = ~pa0 & new_n5386;
  assign new_n5388 = ~pb0 & new_n5387;
  assign new_n5389 = ~pc0 & new_n5388;
  assign new_n5390 = pd0 & new_n5389;
  assign new_n5391 = ~px & new_n5390;
  assign new_n5392 = ~py & new_n5391;
  assign new_n5393 = ~pu & new_n5392;
  assign new_n5394 = ~pq & new_n5393;
  assign new_n5395 = ~pr & new_n5394;
  assign new_n5396 = ~pj & new_n5395;
  assign new_n5397 = pn & new_n5396;
  assign new_n5398 = pi0 & new_n441;
  assign new_n5399 = ~pb & new_n5398;
  assign new_n5400 = pl0 & new_n5399;
  assign new_n5401 = ~pg0 & new_n5400;
  assign new_n5402 = ~pj0 & new_n5401;
  assign new_n5403 = ~pc & new_n5402;
  assign new_n5404 = ~pd0 & new_n5403;
  assign new_n5405 = ~ph0 & new_n5404;
  assign new_n5406 = ~pc0 & new_n5405;
  assign new_n5407 = ~py & new_n5406;
  assign new_n5408 = ~pb0 & new_n5407;
  assign new_n5409 = ~pr & new_n5408;
  assign new_n5410 = ~px & new_n5409;
  assign new_n5411 = ~pb0 & new_n5273;
  assign new_n5412 = ~pc0 & new_n5411;
  assign new_n5413 = pd0 & new_n5412;
  assign new_n5414 = pl0 & new_n5413;
  assign new_n5415 = ~py & new_n5414;
  assign new_n5416 = ~pa0 & new_n5415;
  assign new_n5417 = ~px & new_n5416;
  assign new_n5418 = ~pr & new_n5417;
  assign new_n5419 = ~pu & new_n5418;
  assign new_n5420 = ~pi & new_n5419;
  assign new_n5421 = ~pq & new_n5420;
  assign new_n5422 = pl0 & new_n4666;
  assign new_n5423 = ~pg0 & new_n5422;
  assign new_n5424 = pj0 & new_n5423;
  assign new_n5425 = ~po & new_n5424;
  assign new_n5426 = ~pc0 & new_n5425;
  assign new_n5427 = ~pd0 & new_n5426;
  assign new_n5428 = ~pb0 & new_n5427;
  assign new_n5429 = ~pr & new_n5428;
  assign new_n5430 = ~px & new_n5429;
  assign new_n5431 = pn & new_n5430;
  assign new_n5432 = ~pq & new_n5431;
  assign new_n5433 = pl0 & new_n4829;
  assign new_n5434 = pj0 & new_n5433;
  assign new_n5435 = ~pc & new_n5434;
  assign new_n5436 = ~pi0 & new_n5435;
  assign new_n5437 = ~pd0 & new_n5436;
  assign new_n5438 = ~ph0 & new_n5437;
  assign new_n5439 = ~pc0 & new_n5438;
  assign new_n5440 = ~px & new_n5439;
  assign new_n5441 = ~pb0 & new_n5440;
  assign new_n5442 = ~pn & new_n5441;
  assign new_n5443 = ~pq & new_n5442;
  assign new_n5444 = pd0 & new_n5307;
  assign new_n5445 = pl0 & new_n5444;
  assign new_n5446 = ~pg0 & new_n5445;
  assign new_n5447 = ~po & new_n5446;
  assign new_n5448 = ~pb0 & new_n5447;
  assign new_n5449 = ~pc0 & new_n5448;
  assign new_n5450 = ~pa0 & new_n5449;
  assign new_n5451 = ~px & new_n5450;
  assign new_n5452 = ~py & new_n5451;
  assign new_n5453 = ~pq & new_n5452;
  assign new_n5454 = ~pu & new_n5453;
  assign new_n5455 = ~new_n752 & ~new_n5454;
  assign new_n5456 = ~new_n5432 & ~new_n5443;
  assign new_n5457 = new_n5455 & new_n5456;
  assign new_n5458 = ~new_n5410 & ~new_n5421;
  assign new_n5459 = ~new_n5385 & ~new_n5397;
  assign new_n5460 = new_n5458 & new_n5459;
  assign new_n5461 = new_n5457 & new_n5460;
  assign new_n5462 = ~new_n5360 & ~new_n5373;
  assign new_n5463 = ~new_n5330 & ~new_n5345;
  assign new_n5464 = new_n5462 & new_n5463;
  assign new_n5465 = ~new_n1252 & ~new_n5318;
  assign new_n5466 = ~new_n5295 & ~new_n5306;
  assign new_n5467 = new_n5465 & new_n5466;
  assign new_n5468 = new_n5464 & new_n5467;
  assign new_n5469 = new_n5461 & new_n5468;
  assign new_n5470 = ~new_n5271 & ~new_n5284;
  assign new_n5471 = ~new_n5244 & ~new_n5258;
  assign new_n5472 = new_n5470 & new_n5471;
  assign new_n5473 = ~new_n5219 & ~new_n5233;
  assign new_n5474 = ~new_n5189 & ~new_n5204;
  assign new_n5475 = new_n5473 & new_n5474;
  assign new_n5476 = new_n5472 & new_n5475;
  assign new_n5477 = ~new_n836 & ~new_n5173;
  assign new_n5478 = ~new_n5146 & ~new_n5158;
  assign new_n5479 = new_n5477 & new_n5478;
  assign new_n5480 = ~new_n5125 & ~new_n5138;
  assign new_n5481 = ~new_n5089 & ~new_n5100;
  assign new_n5482 = ~new_n5113 & new_n5481;
  assign new_n5483 = new_n5480 & new_n5482;
  assign new_n5484 = new_n5479 & new_n5483;
  assign new_n5485 = new_n5476 & new_n5484;
  assign new_n5486 = new_n5469 & new_n5485;
  assign new_n5487 = ~new_n5060 & ~new_n5075;
  assign new_n5488 = ~new_n5032 & ~new_n5045;
  assign new_n5489 = new_n5487 & new_n5488;
  assign new_n5490 = ~new_n796 & ~new_n5016;
  assign new_n5491 = ~new_n4997 & ~new_n5006;
  assign new_n5492 = new_n5490 & new_n5491;
  assign new_n5493 = new_n5489 & new_n5492;
  assign new_n5494 = ~new_n4973 & ~new_n4986;
  assign new_n5495 = ~new_n4947 & ~new_n4960;
  assign new_n5496 = new_n5494 & new_n5495;
  assign new_n5497 = ~new_n4920 & ~new_n4935;
  assign new_n5498 = ~new_n4889 & ~new_n4905;
  assign new_n5499 = new_n5497 & new_n5498;
  assign new_n5500 = new_n5496 & new_n5499;
  assign new_n5501 = new_n5493 & new_n5500;
  assign new_n5502 = ~new_n4862 & ~new_n4875;
  assign new_n5503 = ~new_n4840 & ~new_n4851;
  assign new_n5504 = new_n5502 & new_n5503;
  assign new_n5505 = ~new_n4816 & ~new_n4828;
  assign new_n5506 = ~new_n4790 & ~new_n4802;
  assign new_n5507 = new_n5505 & new_n5506;
  assign new_n5508 = new_n5504 & new_n5507;
  assign new_n5509 = ~new_n4760 & ~new_n4775;
  assign new_n5510 = ~new_n870 & ~new_n4749;
  assign new_n5511 = new_n5509 & new_n5510;
  assign new_n5512 = ~new_n4727 & ~new_n4738;
  assign new_n5513 = ~new_n4692 & ~new_n4704;
  assign new_n5514 = ~new_n4716 & new_n5513;
  assign new_n5515 = new_n5512 & new_n5514;
  assign new_n5516 = new_n5511 & new_n5515;
  assign new_n5517 = new_n5508 & new_n5516;
  assign new_n5518 = new_n5501 & new_n5517;
  assign new_n5519 = new_n5486 & new_n5518;
  assign new_n5520 = ~new_n4665 & ~new_n4678;
  assign new_n5521 = ~new_n4635 & ~new_n4650;
  assign new_n5522 = new_n5520 & new_n5521;
  assign new_n5523 = ~new_n4610 & ~new_n4621;
  assign new_n5524 = ~new_n4591 & ~new_n4602;
  assign new_n5525 = new_n5523 & new_n5524;
  assign new_n5526 = new_n5522 & new_n5525;
  assign new_n5527 = ~new_n4567 & ~new_n4580;
  assign new_n5528 = ~new_n4541 & ~new_n4554;
  assign new_n5529 = new_n5527 & new_n5528;
  assign new_n5530 = ~new_n4511 & ~new_n4526;
  assign new_n5531 = ~new_n4487 & ~new_n4498;
  assign new_n5532 = new_n5530 & new_n5531;
  assign new_n5533 = new_n5529 & new_n5532;
  assign new_n5534 = new_n5526 & new_n5533;
  assign new_n5535 = ~new_n4465 & ~new_n4476;
  assign new_n5536 = ~new_n4442 & ~new_n4454;
  assign new_n5537 = new_n5535 & new_n5536;
  assign new_n5538 = ~new_n4415 & ~new_n4429;
  assign new_n5539 = ~new_n4385 & ~new_n4400;
  assign new_n5540 = new_n5538 & new_n5539;
  assign new_n5541 = new_n5537 & new_n5540;
  assign new_n5542 = ~new_n4365 & ~new_n4370;
  assign new_n5543 = ~new_n4353 & ~new_n4358;
  assign new_n5544 = new_n5542 & new_n5543;
  assign new_n5545 = ~new_n4340 & ~new_n4347;
  assign new_n5546 = ~new_n4305 & ~new_n4320;
  assign new_n5547 = ~new_n4331 & new_n5546;
  assign new_n5548 = new_n5545 & new_n5547;
  assign new_n5549 = new_n5544 & new_n5548;
  assign new_n5550 = new_n5541 & new_n5549;
  assign new_n5551 = new_n5534 & new_n5550;
  assign new_n5552 = ~new_n4279 & ~new_n4293;
  assign new_n5553 = ~new_n4267 & ~new_n4274;
  assign new_n5554 = new_n5552 & new_n5553;
  assign new_n5555 = ~new_n4253 & ~new_n4262;
  assign new_n5556 = ~new_n4235 & ~new_n4244;
  assign new_n5557 = new_n5555 & new_n5556;
  assign new_n5558 = new_n5554 & new_n5557;
  assign new_n5559 = ~new_n4212 & ~new_n4224;
  assign new_n5560 = ~new_n4186 & ~new_n4199;
  assign new_n5561 = new_n5559 & new_n5560;
  assign new_n5562 = ~new_n4177 & ~new_n4181;
  assign new_n5563 = ~new_n4163 & ~new_n4170;
  assign new_n5564 = new_n5562 & new_n5563;
  assign new_n5565 = new_n5561 & new_n5564;
  assign new_n5566 = new_n5558 & new_n5565;
  assign new_n5567 = ~new_n4143 & ~new_n4152;
  assign new_n5568 = ~new_n4118 & ~new_n4130;
  assign new_n5569 = new_n5567 & new_n5568;
  assign new_n5570 = ~new_n4092 & ~new_n4107;
  assign new_n5571 = ~new_n4083 & ~new_n4087;
  assign new_n5572 = new_n5570 & new_n5571;
  assign new_n5573 = new_n5569 & new_n5572;
  assign new_n5574 = ~new_n4069 & ~new_n4075;
  assign new_n5575 = ~new_n4051 & ~new_n4060;
  assign new_n5576 = new_n5574 & new_n5575;
  assign new_n5577 = ~new_n4026 & ~new_n4038;
  assign new_n5578 = ~new_n590 & ~new_n4000;
  assign new_n5579 = ~new_n4015 & new_n5578;
  assign new_n5580 = new_n5577 & new_n5579;
  assign new_n5581 = new_n5576 & new_n5580;
  assign new_n5582 = new_n5573 & new_n5581;
  assign new_n5583 = new_n5566 & new_n5582;
  assign new_n5584 = new_n5551 & new_n5583;
  assign new_n5585 = new_n5519 & new_n5584;
  assign new_n5586 = ~new_n3986 & ~new_n3991;
  assign new_n5587 = ~new_n3970 & ~new_n3979;
  assign new_n5588 = new_n5586 & new_n5587;
  assign new_n5589 = ~new_n3950 & ~new_n3962;
  assign new_n5590 = ~new_n3924 & ~new_n3937;
  assign new_n5591 = new_n5589 & new_n5590;
  assign new_n5592 = new_n5588 & new_n5591;
  assign new_n5593 = ~new_n3899 & ~new_n3911;
  assign new_n5594 = ~new_n533 & ~new_n539;
  assign new_n5595 = new_n5593 & new_n5594;
  assign new_n5596 = ~new_n3873 & ~new_n3883;
  assign new_n5597 = ~new_n3862 & ~new_n3866;
  assign new_n5598 = new_n5596 & new_n5597;
  assign new_n5599 = new_n5595 & new_n5598;
  assign new_n5600 = new_n5592 & new_n5599;
  assign new_n5601 = ~new_n3848 & ~new_n3856;
  assign new_n5602 = ~new_n3824 & ~new_n3837;
  assign new_n5603 = new_n5601 & new_n5602;
  assign new_n5604 = ~new_n3797 & ~new_n3811;
  assign new_n5605 = ~new_n3785 & ~new_n3790;
  assign new_n5606 = new_n5604 & new_n5605;
  assign new_n5607 = new_n5603 & new_n5606;
  assign new_n5608 = ~new_n3767 & ~new_n3776;
  assign new_n5609 = ~new_n3748 & ~new_n3757;
  assign new_n5610 = new_n5608 & new_n5609;
  assign new_n5611 = ~new_n3727 & ~new_n3740;
  assign new_n5612 = ~new_n3688 & ~new_n3702;
  assign new_n5613 = ~new_n3715 & new_n5612;
  assign new_n5614 = new_n5611 & new_n5613;
  assign new_n5615 = new_n5610 & new_n5614;
  assign new_n5616 = new_n5607 & new_n5615;
  assign new_n5617 = new_n5600 & new_n5616;
  assign new_n5618 = ~new_n3676 & ~new_n3682;
  assign new_n5619 = ~new_n3664 & ~new_n3669;
  assign new_n5620 = new_n5618 & new_n5619;
  assign new_n5621 = ~new_n3647 & ~new_n3655;
  assign new_n5622 = ~new_n3625 & ~new_n3636;
  assign new_n5623 = new_n5621 & new_n5622;
  assign new_n5624 = new_n5620 & new_n5623;
  assign new_n5625 = ~new_n3599 & ~new_n3612;
  assign new_n5626 = ~new_n969 & ~new_n3586;
  assign new_n5627 = new_n5625 & new_n5626;
  assign new_n5628 = ~new_n3570 & ~new_n3577;
  assign new_n5629 = ~new_n3557 & ~new_n3562;
  assign new_n5630 = new_n5628 & new_n5629;
  assign new_n5631 = new_n5627 & new_n5630;
  assign new_n5632 = new_n5624 & new_n5631;
  assign new_n5633 = ~new_n660 & ~new_n1054;
  assign new_n5634 = ~new_n3539 & ~new_n3547;
  assign new_n5635 = new_n5633 & new_n5634;
  assign new_n5636 = ~new_n3525 & ~new_n3530;
  assign new_n5637 = ~new_n599 & ~new_n700;
  assign new_n5638 = new_n5636 & new_n5637;
  assign new_n5639 = new_n5635 & new_n5638;
  assign new_n5640 = ~new_n3512 & ~new_n3518;
  assign new_n5641 = ~new_n3497 & ~new_n3507;
  assign new_n5642 = new_n5640 & new_n5641;
  assign new_n5643 = ~new_n652 & ~new_n3491;
  assign new_n5644 = ~new_n3472 & ~new_n3480;
  assign new_n5645 = ~new_n3484 & new_n5644;
  assign new_n5646 = new_n5643 & new_n5645;
  assign new_n5647 = new_n5642 & new_n5646;
  assign new_n5648 = new_n5639 & new_n5647;
  assign new_n5649 = new_n5632 & new_n5648;
  assign new_n5650 = new_n5617 & new_n5649;
  assign new_n5651 = ~new_n864 & ~new_n3465;
  assign new_n5652 = ~new_n739 & ~new_n3456;
  assign new_n5653 = new_n5651 & new_n5652;
  assign new_n5654 = ~new_n3442 & ~new_n3447;
  assign new_n5655 = ~new_n3425 & ~new_n3435;
  assign new_n5656 = new_n5654 & new_n5655;
  assign new_n5657 = new_n5653 & new_n5656;
  assign new_n5658 = ~new_n747 & ~new_n782;
  assign new_n5659 = ~new_n3412 & ~new_n3418;
  assign new_n5660 = new_n5658 & new_n5659;
  assign new_n5661 = ~new_n3398 & ~new_n3407;
  assign new_n5662 = ~new_n787 & ~new_n3390;
  assign new_n5663 = new_n5661 & new_n5662;
  assign new_n5664 = new_n5660 & new_n5663;
  assign new_n5665 = new_n5657 & new_n5664;
  assign new_n5666 = ~new_n823 & ~new_n3378;
  assign new_n5667 = ~new_n3360 & ~new_n3369;
  assign new_n5668 = new_n5666 & new_n5667;
  assign new_n5669 = ~new_n3338 & ~new_n3350;
  assign new_n5670 = ~new_n859 & ~new_n3327;
  assign new_n5671 = new_n5669 & new_n5670;
  assign new_n5672 = new_n5668 & new_n5671;
  assign new_n5673 = ~new_n3308 & ~new_n3317;
  assign new_n5674 = ~new_n3291 & ~new_n3300;
  assign new_n5675 = new_n5673 & new_n5674;
  assign new_n5676 = ~new_n3268 & ~new_n3279;
  assign new_n5677 = ~new_n3234 & ~new_n3245;
  assign new_n5678 = ~new_n3256 & new_n5677;
  assign new_n5679 = new_n5676 & new_n5678;
  assign new_n5680 = new_n5675 & new_n5679;
  assign new_n5681 = new_n5672 & new_n5680;
  assign new_n5682 = new_n5665 & new_n5681;
  assign new_n5683 = ~new_n3050 & ~new_n3064;
  assign new_n5684 = ~new_n241 & ~new_n3035;
  assign new_n5685 = new_n5683 & new_n5684;
  assign new_n5686 = ~new_n3010 & ~new_n3019;
  assign new_n5687 = ~new_n2986 & ~new_n3000;
  assign new_n5688 = new_n5686 & new_n5687;
  assign new_n5689 = new_n5685 & new_n5688;
  assign new_n5690 = ~new_n1153 & ~new_n2972;
  assign new_n5691 = ~new_n2943 & ~new_n2957;
  assign new_n5692 = new_n5690 & new_n5691;
  assign new_n5693 = ~new_n101 & ~new_n2929;
  assign new_n5694 = ~new_n2882 & ~new_n2896;
  assign new_n5695 = ~new_n2914 & new_n5694;
  assign new_n5696 = new_n5693 & new_n5695;
  assign new_n5697 = new_n5692 & new_n5696;
  assign new_n5698 = new_n5689 & new_n5697;
  assign new_n5699 = ~new_n3209 & ~new_n3222;
  assign new_n5700 = ~new_n3190 & ~new_n3202;
  assign new_n5701 = new_n5699 & new_n5700;
  assign new_n5702 = ~new_n406 & ~new_n3177;
  assign new_n5703 = ~new_n3156 & ~new_n3168;
  assign new_n5704 = new_n5702 & new_n5703;
  assign new_n5705 = new_n5701 & new_n5704;
  assign new_n5706 = ~new_n3131 & ~new_n3145;
  assign new_n5707 = ~new_n3109 & ~new_n3118;
  assign new_n5708 = new_n5706 & new_n5707;
  assign new_n5709 = ~new_n3071 & ~new_n3080;
  assign new_n5710 = ~new_n310 & ~new_n3095;
  assign new_n5711 = new_n5709 & new_n5710;
  assign new_n5712 = new_n5708 & new_n5711;
  assign new_n5713 = new_n5705 & new_n5712;
  assign new_n5714 = new_n5698 & new_n5713;
  assign new_n5715 = new_n5682 & new_n5714;
  assign new_n5716 = new_n5650 & new_n5715;
  assign po0 = ~new_n5585 | ~new_n5716;
  assign new_n5718 = ~py & ~pz;
  assign new_n5719 = pj & new_n5718;
  assign new_n5720 = ~pn & new_n5719;
  assign new_n5721 = ~pc & new_n5720;
  assign new_n5722 = ~pm & new_n5721;
  assign new_n5723 = pt & new_n5722;
  assign new_n5724 = ~pd0 & new_n5723;
  assign new_n5725 = pi0 & new_n5724;
  assign new_n5726 = ~pd & new_n5725;
  assign new_n5727 = ~pg & new_n5726;
  assign new_n5728 = ~pi & new_n5727;
  assign new_n5729 = ~pf & new_n5728;
  assign new_n5730 = pm0 & new_n5729;
  assign new_n5731 = ~pe & new_n5730;
  assign new_n5732 = ~pc0 & new_n5731;
  assign new_n5733 = ~pj0 & new_n5732;
  assign new_n5734 = ~py & ~pn;
  assign new_n5735 = pj & new_n5734;
  assign new_n5736 = pl & new_n5735;
  assign new_n5737 = ~pc & new_n5736;
  assign new_n5738 = ~pm & new_n5737;
  assign new_n5739 = ~pg & new_n5738;
  assign new_n5740 = ~pi & new_n5739;
  assign new_n5741 = ~pd0 & new_n5740;
  assign new_n5742 = ~pd & new_n5741;
  assign new_n5743 = ~pe & new_n5742;
  assign new_n5744 = ~pf & new_n5743;
  assign new_n5745 = ~ph0 & new_n5744;
  assign new_n5746 = ~pj0 & new_n5745;
  assign new_n5747 = pm0 & new_n5746;
  assign new_n5748 = ~pa0 & new_n5747;
  assign new_n5749 = ~pc0 & new_n5748;
  assign new_n5750 = ps & ~pw;
  assign new_n5751 = pj & new_n5750;
  assign new_n5752 = ~pn & new_n5751;
  assign new_n5753 = ~pc & new_n5752;
  assign new_n5754 = ~pm & new_n5753;
  assign new_n5755 = ~pe & new_n5754;
  assign new_n5756 = ~pf & new_n5755;
  assign new_n5757 = ~pg & new_n5756;
  assign new_n5758 = pt & new_n5757;
  assign new_n5759 = ~pj0 & new_n5758;
  assign new_n5760 = pm0 & new_n5759;
  assign new_n5761 = ~pg0 & new_n5760;
  assign new_n5762 = ~pa0 & new_n5761;
  assign new_n5763 = ~pc0 & new_n5762;
  assign new_n5764 = ~py & new_n5763;
  assign new_n5765 = ~pz & new_n5764;
  assign new_n5766 = ~pd & new_n5737;
  assign new_n5767 = ~pg & new_n5766;
  assign new_n5768 = ~pd0 & new_n5767;
  assign new_n5769 = pi0 & new_n5768;
  assign new_n5770 = ~pb & new_n5769;
  assign new_n5771 = ~pe & new_n5770;
  assign new_n5772 = ~pf & new_n5771;
  assign new_n5773 = ~ph0 & new_n5772;
  assign new_n5774 = ~pj0 & new_n5773;
  assign new_n5775 = pm0 & new_n5774;
  assign new_n5776 = ~pc0 & new_n5775;
  assign new_n5777 = ~pg0 & new_n5776;
  assign new_n5778 = ~pw & ~py;
  assign new_n5779 = pj & new_n5778;
  assign new_n5780 = ~pn & new_n5779;
  assign new_n5781 = ~pc & new_n5780;
  assign new_n5782 = ~pd & new_n5781;
  assign new_n5783 = ~pg & new_n5782;
  assign new_n5784 = ~pi & new_n5783;
  assign new_n5785 = pt & new_n5784;
  assign new_n5786 = ~pb & new_n5785;
  assign new_n5787 = ~pe & new_n5786;
  assign new_n5788 = ~pf & new_n5787;
  assign new_n5789 = pm0 & new_n5788;
  assign new_n5790 = ~pc0 & new_n5789;
  assign new_n5791 = ~pj0 & new_n5790;
  assign new_n5792 = ~pz & new_n5791;
  assign new_n5793 = ~pa0 & new_n5792;
  assign new_n5794 = ps & ~pn;
  assign new_n5795 = pj & new_n5794;
  assign new_n5796 = pl & new_n5795;
  assign new_n5797 = ~pc & new_n5796;
  assign new_n5798 = ~pb & new_n5797;
  assign new_n5799 = ~pg & new_n5798;
  assign new_n5800 = ~pi & new_n5799;
  assign new_n5801 = ~pd0 & new_n5800;
  assign new_n5802 = pi0 & new_n5801;
  assign new_n5803 = ~pe & new_n5802;
  assign new_n5804 = ~pf & new_n5803;
  assign new_n5805 = ~ph0 & new_n5804;
  assign new_n5806 = ~pj0 & new_n5805;
  assign new_n5807 = pm0 & new_n5806;
  assign new_n5808 = ~py & new_n5807;
  assign new_n5809 = ~pc0 & new_n5808;
  assign new_n5810 = ~pe & new_n5798;
  assign new_n5811 = ~pf & new_n5810;
  assign new_n5812 = ~pg & new_n5811;
  assign new_n5813 = ~pd0 & new_n5812;
  assign new_n5814 = ~pj0 & new_n5813;
  assign new_n5815 = pm0 & new_n5814;
  assign new_n5816 = ~pg0 & new_n5815;
  assign new_n5817 = ~pa0 & new_n5816;
  assign new_n5818 = ~pc0 & new_n5817;
  assign new_n5819 = ~py & new_n5818;
  assign new_n5820 = ~pz & new_n5819;
  assign new_n5821 = ~pc0 & ~py;
  assign new_n5822 = ~pj & new_n5821;
  assign new_n5823 = ~ps & new_n5822;
  assign new_n5824 = ~pc & new_n5823;
  assign new_n5825 = ~pg & new_n5824;
  assign new_n5826 = ~pd0 & new_n5825;
  assign new_n5827 = pi0 & new_n5826;
  assign new_n5828 = pd & new_n5827;
  assign new_n5829 = ~pe & new_n5828;
  assign new_n5830 = ~pf & new_n5829;
  assign new_n5831 = ~ph0 & new_n5830;
  assign new_n5832 = pm0 & new_n5831;
  assign new_n5833 = ~pf0 & new_n5832;
  assign new_n5834 = ~pg0 & new_n5833;
  assign new_n5835 = ~pj0 & new_n5834;
  assign new_n5836 = ~pj & new_n5718;
  assign new_n5837 = ~pl & new_n5836;
  assign new_n5838 = ~pc & new_n5837;
  assign new_n5839 = ~pi & new_n5838;
  assign new_n5840 = ~pt & new_n5839;
  assign new_n5841 = ~pd0 & new_n5840;
  assign new_n5842 = pi0 & new_n5841;
  assign new_n5843 = ~pf & new_n5842;
  assign new_n5844 = ~pg & new_n5843;
  assign new_n5845 = ~pe & new_n5844;
  assign new_n5846 = pm0 & new_n5845;
  assign new_n5847 = ~pf0 & new_n5846;
  assign new_n5848 = ~pc0 & new_n5847;
  assign new_n5849 = ~pj0 & new_n5848;
  assign new_n5850 = pj & new_n1763;
  assign new_n5851 = ~py & new_n5850;
  assign new_n5852 = ~pc & new_n5851;
  assign new_n5853 = pi0 & new_n5852;
  assign new_n5854 = ~pm & new_n5853;
  assign new_n5855 = ~pk & new_n5854;
  assign new_n5856 = ~pi & new_n5855;
  assign new_n5857 = ~pd0 & new_n5856;
  assign new_n5858 = ~pg & new_n5857;
  assign new_n5859 = ~pe & new_n5858;
  assign new_n5860 = ~pf & new_n5859;
  assign new_n5861 = pm0 & new_n5860;
  assign new_n5862 = ~ph0 & new_n5861;
  assign new_n5863 = ~pw & new_n5719;
  assign new_n5864 = ~pc & new_n5863;
  assign new_n5865 = ~pg & new_n5864;
  assign new_n5866 = ~pm & new_n5865;
  assign new_n5867 = ~pk & new_n5866;
  assign new_n5868 = ~pe & new_n5867;
  assign new_n5869 = ~pf & new_n5868;
  assign new_n5870 = pm0 & new_n5869;
  assign new_n5871 = ~pg0 & new_n5870;
  assign new_n5872 = ~pj0 & new_n5871;
  assign new_n5873 = ~pa0 & new_n5872;
  assign new_n5874 = ~pc0 & new_n5873;
  assign new_n5875 = ~pc0 & ~pz;
  assign new_n5876 = ~pj & new_n5875;
  assign new_n5877 = ~ps & new_n5876;
  assign new_n5878 = ~pc & new_n5877;
  assign new_n5879 = ~pd0 & new_n5878;
  assign new_n5880 = ~pi0 & new_n5879;
  assign new_n5881 = pd & new_n5880;
  assign new_n5882 = ~ph & new_n5881;
  assign new_n5883 = ~pi & new_n5882;
  assign new_n5884 = ~pg & new_n5883;
  assign new_n5885 = ~pe & new_n5884;
  assign new_n5886 = ~pf & new_n5885;
  assign new_n5887 = pj0 & new_n5886;
  assign new_n5888 = pm0 & new_n5887;
  assign new_n5889 = ~pj & new_n5778;
  assign new_n5890 = ~ps & new_n5889;
  assign new_n5891 = ~pc & new_n5890;
  assign new_n5892 = ~ph & new_n5891;
  assign new_n5893 = ~pi & new_n5892;
  assign new_n5894 = pd & new_n5893;
  assign new_n5895 = ~pf & new_n5894;
  assign new_n5896 = ~pg & new_n5895;
  assign new_n5897 = ~pe & new_n5896;
  assign new_n5898 = pm0 & new_n5897;
  assign new_n5899 = ~ph0 & new_n5898;
  assign new_n5900 = ~pa0 & new_n5899;
  assign new_n5901 = ~pc0 & new_n5900;
  assign new_n5902 = ~pt & new_n5838;
  assign new_n5903 = ~pd0 & new_n5902;
  assign new_n5904 = pi0 & new_n5903;
  assign new_n5905 = ~pg & new_n5904;
  assign new_n5906 = ~ph & new_n5905;
  assign new_n5907 = ~pf & new_n5906;
  assign new_n5908 = pm0 & new_n5907;
  assign new_n5909 = ~pe & new_n5908;
  assign new_n5910 = ~pc0 & new_n5909;
  assign new_n5911 = ~pg0 & new_n5910;
  assign new_n5912 = ~pj & new_n3448;
  assign new_n5913 = pn & new_n5912;
  assign new_n5914 = ~pc & new_n5913;
  assign new_n5915 = ~pf & new_n5914;
  assign new_n5916 = ~pg & new_n5915;
  assign new_n5917 = ~pd0 & new_n5916;
  assign new_n5918 = ~ph0 & new_n5917;
  assign new_n5919 = ~pe & new_n5918;
  assign new_n5920 = ~pf0 & new_n5919;
  assign new_n5921 = ~pj0 & new_n5920;
  assign new_n5922 = pm0 & new_n5921;
  assign new_n5923 = ~pc0 & new_n5922;
  assign new_n5924 = ~pg0 & new_n5923;
  assign new_n5925 = ~pc0 & pj0;
  assign new_n5926 = ~pj & new_n5925;
  assign new_n5927 = ~pz & new_n5926;
  assign new_n5928 = ~pc & new_n5927;
  assign new_n5929 = ~pi0 & new_n5928;
  assign new_n5930 = ~pk & new_n5929;
  assign new_n5931 = ~pi & new_n5930;
  assign new_n5932 = ~pd0 & new_n5931;
  assign new_n5933 = ~ph & new_n5932;
  assign new_n5934 = ~pf & new_n5933;
  assign new_n5935 = ~pg & new_n5934;
  assign new_n5936 = pm0 & new_n5935;
  assign new_n5937 = ~pe & new_n5936;
  assign new_n5938 = ~pw & new_n5912;
  assign new_n5939 = ~pc & new_n5938;
  assign new_n5940 = ~pi & new_n5939;
  assign new_n5941 = ~pk & new_n5940;
  assign new_n5942 = ~pg & new_n5941;
  assign new_n5943 = ~ph & new_n5942;
  assign new_n5944 = ~pf & new_n5943;
  assign new_n5945 = ~ph0 & new_n5944;
  assign new_n5946 = ~pe & new_n5945;
  assign new_n5947 = ~pc0 & new_n5946;
  assign new_n5948 = pm0 & new_n5947;
  assign new_n5949 = pn & new_n5836;
  assign new_n5950 = ~pc & new_n5949;
  assign new_n5951 = ~pd0 & new_n5950;
  assign new_n5952 = pi0 & new_n5951;
  assign new_n5953 = ~pg & new_n5952;
  assign new_n5954 = ~ph & new_n5953;
  assign new_n5955 = ~pf & new_n5954;
  assign new_n5956 = pm0 & new_n5955;
  assign new_n5957 = ~pe & new_n5956;
  assign new_n5958 = ~pc0 & new_n5957;
  assign new_n5959 = ~pg0 & new_n5958;
  assign new_n5960 = ~ph0 & new_n5797;
  assign new_n5961 = ~pi & new_n5960;
  assign new_n5962 = ~pj0 & new_n5961;
  assign new_n5963 = pm0 & new_n5962;
  assign new_n5964 = ~pe0 & new_n5963;
  assign new_n5965 = ~pa0 & new_n5964;
  assign new_n5966 = ~pc0 & new_n5965;
  assign new_n5967 = ~pw & new_n5966;
  assign new_n5968 = ~py & new_n5967;
  assign new_n5969 = ~pc0 & pm0;
  assign new_n5970 = ~py & new_n5969;
  assign new_n5971 = ~pz & new_n5970;
  assign new_n5972 = ~pc & new_n5971;
  assign new_n5973 = ~pm & new_n5972;
  assign new_n5974 = ~pd0 & new_n5973;
  assign new_n5975 = pi0 & new_n5974;
  assign new_n5976 = ~pi & new_n5975;
  assign new_n5977 = ~pg & new_n5976;
  assign new_n5978 = ~ph & new_n5977;
  assign new_n5979 = ~pe & new_n5978;
  assign new_n5980 = ~pf & new_n5979;
  assign new_n5981 = pj & new_n5821;
  assign new_n5982 = ~pn & new_n5981;
  assign new_n5983 = ~pc & new_n5982;
  assign new_n5984 = ~pm & new_n5983;
  assign new_n5985 = pt & new_n5984;
  assign new_n5986 = ~pd0 & new_n5985;
  assign new_n5987 = pi0 & new_n5986;
  assign new_n5988 = ~pd & new_n5987;
  assign new_n5989 = ~pf & new_n5988;
  assign new_n5990 = ~pg & new_n5989;
  assign new_n5991 = ~pe & new_n5990;
  assign new_n5992 = pm0 & new_n5991;
  assign new_n5993 = ~ph0 & new_n5992;
  assign new_n5994 = ~pg0 & new_n5993;
  assign new_n5995 = ~pj0 & new_n5994;
  assign new_n5996 = ~pg & new_n5722;
  assign new_n5997 = pt & new_n5996;
  assign new_n5998 = ~pd0 & new_n5997;
  assign new_n5999 = ~pd & new_n5998;
  assign new_n6000 = ~pe & new_n5999;
  assign new_n6001 = ~pf & new_n6000;
  assign new_n6002 = pm0 & new_n6001;
  assign new_n6003 = ~pg0 & new_n6002;
  assign new_n6004 = ~pj0 & new_n6003;
  assign new_n6005 = ~pa0 & new_n6004;
  assign new_n6006 = ~pc0 & new_n6005;
  assign new_n6007 = ps & ~py;
  assign new_n6008 = pj & new_n6007;
  assign new_n6009 = ~pn & new_n6008;
  assign new_n6010 = ~pc & new_n6009;
  assign new_n6011 = ~pm & new_n6010;
  assign new_n6012 = ~pg & new_n6011;
  assign new_n6013 = ~pi & new_n6012;
  assign new_n6014 = pt & new_n6013;
  assign new_n6015 = ~pd0 & new_n6014;
  assign new_n6016 = ~pe & new_n6015;
  assign new_n6017 = ~pf & new_n6016;
  assign new_n6018 = pm0 & new_n6017;
  assign new_n6019 = ~pc0 & new_n6018;
  assign new_n6020 = ~pj0 & new_n6019;
  assign new_n6021 = ~pz & new_n6020;
  assign new_n6022 = ~pa0 & new_n6021;
  assign new_n6023 = pm0 & new_n5772;
  assign new_n6024 = ~pg0 & new_n6023;
  assign new_n6025 = ~pj0 & new_n6024;
  assign new_n6026 = ~pz & new_n6025;
  assign new_n6027 = ~pc0 & new_n6026;
  assign new_n6028 = ~ph0 & new_n5788;
  assign new_n6029 = ~pj0 & new_n6028;
  assign new_n6030 = pm0 & new_n6029;
  assign new_n6031 = ~pa0 & new_n6030;
  assign new_n6032 = ~pc0 & new_n6031;
  assign new_n6033 = pm0 & new_n5804;
  assign new_n6034 = ~pc0 & new_n6033;
  assign new_n6035 = ~pj0 & new_n6034;
  assign new_n6036 = ~py & new_n6035;
  assign new_n6037 = ~pz & new_n6036;
  assign new_n6038 = pm0 & new_n5813;
  assign new_n6039 = ~ph0 & new_n6038;
  assign new_n6040 = ~pj0 & new_n6039;
  assign new_n6041 = ~pc0 & new_n6040;
  assign new_n6042 = ~pg0 & new_n6041;
  assign new_n6043 = ~py & new_n6042;
  assign new_n6044 = ~pa0 & new_n6043;
  assign new_n6045 = ~ps & new_n5836;
  assign new_n6046 = ~pc & new_n6045;
  assign new_n6047 = ~pg & new_n6046;
  assign new_n6048 = ~pd0 & new_n6047;
  assign new_n6049 = pi0 & new_n6048;
  assign new_n6050 = pd & new_n6049;
  assign new_n6051 = ~pe & new_n6050;
  assign new_n6052 = ~pf & new_n6051;
  assign new_n6053 = ~pf0 & new_n6052;
  assign new_n6054 = ~pj0 & new_n6053;
  assign new_n6055 = pm0 & new_n6054;
  assign new_n6056 = ~pc0 & new_n6055;
  assign new_n6057 = ~pg0 & new_n6056;
  assign new_n6058 = ~pl & new_n5822;
  assign new_n6059 = ~pc & new_n6058;
  assign new_n6060 = ~pi & new_n6059;
  assign new_n6061 = ~pt & new_n6060;
  assign new_n6062 = ~pd0 & new_n6061;
  assign new_n6063 = pi0 & new_n6062;
  assign new_n6064 = ~pf & new_n6063;
  assign new_n6065 = ~pg & new_n6064;
  assign new_n6066 = ~pe & new_n6065;
  assign new_n6067 = ~pf0 & new_n6066;
  assign new_n6068 = ~ph0 & new_n6067;
  assign new_n6069 = ~pj0 & new_n6068;
  assign new_n6070 = pm0 & new_n6069;
  assign new_n6071 = pj & new_n5875;
  assign new_n6072 = ~py & new_n6071;
  assign new_n6073 = ~pc & new_n6072;
  assign new_n6074 = pi0 & new_n6073;
  assign new_n6075 = ~pm & new_n6074;
  assign new_n6076 = ~pk & new_n6075;
  assign new_n6077 = ~pi & new_n6076;
  assign new_n6078 = ~pd0 & new_n6077;
  assign new_n6079 = ~pg & new_n6078;
  assign new_n6080 = ~pe & new_n6079;
  assign new_n6081 = ~pf & new_n6080;
  assign new_n6082 = ~pj0 & new_n6081;
  assign new_n6083 = pm0 & new_n6082;
  assign new_n6084 = pj & new_n3448;
  assign new_n6085 = ~pw & new_n6084;
  assign new_n6086 = ~pc & new_n6085;
  assign new_n6087 = ~pg & new_n6086;
  assign new_n6088 = ~pm & new_n6087;
  assign new_n6089 = ~pk & new_n6088;
  assign new_n6090 = ~pe & new_n6089;
  assign new_n6091 = ~pf & new_n6090;
  assign new_n6092 = ~ph0 & new_n6091;
  assign new_n6093 = ~pj0 & new_n6092;
  assign new_n6094 = pm0 & new_n6093;
  assign new_n6095 = ~pc0 & new_n6094;
  assign new_n6096 = ~pg0 & new_n6095;
  assign new_n6097 = ~pc0 & ~pg0;
  assign new_n6098 = ~pj & new_n6097;
  assign new_n6099 = ~ps & new_n6098;
  assign new_n6100 = ~pc & new_n6099;
  assign new_n6101 = ~pd0 & new_n6100;
  assign new_n6102 = ~pi0 & new_n6101;
  assign new_n6103 = pd & new_n6102;
  assign new_n6104 = ~pg & new_n6103;
  assign new_n6105 = ~ph & new_n6104;
  assign new_n6106 = ~pf & new_n6105;
  assign new_n6107 = ~ph0 & new_n6106;
  assign new_n6108 = ~pe & new_n6107;
  assign new_n6109 = pj0 & new_n6108;
  assign new_n6110 = pm0 & new_n6109;
  assign new_n6111 = ~ph & new_n6046;
  assign new_n6112 = ~pd0 & new_n6111;
  assign new_n6113 = pd & new_n6112;
  assign new_n6114 = ~pf & new_n6113;
  assign new_n6115 = ~pg & new_n6114;
  assign new_n6116 = ~pe & new_n6115;
  assign new_n6117 = ~pg0 & new_n6116;
  assign new_n6118 = pm0 & new_n6117;
  assign new_n6119 = ~pa0 & new_n6118;
  assign new_n6120 = ~pc0 & new_n6119;
  assign new_n6121 = pn & new_n5822;
  assign new_n6122 = ~pc & new_n6121;
  assign new_n6123 = ~pi & new_n6122;
  assign new_n6124 = ~pd0 & new_n6123;
  assign new_n6125 = pi0 & new_n6124;
  assign new_n6126 = ~pf & new_n6125;
  assign new_n6127 = ~pg & new_n6126;
  assign new_n6128 = ~pe & new_n6127;
  assign new_n6129 = ~pf0 & new_n6128;
  assign new_n6130 = ~ph0 & new_n6129;
  assign new_n6131 = ~pj0 & new_n6130;
  assign new_n6132 = pm0 & new_n6131;
  assign new_n6133 = ~pg & new_n5950;
  assign new_n6134 = ~pi & new_n6133;
  assign new_n6135 = ~pd0 & new_n6134;
  assign new_n6136 = ~pe & new_n6135;
  assign new_n6137 = ~pf & new_n6136;
  assign new_n6138 = ~pf0 & new_n6137;
  assign new_n6139 = ~pj0 & new_n6138;
  assign new_n6140 = pm0 & new_n6139;
  assign new_n6141 = ~pa0 & new_n6140;
  assign new_n6142 = ~pc0 & new_n6141;
  assign new_n6143 = ~pj & new_n685;
  assign new_n6144 = ~pc0 & new_n6143;
  assign new_n6145 = ~pc & new_n6144;
  assign new_n6146 = ~pi0 & new_n6145;
  assign new_n6147 = ~pk & new_n6146;
  assign new_n6148 = ~ph & new_n6147;
  assign new_n6149 = ~pd0 & new_n6148;
  assign new_n6150 = ~pg & new_n6149;
  assign new_n6151 = ~pe & new_n6150;
  assign new_n6152 = ~pf & new_n6151;
  assign new_n6153 = pm0 & new_n6152;
  assign new_n6154 = ~ph0 & new_n6153;
  assign new_n6155 = ~pa0 & ~pz;
  assign new_n6156 = ~pj & new_n6155;
  assign new_n6157 = ~py & new_n6156;
  assign new_n6158 = ~pc & new_n6157;
  assign new_n6159 = ~pd0 & new_n6158;
  assign new_n6160 = ~pk & new_n6159;
  assign new_n6161 = ~pg & new_n6160;
  assign new_n6162 = ~ph & new_n6161;
  assign new_n6163 = ~pf & new_n6162;
  assign new_n6164 = pm0 & new_n6163;
  assign new_n6165 = ~pe & new_n6164;
  assign new_n6166 = ~pc0 & new_n6165;
  assign new_n6167 = ~pg0 & new_n6166;
  assign new_n6168 = ~pw & new_n6155;
  assign new_n6169 = ~py & new_n6168;
  assign new_n6170 = ~pc & new_n6169;
  assign new_n6171 = ~pi & new_n6170;
  assign new_n6172 = ~pb & new_n6171;
  assign new_n6173 = ~pf & new_n6172;
  assign new_n6174 = ~pg & new_n6173;
  assign new_n6175 = ~pe & new_n6174;
  assign new_n6176 = pm0 & new_n6175;
  assign new_n6177 = ~pf0 & new_n6176;
  assign new_n6178 = ~pc0 & new_n6177;
  assign new_n6179 = ~pj0 & new_n6178;
  assign new_n6180 = pm0 & new_n5797;
  assign new_n6181 = ~pi & new_n6180;
  assign new_n6182 = ~pe0 & new_n6181;
  assign new_n6183 = ~pj0 & new_n6182;
  assign new_n6184 = ~pc0 & new_n6183;
  assign new_n6185 = ~pz & new_n6184;
  assign new_n6186 = ~pa0 & new_n6185;
  assign new_n6187 = ~pw & new_n6186;
  assign new_n6188 = ~py & new_n6187;
  assign new_n6189 = ~ph0 & pm0;
  assign new_n6190 = ~py & new_n6189;
  assign new_n6191 = ~pc0 & new_n6190;
  assign new_n6192 = ~pc & new_n6191;
  assign new_n6193 = ~pm & new_n6192;
  assign new_n6194 = ~pd0 & new_n6193;
  assign new_n6195 = pi0 & new_n6194;
  assign new_n6196 = ~pi & new_n6195;
  assign new_n6197 = ~pg & new_n6196;
  assign new_n6198 = ~ph & new_n6197;
  assign new_n6199 = ~pe & new_n6198;
  assign new_n6200 = ~pf & new_n6199;
  assign new_n6201 = ~pn & new_n6084;
  assign new_n6202 = ~pc & new_n6201;
  assign new_n6203 = ~pm & new_n6202;
  assign new_n6204 = ~pg & new_n6203;
  assign new_n6205 = pt & new_n6204;
  assign new_n6206 = ~pd0 & new_n6205;
  assign new_n6207 = ~pd & new_n6206;
  assign new_n6208 = ~pe & new_n6207;
  assign new_n6209 = ~pf & new_n6208;
  assign new_n6210 = ~ph0 & new_n6209;
  assign new_n6211 = ~pj0 & new_n6210;
  assign new_n6212 = pm0 & new_n6211;
  assign new_n6213 = ~pc0 & new_n6212;
  assign new_n6214 = ~pg0 & new_n6213;
  assign new_n6215 = ~pf & new_n6011;
  assign new_n6216 = ~pg & new_n6215;
  assign new_n6217 = pt & new_n6216;
  assign new_n6218 = ~pd0 & new_n6217;
  assign new_n6219 = ~ph0 & new_n6218;
  assign new_n6220 = ~pe & new_n6219;
  assign new_n6221 = pm0 & new_n6220;
  assign new_n6222 = ~pg0 & new_n6221;
  assign new_n6223 = ~pj0 & new_n6222;
  assign new_n6224 = ~pa0 & new_n6223;
  assign new_n6225 = ~pc0 & new_n6224;
  assign new_n6226 = ~pm & new_n5797;
  assign new_n6227 = ~pe & new_n6226;
  assign new_n6228 = ~pf & new_n6227;
  assign new_n6229 = ~pg & new_n6228;
  assign new_n6230 = ~pi & new_n6229;
  assign new_n6231 = ~pj0 & new_n6230;
  assign new_n6232 = pm0 & new_n6231;
  assign new_n6233 = ~pc0 & new_n6232;
  assign new_n6234 = ~pz & new_n6233;
  assign new_n6235 = ~pa0 & new_n6234;
  assign new_n6236 = ~pw & new_n6235;
  assign new_n6237 = ~py & new_n6236;
  assign new_n6238 = ~pf & new_n5766;
  assign new_n6239 = ~pg & new_n6238;
  assign new_n6240 = ~pd0 & new_n6239;
  assign new_n6241 = ~pb & new_n6240;
  assign new_n6242 = pm0 & new_n6241;
  assign new_n6243 = ~pe & new_n6242;
  assign new_n6244 = ~pj0 & new_n6243;
  assign new_n6245 = ~pc0 & new_n6244;
  assign new_n6246 = ~pg0 & new_n6245;
  assign new_n6247 = ~pz & new_n6246;
  assign new_n6248 = ~pa0 & new_n6247;
  assign new_n6249 = ~pf & new_n5798;
  assign new_n6250 = ~pg & new_n6249;
  assign new_n6251 = ~pd0 & new_n6250;
  assign new_n6252 = pi0 & new_n6251;
  assign new_n6253 = ~ph0 & new_n6252;
  assign new_n6254 = ~pe & new_n6253;
  assign new_n6255 = pm0 & new_n6254;
  assign new_n6256 = ~pg0 & new_n6255;
  assign new_n6257 = ~pj0 & new_n6256;
  assign new_n6258 = ~py & new_n6257;
  assign new_n6259 = ~pc0 & new_n6258;
  assign new_n6260 = ~pb & new_n5753;
  assign new_n6261 = ~pf & new_n6260;
  assign new_n6262 = ~pg & new_n6261;
  assign new_n6263 = ~pi & new_n6262;
  assign new_n6264 = pt & new_n6263;
  assign new_n6265 = pm0 & new_n6264;
  assign new_n6266 = ~pe & new_n6265;
  assign new_n6267 = ~pj0 & new_n6266;
  assign new_n6268 = ~pa0 & new_n6267;
  assign new_n6269 = ~pc0 & new_n6268;
  assign new_n6270 = ~py & new_n6269;
  assign new_n6271 = ~pz & new_n6270;
  assign new_n6272 = ~pi & new_n5824;
  assign new_n6273 = ~pd0 & new_n6272;
  assign new_n6274 = pi0 & new_n6273;
  assign new_n6275 = pd & new_n6274;
  assign new_n6276 = ~pf & new_n6275;
  assign new_n6277 = ~pg & new_n6276;
  assign new_n6278 = ~pe & new_n6277;
  assign new_n6279 = ~pf0 & new_n6278;
  assign new_n6280 = ~ph0 & new_n6279;
  assign new_n6281 = ~pj0 & new_n6280;
  assign new_n6282 = pm0 & new_n6281;
  assign new_n6283 = ~pe & new_n5891;
  assign new_n6284 = ~pf & new_n6283;
  assign new_n6285 = ~pg & new_n6284;
  assign new_n6286 = pd & new_n6285;
  assign new_n6287 = pm0 & new_n6286;
  assign new_n6288 = ~pf0 & new_n6287;
  assign new_n6289 = ~pj0 & new_n6288;
  assign new_n6290 = ~pc0 & new_n6289;
  assign new_n6291 = ~pg0 & new_n6290;
  assign new_n6292 = ~pz & new_n6291;
  assign new_n6293 = ~pa0 & new_n6292;
  assign new_n6294 = pj & new_n6097;
  assign new_n6295 = ~py & new_n6294;
  assign new_n6296 = ~pc & new_n6295;
  assign new_n6297 = pi0 & new_n6296;
  assign new_n6298 = ~pm & new_n6297;
  assign new_n6299 = ~pk & new_n6298;
  assign new_n6300 = ~pg & new_n6299;
  assign new_n6301 = ~pd0 & new_n6300;
  assign new_n6302 = ~pf & new_n6301;
  assign new_n6303 = ~ph0 & new_n6302;
  assign new_n6304 = ~pe & new_n6303;
  assign new_n6305 = ~pj0 & new_n6304;
  assign new_n6306 = pm0 & new_n6305;
  assign new_n6307 = ~pg & new_n5881;
  assign new_n6308 = ~ph & new_n6307;
  assign new_n6309 = ~pf & new_n6308;
  assign new_n6310 = pm0 & new_n6309;
  assign new_n6311 = ~pe & new_n6310;
  assign new_n6312 = ~pg0 & new_n6311;
  assign new_n6313 = pj0 & new_n6312;
  assign new_n6314 = ~pg & new_n5891;
  assign new_n6315 = ~ph & new_n6314;
  assign new_n6316 = pd & new_n6315;
  assign new_n6317 = ~pe & new_n6316;
  assign new_n6318 = ~pf & new_n6317;
  assign new_n6319 = ~ph0 & new_n6318;
  assign new_n6320 = ~pg0 & new_n6319;
  assign new_n6321 = pm0 & new_n6320;
  assign new_n6322 = ~pa0 & new_n6321;
  assign new_n6323 = ~pc0 & new_n6322;
  assign new_n6324 = ~ph & new_n5904;
  assign new_n6325 = ~pi & new_n6324;
  assign new_n6326 = ~pg & new_n6325;
  assign new_n6327 = ~pe & new_n6326;
  assign new_n6328 = ~pf & new_n6327;
  assign new_n6329 = ~pc0 & new_n6328;
  assign new_n6330 = pm0 & new_n6329;
  assign new_n6331 = ~pg & new_n5914;
  assign new_n6332 = ~pi & new_n6331;
  assign new_n6333 = ~pd0 & new_n6332;
  assign new_n6334 = ~pe & new_n6333;
  assign new_n6335 = ~pf & new_n6334;
  assign new_n6336 = ~ph0 & new_n6335;
  assign new_n6337 = pm0 & new_n6336;
  assign new_n6338 = ~pf0 & new_n6337;
  assign new_n6339 = ~pc0 & new_n6338;
  assign new_n6340 = ~pj0 & new_n6339;
  assign new_n6341 = ~pz & new_n6098;
  assign new_n6342 = ~pc & new_n6341;
  assign new_n6343 = ~pi0 & new_n6342;
  assign new_n6344 = ~pk & new_n6343;
  assign new_n6345 = ~ph & new_n6344;
  assign new_n6346 = ~pd0 & new_n6345;
  assign new_n6347 = ~pg & new_n6346;
  assign new_n6348 = ~pe & new_n6347;
  assign new_n6349 = ~pf & new_n6348;
  assign new_n6350 = pj0 & new_n6349;
  assign new_n6351 = pm0 & new_n6350;
  assign new_n6352 = ~ph & new_n5939;
  assign new_n6353 = ~pk & new_n6352;
  assign new_n6354 = ~pf & new_n6353;
  assign new_n6355 = ~pg & new_n6354;
  assign new_n6356 = ~pe & new_n6355;
  assign new_n6357 = pm0 & new_n6356;
  assign new_n6358 = ~ph0 & new_n6357;
  assign new_n6359 = ~pc0 & new_n6358;
  assign new_n6360 = ~pg0 & new_n6359;
  assign new_n6361 = ~pw & ~pn;
  assign new_n6362 = pj & new_n6361;
  assign new_n6363 = pl & new_n6362;
  assign new_n6364 = ~pc & new_n6363;
  assign new_n6365 = pm0 & new_n6364;
  assign new_n6366 = ~pd & new_n6365;
  assign new_n6367 = ~pg0 & new_n6366;
  assign new_n6368 = ~pj0 & new_n6367;
  assign new_n6369 = ~pe0 & new_n6368;
  assign new_n6370 = ~pa0 & new_n6369;
  assign new_n6371 = ~pc0 & new_n6370;
  assign new_n6372 = ~py & new_n6371;
  assign new_n6373 = ~pz & new_n6372;
  assign new_n6374 = pn & new_n5889;
  assign new_n6375 = ~pc & new_n6374;
  assign new_n6376 = ~pg & new_n6375;
  assign new_n6377 = ~ph & new_n6376;
  assign new_n6378 = ~pe & new_n6377;
  assign new_n6379 = ~pf & new_n6378;
  assign new_n6380 = ~ph0 & new_n6379;
  assign new_n6381 = ~pg0 & new_n6380;
  assign new_n6382 = pm0 & new_n6381;
  assign new_n6383 = ~pa0 & new_n6382;
  assign new_n6384 = ~pc0 & new_n6383;
  assign new_n6385 = ~py & new_n6097;
  assign new_n6386 = ~pz & new_n6385;
  assign new_n6387 = ~pc & new_n6386;
  assign new_n6388 = ~pm & new_n6387;
  assign new_n6389 = ~pd0 & new_n6388;
  assign new_n6390 = pi0 & new_n6389;
  assign new_n6391 = ~ph & new_n6390;
  assign new_n6392 = ~pf & new_n6391;
  assign new_n6393 = ~pg & new_n6392;
  assign new_n6394 = pm0 & new_n6393;
  assign new_n6395 = ~pe & new_n6394;
  assign new_n6396 = ~pe0 & ~pj0;
  assign new_n6397 = ~pz & new_n6396;
  assign new_n6398 = ~pc0 & new_n6397;
  assign new_n6399 = ~py & new_n6398;
  assign new_n6400 = pi0 & new_n6399;
  assign new_n6401 = ~pi & new_n6400;
  assign new_n6402 = ~pd0 & new_n6401;
  assign new_n6403 = pm0 & new_n6402;
  assign new_n6404 = ~pf0 & new_n6403;
  assign new_n6405 = ~pe0 & new_n6189;
  assign new_n6406 = pj0 & new_n6405;
  assign new_n6407 = ~pc0 & new_n6406;
  assign new_n6408 = ~pd0 & new_n6407;
  assign new_n6409 = ~pi0 & new_n6408;
  assign new_n6410 = ~ph & new_n6409;
  assign new_n6411 = ~pi & new_n6410;
  assign new_n6412 = ~pg & new_n5988;
  assign new_n6413 = ~pi & new_n6412;
  assign new_n6414 = ~pf & new_n6413;
  assign new_n6415 = ~ph0 & new_n6414;
  assign new_n6416 = ~pe & new_n6415;
  assign new_n6417 = ~pj0 & new_n6416;
  assign new_n6418 = pm0 & new_n6417;
  assign new_n6419 = ~pi & new_n5722;
  assign new_n6420 = pt & new_n6419;
  assign new_n6421 = ~pd0 & new_n6420;
  assign new_n6422 = ~pd & new_n6421;
  assign new_n6423 = ~pf & new_n6422;
  assign new_n6424 = ~pg & new_n6423;
  assign new_n6425 = ~pe & new_n6424;
  assign new_n6426 = ~pj0 & new_n6425;
  assign new_n6427 = pm0 & new_n6426;
  assign new_n6428 = ~pa0 & new_n6427;
  assign new_n6429 = ~pc0 & new_n6428;
  assign new_n6430 = pm0 & new_n6218;
  assign new_n6431 = ~pe & new_n6430;
  assign new_n6432 = ~pj0 & new_n6431;
  assign new_n6433 = ~pc0 & new_n6432;
  assign new_n6434 = ~pg0 & new_n6433;
  assign new_n6435 = ~pz & new_n6434;
  assign new_n6436 = ~pa0 & new_n6435;
  assign new_n6437 = pm0 & new_n6230;
  assign new_n6438 = ~ph0 & new_n6437;
  assign new_n6439 = ~pj0 & new_n6438;
  assign new_n6440 = ~pa0 & new_n6439;
  assign new_n6441 = ~pc0 & new_n6440;
  assign new_n6442 = ~pw & new_n6441;
  assign new_n6443 = ~py & new_n6442;
  assign new_n6444 = ~pi & new_n5766;
  assign new_n6445 = ~pd0 & new_n6444;
  assign new_n6446 = pi0 & new_n6445;
  assign new_n6447 = ~pb & new_n6446;
  assign new_n6448 = ~pf & new_n6447;
  assign new_n6449 = ~pg & new_n6448;
  assign new_n6450 = ~pe & new_n6449;
  assign new_n6451 = ~pj0 & new_n6450;
  assign new_n6452 = pm0 & new_n6451;
  assign new_n6453 = ~pz & new_n6452;
  assign new_n6454 = ~pc0 & new_n6453;
  assign new_n6455 = pm0 & new_n6252;
  assign new_n6456 = ~pe & new_n6455;
  assign new_n6457 = ~pj0 & new_n6456;
  assign new_n6458 = ~pc0 & new_n6457;
  assign new_n6459 = ~pg0 & new_n6458;
  assign new_n6460 = ~py & new_n6459;
  assign new_n6461 = ~pz & new_n6460;
  assign new_n6462 = ~ph0 & new_n6264;
  assign new_n6463 = ~pe & new_n6462;
  assign new_n6464 = pm0 & new_n6463;
  assign new_n6465 = ~pc0 & new_n6464;
  assign new_n6466 = ~pj0 & new_n6465;
  assign new_n6467 = ~py & new_n6466;
  assign new_n6468 = ~pa0 & new_n6467;
  assign new_n6469 = ~pi & new_n6046;
  assign new_n6470 = ~pd0 & new_n6469;
  assign new_n6471 = pi0 & new_n6470;
  assign new_n6472 = pd & new_n6471;
  assign new_n6473 = ~pf & new_n6472;
  assign new_n6474 = ~pg & new_n6473;
  assign new_n6475 = ~pe & new_n6474;
  assign new_n6476 = pm0 & new_n6475;
  assign new_n6477 = ~pf0 & new_n6476;
  assign new_n6478 = ~pc0 & new_n6477;
  assign new_n6479 = ~pj0 & new_n6478;
  assign new_n6480 = ~pf0 & new_n6286;
  assign new_n6481 = ~ph0 & new_n6480;
  assign new_n6482 = pm0 & new_n6481;
  assign new_n6483 = ~pg0 & new_n6482;
  assign new_n6484 = ~pj0 & new_n6483;
  assign new_n6485 = ~pa0 & new_n6484;
  assign new_n6486 = ~pc0 & new_n6485;
  assign new_n6487 = ~pb & new_n5853;
  assign new_n6488 = ~pk & new_n6487;
  assign new_n6489 = ~pi & new_n6488;
  assign new_n6490 = ~pd0 & new_n6489;
  assign new_n6491 = ~pg & new_n6490;
  assign new_n6492 = ~pe & new_n6491;
  assign new_n6493 = ~pf & new_n6492;
  assign new_n6494 = pm0 & new_n6493;
  assign new_n6495 = ~ph0 & new_n6494;
  assign new_n6496 = ~pd0 & new_n5824;
  assign new_n6497 = pi0 & new_n6496;
  assign new_n6498 = pd & new_n6497;
  assign new_n6499 = ~ph & new_n6498;
  assign new_n6500 = ~pi & new_n6499;
  assign new_n6501 = ~pg & new_n6500;
  assign new_n6502 = ~pe & new_n6501;
  assign new_n6503 = ~pf & new_n6502;
  assign new_n6504 = pm0 & new_n6503;
  assign new_n6505 = ~ph0 & new_n6504;
  assign new_n6506 = ~pc0 & new_n5897;
  assign new_n6507 = pm0 & new_n6506;
  assign new_n6508 = ~pz & new_n6507;
  assign new_n6509 = ~pa0 & new_n6508;
  assign new_n6510 = ~pt & new_n6059;
  assign new_n6511 = ~pd0 & new_n6510;
  assign new_n6512 = pi0 & new_n6511;
  assign new_n6513 = ~pg & new_n6512;
  assign new_n6514 = ~ph & new_n6513;
  assign new_n6515 = ~pf & new_n6514;
  assign new_n6516 = ~ph0 & new_n6515;
  assign new_n6517 = ~pe & new_n6516;
  assign new_n6518 = ~pg0 & new_n6517;
  assign new_n6519 = pm0 & new_n6518;
  assign new_n6520 = ~ph & new_n5838;
  assign new_n6521 = ~pt & new_n6520;
  assign new_n6522 = ~pd0 & new_n6521;
  assign new_n6523 = ~pf & new_n6522;
  assign new_n6524 = ~pg & new_n6523;
  assign new_n6525 = ~pe & new_n6524;
  assign new_n6526 = ~pg0 & new_n6525;
  assign new_n6527 = pm0 & new_n6526;
  assign new_n6528 = ~pa0 & new_n6527;
  assign new_n6529 = ~pc0 & new_n6528;
  assign new_n6530 = ~pj & new_n5969;
  assign new_n6531 = ~py & new_n6530;
  assign new_n6532 = ~pc & new_n6531;
  assign new_n6533 = pi0 & new_n6532;
  assign new_n6534 = ~pk & new_n6533;
  assign new_n6535 = ~pi & new_n6534;
  assign new_n6536 = ~pd0 & new_n6535;
  assign new_n6537 = ~ph & new_n6536;
  assign new_n6538 = ~pf & new_n6537;
  assign new_n6539 = ~pg & new_n6538;
  assign new_n6540 = ~ph0 & new_n6539;
  assign new_n6541 = ~pe & new_n6540;
  assign new_n6542 = ~pw & new_n5836;
  assign new_n6543 = ~pc & new_n6542;
  assign new_n6544 = ~pi & new_n6543;
  assign new_n6545 = ~pk & new_n6544;
  assign new_n6546 = ~pg & new_n6545;
  assign new_n6547 = ~ph & new_n6546;
  assign new_n6548 = ~pf & new_n6547;
  assign new_n6549 = pm0 & new_n6548;
  assign new_n6550 = ~pe & new_n6549;
  assign new_n6551 = ~pa0 & new_n6550;
  assign new_n6552 = ~pc0 & new_n6551;
  assign new_n6553 = pl & new_n5750;
  assign new_n6554 = ~pn & new_n6553;
  assign new_n6555 = pj & new_n6554;
  assign new_n6556 = ~pi & new_n6555;
  assign new_n6557 = pm & new_n6556;
  assign new_n6558 = ~pj0 & new_n6557;
  assign new_n6559 = pm0 & new_n6558;
  assign new_n6560 = ~pe0 & new_n6559;
  assign new_n6561 = ~pa0 & new_n6560;
  assign new_n6562 = ~pc0 & new_n6561;
  assign new_n6563 = ~py & new_n6562;
  assign new_n6564 = ~pz & new_n6563;
  assign new_n6565 = pm0 & new_n6379;
  assign new_n6566 = ~pc0 & new_n6565;
  assign new_n6567 = ~pg0 & new_n6566;
  assign new_n6568 = ~pz & new_n6567;
  assign new_n6569 = ~pa0 & new_n6568;
  assign new_n6570 = ~pg0 & pm0;
  assign new_n6571 = ~py & new_n6570;
  assign new_n6572 = ~pc0 & new_n6571;
  assign new_n6573 = ~pc & new_n6572;
  assign new_n6574 = ~pm & new_n6573;
  assign new_n6575 = ~pd0 & new_n6574;
  assign new_n6576 = pi0 & new_n6575;
  assign new_n6577 = ~ph & new_n6576;
  assign new_n6578 = ~pf & new_n6577;
  assign new_n6579 = ~pg & new_n6578;
  assign new_n6580 = ~ph0 & new_n6579;
  assign new_n6581 = ~pe & new_n6580;
  assign new_n6582 = ~pg0 & ~pj0;
  assign new_n6583 = ~pc0 & new_n6582;
  assign new_n6584 = ~pe0 & new_n6583;
  assign new_n6585 = ~py & new_n6584;
  assign new_n6586 = pi0 & new_n6585;
  assign new_n6587 = ~ph0 & new_n6586;
  assign new_n6588 = ~pd0 & new_n6587;
  assign new_n6589 = pm0 & new_n6588;
  assign new_n6590 = ~pf0 & new_n6589;
  assign new_n6591 = ~ph & new_n6170;
  assign new_n6592 = ~pg0 & new_n6591;
  assign new_n6593 = pm0 & new_n6592;
  assign new_n6594 = ~pc0 & new_n6593;
  assign new_n6595 = ~pe0 & new_n6594;
  assign new_n6596 = ~pi & new_n6203;
  assign new_n6597 = pt & new_n6596;
  assign new_n6598 = ~pd0 & new_n6597;
  assign new_n6599 = ~pd & new_n6598;
  assign new_n6600 = ~pf & new_n6599;
  assign new_n6601 = ~pg & new_n6600;
  assign new_n6602 = ~pe & new_n6601;
  assign new_n6603 = pm0 & new_n6602;
  assign new_n6604 = ~ph0 & new_n6603;
  assign new_n6605 = ~pc0 & new_n6604;
  assign new_n6606 = ~pj0 & new_n6605;
  assign new_n6607 = ~pf & new_n6226;
  assign new_n6608 = ~pg & new_n6607;
  assign new_n6609 = ~pi & new_n6608;
  assign new_n6610 = ~pd0 & new_n6609;
  assign new_n6611 = ~ph0 & new_n6610;
  assign new_n6612 = ~pe & new_n6611;
  assign new_n6613 = pm0 & new_n6612;
  assign new_n6614 = ~pc0 & new_n6613;
  assign new_n6615 = ~pj0 & new_n6614;
  assign new_n6616 = ~py & new_n6615;
  assign new_n6617 = ~pa0 & new_n6616;
  assign new_n6618 = pm0 & new_n6226;
  assign new_n6619 = ~pe & new_n6618;
  assign new_n6620 = ~pf & new_n6619;
  assign new_n6621 = ~pg & new_n6620;
  assign new_n6622 = ~pg0 & new_n6621;
  assign new_n6623 = ~pj0 & new_n6622;
  assign new_n6624 = ~pc0 & new_n6623;
  assign new_n6625 = ~pz & new_n6624;
  assign new_n6626 = ~pa0 & new_n6625;
  assign new_n6627 = ~pw & new_n6626;
  assign new_n6628 = ~py & new_n6627;
  assign new_n6629 = ~pd & new_n6202;
  assign new_n6630 = ~pg & new_n6629;
  assign new_n6631 = pt & new_n6630;
  assign new_n6632 = ~pd0 & new_n6631;
  assign new_n6633 = ~pb & new_n6632;
  assign new_n6634 = ~pe & new_n6633;
  assign new_n6635 = ~pf & new_n6634;
  assign new_n6636 = ~ph0 & new_n6635;
  assign new_n6637 = ~pj0 & new_n6636;
  assign new_n6638 = pm0 & new_n6637;
  assign new_n6639 = ~pc0 & new_n6638;
  assign new_n6640 = ~pg0 & new_n6639;
  assign new_n6641 = ~pd & new_n6364;
  assign new_n6642 = ~pf & new_n6641;
  assign new_n6643 = ~pg & new_n6642;
  assign new_n6644 = ~pi & new_n6643;
  assign new_n6645 = ~pb & new_n6644;
  assign new_n6646 = pm0 & new_n6645;
  assign new_n6647 = ~pe & new_n6646;
  assign new_n6648 = ~pj0 & new_n6647;
  assign new_n6649 = ~pa0 & new_n6648;
  assign new_n6650 = ~pc0 & new_n6649;
  assign new_n6651 = ~py & new_n6650;
  assign new_n6652 = ~pz & new_n6651;
  assign new_n6653 = ~pb & new_n6010;
  assign new_n6654 = ~pf & new_n6653;
  assign new_n6655 = ~pg & new_n6654;
  assign new_n6656 = pt & new_n6655;
  assign new_n6657 = ~pd0 & new_n6656;
  assign new_n6658 = pm0 & new_n6657;
  assign new_n6659 = ~pe & new_n6658;
  assign new_n6660 = ~pj0 & new_n6659;
  assign new_n6661 = ~pc0 & new_n6660;
  assign new_n6662 = ~pg0 & new_n6661;
  assign new_n6663 = ~pz & new_n6662;
  assign new_n6664 = ~pa0 & new_n6663;
  assign new_n6665 = ~ph0 & new_n5798;
  assign new_n6666 = ~pe & new_n6665;
  assign new_n6667 = ~pf & new_n6666;
  assign new_n6668 = ~pg & new_n6667;
  assign new_n6669 = ~pj0 & new_n6668;
  assign new_n6670 = pm0 & new_n6669;
  assign new_n6671 = ~pg0 & new_n6670;
  assign new_n6672 = ~pa0 & new_n6671;
  assign new_n6673 = ~pc0 & new_n6672;
  assign new_n6674 = ~pw & new_n6673;
  assign new_n6675 = ~py & new_n6674;
  assign new_n6676 = ~pf & new_n5891;
  assign new_n6677 = ~pg & new_n6676;
  assign new_n6678 = ~pi & new_n6677;
  assign new_n6679 = pd & new_n6678;
  assign new_n6680 = ~pf0 & new_n6679;
  assign new_n6681 = ~pe & new_n6680;
  assign new_n6682 = pm0 & new_n6681;
  assign new_n6683 = ~pc0 & new_n6682;
  assign new_n6684 = ~pj0 & new_n6683;
  assign new_n6685 = ~pz & new_n6684;
  assign new_n6686 = ~pa0 & new_n6685;
  assign new_n6687 = ~pb & new_n6074;
  assign new_n6688 = ~pk & new_n6687;
  assign new_n6689 = ~pi & new_n6688;
  assign new_n6690 = ~pd0 & new_n6689;
  assign new_n6691 = ~pg & new_n6690;
  assign new_n6692 = ~pe & new_n6691;
  assign new_n6693 = ~pf & new_n6692;
  assign new_n6694 = ~pj0 & new_n6693;
  assign new_n6695 = pm0 & new_n6694;
  assign new_n6696 = ~pj & new_n1763;
  assign new_n6697 = ~py & new_n6696;
  assign new_n6698 = ~pc & new_n6697;
  assign new_n6699 = ~pd0 & new_n6698;
  assign new_n6700 = pi0 & new_n6699;
  assign new_n6701 = ~pk & new_n6700;
  assign new_n6702 = ~pg & new_n6701;
  assign new_n6703 = ~pi & new_n6702;
  assign new_n6704 = ~pf & new_n6703;
  assign new_n6705 = ~ph0 & new_n6704;
  assign new_n6706 = ~pe & new_n6705;
  assign new_n6707 = pm0 & new_n6706;
  assign new_n6708 = ~pf0 & new_n6707;
  assign new_n6709 = ~pf & new_n6543;
  assign new_n6710 = ~pg & new_n6709;
  assign new_n6711 = ~pk & new_n6710;
  assign new_n6712 = ~pf0 & new_n6711;
  assign new_n6713 = ~pe & new_n6712;
  assign new_n6714 = pm0 & new_n6713;
  assign new_n6715 = ~pg0 & new_n6714;
  assign new_n6716 = ~pj0 & new_n6715;
  assign new_n6717 = ~pa0 & new_n6716;
  assign new_n6718 = ~pc0 & new_n6717;
  assign new_n6719 = ps & new_n3448;
  assign new_n6720 = ~pw & new_n6719;
  assign new_n6721 = ~pn & new_n6720;
  assign new_n6722 = pt & new_n6721;
  assign new_n6723 = pm & new_n6722;
  assign new_n6724 = pk & new_n6723;
  assign new_n6725 = ~pf0 & new_n6724;
  assign new_n6726 = ~ph0 & new_n6725;
  assign new_n6727 = pm0 & new_n6726;
  assign new_n6728 = ~pg0 & new_n6727;
  assign new_n6729 = ~pj0 & new_n6728;
  assign new_n6730 = ~pc0 & new_n6729;
  assign new_n6731 = ~pe0 & new_n6730;
  assign new_n6732 = ~py & new_n5876;
  assign new_n6733 = ~pc & new_n6732;
  assign new_n6734 = pi0 & new_n6733;
  assign new_n6735 = ~pk & new_n6734;
  assign new_n6736 = ~pi & new_n6735;
  assign new_n6737 = ~pd0 & new_n6736;
  assign new_n6738 = ~ph & new_n6737;
  assign new_n6739 = ~pf & new_n6738;
  assign new_n6740 = ~pg & new_n6739;
  assign new_n6741 = pm0 & new_n6740;
  assign new_n6742 = ~pe & new_n6741;
  assign new_n6743 = ~pa0 & ~pc0;
  assign new_n6744 = ~pw & new_n6743;
  assign new_n6745 = ~py & new_n6744;
  assign new_n6746 = ~pn & new_n6745;
  assign new_n6747 = pm & new_n6746;
  assign new_n6748 = pk & new_n6747;
  assign new_n6749 = pt & new_n6748;
  assign new_n6750 = ~pd & new_n6749;
  assign new_n6751 = ~pi & new_n6750;
  assign new_n6752 = ~ph0 & new_n6751;
  assign new_n6753 = ~ph & new_n6752;
  assign new_n6754 = ~pe0 & new_n6753;
  assign new_n6755 = pm0 & new_n6754;
  assign new_n6756 = ~pn & new_n5718;
  assign new_n6757 = ~pw & new_n6756;
  assign new_n6758 = pj & new_n6757;
  assign new_n6759 = ~pd & new_n6758;
  assign new_n6760 = pm & new_n6759;
  assign new_n6761 = pm0 & new_n6760;
  assign new_n6762 = pt & new_n6761;
  assign new_n6763 = ~pj0 & new_n6762;
  assign new_n6764 = ~pe0 & new_n6763;
  assign new_n6765 = ~pg0 & new_n6764;
  assign new_n6766 = ~pa0 & new_n6765;
  assign new_n6767 = ~pc0 & new_n6766;
  assign new_n6768 = ~ph0 & new_n6180;
  assign new_n6769 = ~pg0 & new_n6768;
  assign new_n6770 = ~pj0 & new_n6769;
  assign new_n6771 = ~pe0 & new_n6770;
  assign new_n6772 = ~pa0 & new_n6771;
  assign new_n6773 = ~pc0 & new_n6772;
  assign new_n6774 = ~pw & new_n6773;
  assign new_n6775 = ~py & new_n6774;
  assign new_n6776 = ~py & new_n6743;
  assign new_n6777 = ~pz & new_n6776;
  assign new_n6778 = ~pc & new_n6777;
  assign new_n6779 = ~pm & new_n6778;
  assign new_n6780 = ~pi & new_n6779;
  assign new_n6781 = ~pd0 & new_n6780;
  assign new_n6782 = ~ph & new_n6781;
  assign new_n6783 = ~pf & new_n6782;
  assign new_n6784 = ~pg & new_n6783;
  assign new_n6785 = pm0 & new_n6784;
  assign new_n6786 = ~pe & new_n6785;
  assign new_n6787 = ~pe0 & ~pg0;
  assign new_n6788 = ~pz & new_n6787;
  assign new_n6789 = ~pc0 & new_n6788;
  assign new_n6790 = ~py & new_n6789;
  assign new_n6791 = pi0 & new_n6790;
  assign new_n6792 = ~pf0 & new_n6791;
  assign new_n6793 = ~pd0 & new_n6792;
  assign new_n6794 = ~pj0 & new_n6793;
  assign new_n6795 = pm0 & new_n6794;
  assign new_n6796 = pj0 & pm0;
  assign new_n6797 = ~pe0 & new_n6796;
  assign new_n6798 = ~pg0 & new_n6797;
  assign new_n6799 = ~pc0 & new_n6798;
  assign new_n6800 = ~pd0 & new_n6799;
  assign new_n6801 = ~pi0 & new_n6800;
  assign new_n6802 = ~ph0 & new_n6801;
  assign new_n6803 = ~ph & new_n6802;
  assign new_n6804 = ~pd0 & new_n5739;
  assign new_n6805 = pi0 & new_n6804;
  assign new_n6806 = ~pd & new_n6805;
  assign new_n6807 = ~pe & new_n6806;
  assign new_n6808 = ~pf & new_n6807;
  assign new_n6809 = pm0 & new_n6808;
  assign new_n6810 = ~pg0 & new_n6809;
  assign new_n6811 = ~pj0 & new_n6810;
  assign new_n6812 = ~pz & new_n6811;
  assign new_n6813 = ~pc0 & new_n6812;
  assign new_n6814 = pm0 & new_n6610;
  assign new_n6815 = ~pe & new_n6814;
  assign new_n6816 = ~pj0 & new_n6815;
  assign new_n6817 = ~pa0 & new_n6816;
  assign new_n6818 = ~pc0 & new_n6817;
  assign new_n6819 = ~py & new_n6818;
  assign new_n6820 = ~pz & new_n6819;
  assign new_n6821 = ~ph0 & new_n6226;
  assign new_n6822 = ~pe & new_n6821;
  assign new_n6823 = ~pf & new_n6822;
  assign new_n6824 = ~pg & new_n6823;
  assign new_n6825 = ~pj0 & new_n6824;
  assign new_n6826 = pm0 & new_n6825;
  assign new_n6827 = ~pg0 & new_n6826;
  assign new_n6828 = ~pa0 & new_n6827;
  assign new_n6829 = ~pc0 & new_n6828;
  assign new_n6830 = ~pw & new_n6829;
  assign new_n6831 = ~py & new_n6830;
  assign new_n6832 = ~pd & new_n5721;
  assign new_n6833 = ~pg & new_n6832;
  assign new_n6834 = pt & new_n6833;
  assign new_n6835 = ~pd0 & new_n6834;
  assign new_n6836 = ~pb & new_n6835;
  assign new_n6837 = ~pe & new_n6836;
  assign new_n6838 = ~pf & new_n6837;
  assign new_n6839 = pm0 & new_n6838;
  assign new_n6840 = ~pg0 & new_n6839;
  assign new_n6841 = ~pj0 & new_n6840;
  assign new_n6842 = ~pa0 & new_n6841;
  assign new_n6843 = ~pc0 & new_n6842;
  assign new_n6844 = ~ph0 & new_n6645;
  assign new_n6845 = ~pe & new_n6844;
  assign new_n6846 = pm0 & new_n6845;
  assign new_n6847 = ~pc0 & new_n6846;
  assign new_n6848 = ~pj0 & new_n6847;
  assign new_n6849 = ~py & new_n6848;
  assign new_n6850 = ~pa0 & new_n6849;
  assign new_n6851 = ~pi & new_n6653;
  assign new_n6852 = pt & new_n6851;
  assign new_n6853 = ~pd0 & new_n6852;
  assign new_n6854 = pi0 & new_n6853;
  assign new_n6855 = ~pf & new_n6854;
  assign new_n6856 = ~pg & new_n6855;
  assign new_n6857 = ~pe & new_n6856;
  assign new_n6858 = ~pj0 & new_n6857;
  assign new_n6859 = pm0 & new_n6858;
  assign new_n6860 = ~pz & new_n6859;
  assign new_n6861 = ~pc0 & new_n6860;
  assign new_n6862 = pm0 & new_n5798;
  assign new_n6863 = ~pe & new_n6862;
  assign new_n6864 = ~pf & new_n6863;
  assign new_n6865 = ~pg & new_n6864;
  assign new_n6866 = ~pg0 & new_n6865;
  assign new_n6867 = ~pj0 & new_n6866;
  assign new_n6868 = ~pc0 & new_n6867;
  assign new_n6869 = ~pz & new_n6868;
  assign new_n6870 = ~pa0 & new_n6869;
  assign new_n6871 = ~pw & new_n6870;
  assign new_n6872 = ~py & new_n6871;
  assign new_n6873 = ~ph0 & new_n6679;
  assign new_n6874 = ~pe & new_n6873;
  assign new_n6875 = ~pf0 & new_n6874;
  assign new_n6876 = ~pj0 & new_n6875;
  assign new_n6877 = pm0 & new_n6876;
  assign new_n6878 = ~pa0 & new_n6877;
  assign new_n6879 = ~pc0 & new_n6878;
  assign new_n6880 = ~pb & new_n6297;
  assign new_n6881 = ~pk & new_n6880;
  assign new_n6882 = ~pg & new_n6881;
  assign new_n6883 = ~pd0 & new_n6882;
  assign new_n6884 = ~pf & new_n6883;
  assign new_n6885 = ~ph0 & new_n6884;
  assign new_n6886 = ~pe & new_n6885;
  assign new_n6887 = ~pj0 & new_n6886;
  assign new_n6888 = pm0 & new_n6887;
  assign new_n6889 = ~pb & new_n5865;
  assign new_n6890 = ~pk & new_n6889;
  assign new_n6891 = ~pe & new_n6890;
  assign new_n6892 = ~pf & new_n6891;
  assign new_n6893 = pm0 & new_n6892;
  assign new_n6894 = ~pg0 & new_n6893;
  assign new_n6895 = ~pj0 & new_n6894;
  assign new_n6896 = ~pa0 & new_n6895;
  assign new_n6897 = ~pc0 & new_n6896;
  assign new_n6898 = ~pd & new_n6746;
  assign new_n6899 = pm & new_n6898;
  assign new_n6900 = pk & new_n6899;
  assign new_n6901 = ~pi & new_n6900;
  assign new_n6902 = pt & new_n6901;
  assign new_n6903 = ~ph0 & new_n6902;
  assign new_n6904 = pm0 & new_n6903;
  assign new_n6905 = ~pf0 & new_n6904;
  assign new_n6906 = ~pe0 & new_n6905;
  assign new_n6907 = ~pj0 & new_n6906;
  assign new_n6908 = ps & new_n5718;
  assign new_n6909 = ~pw & new_n6908;
  assign new_n6910 = ~pn & new_n6909;
  assign new_n6911 = pt & new_n6910;
  assign new_n6912 = pm & new_n6911;
  assign new_n6913 = pk & new_n6912;
  assign new_n6914 = ~pf0 & new_n6913;
  assign new_n6915 = ~pi & new_n6914;
  assign new_n6916 = pm0 & new_n6915;
  assign new_n6917 = ~pe0 & new_n6916;
  assign new_n6918 = ~pj0 & new_n6917;
  assign new_n6919 = ~pa0 & new_n6918;
  assign new_n6920 = ~pc0 & new_n6919;
  assign new_n6921 = ~py & new_n6098;
  assign new_n6922 = ~pc & new_n6921;
  assign new_n6923 = pi0 & new_n6922;
  assign new_n6924 = ~pk & new_n6923;
  assign new_n6925 = ~ph & new_n6924;
  assign new_n6926 = ~pd0 & new_n6925;
  assign new_n6927 = ~pg & new_n6926;
  assign new_n6928 = ~pe & new_n6927;
  assign new_n6929 = ~pf & new_n6928;
  assign new_n6930 = pm0 & new_n6929;
  assign new_n6931 = ~ph0 & new_n6930;
  assign new_n6932 = ~ph & new_n6543;
  assign new_n6933 = ~pk & new_n6932;
  assign new_n6934 = ~pf & new_n6933;
  assign new_n6935 = ~pg & new_n6934;
  assign new_n6936 = ~pe & new_n6935;
  assign new_n6937 = ~pg0 & new_n6936;
  assign new_n6938 = pm0 & new_n6937;
  assign new_n6939 = ~pa0 & new_n6938;
  assign new_n6940 = ~pc0 & new_n6939;
  assign new_n6941 = ~pd0 & new_n6778;
  assign new_n6942 = ~pm & new_n6941;
  assign new_n6943 = ~pg & new_n6942;
  assign new_n6944 = ~pi & new_n6943;
  assign new_n6945 = ~pf & new_n6944;
  assign new_n6946 = ~pf0 & new_n6945;
  assign new_n6947 = ~pe & new_n6946;
  assign new_n6948 = ~pj0 & new_n6947;
  assign new_n6949 = pm0 & new_n6948;
  assign new_n6950 = ~pj0 & new_n5797;
  assign new_n6951 = pm0 & new_n6950;
  assign new_n6952 = ~pe0 & new_n6951;
  assign new_n6953 = ~pg0 & new_n6952;
  assign new_n6954 = ~pc0 & new_n6953;
  assign new_n6955 = ~pz & new_n6954;
  assign new_n6956 = ~pa0 & new_n6955;
  assign new_n6957 = ~pw & new_n6956;
  assign new_n6958 = ~py & new_n6957;
  assign new_n6959 = ~pa0 & new_n5970;
  assign new_n6960 = ~pc & new_n6959;
  assign new_n6961 = ~pm & new_n6960;
  assign new_n6962 = ~pi & new_n6961;
  assign new_n6963 = ~pd0 & new_n6962;
  assign new_n6964 = ~ph & new_n6963;
  assign new_n6965 = ~pf & new_n6964;
  assign new_n6966 = ~pg & new_n6965;
  assign new_n6967 = ~ph0 & new_n6966;
  assign new_n6968 = ~pe & new_n6967;
  assign new_n6969 = ~pa0 & new_n6396;
  assign new_n6970 = ~pc0 & new_n6969;
  assign new_n6971 = ~py & new_n6970;
  assign new_n6972 = ~pd0 & new_n6971;
  assign new_n6973 = ~ph0 & new_n6972;
  assign new_n6974 = ~pi & new_n6973;
  assign new_n6975 = pm0 & new_n6974;
  assign new_n6976 = ~pf0 & new_n6975;
  assign new_n6977 = ~pc0 & new_n6796;
  assign new_n6978 = ~pe0 & new_n6977;
  assign new_n6979 = ~pz & new_n6978;
  assign new_n6980 = ~pd0 & new_n6979;
  assign new_n6981 = ~pi0 & new_n6980;
  assign new_n6982 = ~ph & new_n6981;
  assign new_n6983 = ~pi & new_n6982;
  assign new_n6984 = ~ph0 & new_n6808;
  assign new_n6985 = ~pj0 & new_n6984;
  assign new_n6986 = pm0 & new_n6985;
  assign new_n6987 = ~pc0 & new_n6986;
  assign new_n6988 = ~pg0 & new_n6987;
  assign new_n6989 = ~pd0 & new_n6229;
  assign new_n6990 = pm0 & new_n6989;
  assign new_n6991 = ~ph0 & new_n6990;
  assign new_n6992 = ~pj0 & new_n6991;
  assign new_n6993 = ~pc0 & new_n6992;
  assign new_n6994 = ~pg0 & new_n6993;
  assign new_n6995 = ~py & new_n6994;
  assign new_n6996 = ~pa0 & new_n6995;
  assign new_n6997 = pt & new_n6832;
  assign new_n6998 = ~pd0 & new_n6997;
  assign new_n6999 = pi0 & new_n6998;
  assign new_n7000 = ~pb & new_n6999;
  assign new_n7001 = ~pg & new_n7000;
  assign new_n7002 = ~pi & new_n7001;
  assign new_n7003 = ~pf & new_n7002;
  assign new_n7004 = pm0 & new_n7003;
  assign new_n7005 = ~pe & new_n7004;
  assign new_n7006 = ~pc0 & new_n7005;
  assign new_n7007 = ~pj0 & new_n7006;
  assign new_n7008 = ~pi & new_n6629;
  assign new_n7009 = pt & new_n7008;
  assign new_n7010 = ~pd0 & new_n7009;
  assign new_n7011 = ~pb & new_n7010;
  assign new_n7012 = ~pf & new_n7011;
  assign new_n7013 = ~pg & new_n7012;
  assign new_n7014 = ~pe & new_n7013;
  assign new_n7015 = pm0 & new_n7014;
  assign new_n7016 = ~ph0 & new_n7015;
  assign new_n7017 = ~pc0 & new_n7016;
  assign new_n7018 = ~pj0 & new_n7017;
  assign new_n7019 = ~pf & new_n5782;
  assign new_n7020 = ~pg & new_n7019;
  assign new_n7021 = pt & new_n7020;
  assign new_n7022 = ~pb & new_n7021;
  assign new_n7023 = pm0 & new_n7022;
  assign new_n7024 = ~pe & new_n7023;
  assign new_n7025 = ~pj0 & new_n7024;
  assign new_n7026 = ~pc0 & new_n7025;
  assign new_n7027 = ~pg0 & new_n7026;
  assign new_n7028 = ~pz & new_n7027;
  assign new_n7029 = ~pa0 & new_n7028;
  assign new_n7030 = ~pg & new_n6653;
  assign new_n7031 = pt & new_n7030;
  assign new_n7032 = ~pd0 & new_n7031;
  assign new_n7033 = pi0 & new_n7032;
  assign new_n7034 = ~pe & new_n7033;
  assign new_n7035 = ~pf & new_n7034;
  assign new_n7036 = ~ph0 & new_n7035;
  assign new_n7037 = ~pj0 & new_n7036;
  assign new_n7038 = pm0 & new_n7037;
  assign new_n7039 = ~pc0 & new_n7038;
  assign new_n7040 = ~pg0 & new_n7039;
  assign new_n7041 = ~pi & new_n6250;
  assign new_n7042 = ~pd0 & new_n7041;
  assign new_n7043 = pm0 & new_n7042;
  assign new_n7044 = ~pe & new_n7043;
  assign new_n7045 = ~pj0 & new_n7044;
  assign new_n7046 = ~pa0 & new_n7045;
  assign new_n7047 = ~pc0 & new_n7046;
  assign new_n7048 = ~py & new_n7047;
  assign new_n7049 = ~pz & new_n7048;
  assign new_n7050 = ~pf & new_n6046;
  assign new_n7051 = ~pg & new_n7050;
  assign new_n7052 = ~pd0 & new_n7051;
  assign new_n7053 = pd & new_n7052;
  assign new_n7054 = ~pf0 & new_n7053;
  assign new_n7055 = ~pe & new_n7054;
  assign new_n7056 = pm0 & new_n7055;
  assign new_n7057 = ~pg0 & new_n7056;
  assign new_n7058 = ~pj0 & new_n7057;
  assign new_n7059 = ~pa0 & new_n7058;
  assign new_n7060 = ~pc0 & new_n7059;
  assign new_n7061 = ~pg & new_n6688;
  assign new_n7062 = ~pd0 & new_n7061;
  assign new_n7063 = ~pf & new_n7062;
  assign new_n7064 = pm0 & new_n7063;
  assign new_n7065 = ~pe & new_n7064;
  assign new_n7066 = ~pg0 & new_n7065;
  assign new_n7067 = ~pj0 & new_n7066;
  assign new_n7068 = ~pd0 & new_n6922;
  assign new_n7069 = pi0 & new_n7068;
  assign new_n7070 = ~pk & new_n7069;
  assign new_n7071 = ~pf & new_n7070;
  assign new_n7072 = ~pg & new_n7071;
  assign new_n7073 = ~pe & new_n7072;
  assign new_n7074 = ~pf0 & new_n7073;
  assign new_n7075 = ~ph0 & new_n7074;
  assign new_n7076 = ~pj0 & new_n7075;
  assign new_n7077 = pm0 & new_n7076;
  assign new_n7078 = ~pg & new_n6543;
  assign new_n7079 = ~pi & new_n7078;
  assign new_n7080 = ~pk & new_n7079;
  assign new_n7081 = ~pe & new_n7080;
  assign new_n7082 = ~pf & new_n7081;
  assign new_n7083 = ~pf0 & new_n7082;
  assign new_n7084 = ~pj0 & new_n7083;
  assign new_n7085 = pm0 & new_n7084;
  assign new_n7086 = ~pa0 & new_n7085;
  assign new_n7087 = ~pc0 & new_n7086;
  assign new_n7088 = ~ph0 & new_n6724;
  assign new_n7089 = ~pi & new_n7088;
  assign new_n7090 = ~pf0 & new_n7089;
  assign new_n7091 = ~pj0 & new_n7090;
  assign new_n7092 = pm0 & new_n7091;
  assign new_n7093 = ~pc0 & new_n7092;
  assign new_n7094 = ~pe0 & new_n7093;
  assign new_n7095 = pm & new_n6910;
  assign new_n7096 = pk & new_n7095;
  assign new_n7097 = ~ph & new_n7096;
  assign new_n7098 = pt & new_n7097;
  assign new_n7099 = pm0 & new_n7098;
  assign new_n7100 = ~pe0 & new_n7099;
  assign new_n7101 = ~pg0 & new_n7100;
  assign new_n7102 = ~pa0 & new_n7101;
  assign new_n7103 = ~pc0 & new_n7102;
  assign new_n7104 = ~pc0 & new_n6189;
  assign new_n7105 = pj0 & new_n7104;
  assign new_n7106 = ~pc & new_n7105;
  assign new_n7107 = ~pm & new_n7106;
  assign new_n7108 = ~pd0 & new_n7107;
  assign new_n7109 = ~pi0 & new_n7108;
  assign new_n7110 = ~pi & new_n7109;
  assign new_n7111 = ~pg & new_n7110;
  assign new_n7112 = ~ph & new_n7111;
  assign new_n7113 = ~pe & new_n7112;
  assign new_n7114 = ~pf & new_n7113;
  assign new_n7115 = ~ph & new_n6779;
  assign new_n7116 = ~pd0 & new_n7115;
  assign new_n7117 = ~pg & new_n7116;
  assign new_n7118 = ~pe & new_n7117;
  assign new_n7119 = ~pf & new_n7118;
  assign new_n7120 = ~pg0 & new_n7119;
  assign new_n7121 = pm0 & new_n7120;
  assign new_n7122 = ~pc0 & ~pe0;
  assign new_n7123 = ~pz & new_n7122;
  assign new_n7124 = ~pa0 & new_n7123;
  assign new_n7125 = ~py & new_n7124;
  assign new_n7126 = ~pd0 & new_n7125;
  assign new_n7127 = ~pf0 & new_n7126;
  assign new_n7128 = ~pi & new_n7127;
  assign new_n7129 = ~pj0 & new_n7128;
  assign new_n7130 = pm0 & new_n7129;
  assign new_n7131 = ~pe0 & new_n7104;
  assign new_n7132 = ~py & new_n7131;
  assign new_n7133 = ~pd0 & new_n7132;
  assign new_n7134 = pi0 & new_n7133;
  assign new_n7135 = ~ph & new_n7134;
  assign new_n7136 = ~pi & new_n7135;
  assign new_n7137 = ~pi & new_n5738;
  assign new_n7138 = ~pd0 & new_n7137;
  assign new_n7139 = pi0 & new_n7138;
  assign new_n7140 = ~pd & new_n7139;
  assign new_n7141 = ~pf & new_n7140;
  assign new_n7142 = ~pg & new_n7141;
  assign new_n7143 = ~pe & new_n7142;
  assign new_n7144 = ~pj0 & new_n7143;
  assign new_n7145 = pm0 & new_n7144;
  assign new_n7146 = ~pz & new_n7145;
  assign new_n7147 = ~pc0 & new_n7146;
  assign new_n7148 = ~pj0 & new_n6989;
  assign new_n7149 = pm0 & new_n7148;
  assign new_n7150 = ~pg0 & new_n7149;
  assign new_n7151 = ~pa0 & new_n7150;
  assign new_n7152 = ~pc0 & new_n7151;
  assign new_n7153 = ~py & new_n7152;
  assign new_n7154 = ~pz & new_n7153;
  assign new_n7155 = ~pd & new_n5983;
  assign new_n7156 = pt & new_n7155;
  assign new_n7157 = ~pd0 & new_n7156;
  assign new_n7158 = pi0 & new_n7157;
  assign new_n7159 = ~pb & new_n7158;
  assign new_n7160 = ~pg & new_n7159;
  assign new_n7161 = ~pi & new_n7160;
  assign new_n7162 = ~pf & new_n7161;
  assign new_n7163 = ~ph0 & new_n7162;
  assign new_n7164 = ~pe & new_n7163;
  assign new_n7165 = ~pj0 & new_n7164;
  assign new_n7166 = pm0 & new_n7165;
  assign new_n7167 = ~pi & new_n6832;
  assign new_n7168 = pt & new_n7167;
  assign new_n7169 = ~pd0 & new_n7168;
  assign new_n7170 = ~pb & new_n7169;
  assign new_n7171 = ~pf & new_n7170;
  assign new_n7172 = ~pg & new_n7171;
  assign new_n7173 = ~pe & new_n7172;
  assign new_n7174 = ~pj0 & new_n7173;
  assign new_n7175 = pm0 & new_n7174;
  assign new_n7176 = ~pa0 & new_n7175;
  assign new_n7177 = ~pc0 & new_n7176;
  assign new_n7178 = ~ph0 & new_n7022;
  assign new_n7179 = ~pe & new_n7178;
  assign new_n7180 = pm0 & new_n7179;
  assign new_n7181 = ~pg0 & new_n7180;
  assign new_n7182 = ~pj0 & new_n7181;
  assign new_n7183 = ~pa0 & new_n7182;
  assign new_n7184 = ~pc0 & new_n7183;
  assign new_n7185 = pm0 & new_n7035;
  assign new_n7186 = ~pg0 & new_n7185;
  assign new_n7187 = ~pj0 & new_n7186;
  assign new_n7188 = ~pz & new_n7187;
  assign new_n7189 = ~pc0 & new_n7188;
  assign new_n7190 = ~ph0 & new_n7042;
  assign new_n7191 = ~pe & new_n7190;
  assign new_n7192 = pm0 & new_n7191;
  assign new_n7193 = ~pc0 & new_n7192;
  assign new_n7194 = ~pj0 & new_n7193;
  assign new_n7195 = ~py & new_n7194;
  assign new_n7196 = ~pa0 & new_n7195;
  assign new_n7197 = ~pi & new_n5812;
  assign new_n7198 = ~pj0 & new_n7197;
  assign new_n7199 = pm0 & new_n7198;
  assign new_n7200 = ~pc0 & new_n7199;
  assign new_n7201 = ~pz & new_n7200;
  assign new_n7202 = ~pa0 & new_n7201;
  assign new_n7203 = ~pw & new_n7202;
  assign new_n7204 = ~py & new_n7203;
  assign new_n7205 = pj & new_n6743;
  assign new_n7206 = ~py & new_n7205;
  assign new_n7207 = ~pc & new_n7206;
  assign new_n7208 = ~pd0 & new_n7207;
  assign new_n7209 = ~pb & new_n7208;
  assign new_n7210 = ~pk & new_n7209;
  assign new_n7211 = ~pg & new_n7210;
  assign new_n7212 = ~pi & new_n7211;
  assign new_n7213 = ~pf & new_n7212;
  assign new_n7214 = ~ph0 & new_n7213;
  assign new_n7215 = ~pe & new_n7214;
  assign new_n7216 = ~pj0 & new_n7215;
  assign new_n7217 = pm0 & new_n7216;
  assign new_n7218 = ~pd0 & new_n6733;
  assign new_n7219 = pi0 & new_n7218;
  assign new_n7220 = ~pk & new_n7219;
  assign new_n7221 = ~pg & new_n7220;
  assign new_n7222 = ~pi & new_n7221;
  assign new_n7223 = ~pf & new_n7222;
  assign new_n7224 = ~pf0 & new_n7223;
  assign new_n7225 = ~pe & new_n7224;
  assign new_n7226 = ~pj0 & new_n7225;
  assign new_n7227 = pm0 & new_n7226;
  assign new_n7228 = ~pf & new_n5939;
  assign new_n7229 = ~pg & new_n7228;
  assign new_n7230 = ~pk & new_n7229;
  assign new_n7231 = ~ph0 & new_n7230;
  assign new_n7232 = ~pe & new_n7231;
  assign new_n7233 = ~pf0 & new_n7232;
  assign new_n7234 = ~pj0 & new_n7233;
  assign new_n7235 = pm0 & new_n7234;
  assign new_n7236 = ~pc0 & new_n7235;
  assign new_n7237 = ~pg0 & new_n7236;
  assign new_n7238 = pl & new_n6757;
  assign new_n7239 = ~pd & new_n7238;
  assign new_n7240 = pm & new_n7239;
  assign new_n7241 = pk & new_n7240;
  assign new_n7242 = pm0 & new_n7241;
  assign new_n7243 = ~pf0 & new_n7242;
  assign new_n7244 = ~pj0 & new_n7243;
  assign new_n7245 = ~pe0 & new_n7244;
  assign new_n7246 = ~pg0 & new_n7245;
  assign new_n7247 = ~pa0 & new_n7246;
  assign new_n7248 = ~pc0 & new_n7247;
  assign new_n7249 = ~pn & new_n6169;
  assign new_n7250 = pm & new_n7249;
  assign new_n7251 = pk & new_n7250;
  assign new_n7252 = pt & new_n7251;
  assign new_n7253 = ~pd & new_n7252;
  assign new_n7254 = ~pi & new_n7253;
  assign new_n7255 = pm0 & new_n7254;
  assign new_n7256 = ~ph & new_n7255;
  assign new_n7257 = ~pc0 & new_n7256;
  assign new_n7258 = ~pe0 & new_n7257;
  assign new_n7259 = ~pz & new_n6796;
  assign new_n7260 = ~pc0 & new_n7259;
  assign new_n7261 = ~pc & new_n7260;
  assign new_n7262 = ~pm & new_n7261;
  assign new_n7263 = ~pd0 & new_n7262;
  assign new_n7264 = ~pi0 & new_n7263;
  assign new_n7265 = ~pi & new_n7264;
  assign new_n7266 = ~pg & new_n7265;
  assign new_n7267 = ~ph & new_n7266;
  assign new_n7268 = ~pe & new_n7267;
  assign new_n7269 = ~pf & new_n7268;
  assign new_n7270 = ~pa0 & new_n6385;
  assign new_n7271 = ~pc & new_n7270;
  assign new_n7272 = ~pm & new_n7271;
  assign new_n7273 = ~ph & new_n7272;
  assign new_n7274 = ~pd0 & new_n7273;
  assign new_n7275 = ~pg & new_n7274;
  assign new_n7276 = ~pe & new_n7275;
  assign new_n7277 = ~pf & new_n7276;
  assign new_n7278 = pm0 & new_n7277;
  assign new_n7279 = ~ph0 & new_n7278;
  assign new_n7280 = ~pa0 & new_n6787;
  assign new_n7281 = ~pc0 & new_n7280;
  assign new_n7282 = ~py & new_n7281;
  assign new_n7283 = ~pd0 & new_n7282;
  assign new_n7284 = ~pf0 & new_n7283;
  assign new_n7285 = ~ph0 & new_n7284;
  assign new_n7286 = ~pj0 & new_n7285;
  assign new_n7287 = pm0 & new_n7286;
  assign new_n7288 = ~pe0 & new_n3791;
  assign new_n7289 = ~pz & new_n7288;
  assign new_n7290 = ~pd0 & new_n7289;
  assign new_n7291 = ~pi0 & new_n7290;
  assign new_n7292 = pm0 & new_n7291;
  assign new_n7293 = ~ph & new_n7292;
  assign new_n7294 = pm0 & new_n7143;
  assign new_n7295 = ~ph0 & new_n7294;
  assign new_n7296 = ~pc0 & new_n7295;
  assign new_n7297 = ~pj0 & new_n7296;
  assign new_n7298 = ~pg0 & new_n6977;
  assign new_n7299 = ~pc & new_n7298;
  assign new_n7300 = ~pm & new_n7299;
  assign new_n7301 = ~pd0 & new_n7300;
  assign new_n7302 = ~pi0 & new_n7301;
  assign new_n7303 = ~ph & new_n7302;
  assign new_n7304 = ~pf & new_n7303;
  assign new_n7305 = ~pg & new_n7304;
  assign new_n7306 = ~ph0 & new_n7305;
  assign new_n7307 = ~pe & new_n7306;
  assign new_n7308 = pm0 & new_n7126;
  assign new_n7309 = ~pf0 & new_n7308;
  assign new_n7310 = ~pg0 & new_n7309;
  assign new_n7311 = ~pj0 & new_n7310;
  assign new_n7312 = ~pc0 & new_n6570;
  assign new_n7313 = ~pe0 & new_n7312;
  assign new_n7314 = ~py & new_n7313;
  assign new_n7315 = ~pd0 & new_n7314;
  assign new_n7316 = pi0 & new_n7315;
  assign new_n7317 = ~ph0 & new_n7316;
  assign new_n7318 = ~ph & new_n7317;
  assign new_n7319 = ~pd0 & ~pi0;
  assign new_n7320 = pg0 & new_n7319;
  assign new_n7321 = pj0 & new_n7320;
  assign new_n7322 = ~pc0 & new_n7321;
  assign new_n7323 = pq & new_n7322;
  assign new_n7324 = ~pw & new_n818;
  assign new_n7325 = pq & new_n7324;
  assign new_n7326 = ~pc0 & pg0;
  assign new_n7327 = ~py & new_n7326;
  assign new_n7328 = ~pa0 & new_n7327;
  assign new_n7329 = pn & new_n7328;
  assign new_n7330 = po & new_n7329;
  assign new_n7331 = pf0 & px;
  assign new_n7332 = ~pa0 & new_n7331;
  assign new_n7333 = ~pc0 & new_n7332;
  assign new_n7334 = ~py & new_n7333;
  assign new_n7335 = ~pf & new_n5726;
  assign new_n7336 = ~pg & new_n7335;
  assign new_n7337 = ~pe & new_n7336;
  assign new_n7338 = ~pj0 & new_n7337;
  assign new_n7339 = pm0 & new_n7338;
  assign new_n7340 = ~pc0 & new_n7339;
  assign new_n7341 = ~pg0 & new_n7340;
  assign new_n7342 = ~pc & new_n6745;
  assign new_n7343 = ~pm & new_n7342;
  assign new_n7344 = ~ph & new_n7343;
  assign new_n7345 = ~pi & new_n7344;
  assign new_n7346 = ~pg & new_n7345;
  assign new_n7347 = ~pe & new_n7346;
  assign new_n7348 = ~pf & new_n7347;
  assign new_n7349 = pm0 & new_n7348;
  assign new_n7350 = ~ph0 & new_n7349;
  assign new_n7351 = ~pi & new_n7342;
  assign new_n7352 = ~ph0 & new_n7351;
  assign new_n7353 = ~ph & new_n7352;
  assign new_n7354 = ~pe0 & new_n7353;
  assign new_n7355 = pm0 & new_n7354;
  assign new_n7356 = ~pe0 & pm0;
  assign new_n7357 = ~pz & new_n7356;
  assign new_n7358 = ~pc0 & new_n7357;
  assign new_n7359 = ~py & new_n7358;
  assign new_n7360 = ~pd0 & new_n7359;
  assign new_n7361 = pi0 & new_n7360;
  assign new_n7362 = ~ph & new_n7361;
  assign new_n7363 = ~pi & new_n7362;
  assign new_n7364 = pe0 & new_n7319;
  assign new_n7365 = pj0 & new_n7364;
  assign new_n7366 = ~pc0 & new_n7365;
  assign new_n7367 = pq & new_n7366;
  assign new_n7368 = pe0 & pi0;
  assign new_n7369 = ~py & new_n7368;
  assign new_n7370 = ~pc0 & new_n7369;
  assign new_n7371 = pw & new_n7370;
  assign new_n7372 = pq & new_n7371;
  assign new_n7373 = ~pc0 & pe0;
  assign new_n7374 = ~py & new_n7373;
  assign new_n7375 = ~pa0 & new_n7374;
  assign new_n7376 = pn & new_n7375;
  assign new_n7377 = po & new_n7376;
  assign new_n7378 = ph0 & po;
  assign new_n7379 = ~pa0 & new_n7378;
  assign new_n7380 = ~pc0 & new_n7379;
  assign new_n7381 = ~py & new_n7380;
  assign new_n7382 = pm0 & new_n6171;
  assign new_n7383 = ~ph & new_n7382;
  assign new_n7384 = ~pc0 & new_n7383;
  assign new_n7385 = ~pe0 & new_n7384;
  assign new_n7386 = ~pa0 & new_n7356;
  assign new_n7387 = ~pc0 & new_n7386;
  assign new_n7388 = ~py & new_n7387;
  assign new_n7389 = ~pi & new_n7388;
  assign new_n7390 = ~pd0 & new_n7389;
  assign new_n7391 = ~ph0 & new_n7390;
  assign new_n7392 = ~ph & new_n7391;
  assign new_n7393 = ~pc0 & new_n1041;
  assign new_n7394 = pf0 & new_n7393;
  assign new_n7395 = ~py & new_n7394;
  assign new_n7396 = pm & new_n7395;
  assign new_n7397 = pr & new_n7396;
  assign new_n7398 = pf0 & ~pi0;
  assign new_n7399 = ~pc0 & new_n7398;
  assign new_n7400 = pj0 & new_n7399;
  assign new_n7401 = pw & new_n7400;
  assign new_n7402 = pq & new_n7401;
  assign new_n7403 = ~pd0 & px;
  assign new_n7404 = pg0 & new_n7403;
  assign new_n7405 = pj0 & new_n7404;
  assign new_n7406 = ~pc0 & new_n7405;
  assign new_n7407 = ~pi0 & new_n7406;
  assign new_n7408 = ~pc0 & px;
  assign new_n7409 = ~py & new_n7408;
  assign new_n7410 = ~pa0 & new_n7409;
  assign new_n7411 = ~pw & new_n7410;
  assign new_n7412 = pd0 & new_n7411;
  assign new_n7413 = px & pi0;
  assign new_n7414 = ~py & new_n7413;
  assign new_n7415 = ~pc0 & new_n7414;
  assign new_n7416 = pw & new_n7415;
  assign new_n7417 = ~ph & new_n7342;
  assign new_n7418 = pm0 & new_n7417;
  assign new_n7419 = ~ph0 & new_n7418;
  assign new_n7420 = ~pe0 & new_n7419;
  assign new_n7421 = ~pg0 & new_n7420;
  assign new_n7422 = ~pd0 & new_n6790;
  assign new_n7423 = pi0 & new_n7422;
  assign new_n7424 = pm0 & new_n7423;
  assign new_n7425 = ~ph & new_n7424;
  assign new_n7426 = pe0 & new_n637;
  assign new_n7427 = pw & new_n7426;
  assign new_n7428 = pm & new_n7427;
  assign new_n7429 = pr & new_n7428;
  assign new_n7430 = pg0 & new_n637;
  assign new_n7431 = pw & new_n7430;
  assign new_n7432 = pq & new_n7431;
  assign new_n7433 = ~pd0 & pf0;
  assign new_n7434 = pj0 & new_n7433;
  assign new_n7435 = px & new_n7434;
  assign new_n7436 = ~pc0 & new_n7435;
  assign new_n7437 = ~pi0 & new_n7436;
  assign new_n7438 = ~pc0 & pf0;
  assign new_n7439 = ~py & new_n7438;
  assign new_n7440 = ~pa0 & new_n7439;
  assign new_n7441 = pn & new_n7440;
  assign new_n7442 = po & new_n7441;
  assign new_n7443 = px & new_n7393;
  assign new_n7444 = ~py & new_n7443;
  assign new_n7445 = pj0 & po;
  assign new_n7446 = ~pc0 & new_n7445;
  assign new_n7447 = pe0 & new_n7446;
  assign new_n7448 = pn & new_n7447;
  assign new_n7449 = ~pd0 & new_n7448;
  assign new_n7450 = ~pi0 & new_n7449;
  assign new_n7451 = pd0 & ~pi0;
  assign new_n7452 = ~pc0 & new_n7451;
  assign new_n7453 = pj0 & new_n7452;
  assign new_n7454 = ~pw & new_n7453;
  assign new_n7455 = pv & new_n7454;
  assign new_n7456 = pq & new_n7427;
  assign new_n7457 = ~pc0 & new_n7378;
  assign new_n7458 = pj0 & new_n7457;
  assign new_n7459 = pw & new_n7458;
  assign new_n7460 = ~pi0 & new_n7459;
  assign new_n7461 = pb0 & pe0;
  assign new_n7462 = ~pa0 & new_n7461;
  assign new_n7463 = ~pc0 & new_n7462;
  assign new_n7464 = ~py & new_n7463;
  assign new_n7465 = pf0 & pj0;
  assign new_n7466 = pw & new_n7465;
  assign new_n7467 = ~pc0 & new_n7466;
  assign new_n7468 = pn & new_n7467;
  assign new_n7469 = po & new_n7468;
  assign new_n7470 = ~pi0 & new_n7469;
  assign new_n7471 = pn & new_n6745;
  assign new_n7472 = po & new_n7471;
  assign new_n7473 = pd0 & new_n7472;
  assign new_n7474 = pq & new_n7395;
  assign new_n7475 = pe0 & new_n7403;
  assign new_n7476 = pj0 & new_n7475;
  assign new_n7477 = ~pc0 & new_n7476;
  assign new_n7478 = ~pi0 & new_n7477;
  assign new_n7479 = pq & pf0;
  assign new_n7480 = ~pa0 & new_n7479;
  assign new_n7481 = ~pc0 & new_n7480;
  assign new_n7482 = ~py & new_n7481;
  assign new_n7483 = pb0 & new_n7366;
  assign new_n7484 = pj0 & new_n7319;
  assign new_n7485 = pf0 & new_n7484;
  assign new_n7486 = ~pc0 & new_n7485;
  assign new_n7487 = pq & new_n7486;
  assign new_n7488 = pg0 & new_n7393;
  assign new_n7489 = ~py & new_n7488;
  assign new_n7490 = pq & new_n7489;
  assign new_n7491 = px & pj0;
  assign new_n7492 = ~pc0 & new_n7491;
  assign new_n7493 = pg0 & new_n7492;
  assign new_n7494 = pw & new_n7493;
  assign new_n7495 = ~pi0 & new_n7494;
  assign new_n7496 = pb0 & pf0;
  assign new_n7497 = ~pa0 & new_n7496;
  assign new_n7498 = ~pc0 & new_n7497;
  assign new_n7499 = ~py & new_n7498;
  assign new_n7500 = pe0 & px;
  assign new_n7501 = ~pa0 & new_n7500;
  assign new_n7502 = ~pc0 & new_n7501;
  assign new_n7503 = ~py & new_n7502;
  assign new_n7504 = pb0 & new_n7401;
  assign new_n7505 = pb0 & new_n7324;
  assign new_n7506 = pe0 & new_n7393;
  assign new_n7507 = ~py & new_n7506;
  assign new_n7508 = pq & new_n7507;
  assign new_n7509 = ~pc0 & new_n7331;
  assign new_n7510 = pj0 & new_n7509;
  assign new_n7511 = pw & new_n7510;
  assign new_n7512 = ~pi0 & new_n7511;
  assign new_n7513 = pb0 & pg0;
  assign new_n7514 = ~pa0 & new_n7513;
  assign new_n7515 = ~pc0 & new_n7514;
  assign new_n7516 = ~py & new_n7515;
  assign new_n7517 = pg0 & px;
  assign new_n7518 = ~pa0 & new_n7517;
  assign new_n7519 = ~pc0 & new_n7518;
  assign new_n7520 = ~py & new_n7519;
  assign new_n7521 = pm & new_n6721;
  assign new_n7522 = pk & new_n7521;
  assign new_n7523 = ~ph & new_n7522;
  assign new_n7524 = pt & new_n7523;
  assign new_n7525 = ~ph0 & new_n7524;
  assign new_n7526 = ~pg0 & new_n7525;
  assign new_n7527 = pm0 & new_n7526;
  assign new_n7528 = ~pc0 & new_n7527;
  assign new_n7529 = ~pe0 & new_n7528;
  assign new_n7530 = ~pn & new_n5875;
  assign new_n7531 = ~py & new_n7530;
  assign new_n7532 = pj & new_n7531;
  assign new_n7533 = ~pd & new_n7532;
  assign new_n7534 = ~pd0 & new_n7533;
  assign new_n7535 = pi0 & new_n7534;
  assign new_n7536 = pt & new_n7535;
  assign new_n7537 = ~pj0 & new_n7536;
  assign new_n7538 = pm0 & new_n7537;
  assign new_n7539 = ~pe0 & new_n7538;
  assign new_n7540 = ~pg0 & new_n7539;
  assign new_n7541 = pl & new_n3448;
  assign new_n7542 = ~pn & new_n7541;
  assign new_n7543 = pj & new_n7542;
  assign new_n7544 = ~pd & new_n7543;
  assign new_n7545 = ~ph0 & new_n7544;
  assign new_n7546 = ~pd0 & new_n7545;
  assign new_n7547 = pm0 & new_n7546;
  assign new_n7548 = ~pg0 & new_n7547;
  assign new_n7549 = ~pj0 & new_n7548;
  assign new_n7550 = ~pc0 & new_n7549;
  assign new_n7551 = ~pe0 & new_n7550;
  assign new_n7552 = ~pb & new_n6778;
  assign new_n7553 = ~pi & new_n7552;
  assign new_n7554 = ~pd0 & new_n7553;
  assign new_n7555 = ~ph & new_n7554;
  assign new_n7556 = ~pf & new_n7555;
  assign new_n7557 = ~pg & new_n7556;
  assign new_n7558 = pm0 & new_n7557;
  assign new_n7559 = ~pe & new_n7558;
  assign new_n7560 = pl & new_n6007;
  assign new_n7561 = ~pn & new_n7560;
  assign new_n7562 = pj & new_n7561;
  assign new_n7563 = pi0 & new_n7562;
  assign new_n7564 = ~pi & new_n7563;
  assign new_n7565 = ~pd0 & new_n7564;
  assign new_n7566 = ~ph0 & new_n7565;
  assign new_n7567 = ~pj0 & new_n7566;
  assign new_n7568 = pm0 & new_n7567;
  assign new_n7569 = ~pc0 & new_n7568;
  assign new_n7570 = ~pe0 & new_n7569;
  assign new_n7571 = pm & new_n7486;
  assign new_n7572 = pr & new_n7571;
  assign new_n7573 = pm & new_n7371;
  assign new_n7574 = pr & new_n7573;
  assign new_n7575 = pw & new_n7438;
  assign new_n7576 = ~py & new_n7575;
  assign new_n7577 = pn & new_n7576;
  assign new_n7578 = po & new_n7577;
  assign new_n7579 = pi0 & new_n7578;
  assign new_n7580 = pb0 & new_n7486;
  assign new_n7581 = pb0 & new_n7371;
  assign new_n7582 = pf0 & pi0;
  assign new_n7583 = ~py & new_n7582;
  assign new_n7584 = ~pc0 & new_n7583;
  assign new_n7585 = pw & new_n7584;
  assign new_n7586 = pq & new_n7585;
  assign new_n7587 = ~py & new_n7378;
  assign new_n7588 = ~pc0 & new_n7587;
  assign new_n7589 = pw & new_n7588;
  assign new_n7590 = pi0 & new_n7589;
  assign new_n7591 = ~py & new_n1763;
  assign new_n7592 = ~pa0 & new_n7591;
  assign new_n7593 = ~pc & new_n7592;
  assign new_n7594 = ~pd0 & new_n7593;
  assign new_n7595 = ~pm & new_n7594;
  assign new_n7596 = ~pg & new_n7595;
  assign new_n7597 = ~pi & new_n7596;
  assign new_n7598 = ~pf & new_n7597;
  assign new_n7599 = ~ph0 & new_n7598;
  assign new_n7600 = ~pe & new_n7599;
  assign new_n7601 = pm0 & new_n7600;
  assign new_n7602 = ~pf0 & new_n7601;
  assign new_n7603 = pl & new_n5821;
  assign new_n7604 = ~pn & new_n7603;
  assign new_n7605 = pj & new_n7604;
  assign new_n7606 = ~pd & new_n7605;
  assign new_n7607 = ~pd0 & new_n7606;
  assign new_n7608 = pi0 & new_n7607;
  assign new_n7609 = ~pi & new_n7608;
  assign new_n7610 = pm0 & new_n7609;
  assign new_n7611 = ~ph0 & new_n7610;
  assign new_n7612 = ~pe0 & new_n7611;
  assign new_n7613 = ~pj0 & new_n7612;
  assign new_n7614 = pl & new_n5718;
  assign new_n7615 = ~pn & new_n7614;
  assign new_n7616 = pj & new_n7615;
  assign new_n7617 = ~pd & new_n7616;
  assign new_n7618 = ~pi & new_n7617;
  assign new_n7619 = ~pd0 & new_n7618;
  assign new_n7620 = pm0 & new_n7619;
  assign new_n7621 = ~pe0 & new_n7620;
  assign new_n7622 = ~pj0 & new_n7621;
  assign new_n7623 = ~pa0 & new_n7622;
  assign new_n7624 = ~pc0 & new_n7623;
  assign new_n7625 = ~pb & new_n7271;
  assign new_n7626 = ~ph & new_n7625;
  assign new_n7627 = ~pd0 & new_n7626;
  assign new_n7628 = ~pg & new_n7627;
  assign new_n7629 = ~pe & new_n7628;
  assign new_n7630 = ~pf & new_n7629;
  assign new_n7631 = pm0 & new_n7630;
  assign new_n7632 = ~ph0 & new_n7631;
  assign new_n7633 = ps & new_n6756;
  assign new_n7634 = pj & new_n7633;
  assign new_n7635 = pi0 & new_n7634;
  assign new_n7636 = pt & new_n7635;
  assign new_n7637 = ~pd0 & new_n7636;
  assign new_n7638 = pm0 & new_n7637;
  assign new_n7639 = ~pg0 & new_n7638;
  assign new_n7640 = ~pj0 & new_n7639;
  assign new_n7641 = ~pc0 & new_n7640;
  assign new_n7642 = ~pe0 & new_n7641;
  assign new_n7643 = ~ph & new_n7125;
  assign new_n7644 = ~pd0 & new_n7643;
  assign new_n7645 = ~pg0 & new_n7644;
  assign new_n7646 = pm0 & new_n7645;
  assign new_n7647 = pm & new_n7324;
  assign new_n7648 = pr & new_n7647;
  assign new_n7649 = pe0 & po;
  assign new_n7650 = ~py & new_n7649;
  assign new_n7651 = ~pc0 & new_n7650;
  assign new_n7652 = pn & new_n7651;
  assign new_n7653 = ~pd0 & new_n7652;
  assign new_n7654 = pi0 & new_n7653;
  assign new_n7655 = pb0 & new_n7322;
  assign new_n7656 = pg0 & pi0;
  assign new_n7657 = ~py & new_n7656;
  assign new_n7658 = ~pc0 & new_n7657;
  assign new_n7659 = pw & new_n7658;
  assign new_n7660 = pb0 & new_n7659;
  assign new_n7661 = pq & new_n7659;
  assign new_n7662 = pe0 & new_n7492;
  assign new_n7663 = pw & new_n7662;
  assign new_n7664 = ~pi0 & new_n7663;
  assign new_n7665 = ~pn & new_n3448;
  assign new_n7666 = ~pw & new_n7665;
  assign new_n7667 = pj & new_n7666;
  assign new_n7668 = ~pd & new_n7667;
  assign new_n7669 = pm & new_n7668;
  assign new_n7670 = ~ph0 & new_n7669;
  assign new_n7671 = pt & new_n7670;
  assign new_n7672 = pm0 & new_n7671;
  assign new_n7673 = ~pg0 & new_n7672;
  assign new_n7674 = ~pj0 & new_n7673;
  assign new_n7675 = ~pc0 & new_n7674;
  assign new_n7676 = ~pe0 & new_n7675;
  assign new_n7677 = ~pd0 & new_n7617;
  assign new_n7678 = pi0 & new_n7677;
  assign new_n7679 = ~pi & new_n7678;
  assign new_n7680 = ~pj0 & new_n7679;
  assign new_n7681 = pm0 & new_n7680;
  assign new_n7682 = ~pc0 & new_n7681;
  assign new_n7683 = ~pe0 & new_n7682;
  assign new_n7684 = ~pb & new_n7106;
  assign new_n7685 = ~pd0 & new_n7684;
  assign new_n7686 = ~pi0 & new_n7685;
  assign new_n7687 = ~pi & new_n7686;
  assign new_n7688 = ~pg & new_n7687;
  assign new_n7689 = ~ph & new_n7688;
  assign new_n7690 = ~pe & new_n7689;
  assign new_n7691 = ~pf & new_n7690;
  assign new_n7692 = ~pb & new_n6387;
  assign new_n7693 = ~pd0 & new_n7692;
  assign new_n7694 = pi0 & new_n7693;
  assign new_n7695 = ~ph & new_n7694;
  assign new_n7696 = ~pf & new_n7695;
  assign new_n7697 = ~pg & new_n7696;
  assign new_n7698 = pm0 & new_n7697;
  assign new_n7699 = ~pe & new_n7698;
  assign new_n7700 = ~pn & new_n5821;
  assign new_n7701 = ps & new_n7700;
  assign new_n7702 = pj & new_n7701;
  assign new_n7703 = pi0 & new_n7702;
  assign new_n7704 = pt & new_n7703;
  assign new_n7705 = ~pd0 & new_n7704;
  assign new_n7706 = ~ph0 & new_n7705;
  assign new_n7707 = ~pj0 & new_n7706;
  assign new_n7708 = pm0 & new_n7707;
  assign new_n7709 = ~pe0 & new_n7708;
  assign new_n7710 = ~pg0 & new_n7709;
  assign new_n7711 = ~ph & new_n7282;
  assign new_n7712 = ~pd0 & new_n7711;
  assign new_n7713 = pm0 & new_n7712;
  assign new_n7714 = ~ph0 & new_n7713;
  assign new_n7715 = pf0 & po;
  assign new_n7716 = ~pc0 & new_n7715;
  assign new_n7717 = pj0 & new_n7716;
  assign new_n7718 = pn & new_n7717;
  assign new_n7719 = ~pd0 & new_n7718;
  assign new_n7720 = ~pi0 & new_n7719;
  assign new_n7721 = pw & new_n7373;
  assign new_n7722 = ~py & new_n7721;
  assign new_n7723 = pn & new_n7722;
  assign new_n7724 = po & new_n7723;
  assign new_n7725 = pi0 & new_n7724;
  assign new_n7726 = pg0 & pm;
  assign new_n7727 = ~pa0 & new_n7726;
  assign new_n7728 = ~pc0 & new_n7727;
  assign new_n7729 = ~py & new_n7728;
  assign new_n7730 = pr & new_n7729;
  assign new_n7731 = pb0 & new_n7585;
  assign new_n7732 = pq & pg0;
  assign new_n7733 = ~pa0 & new_n7732;
  assign new_n7734 = ~pc0 & new_n7733;
  assign new_n7735 = ~py & new_n7734;
  assign new_n7736 = pm0 & new_n6557;
  assign new_n7737 = ~ph0 & new_n7736;
  assign new_n7738 = ~pj0 & new_n7737;
  assign new_n7739 = ~pc0 & new_n7738;
  assign new_n7740 = ~pe0 & new_n7739;
  assign new_n7741 = ~py & new_n7740;
  assign new_n7742 = ~pa0 & new_n7741;
  assign new_n7743 = ~ph0 & new_n7608;
  assign new_n7744 = ~pj0 & new_n7743;
  assign new_n7745 = pm0 & new_n7744;
  assign new_n7746 = ~pe0 & new_n7745;
  assign new_n7747 = ~pg0 & new_n7746;
  assign new_n7748 = pm0 & new_n7617;
  assign new_n7749 = ~pd0 & new_n7748;
  assign new_n7750 = ~pj0 & new_n7749;
  assign new_n7751 = ~pe0 & new_n7750;
  assign new_n7752 = ~pg0 & new_n7751;
  assign new_n7753 = ~pa0 & new_n7752;
  assign new_n7754 = ~pc0 & new_n7753;
  assign new_n7755 = ~pb & new_n6960;
  assign new_n7756 = ~pi & new_n7755;
  assign new_n7757 = ~pd0 & new_n7756;
  assign new_n7758 = ~ph & new_n7757;
  assign new_n7759 = ~pf & new_n7758;
  assign new_n7760 = ~pg & new_n7759;
  assign new_n7761 = ~ph0 & new_n7760;
  assign new_n7762 = ~pe & new_n7761;
  assign new_n7763 = ~pi & new_n7637;
  assign new_n7764 = ~pj0 & new_n7763;
  assign new_n7765 = pm0 & new_n7764;
  assign new_n7766 = ~pc0 & new_n7765;
  assign new_n7767 = ~pe0 & new_n7766;
  assign new_n7768 = ~pi & new_n7125;
  assign new_n7769 = ~pd0 & new_n7768;
  assign new_n7770 = pm0 & new_n7769;
  assign new_n7771 = ~ph & new_n7770;
  assign new_n7772 = pg0 & new_n7446;
  assign new_n7773 = pn & new_n7772;
  assign new_n7774 = ~pd0 & new_n7773;
  assign new_n7775 = ~pi0 & new_n7774;
  assign new_n7776 = pw & new_n7326;
  assign new_n7777 = ~py & new_n7776;
  assign new_n7778 = pn & new_n7777;
  assign new_n7779 = po & new_n7778;
  assign new_n7780 = pi0 & new_n7779;
  assign new_n7781 = pe0 & pm;
  assign new_n7782 = ~pa0 & new_n7781;
  assign new_n7783 = ~pc0 & new_n7782;
  assign new_n7784 = ~py & new_n7783;
  assign new_n7785 = pr & new_n7784;
  assign new_n7786 = pb0 & new_n7507;
  assign new_n7787 = pq & pe0;
  assign new_n7788 = ~pa0 & new_n7787;
  assign new_n7789 = ~pc0 & new_n7788;
  assign new_n7790 = ~py & new_n7789;
  assign new_n7791 = ~ph0 & new_n6364;
  assign new_n7792 = ~pd & new_n7791;
  assign new_n7793 = ~pj0 & new_n7792;
  assign new_n7794 = pm0 & new_n7793;
  assign new_n7795 = ~pg0 & new_n7794;
  assign new_n7796 = ~pc0 & new_n7795;
  assign new_n7797 = ~pe0 & new_n7796;
  assign new_n7798 = ~py & new_n7797;
  assign new_n7799 = ~pa0 & new_n7798;
  assign new_n7800 = ~pd0 & new_n7634;
  assign new_n7801 = pm0 & new_n7800;
  assign new_n7802 = pt & new_n7801;
  assign new_n7803 = ~pj0 & new_n7802;
  assign new_n7804 = ~pe0 & new_n7803;
  assign new_n7805 = ~pg0 & new_n7804;
  assign new_n7806 = ~pa0 & new_n7805;
  assign new_n7807 = ~pc0 & new_n7806;
  assign new_n7808 = ~ph0 & new_n6086;
  assign new_n7809 = ~pk & new_n7808;
  assign new_n7810 = pm0 & new_n7809;
  assign new_n7811 = ~pg0 & new_n7810;
  assign new_n7812 = ~pj0 & new_n7811;
  assign new_n7813 = ~pc0 & new_n7812;
  assign new_n7814 = ~pe0 & new_n7813;
  assign new_n7815 = pj & new_n6777;
  assign new_n7816 = ~pk & new_n7815;
  assign new_n7817 = ~pd0 & new_n7816;
  assign new_n7818 = pm0 & new_n7817;
  assign new_n7819 = ~pi & new_n7818;
  assign new_n7820 = ~pe0 & new_n7819;
  assign new_n7821 = ~pj0 & new_n7820;
  assign new_n7822 = ~pj0 & pm0;
  assign new_n7823 = ~pc0 & new_n7822;
  assign new_n7824 = ~pe0 & new_n7823;
  assign new_n7825 = ~py & new_n7824;
  assign new_n7826 = pi0 & new_n7825;
  assign new_n7827 = ~pi & new_n7826;
  assign new_n7828 = ~pd0 & new_n7827;
  assign new_n7829 = ~pf0 & new_n7828;
  assign new_n7830 = ~ph0 & new_n7829;
  assign new_n7831 = pm & new_n7431;
  assign new_n7832 = pr & new_n7831;
  assign new_n7833 = pm & new_n7489;
  assign new_n7834 = pr & new_n7833;
  assign new_n7835 = pe0 & pj0;
  assign new_n7836 = pw & new_n7835;
  assign new_n7837 = ~pc0 & new_n7836;
  assign new_n7838 = pn & new_n7837;
  assign new_n7839 = po & new_n7838;
  assign new_n7840 = ~pi0 & new_n7839;
  assign new_n7841 = pd0 & pi0;
  assign new_n7842 = ~py & new_n7841;
  assign new_n7843 = ~pc0 & new_n7842;
  assign new_n7844 = ~pw & new_n7843;
  assign new_n7845 = pu & new_n7844;
  assign new_n7846 = pb0 & new_n7489;
  assign new_n7847 = ~pb & new_n7351;
  assign new_n7848 = ~pf & new_n7847;
  assign new_n7849 = ~pg & new_n7848;
  assign new_n7850 = ~pe & new_n7849;
  assign new_n7851 = ~pf0 & new_n7850;
  assign new_n7852 = ~ph0 & new_n7851;
  assign new_n7853 = ~pj0 & new_n7852;
  assign new_n7854 = pm0 & new_n7853;
  assign new_n7855 = ~pd0 & new_n7562;
  assign new_n7856 = ~ph0 & new_n7855;
  assign new_n7857 = ~pi & new_n7856;
  assign new_n7858 = pm0 & new_n7857;
  assign new_n7859 = ~pe0 & new_n7858;
  assign new_n7860 = ~pj0 & new_n7859;
  assign new_n7861 = ~pa0 & new_n7860;
  assign new_n7862 = ~pc0 & new_n7861;
  assign new_n7863 = ~pi & new_n5864;
  assign new_n7864 = ~pk & new_n7863;
  assign new_n7865 = pm0 & new_n7864;
  assign new_n7866 = ~pe0 & new_n7865;
  assign new_n7867 = ~pj0 & new_n7866;
  assign new_n7868 = ~pa0 & new_n7867;
  assign new_n7869 = ~pc0 & new_n7868;
  assign new_n7870 = ~py & new_n7122;
  assign new_n7871 = ~pa0 & new_n7870;
  assign new_n7872 = pj & new_n7871;
  assign new_n7873 = ~pk & new_n7872;
  assign new_n7874 = ~pd0 & new_n7873;
  assign new_n7875 = pm0 & new_n7874;
  assign new_n7876 = ~ph0 & new_n7875;
  assign new_n7877 = ~pg0 & new_n7876;
  assign new_n7878 = ~pj0 & new_n7877;
  assign new_n7879 = ~pf0 & new_n6170;
  assign new_n7880 = pm0 & new_n7879;
  assign new_n7881 = ~pg0 & new_n7880;
  assign new_n7882 = ~pj0 & new_n7881;
  assign new_n7883 = ~pc0 & new_n7882;
  assign new_n7884 = ~pe0 & new_n7883;
  assign new_n7885 = pm & new_n7401;
  assign new_n7886 = pr & new_n7885;
  assign new_n7887 = pm & new_n7507;
  assign new_n7888 = pr & new_n7887;
  assign new_n7889 = pg0 & pj0;
  assign new_n7890 = pw & new_n7889;
  assign new_n7891 = ~pc0 & new_n7890;
  assign new_n7892 = pn & new_n7891;
  assign new_n7893 = po & new_n7892;
  assign new_n7894 = ~pi0 & new_n7893;
  assign new_n7895 = pf0 & pm;
  assign new_n7896 = ~pa0 & new_n7895;
  assign new_n7897 = ~pc0 & new_n7896;
  assign new_n7898 = ~py & new_n7897;
  assign new_n7899 = pr & new_n7898;
  assign new_n7900 = pb0 & new_n7395;
  assign new_n7901 = pm0 & new_n5744;
  assign new_n7902 = ~pc0 & new_n7901;
  assign new_n7903 = ~pj0 & new_n7902;
  assign new_n7904 = ~pz & new_n7903;
  assign new_n7905 = ~pa0 & new_n7904;
  assign new_n7906 = ~pi & new_n6011;
  assign new_n7907 = pt & new_n7906;
  assign new_n7908 = ~pd0 & new_n7907;
  assign new_n7909 = pi0 & new_n7908;
  assign new_n7910 = ~pf & new_n7909;
  assign new_n7911 = ~pg & new_n7910;
  assign new_n7912 = ~pe & new_n7911;
  assign new_n7913 = pm0 & new_n7912;
  assign new_n7914 = ~ph0 & new_n7913;
  assign new_n7915 = ~pc0 & new_n7914;
  assign new_n7916 = ~pj0 & new_n7915;
  assign new_n7917 = ~pd0 & new_n6122;
  assign new_n7918 = pi0 & new_n7917;
  assign new_n7919 = ~pg & new_n7918;
  assign new_n7920 = ~ph & new_n7919;
  assign new_n7921 = ~pf & new_n7920;
  assign new_n7922 = ~ph0 & new_n7921;
  assign new_n7923 = ~pe & new_n7922;
  assign new_n7924 = ~pg0 & new_n7923;
  assign new_n7925 = pm0 & new_n7924;
  assign new_n7926 = pm0 & new_n7855;
  assign new_n7927 = ~pi & new_n7926;
  assign new_n7928 = ~pj0 & new_n7927;
  assign new_n7929 = ~pc0 & new_n7928;
  assign new_n7930 = ~pe0 & new_n7929;
  assign new_n7931 = ~pz & new_n7930;
  assign new_n7932 = ~pa0 & new_n7931;
  assign new_n7933 = pj & new_n6745;
  assign new_n7934 = ~pi & new_n7933;
  assign new_n7935 = pm & new_n7934;
  assign new_n7936 = ~ph0 & new_n7935;
  assign new_n7937 = pm0 & new_n7936;
  assign new_n7938 = ~pf0 & new_n7937;
  assign new_n7939 = ~pe0 & new_n7938;
  assign new_n7940 = ~pj0 & new_n7939;
  assign new_n7941 = ~pz & new_n7870;
  assign new_n7942 = pj & new_n7941;
  assign new_n7943 = ~pk & new_n7942;
  assign new_n7944 = pi0 & new_n7943;
  assign new_n7945 = pm0 & new_n7944;
  assign new_n7946 = ~pd0 & new_n7945;
  assign new_n7947 = ~pg0 & new_n7946;
  assign new_n7948 = ~pj0 & new_n7947;
  assign new_n7949 = ~ph0 & new_n7342;
  assign new_n7950 = ~pf0 & new_n7949;
  assign new_n7951 = ~pj0 & new_n7950;
  assign new_n7952 = pm0 & new_n7951;
  assign new_n7953 = ~pe0 & new_n7952;
  assign new_n7954 = ~pg0 & new_n7953;
  assign new_n7955 = pm & new_n7366;
  assign new_n7956 = pr & new_n7955;
  assign new_n7957 = pm & new_n7585;
  assign new_n7958 = pr & new_n7957;
  assign new_n7959 = pg0 & po;
  assign new_n7960 = ~py & new_n7959;
  assign new_n7961 = ~pc0 & new_n7960;
  assign new_n7962 = pn & new_n7961;
  assign new_n7963 = ~pd0 & new_n7962;
  assign new_n7964 = pi0 & new_n7963;
  assign new_n7965 = pv & new_n7844;
  assign new_n7966 = pb0 & new_n7427;
  assign new_n7967 = ~pf & new_n5738;
  assign new_n7968 = ~pg & new_n7967;
  assign new_n7969 = ~pd0 & new_n7968;
  assign new_n7970 = ~pd & new_n7969;
  assign new_n7971 = ~ph0 & new_n7970;
  assign new_n7972 = ~pe & new_n7971;
  assign new_n7973 = pm0 & new_n7972;
  assign new_n7974 = ~pg0 & new_n7973;
  assign new_n7975 = ~pj0 & new_n7974;
  assign new_n7976 = ~pa0 & new_n7975;
  assign new_n7977 = ~pc0 & new_n7976;
  assign new_n7978 = ~pm & new_n6364;
  assign new_n7979 = ~pe & new_n7978;
  assign new_n7980 = ~pf & new_n7979;
  assign new_n7981 = ~pg & new_n7980;
  assign new_n7982 = ~pd & new_n7981;
  assign new_n7983 = ~pj0 & new_n7982;
  assign new_n7984 = pm0 & new_n7983;
  assign new_n7985 = ~pg0 & new_n7984;
  assign new_n7986 = ~pa0 & new_n7985;
  assign new_n7987 = ~pc0 & new_n7986;
  assign new_n7988 = ~py & new_n7987;
  assign new_n7989 = ~pz & new_n7988;
  assign new_n7990 = ~ph & new_n6375;
  assign new_n7991 = ~pi & new_n7990;
  assign new_n7992 = ~pf & new_n7991;
  assign new_n7993 = ~pg & new_n7992;
  assign new_n7994 = ~pe & new_n7993;
  assign new_n7995 = pm0 & new_n7994;
  assign new_n7996 = ~ph0 & new_n7995;
  assign new_n7997 = ~pa0 & new_n7996;
  assign new_n7998 = ~pc0 & new_n7997;
  assign new_n7999 = ~ph0 & new_n7926;
  assign new_n8000 = ~pj0 & new_n7999;
  assign new_n8001 = ~pe0 & new_n8000;
  assign new_n8002 = ~pg0 & new_n8001;
  assign new_n8003 = ~pa0 & new_n8002;
  assign new_n8004 = ~pc0 & new_n8003;
  assign new_n8005 = pm0 & new_n5864;
  assign new_n8006 = ~pk & new_n8005;
  assign new_n8007 = ~pj0 & new_n8006;
  assign new_n8008 = ~pe0 & new_n8007;
  assign new_n8009 = ~pg0 & new_n8008;
  assign new_n8010 = ~pa0 & new_n8009;
  assign new_n8011 = ~pc0 & new_n8010;
  assign new_n8012 = ~ph0 & new_n7874;
  assign new_n8013 = ~pi & new_n8012;
  assign new_n8014 = ~pj0 & new_n8013;
  assign new_n8015 = pm0 & new_n8014;
  assign new_n8016 = ~pf0 & new_n6171;
  assign new_n8017 = ~pj0 & new_n8016;
  assign new_n8018 = pm0 & new_n8017;
  assign new_n8019 = ~pc0 & new_n8018;
  assign new_n8020 = ~pe0 & new_n8019;
  assign new_n8021 = pm & new_n7322;
  assign new_n8022 = pr & new_n8021;
  assign new_n8023 = pm & new_n7659;
  assign new_n8024 = pr & new_n8023;
  assign new_n8025 = ~py & new_n7715;
  assign new_n8026 = ~pc0 & new_n8025;
  assign new_n8027 = pn & new_n8026;
  assign new_n8028 = ~pd0 & new_n8027;
  assign new_n8029 = pi0 & new_n8028;
  assign new_n8030 = pu & new_n7454;
  assign new_n8031 = pb0 & new_n7431;
  assign new_n8032 = pm0 & new_n7970;
  assign new_n8033 = ~pe & new_n8032;
  assign new_n8034 = ~pj0 & new_n8033;
  assign new_n8035 = ~pc0 & new_n8034;
  assign new_n8036 = ~pg0 & new_n8035;
  assign new_n8037 = ~pz & new_n8036;
  assign new_n8038 = ~pa0 & new_n8037;
  assign new_n8039 = pt & new_n6012;
  assign new_n8040 = ~pd0 & new_n8039;
  assign new_n8041 = pi0 & new_n8040;
  assign new_n8042 = ~pe & new_n8041;
  assign new_n8043 = ~pf & new_n8042;
  assign new_n8044 = ~ph0 & new_n8043;
  assign new_n8045 = ~pj0 & new_n8044;
  assign new_n8046 = pm0 & new_n8045;
  assign new_n8047 = ~pc0 & new_n8046;
  assign new_n8048 = ~pg0 & new_n8047;
  assign new_n8049 = ~pf & new_n5754;
  assign new_n8050 = ~pg & new_n8049;
  assign new_n8051 = ~pi & new_n8050;
  assign new_n8052 = pt & new_n8051;
  assign new_n8053 = ~ph0 & new_n8052;
  assign new_n8054 = ~pe & new_n8053;
  assign new_n8055 = pm0 & new_n8054;
  assign new_n8056 = ~pc0 & new_n8055;
  assign new_n8057 = ~pj0 & new_n8056;
  assign new_n8058 = ~py & new_n8057;
  assign new_n8059 = ~pa0 & new_n8058;
  assign new_n8060 = ~pf & new_n7000;
  assign new_n8061 = ~pg & new_n8060;
  assign new_n8062 = ~pe & new_n8061;
  assign new_n8063 = ~pj0 & new_n8062;
  assign new_n8064 = pm0 & new_n8063;
  assign new_n8065 = ~pc0 & new_n8064;
  assign new_n8066 = ~pg0 & new_n8065;
  assign new_n8067 = ~ph0 & new_n6241;
  assign new_n8068 = ~pe & new_n8067;
  assign new_n8069 = pm0 & new_n8068;
  assign new_n8070 = ~pg0 & new_n8069;
  assign new_n8071 = ~pj0 & new_n8070;
  assign new_n8072 = ~pa0 & new_n8071;
  assign new_n8073 = ~pc0 & new_n8072;
  assign new_n8074 = ~pg & new_n6076;
  assign new_n8075 = ~pd0 & new_n8074;
  assign new_n8076 = ~pf & new_n8075;
  assign new_n8077 = pm0 & new_n8076;
  assign new_n8078 = ~pe & new_n8077;
  assign new_n8079 = ~pg0 & new_n8078;
  assign new_n8080 = ~pj0 & new_n8079;
  assign new_n8081 = pj & new_n6155;
  assign new_n8082 = ~py & new_n8081;
  assign new_n8083 = ~pc & new_n8082;
  assign new_n8084 = ~pd0 & new_n8083;
  assign new_n8085 = ~pb & new_n8084;
  assign new_n8086 = ~pk & new_n8085;
  assign new_n8087 = ~pg & new_n8086;
  assign new_n8088 = ~pi & new_n8087;
  assign new_n8089 = ~pf & new_n8088;
  assign new_n8090 = pm0 & new_n8089;
  assign new_n8091 = ~pe & new_n8090;
  assign new_n8092 = ~pc0 & new_n8091;
  assign new_n8093 = ~pj0 & new_n8092;
  assign new_n8094 = ~pj & new_n6743;
  assign new_n8095 = ~py & new_n8094;
  assign new_n8096 = ~pc & new_n8095;
  assign new_n8097 = ~pi & new_n8096;
  assign new_n8098 = ~pd0 & new_n8097;
  assign new_n8099 = ~pk & new_n8098;
  assign new_n8100 = ~pf & new_n8099;
  assign new_n8101 = ~pg & new_n8100;
  assign new_n8102 = ~pe & new_n8101;
  assign new_n8103 = ~pf0 & new_n8102;
  assign new_n8104 = ~ph0 & new_n8103;
  assign new_n8105 = ~pj0 & new_n8104;
  assign new_n8106 = pm0 & new_n8105;
  assign new_n8107 = ~pd & new_n7249;
  assign new_n8108 = pm & new_n8107;
  assign new_n8109 = pk & new_n8108;
  assign new_n8110 = ~pf0 & new_n8109;
  assign new_n8111 = pt & new_n8110;
  assign new_n8112 = pm0 & new_n8111;
  assign new_n8113 = ~pg0 & new_n8112;
  assign new_n8114 = ~pj0 & new_n8113;
  assign new_n8115 = ~pc0 & new_n8114;
  assign new_n8116 = ~pe0 & new_n8115;
  assign new_n8117 = ~pn & new_n5778;
  assign new_n8118 = ps & new_n8117;
  assign new_n8119 = pl & new_n8118;
  assign new_n8120 = ~ph0 & new_n8119;
  assign new_n8121 = pm & new_n8120;
  assign new_n8122 = pk & new_n8121;
  assign new_n8123 = pm0 & new_n8122;
  assign new_n8124 = ~pf0 & new_n8123;
  assign new_n8125 = ~pj0 & new_n8124;
  assign new_n8126 = ~pe0 & new_n8125;
  assign new_n8127 = ~pg0 & new_n8126;
  assign new_n8128 = ~pa0 & new_n8127;
  assign new_n8129 = ~pc0 & new_n8128;
  assign new_n8130 = pd & new_n6470;
  assign new_n8131 = ~pg & new_n8130;
  assign new_n8132 = ~ph & new_n8131;
  assign new_n8133 = ~pf & new_n8132;
  assign new_n8134 = pm0 & new_n8133;
  assign new_n8135 = ~pe & new_n8134;
  assign new_n8136 = ~pa0 & new_n8135;
  assign new_n8137 = ~pc0 & new_n8136;
  assign new_n8138 = ~ph & new_n6512;
  assign new_n8139 = ~pi & new_n8138;
  assign new_n8140 = ~pg & new_n8139;
  assign new_n8141 = ~pe & new_n8140;
  assign new_n8142 = ~pf & new_n8141;
  assign new_n8143 = pm0 & new_n8142;
  assign new_n8144 = ~ph0 & new_n8143;
  assign new_n8145 = ~ph & new_n6750;
  assign new_n8146 = pm0 & new_n8145;
  assign new_n8147 = ~ph0 & new_n8146;
  assign new_n8148 = ~pe0 & new_n8147;
  assign new_n8149 = ~pg0 & new_n8148;
  assign new_n8150 = pm & new_n8119;
  assign new_n8151 = pk & new_n8150;
  assign new_n8152 = ~ph & new_n8151;
  assign new_n8153 = ~pi & new_n8152;
  assign new_n8154 = pm0 & new_n8153;
  assign new_n8155 = ~pc0 & new_n8154;
  assign new_n8156 = ~pe0 & new_n8155;
  assign new_n8157 = ~pz & new_n8156;
  assign new_n8158 = ~pa0 & new_n8157;
  assign new_n8159 = ~pm & new_n7351;
  assign new_n8160 = ~pf & new_n8159;
  assign new_n8161 = ~pg & new_n8160;
  assign new_n8162 = ~pe & new_n8161;
  assign new_n8163 = ~pf0 & new_n8162;
  assign new_n8164 = ~ph0 & new_n8163;
  assign new_n8165 = ~pj0 & new_n8164;
  assign new_n8166 = pm0 & new_n8165;
  assign new_n8167 = pl & new_n5778;
  assign new_n8168 = ~pn & new_n8167;
  assign new_n8169 = pj & new_n8168;
  assign new_n8170 = ~pd & new_n8169;
  assign new_n8171 = pm & new_n8170;
  assign new_n8172 = ~pj0 & new_n8171;
  assign new_n8173 = pm0 & new_n8172;
  assign new_n8174 = ~pg0 & new_n8173;
  assign new_n8175 = ~pc0 & new_n8174;
  assign new_n8176 = ~pe0 & new_n8175;
  assign new_n8177 = ~pz & new_n8176;
  assign new_n8178 = ~pa0 & new_n8177;
  assign new_n8179 = pt & new_n5781;
  assign new_n8180 = ~pd & new_n8179;
  assign new_n8181 = pm0 & new_n8180;
  assign new_n8182 = ~ph0 & new_n8181;
  assign new_n8183 = ~pj0 & new_n8182;
  assign new_n8184 = ~pe0 & new_n8183;
  assign new_n8185 = ~pg0 & new_n8184;
  assign new_n8186 = ~pa0 & new_n8185;
  assign new_n8187 = ~pc0 & new_n8186;
  assign new_n8188 = ~pb & new_n6941;
  assign new_n8189 = ~pg & new_n8188;
  assign new_n8190 = ~pi & new_n8189;
  assign new_n8191 = ~pf & new_n8190;
  assign new_n8192 = ~pf0 & new_n8191;
  assign new_n8193 = ~pe & new_n8192;
  assign new_n8194 = ~pj0 & new_n8193;
  assign new_n8195 = pm0 & new_n8194;
  assign new_n8196 = ~ph & new_n7918;
  assign new_n8197 = ~pi & new_n8196;
  assign new_n8198 = ~pg & new_n8197;
  assign new_n8199 = ~pe & new_n8198;
  assign new_n8200 = ~pf & new_n8199;
  assign new_n8201 = pm0 & new_n8200;
  assign new_n8202 = ~ph0 & new_n8201;
  assign new_n8203 = pm0 & new_n5753;
  assign new_n8204 = pt & new_n8203;
  assign new_n8205 = ~pg0 & new_n8204;
  assign new_n8206 = ~pj0 & new_n8205;
  assign new_n8207 = ~pe0 & new_n8206;
  assign new_n8208 = ~pa0 & new_n8207;
  assign new_n8209 = ~pc0 & new_n8208;
  assign new_n8210 = ~py & new_n8209;
  assign new_n8211 = ~pz & new_n8210;
  assign new_n8212 = ~pb & new_n7261;
  assign new_n8213 = ~pd0 & new_n8212;
  assign new_n8214 = ~pi0 & new_n8213;
  assign new_n8215 = ~pi & new_n8214;
  assign new_n8216 = ~pg & new_n8215;
  assign new_n8217 = ~ph & new_n8216;
  assign new_n8218 = ~pe & new_n8217;
  assign new_n8219 = ~pf & new_n8218;
  assign new_n8220 = ~pb & new_n7342;
  assign new_n8221 = ~ph & new_n8220;
  assign new_n8222 = ~pi & new_n8221;
  assign new_n8223 = ~pg & new_n8222;
  assign new_n8224 = ~pe & new_n8223;
  assign new_n8225 = ~pf & new_n8224;
  assign new_n8226 = pm0 & new_n8225;
  assign new_n8227 = ~ph0 & new_n8226;
  assign new_n8228 = pm0 & new_n7563;
  assign new_n8229 = ~pd0 & new_n8228;
  assign new_n8230 = ~pj0 & new_n8229;
  assign new_n8231 = ~pe0 & new_n8230;
  assign new_n8232 = ~pg0 & new_n8231;
  assign new_n8233 = ~pz & new_n8232;
  assign new_n8234 = ~pc0 & new_n8233;
  assign new_n8235 = pm & new_n7933;
  assign new_n8236 = ~pk & new_n8235;
  assign new_n8237 = ~ph0 & new_n8236;
  assign new_n8238 = ~pj0 & new_n8237;
  assign new_n8239 = pm0 & new_n8238;
  assign new_n8240 = ~pe0 & new_n8239;
  assign new_n8241 = ~pg0 & new_n8240;
  assign new_n8242 = ~pi & new_n7944;
  assign new_n8243 = ~pd0 & new_n8242;
  assign new_n8244 = ~pj0 & new_n8243;
  assign new_n8245 = pm0 & new_n8244;
  assign new_n8246 = pm0 & new_n7352;
  assign new_n8247 = ~pf0 & new_n8246;
  assign new_n8248 = ~pe0 & new_n8247;
  assign new_n8249 = ~pj0 & new_n8248;
  assign new_n8250 = ~pm & new_n5781;
  assign new_n8251 = ~pg & new_n8250;
  assign new_n8252 = ~pi & new_n8251;
  assign new_n8253 = pt & new_n8252;
  assign new_n8254 = ~pd & new_n8253;
  assign new_n8255 = ~pe & new_n8254;
  assign new_n8256 = ~pf & new_n8255;
  assign new_n8257 = ~ph0 & new_n8256;
  assign new_n8258 = ~pj0 & new_n8257;
  assign new_n8259 = pm0 & new_n8258;
  assign new_n8260 = ~pa0 & new_n8259;
  assign new_n8261 = ~pc0 & new_n8260;
  assign new_n8262 = ~pj0 & new_n7912;
  assign new_n8263 = pm0 & new_n8262;
  assign new_n8264 = ~pz & new_n8263;
  assign new_n8265 = ~pc0 & new_n8264;
  assign new_n8266 = pm0 & new_n8052;
  assign new_n8267 = ~pe & new_n8266;
  assign new_n8268 = ~pj0 & new_n8267;
  assign new_n8269 = ~pa0 & new_n8268;
  assign new_n8270 = ~pc0 & new_n8269;
  assign new_n8271 = ~py & new_n8270;
  assign new_n8272 = ~pz & new_n8271;
  assign new_n8273 = ~pf & new_n7159;
  assign new_n8274 = ~pg & new_n8273;
  assign new_n8275 = ~pe & new_n8274;
  assign new_n8276 = pm0 & new_n8275;
  assign new_n8277 = ~ph0 & new_n8276;
  assign new_n8278 = ~pg0 & new_n8277;
  assign new_n8279 = ~pj0 & new_n8278;
  assign new_n8280 = pm0 & new_n6857;
  assign new_n8281 = ~ph0 & new_n8280;
  assign new_n8282 = ~pc0 & new_n8281;
  assign new_n8283 = ~pj0 & new_n8282;
  assign new_n8284 = ~pg & new_n5838;
  assign new_n8285 = ~pi & new_n8284;
  assign new_n8286 = ~pt & new_n8285;
  assign new_n8287 = ~pd0 & new_n8286;
  assign new_n8288 = ~pe & new_n8287;
  assign new_n8289 = ~pf & new_n8288;
  assign new_n8290 = ~pf0 & new_n8289;
  assign new_n8291 = ~pj0 & new_n8290;
  assign new_n8292 = pm0 & new_n8291;
  assign new_n8293 = ~pa0 & new_n8292;
  assign new_n8294 = ~pc0 & new_n8293;
  assign new_n8295 = ~pf & new_n7210;
  assign new_n8296 = ~pg & new_n8295;
  assign new_n8297 = ~pe & new_n8296;
  assign new_n8298 = pm0 & new_n8297;
  assign new_n8299 = ~ph0 & new_n8298;
  assign new_n8300 = ~pg0 & new_n8299;
  assign new_n8301 = ~pj0 & new_n8300;
  assign new_n8302 = ~pf & new_n7220;
  assign new_n8303 = ~pg & new_n8302;
  assign new_n8304 = ~pe & new_n8303;
  assign new_n8305 = pm0 & new_n8304;
  assign new_n8306 = ~pf0 & new_n8305;
  assign new_n8307 = ~pg0 & new_n8306;
  assign new_n8308 = ~pj0 & new_n8307;
  assign new_n8309 = pl & new_n7666;
  assign new_n8310 = ~pd & new_n8309;
  assign new_n8311 = pm & new_n8310;
  assign new_n8312 = pk & new_n8311;
  assign new_n8313 = ~ph0 & new_n8312;
  assign new_n8314 = ~pi & new_n8313;
  assign new_n8315 = ~pf0 & new_n8314;
  assign new_n8316 = ~pj0 & new_n8315;
  assign new_n8317 = pm0 & new_n8316;
  assign new_n8318 = ~pc0 & new_n8317;
  assign new_n8319 = ~pe0 & new_n8318;
  assign new_n8320 = ~pi & new_n8119;
  assign new_n8321 = pm & new_n8320;
  assign new_n8322 = pk & new_n8321;
  assign new_n8323 = pm0 & new_n8322;
  assign new_n8324 = ~pf0 & new_n8323;
  assign new_n8325 = ~pj0 & new_n8324;
  assign new_n8326 = ~pc0 & new_n8325;
  assign new_n8327 = ~pe0 & new_n8326;
  assign new_n8328 = ~pz & new_n8327;
  assign new_n8329 = ~pa0 & new_n8328;
  assign new_n8330 = ~ps & new_n5912;
  assign new_n8331 = ~pc & new_n8330;
  assign new_n8332 = ~ph & new_n8331;
  assign new_n8333 = ~pd0 & new_n8332;
  assign new_n8334 = pd & new_n8333;
  assign new_n8335 = ~pf & new_n8334;
  assign new_n8336 = ~pg & new_n8335;
  assign new_n8337 = ~pe & new_n8336;
  assign new_n8338 = pm0 & new_n8337;
  assign new_n8339 = ~ph0 & new_n8338;
  assign new_n8340 = ~pc0 & new_n8339;
  assign new_n8341 = ~pg0 & new_n8340;
  assign new_n8342 = ~pl & new_n5876;
  assign new_n8343 = ~pc & new_n8342;
  assign new_n8344 = ~pt & new_n8343;
  assign new_n8345 = ~pd0 & new_n8344;
  assign new_n8346 = ~pi0 & new_n8345;
  assign new_n8347 = ~pg & new_n8346;
  assign new_n8348 = ~ph & new_n8347;
  assign new_n8349 = ~pf & new_n8348;
  assign new_n8350 = pm0 & new_n8349;
  assign new_n8351 = ~pe & new_n8350;
  assign new_n8352 = ~pg0 & new_n8351;
  assign new_n8353 = pj0 & new_n8352;
  assign new_n8354 = ~ph & new_n7253;
  assign new_n8355 = ~pg0 & new_n8354;
  assign new_n8356 = pm0 & new_n8355;
  assign new_n8357 = ~pc0 & new_n8356;
  assign new_n8358 = ~pe0 & new_n8357;
  assign new_n8359 = ~ph0 & new_n8153;
  assign new_n8360 = ~pe0 & new_n8359;
  assign new_n8361 = pm0 & new_n8360;
  assign new_n8362 = ~pa0 & new_n8361;
  assign new_n8363 = ~pc0 & new_n8362;
  assign new_n8364 = ~pm & new_n6171;
  assign new_n8365 = ~pf & new_n8364;
  assign new_n8366 = ~pg & new_n8365;
  assign new_n8367 = ~pe & new_n8366;
  assign new_n8368 = pm0 & new_n8367;
  assign new_n8369 = ~pf0 & new_n8368;
  assign new_n8370 = ~pc0 & new_n8369;
  assign new_n8371 = ~pj0 & new_n8370;
  assign new_n8372 = pm0 & new_n8171;
  assign new_n8373 = ~ph0 & new_n8372;
  assign new_n8374 = ~pj0 & new_n8373;
  assign new_n8375 = ~pe0 & new_n8374;
  assign new_n8376 = ~pg0 & new_n8375;
  assign new_n8377 = ~pa0 & new_n8376;
  assign new_n8378 = ~pc0 & new_n8377;
  assign new_n8379 = ~pj0 & new_n8180;
  assign new_n8380 = pm0 & new_n8379;
  assign new_n8381 = ~pg0 & new_n8380;
  assign new_n8382 = ~pc0 & new_n8381;
  assign new_n8383 = ~pe0 & new_n8382;
  assign new_n8384 = ~pz & new_n8383;
  assign new_n8385 = ~pa0 & new_n8384;
  assign new_n8386 = ~pb & new_n7594;
  assign new_n8387 = ~pg & new_n8386;
  assign new_n8388 = ~pi & new_n8387;
  assign new_n8389 = ~pf & new_n8388;
  assign new_n8390 = ~ph0 & new_n8389;
  assign new_n8391 = ~pe & new_n8390;
  assign new_n8392 = pm0 & new_n8391;
  assign new_n8393 = ~pf0 & new_n8392;
  assign new_n8394 = ~ph & new_n5952;
  assign new_n8395 = ~pi & new_n8394;
  assign new_n8396 = ~pg & new_n8395;
  assign new_n8397 = ~pe & new_n8396;
  assign new_n8398 = ~pf & new_n8397;
  assign new_n8399 = ~pc0 & new_n8398;
  assign new_n8400 = pm0 & new_n8399;
  assign new_n8401 = ~ph0 & new_n5753;
  assign new_n8402 = pt & new_n8401;
  assign new_n8403 = ~pj0 & new_n8402;
  assign new_n8404 = pm0 & new_n8403;
  assign new_n8405 = ~pg0 & new_n8404;
  assign new_n8406 = ~pc0 & new_n8405;
  assign new_n8407 = ~pe0 & new_n8406;
  assign new_n8408 = ~py & new_n8407;
  assign new_n8409 = ~pa0 & new_n8408;
  assign new_n8410 = ~pb & new_n7299;
  assign new_n8411 = ~pd0 & new_n8410;
  assign new_n8412 = ~pi0 & new_n8411;
  assign new_n8413 = ~ph & new_n8412;
  assign new_n8414 = ~pf & new_n8413;
  assign new_n8415 = ~pg & new_n8414;
  assign new_n8416 = ~ph0 & new_n8415;
  assign new_n8417 = ~pe & new_n8416;
  assign new_n8418 = ~ph & new_n7552;
  assign new_n8419 = ~pd0 & new_n8418;
  assign new_n8420 = ~pg & new_n8419;
  assign new_n8421 = ~pe & new_n8420;
  assign new_n8422 = ~pf & new_n8421;
  assign new_n8423 = ~pg0 & new_n8422;
  assign new_n8424 = pm0 & new_n8423;
  assign new_n8425 = ps & new_n7665;
  assign new_n8426 = pj & new_n8425;
  assign new_n8427 = ~pd0 & new_n8426;
  assign new_n8428 = ~pi & new_n8427;
  assign new_n8429 = pt & new_n8428;
  assign new_n8430 = ~ph0 & new_n8429;
  assign new_n8431 = ~pj0 & new_n8430;
  assign new_n8432 = pm0 & new_n8431;
  assign new_n8433 = ~pc0 & new_n8432;
  assign new_n8434 = ~pe0 & new_n8433;
  assign new_n8435 = pj & new_n6169;
  assign new_n8436 = pm & new_n8435;
  assign new_n8437 = ~pk & new_n8436;
  assign new_n8438 = ~pi & new_n8437;
  assign new_n8439 = ~pj0 & new_n8438;
  assign new_n8440 = pm0 & new_n8439;
  assign new_n8441 = ~pc0 & new_n8440;
  assign new_n8442 = ~pe0 & new_n8441;
  assign new_n8443 = ~py & new_n6787;
  assign new_n8444 = ~pc0 & new_n8443;
  assign new_n8445 = pj & new_n8444;
  assign new_n8446 = ~pk & new_n8445;
  assign new_n8447 = pi0 & new_n8446;
  assign new_n8448 = ~ph0 & new_n8447;
  assign new_n8449 = ~pd0 & new_n8448;
  assign new_n8450 = ~pj0 & new_n8449;
  assign new_n8451 = pm0 & new_n8450;
  assign new_n8452 = ~ph & new_n8436;
  assign new_n8453 = ~pg0 & new_n8452;
  assign new_n8454 = pm0 & new_n8453;
  assign new_n8455 = ~pc0 & new_n8454;
  assign new_n8456 = ~pe0 & new_n8455;
  assign new_n8457 = pm0 & new_n8256;
  assign new_n8458 = ~pc0 & new_n8457;
  assign new_n8459 = ~pj0 & new_n8458;
  assign new_n8460 = ~pz & new_n8459;
  assign new_n8461 = ~pa0 & new_n8460;
  assign new_n8462 = ~pg & new_n6226;
  assign new_n8463 = ~pi & new_n8462;
  assign new_n8464 = ~pd0 & new_n8463;
  assign new_n8465 = pi0 & new_n8464;
  assign new_n8466 = ~pe & new_n8465;
  assign new_n8467 = ~pf & new_n8466;
  assign new_n8468 = ~ph0 & new_n8467;
  assign new_n8469 = ~pj0 & new_n8468;
  assign new_n8470 = pm0 & new_n8469;
  assign new_n8471 = ~py & new_n8470;
  assign new_n8472 = ~pc0 & new_n8471;
  assign new_n8473 = pm0 & new_n5758;
  assign new_n8474 = ~ph0 & new_n8473;
  assign new_n8475 = ~pj0 & new_n8474;
  assign new_n8476 = ~pc0 & new_n8475;
  assign new_n8477 = ~pg0 & new_n8476;
  assign new_n8478 = ~py & new_n8477;
  assign new_n8479 = ~pa0 & new_n8478;
  assign new_n8480 = ~pi & new_n5767;
  assign new_n8481 = ~pd0 & new_n8480;
  assign new_n8482 = ~pb & new_n8481;
  assign new_n8483 = ~pe & new_n8482;
  assign new_n8484 = ~pf & new_n8483;
  assign new_n8485 = ~ph0 & new_n8484;
  assign new_n8486 = ~pj0 & new_n8485;
  assign new_n8487 = pm0 & new_n8486;
  assign new_n8488 = ~pa0 & new_n8487;
  assign new_n8489 = ~pc0 & new_n8488;
  assign new_n8490 = ~pe & new_n6641;
  assign new_n8491 = ~pf & new_n8490;
  assign new_n8492 = ~pg & new_n8491;
  assign new_n8493 = ~pb & new_n8492;
  assign new_n8494 = ~pj0 & new_n8493;
  assign new_n8495 = pm0 & new_n8494;
  assign new_n8496 = ~pg0 & new_n8495;
  assign new_n8497 = ~pa0 & new_n8496;
  assign new_n8498 = ~pc0 & new_n8497;
  assign new_n8499 = ~py & new_n8498;
  assign new_n8500 = ~pz & new_n8499;
  assign new_n8501 = ~pl & new_n5912;
  assign new_n8502 = ~pc & new_n8501;
  assign new_n8503 = ~pf & new_n8502;
  assign new_n8504 = ~pg & new_n8503;
  assign new_n8505 = ~pt & new_n8504;
  assign new_n8506 = ~pd0 & new_n8505;
  assign new_n8507 = ~ph0 & new_n8506;
  assign new_n8508 = ~pe & new_n8507;
  assign new_n8509 = ~pf0 & new_n8508;
  assign new_n8510 = ~pj0 & new_n8509;
  assign new_n8511 = pm0 & new_n8510;
  assign new_n8512 = ~pc0 & new_n8511;
  assign new_n8513 = ~pg0 & new_n8512;
  assign new_n8514 = ~pm & new_n8084;
  assign new_n8515 = ~pk & new_n8514;
  assign new_n8516 = ~pg & new_n8515;
  assign new_n8517 = ~pi & new_n8516;
  assign new_n8518 = ~pf & new_n8517;
  assign new_n8519 = pm0 & new_n8518;
  assign new_n8520 = ~pe & new_n8519;
  assign new_n8521 = ~pc0 & new_n8520;
  assign new_n8522 = ~pj0 & new_n8521;
  assign new_n8523 = ~pf & new_n8086;
  assign new_n8524 = ~pg & new_n8523;
  assign new_n8525 = ~pe & new_n8524;
  assign new_n8526 = ~pj0 & new_n8525;
  assign new_n8527 = pm0 & new_n8526;
  assign new_n8528 = ~pc0 & new_n8527;
  assign new_n8529 = ~pg0 & new_n8528;
  assign new_n8530 = ~pg & new_n8096;
  assign new_n8531 = ~pd0 & new_n8530;
  assign new_n8532 = ~pk & new_n8531;
  assign new_n8533 = ~pe & new_n8532;
  assign new_n8534 = ~pf & new_n8533;
  assign new_n8535 = ~ph0 & new_n8534;
  assign new_n8536 = pm0 & new_n8535;
  assign new_n8537 = ~pf0 & new_n8536;
  assign new_n8538 = ~pg0 & new_n8537;
  assign new_n8539 = ~pj0 & new_n8538;
  assign new_n8540 = ~pi & new_n8109;
  assign new_n8541 = pt & new_n8540;
  assign new_n8542 = ~pf0 & new_n8541;
  assign new_n8543 = ~pj0 & new_n8542;
  assign new_n8544 = pm0 & new_n8543;
  assign new_n8545 = ~pc0 & new_n8544;
  assign new_n8546 = ~pe0 & new_n8545;
  assign new_n8547 = ~pf0 & new_n8322;
  assign new_n8548 = ~ph0 & new_n8547;
  assign new_n8549 = pm0 & new_n8548;
  assign new_n8550 = ~pe0 & new_n8549;
  assign new_n8551 = ~pj0 & new_n8550;
  assign new_n8552 = ~pa0 & new_n8551;
  assign new_n8553 = ~pc0 & new_n8552;
  assign new_n8554 = ~pg & new_n5841;
  assign new_n8555 = ~ph & new_n8554;
  assign new_n8556 = ~pf & new_n8555;
  assign new_n8557 = pm0 & new_n8556;
  assign new_n8558 = ~pe & new_n8557;
  assign new_n8559 = ~pa0 & new_n8558;
  assign new_n8560 = ~pc0 & new_n8559;
  assign new_n8561 = ~pf & new_n6375;
  assign new_n8562 = ~pg & new_n8561;
  assign new_n8563 = ~pi & new_n8562;
  assign new_n8564 = ~ph0 & new_n8563;
  assign new_n8565 = ~pe & new_n8564;
  assign new_n8566 = ~pf0 & new_n8565;
  assign new_n8567 = ~pj0 & new_n8566;
  assign new_n8568 = pm0 & new_n8567;
  assign new_n8569 = ~pa0 & new_n8568;
  assign new_n8570 = ~pc0 & new_n8569;
  assign new_n8571 = pm & new_n8309;
  assign new_n8572 = pk & new_n8571;
  assign new_n8573 = ~pi & new_n8572;
  assign new_n8574 = ~pd & new_n8573;
  assign new_n8575 = ~ph & new_n8574;
  assign new_n8576 = pm0 & new_n8575;
  assign new_n8577 = ~ph0 & new_n8576;
  assign new_n8578 = ~pc0 & new_n8577;
  assign new_n8579 = ~pe0 & new_n8578;
  assign new_n8580 = pm0 & new_n8151;
  assign new_n8581 = ~ph & new_n8580;
  assign new_n8582 = ~pg0 & new_n8581;
  assign new_n8583 = ~pc0 & new_n8582;
  assign new_n8584 = ~pe0 & new_n8583;
  assign new_n8585 = ~pz & new_n8584;
  assign new_n8586 = ~pa0 & new_n8585;
  assign new_n8587 = ~pd0 & new_n7271;
  assign new_n8588 = ~pm & new_n8587;
  assign new_n8589 = ~pf & new_n8588;
  assign new_n8590 = ~pg & new_n8589;
  assign new_n8591 = ~pe & new_n8590;
  assign new_n8592 = ~pf0 & new_n8591;
  assign new_n8593 = ~ph0 & new_n8592;
  assign new_n8594 = ~pj0 & new_n8593;
  assign new_n8595 = pm0 & new_n8594;
  assign new_n8596 = ~pi & new_n8372;
  assign new_n8597 = ~pj0 & new_n8596;
  assign new_n8598 = ~pc0 & new_n8597;
  assign new_n8599 = ~pe0 & new_n8598;
  assign new_n8600 = ~pz & new_n8599;
  assign new_n8601 = ~pa0 & new_n8600;
  assign new_n8602 = ~pi & new_n6364;
  assign new_n8603 = ~pd & new_n8602;
  assign new_n8604 = pm0 & new_n8603;
  assign new_n8605 = ~ph0 & new_n8604;
  assign new_n8606 = ~pj0 & new_n8605;
  assign new_n8607 = ~pc0 & new_n8606;
  assign new_n8608 = ~pe0 & new_n8607;
  assign new_n8609 = ~py & new_n8608;
  assign new_n8610 = ~pa0 & new_n8609;
  assign new_n8611 = ~pf & new_n8188;
  assign new_n8612 = ~pg & new_n8611;
  assign new_n8613 = ~pe & new_n8612;
  assign new_n8614 = pm0 & new_n8613;
  assign new_n8615 = ~pf0 & new_n8614;
  assign new_n8616 = ~pg0 & new_n8615;
  assign new_n8617 = ~pj0 & new_n8616;
  assign new_n8618 = pn & new_n6098;
  assign new_n8619 = ~pc & new_n8618;
  assign new_n8620 = ~pd0 & new_n8619;
  assign new_n8621 = ~pi0 & new_n8620;
  assign new_n8622 = ~pg & new_n8621;
  assign new_n8623 = ~ph & new_n8622;
  assign new_n8624 = ~pf & new_n8623;
  assign new_n8625 = ~ph0 & new_n8624;
  assign new_n8626 = ~pe & new_n8625;
  assign new_n8627 = pj0 & new_n8626;
  assign new_n8628 = pm0 & new_n8627;
  assign new_n8629 = ~pi & new_n5753;
  assign new_n8630 = pt & new_n8629;
  assign new_n8631 = ~pj0 & new_n8630;
  assign new_n8632 = pm0 & new_n8631;
  assign new_n8633 = ~pe0 & new_n8632;
  assign new_n8634 = ~pa0 & new_n8633;
  assign new_n8635 = ~pc0 & new_n8634;
  assign new_n8636 = ~py & new_n8635;
  assign new_n8637 = ~pz & new_n8636;
  assign new_n8638 = ~pm & new_n6170;
  assign new_n8639 = ~ph & new_n8638;
  assign new_n8640 = ~pi & new_n8639;
  assign new_n8641 = ~pg & new_n8640;
  assign new_n8642 = ~pe & new_n8641;
  assign new_n8643 = ~pf & new_n8642;
  assign new_n8644 = ~pc0 & new_n8643;
  assign new_n8645 = pm0 & new_n8644;
  assign new_n8646 = ~pn & new_n6743;
  assign new_n8647 = ~py & new_n8646;
  assign new_n8648 = pj & new_n8647;
  assign new_n8649 = ~pd & new_n8648;
  assign new_n8650 = pt & new_n8649;
  assign new_n8651 = ~pd0 & new_n8650;
  assign new_n8652 = ~pi & new_n8651;
  assign new_n8653 = pm0 & new_n8652;
  assign new_n8654 = ~ph0 & new_n8653;
  assign new_n8655 = ~pe0 & new_n8654;
  assign new_n8656 = ~pj0 & new_n8655;
  assign new_n8657 = ~pi & new_n7800;
  assign new_n8658 = pt & new_n8657;
  assign new_n8659 = pm0 & new_n8658;
  assign new_n8660 = ~pe0 & new_n8659;
  assign new_n8661 = ~pj0 & new_n8660;
  assign new_n8662 = ~pa0 & new_n8661;
  assign new_n8663 = ~pc0 & new_n8662;
  assign new_n8664 = ~pi & new_n6086;
  assign new_n8665 = ~pk & new_n8664;
  assign new_n8666 = ~ph0 & new_n8665;
  assign new_n8667 = ~pj0 & new_n8666;
  assign new_n8668 = pm0 & new_n8667;
  assign new_n8669 = ~pc0 & new_n8668;
  assign new_n8670 = ~pe0 & new_n8669;
  assign new_n8671 = ~pf0 & new_n8435;
  assign new_n8672 = pm & new_n8671;
  assign new_n8673 = pm0 & new_n8672;
  assign new_n8674 = ~pg0 & new_n8673;
  assign new_n8675 = ~pj0 & new_n8674;
  assign new_n8676 = ~pc0 & new_n8675;
  assign new_n8677 = ~pe0 & new_n8676;
  assign new_n8678 = ~ph & new_n8235;
  assign new_n8679 = pm0 & new_n8678;
  assign new_n8680 = ~ph0 & new_n8679;
  assign new_n8681 = ~pe0 & new_n8680;
  assign new_n8682 = ~pg0 & new_n8681;
  assign new_n8683 = ~pf & new_n8250;
  assign new_n8684 = ~pg & new_n8683;
  assign new_n8685 = pt & new_n8684;
  assign new_n8686 = ~pd & new_n8685;
  assign new_n8687 = ~ph0 & new_n8686;
  assign new_n8688 = ~pe & new_n8687;
  assign new_n8689 = pm0 & new_n8688;
  assign new_n8690 = ~pg0 & new_n8689;
  assign new_n8691 = ~pj0 & new_n8690;
  assign new_n8692 = ~pa0 & new_n8691;
  assign new_n8693 = ~pc0 & new_n8692;
  assign new_n8694 = pm0 & new_n8043;
  assign new_n8695 = ~pg0 & new_n8694;
  assign new_n8696 = ~pj0 & new_n8695;
  assign new_n8697 = ~pz & new_n8696;
  assign new_n8698 = ~pc0 & new_n8697;
  assign new_n8699 = pm0 & new_n6450;
  assign new_n8700 = ~ph0 & new_n8699;
  assign new_n8701 = ~pc0 & new_n8700;
  assign new_n8702 = ~pj0 & new_n8701;
  assign new_n8703 = pm0 & new_n8484;
  assign new_n8704 = ~pc0 & new_n8703;
  assign new_n8705 = ~pj0 & new_n8704;
  assign new_n8706 = ~pz & new_n8705;
  assign new_n8707 = ~pa0 & new_n8706;
  assign new_n8708 = pm0 & new_n8493;
  assign new_n8709 = ~ph0 & new_n8708;
  assign new_n8710 = ~pj0 & new_n8709;
  assign new_n8711 = ~pc0 & new_n8710;
  assign new_n8712 = ~pg0 & new_n8711;
  assign new_n8713 = ~py & new_n8712;
  assign new_n8714 = ~pa0 & new_n8713;
  assign new_n8715 = ~pf & new_n5838;
  assign new_n8716 = ~pg & new_n8715;
  assign new_n8717 = ~pt & new_n8716;
  assign new_n8718 = ~pd0 & new_n8717;
  assign new_n8719 = ~pf0 & new_n8718;
  assign new_n8720 = ~pe & new_n8719;
  assign new_n8721 = pm0 & new_n8720;
  assign new_n8722 = ~pg0 & new_n8721;
  assign new_n8723 = ~pj0 & new_n8722;
  assign new_n8724 = ~pa0 & new_n8723;
  assign new_n8725 = ~pc0 & new_n8724;
  assign new_n8726 = ~pm & new_n7208;
  assign new_n8727 = ~pk & new_n8726;
  assign new_n8728 = ~pg & new_n8727;
  assign new_n8729 = ~pi & new_n8728;
  assign new_n8730 = ~pf & new_n8729;
  assign new_n8731 = ~ph0 & new_n8730;
  assign new_n8732 = ~pe & new_n8731;
  assign new_n8733 = ~pj0 & new_n8732;
  assign new_n8734 = pm0 & new_n8733;
  assign new_n8735 = ~pb & new_n8664;
  assign new_n8736 = ~pk & new_n8735;
  assign new_n8737 = ~pf & new_n8736;
  assign new_n8738 = ~pg & new_n8737;
  assign new_n8739 = ~pe & new_n8738;
  assign new_n8740 = pm0 & new_n8739;
  assign new_n8741 = ~ph0 & new_n8740;
  assign new_n8742 = ~pc0 & new_n8741;
  assign new_n8743 = ~pj0 & new_n8742;
  assign new_n8744 = ~pi & new_n6158;
  assign new_n8745 = ~pd0 & new_n8744;
  assign new_n8746 = ~pk & new_n8745;
  assign new_n8747 = ~pf & new_n8746;
  assign new_n8748 = ~pg & new_n8747;
  assign new_n8749 = ~pe & new_n8748;
  assign new_n8750 = pm0 & new_n8749;
  assign new_n8751 = ~pf0 & new_n8750;
  assign new_n8752 = ~pc0 & new_n8751;
  assign new_n8753 = ~pj0 & new_n8752;
  assign new_n8754 = ~ph0 & new_n6900;
  assign new_n8755 = pt & new_n8754;
  assign new_n8756 = ~pf0 & new_n8755;
  assign new_n8757 = ~pj0 & new_n8756;
  assign new_n8758 = pm0 & new_n8757;
  assign new_n8759 = ~pe0 & new_n8758;
  assign new_n8760 = ~pg0 & new_n8759;
  assign new_n8761 = pm0 & new_n6913;
  assign new_n8762 = ~pf0 & new_n8761;
  assign new_n8763 = ~pj0 & new_n8762;
  assign new_n8764 = ~pe0 & new_n8763;
  assign new_n8765 = ~pg0 & new_n8764;
  assign new_n8766 = ~pa0 & new_n8765;
  assign new_n8767 = ~pc0 & new_n8766;
  assign new_n8768 = ~ph & new_n8502;
  assign new_n8769 = ~pt & new_n8768;
  assign new_n8770 = ~pd0 & new_n8769;
  assign new_n8771 = ~pf & new_n8770;
  assign new_n8772 = ~pg & new_n8771;
  assign new_n8773 = ~pe & new_n8772;
  assign new_n8774 = pm0 & new_n8773;
  assign new_n8775 = ~ph0 & new_n8774;
  assign new_n8776 = ~pc0 & new_n8775;
  assign new_n8777 = ~pg0 & new_n8776;
  assign new_n8778 = ~pl & new_n5889;
  assign new_n8779 = ~pc & new_n8778;
  assign new_n8780 = ~pg & new_n8779;
  assign new_n8781 = ~ph & new_n8780;
  assign new_n8782 = ~pt & new_n8781;
  assign new_n8783 = ~pe & new_n8782;
  assign new_n8784 = ~pf & new_n8783;
  assign new_n8785 = pm0 & new_n8784;
  assign new_n8786 = ~pc0 & new_n8785;
  assign new_n8787 = ~pg0 & new_n8786;
  assign new_n8788 = ~pz & new_n8787;
  assign new_n8789 = ~pa0 & new_n8788;
  assign new_n8790 = pm & new_n7238;
  assign new_n8791 = pk & new_n8790;
  assign new_n8792 = ~pi & new_n8791;
  assign new_n8793 = ~pd & new_n8792;
  assign new_n8794 = ~ph & new_n8793;
  assign new_n8795 = ~pe0 & new_n8794;
  assign new_n8796 = pm0 & new_n8795;
  assign new_n8797 = ~pa0 & new_n8796;
  assign new_n8798 = ~pc0 & new_n8797;
  assign new_n8799 = ~ph0 & new_n8151;
  assign new_n8800 = ~ph & new_n8799;
  assign new_n8801 = pm0 & new_n8800;
  assign new_n8802 = ~pe0 & new_n8801;
  assign new_n8803 = ~pg0 & new_n8802;
  assign new_n8804 = ~pa0 & new_n8803;
  assign new_n8805 = ~pc0 & new_n8804;
  assign new_n8806 = ~pf & new_n6942;
  assign new_n8807 = ~pg & new_n8806;
  assign new_n8808 = ~pe & new_n8807;
  assign new_n8809 = pm0 & new_n8808;
  assign new_n8810 = ~pf0 & new_n8809;
  assign new_n8811 = ~pg0 & new_n8810;
  assign new_n8812 = ~pj0 & new_n8811;
  assign new_n8813 = ~ph0 & new_n8171;
  assign new_n8814 = ~pi & new_n8813;
  assign new_n8815 = pm0 & new_n8814;
  assign new_n8816 = ~pe0 & new_n8815;
  assign new_n8817 = ~pj0 & new_n8816;
  assign new_n8818 = ~pa0 & new_n8817;
  assign new_n8819 = ~pc0 & new_n8818;
  assign new_n8820 = ~pj0 & new_n8603;
  assign new_n8821 = pm0 & new_n8820;
  assign new_n8822 = ~pe0 & new_n8821;
  assign new_n8823 = ~pa0 & new_n8822;
  assign new_n8824 = ~pc0 & new_n8823;
  assign new_n8825 = ~py & new_n8824;
  assign new_n8826 = ~pz & new_n8825;
  assign new_n8827 = ~pb & new_n8587;
  assign new_n8828 = ~pf & new_n8827;
  assign new_n8829 = ~pg & new_n8828;
  assign new_n8830 = ~pe & new_n8829;
  assign new_n8831 = ~pf0 & new_n8830;
  assign new_n8832 = ~ph0 & new_n8831;
  assign new_n8833 = ~pj0 & new_n8832;
  assign new_n8834 = pm0 & new_n8833;
  assign new_n8835 = pn & new_n5876;
  assign new_n8836 = ~pc & new_n8835;
  assign new_n8837 = ~pd0 & new_n8836;
  assign new_n8838 = ~pi0 & new_n8837;
  assign new_n8839 = ~pg & new_n8838;
  assign new_n8840 = ~ph & new_n8839;
  assign new_n8841 = ~pf & new_n8840;
  assign new_n8842 = pm0 & new_n8841;
  assign new_n8843 = ~pe & new_n8842;
  assign new_n8844 = ~pg0 & new_n8843;
  assign new_n8845 = pj0 & new_n8844;
  assign new_n8846 = pm0 & new_n8630;
  assign new_n8847 = ~ph0 & new_n8846;
  assign new_n8848 = ~pj0 & new_n8847;
  assign new_n8849 = ~pc0 & new_n8848;
  assign new_n8850 = ~pe0 & new_n8849;
  assign new_n8851 = ~py & new_n8850;
  assign new_n8852 = ~pa0 & new_n8851;
  assign new_n8853 = ~pg & new_n7343;
  assign new_n8854 = ~ph & new_n8853;
  assign new_n8855 = ~pf & new_n8854;
  assign new_n8856 = ~ph0 & new_n8855;
  assign new_n8857 = ~pe & new_n8856;
  assign new_n8858 = ~pg0 & new_n8857;
  assign new_n8859 = pm0 & new_n8858;
  assign new_n8860 = pm0 & new_n7678;
  assign new_n8861 = ~pg0 & new_n8860;
  assign new_n8862 = ~pj0 & new_n8861;
  assign new_n8863 = ~pc0 & new_n8862;
  assign new_n8864 = ~pe0 & new_n8863;
  assign new_n8865 = ~ph0 & new_n8427;
  assign new_n8866 = pt & new_n8865;
  assign new_n8867 = pm0 & new_n8866;
  assign new_n8868 = ~pg0 & new_n8867;
  assign new_n8869 = ~pj0 & new_n8868;
  assign new_n8870 = ~pc0 & new_n8869;
  assign new_n8871 = ~pe0 & new_n8870;
  assign new_n8872 = pm0 & new_n8437;
  assign new_n8873 = ~pg0 & new_n8872;
  assign new_n8874 = ~pj0 & new_n8873;
  assign new_n8875 = ~pc0 & new_n8874;
  assign new_n8876 = ~pe0 & new_n8875;
  assign new_n8877 = ~py & new_n6396;
  assign new_n8878 = ~pc0 & new_n8877;
  assign new_n8879 = pj & new_n8878;
  assign new_n8880 = ~pk & new_n8879;
  assign new_n8881 = pi0 & new_n8880;
  assign new_n8882 = ~pi & new_n8881;
  assign new_n8883 = ~pd0 & new_n8882;
  assign new_n8884 = pm0 & new_n8883;
  assign new_n8885 = ~ph0 & new_n8884;
  assign new_n8886 = ~pi & new_n8436;
  assign new_n8887 = pm0 & new_n8886;
  assign new_n8888 = ~ph & new_n8887;
  assign new_n8889 = ~pc0 & new_n8888;
  assign new_n8890 = ~pe0 & new_n8889;
  assign new_n8891 = pm0 & new_n8686;
  assign new_n8892 = ~pe & new_n8891;
  assign new_n8893 = ~pj0 & new_n8892;
  assign new_n8894 = ~pc0 & new_n8893;
  assign new_n8895 = ~pg0 & new_n8894;
  assign new_n8896 = ~pz & new_n8895;
  assign new_n8897 = ~pa0 & new_n8896;
  assign new_n8898 = ~pd0 & new_n6608;
  assign new_n8899 = pi0 & new_n8898;
  assign new_n8900 = ~ph0 & new_n8899;
  assign new_n8901 = ~pe & new_n8900;
  assign new_n8902 = pm0 & new_n8901;
  assign new_n8903 = ~pg0 & new_n8902;
  assign new_n8904 = ~pj0 & new_n8903;
  assign new_n8905 = ~py & new_n8904;
  assign new_n8906 = ~pc0 & new_n8905;
  assign new_n8907 = ~pi & new_n7030;
  assign new_n8908 = pt & new_n8907;
  assign new_n8909 = ~pd0 & new_n8908;
  assign new_n8910 = ~pe & new_n8909;
  assign new_n8911 = ~pf & new_n8910;
  assign new_n8912 = ~ph0 & new_n8911;
  assign new_n8913 = ~pj0 & new_n8912;
  assign new_n8914 = pm0 & new_n8913;
  assign new_n8915 = ~pa0 & new_n8914;
  assign new_n8916 = ~pc0 & new_n8915;
  assign new_n8917 = ~pe & new_n6260;
  assign new_n8918 = ~pf & new_n8917;
  assign new_n8919 = ~pg & new_n8918;
  assign new_n8920 = pt & new_n8919;
  assign new_n8921 = ~pj0 & new_n8920;
  assign new_n8922 = pm0 & new_n8921;
  assign new_n8923 = ~pg0 & new_n8922;
  assign new_n8924 = ~pa0 & new_n8923;
  assign new_n8925 = ~pc0 & new_n8924;
  assign new_n8926 = ~py & new_n8925;
  assign new_n8927 = ~pz & new_n8926;
  assign new_n8928 = ~pf & new_n8331;
  assign new_n8929 = ~pg & new_n8928;
  assign new_n8930 = ~pd0 & new_n8929;
  assign new_n8931 = pd & new_n8930;
  assign new_n8932 = ~ph0 & new_n8931;
  assign new_n8933 = ~pe & new_n8932;
  assign new_n8934 = ~pf0 & new_n8933;
  assign new_n8935 = ~pj0 & new_n8934;
  assign new_n8936 = pm0 & new_n8935;
  assign new_n8937 = ~pc0 & new_n8936;
  assign new_n8938 = ~pg0 & new_n8937;
  assign new_n8939 = ~pf & new_n8779;
  assign new_n8940 = ~pg & new_n8939;
  assign new_n8941 = ~pi & new_n8940;
  assign new_n8942 = ~pt & new_n8941;
  assign new_n8943 = ~ph0 & new_n8942;
  assign new_n8944 = ~pe & new_n8943;
  assign new_n8945 = ~pf0 & new_n8944;
  assign new_n8946 = ~pj0 & new_n8945;
  assign new_n8947 = pm0 & new_n8946;
  assign new_n8948 = ~pa0 & new_n8947;
  assign new_n8949 = ~pc0 & new_n8948;
  assign new_n8950 = ~pf & new_n8515;
  assign new_n8951 = ~pg & new_n8950;
  assign new_n8952 = ~pe & new_n8951;
  assign new_n8953 = ~pj0 & new_n8952;
  assign new_n8954 = pm0 & new_n8953;
  assign new_n8955 = ~pc0 & new_n8954;
  assign new_n8956 = ~pg0 & new_n8955;
  assign new_n8957 = ~pb & new_n7863;
  assign new_n8958 = ~pk & new_n8957;
  assign new_n8959 = ~pf & new_n8958;
  assign new_n8960 = ~pg & new_n8959;
  assign new_n8961 = ~pe & new_n8960;
  assign new_n8962 = ~pj0 & new_n8961;
  assign new_n8963 = pm0 & new_n8962;
  assign new_n8964 = ~pa0 & new_n8963;
  assign new_n8965 = ~pc0 & new_n8964;
  assign new_n8966 = ~pg & new_n5939;
  assign new_n8967 = ~pi & new_n8966;
  assign new_n8968 = ~pk & new_n8967;
  assign new_n8969 = ~pe & new_n8968;
  assign new_n8970 = ~pf & new_n8969;
  assign new_n8971 = ~ph0 & new_n8970;
  assign new_n8972 = pm0 & new_n8971;
  assign new_n8973 = ~pf0 & new_n8972;
  assign new_n8974 = ~pc0 & new_n8973;
  assign new_n8975 = ~pj0 & new_n8974;
  assign new_n8976 = ~pd0 & new_n6046;
  assign new_n8977 = pi0 & new_n8976;
  assign new_n8978 = pd & new_n8977;
  assign new_n8979 = ~ph & new_n8978;
  assign new_n8980 = ~pi & new_n8979;
  assign new_n8981 = ~pg & new_n8980;
  assign new_n8982 = ~pe & new_n8981;
  assign new_n8983 = ~pf & new_n8982;
  assign new_n8984 = ~pc0 & new_n8983;
  assign new_n8985 = pm0 & new_n8984;
  assign new_n8986 = ~pl & new_n5926;
  assign new_n8987 = ~pc & new_n8986;
  assign new_n8988 = ~pt & new_n8987;
  assign new_n8989 = ~pd0 & new_n8988;
  assign new_n8990 = ~pi0 & new_n8989;
  assign new_n8991 = ~ph & new_n8990;
  assign new_n8992 = ~pi & new_n8991;
  assign new_n8993 = ~pg & new_n8992;
  assign new_n8994 = ~pe & new_n8993;
  assign new_n8995 = ~pf & new_n8994;
  assign new_n8996 = pm0 & new_n8995;
  assign new_n8997 = ~ph0 & new_n8996;
  assign new_n8998 = ~pd0 & new_n6133;
  assign new_n8999 = pi0 & new_n8998;
  assign new_n9000 = ~pe & new_n8999;
  assign new_n9001 = ~pf & new_n9000;
  assign new_n9002 = ~pf0 & new_n9001;
  assign new_n9003 = ~pj0 & new_n9002;
  assign new_n9004 = pm0 & new_n9003;
  assign new_n9005 = ~pc0 & new_n9004;
  assign new_n9006 = ~pg0 & new_n9005;
  assign new_n9007 = ~ph0 & new_n8784;
  assign new_n9008 = ~pg0 & new_n9007;
  assign new_n9009 = pm0 & new_n9008;
  assign new_n9010 = ~pa0 & new_n9009;
  assign new_n9011 = ~pc0 & new_n9010;
  assign new_n9012 = ~pf0 & new_n8563;
  assign new_n9013 = ~pe & new_n9012;
  assign new_n9014 = pm0 & new_n9013;
  assign new_n9015 = ~pc0 & new_n9014;
  assign new_n9016 = ~pj0 & new_n9015;
  assign new_n9017 = ~pz & new_n9016;
  assign new_n9018 = ~pa0 & new_n9017;
  assign new_n9019 = ~pd0 & new_n8096;
  assign new_n9020 = ~pk & new_n9019;
  assign new_n9021 = ~ph & new_n9020;
  assign new_n9022 = ~pi & new_n9021;
  assign new_n9023 = ~pg & new_n9022;
  assign new_n9024 = ~pe & new_n9023;
  assign new_n9025 = ~pf & new_n9024;
  assign new_n9026 = pm0 & new_n9025;
  assign new_n9027 = ~ph0 & new_n9026;
  assign new_n9028 = ~ph & new_n8572;
  assign new_n9029 = ~pd & new_n9028;
  assign new_n9030 = ~ph0 & new_n9029;
  assign new_n9031 = ~pg0 & new_n9030;
  assign new_n9032 = pm0 & new_n9031;
  assign new_n9033 = ~pc0 & new_n9032;
  assign new_n9034 = ~pe0 & new_n9033;
  assign new_n9035 = ~pz & new_n7591;
  assign new_n9036 = ~pc & new_n9035;
  assign new_n9037 = pi0 & new_n9036;
  assign new_n9038 = ~pm & new_n9037;
  assign new_n9039 = ~pi & new_n9038;
  assign new_n9040 = ~pd0 & new_n9039;
  assign new_n9041 = ~pg & new_n9040;
  assign new_n9042 = ~pe & new_n9041;
  assign new_n9043 = ~pf & new_n9042;
  assign new_n9044 = pm0 & new_n9043;
  assign new_n9045 = ~pf0 & new_n9044;
  assign new_n9046 = ~pi & new_n7669;
  assign new_n9047 = pt & new_n9046;
  assign new_n9048 = ~ph0 & new_n9047;
  assign new_n9049 = ~pj0 & new_n9048;
  assign new_n9050 = pm0 & new_n9049;
  assign new_n9051 = ~pc0 & new_n9050;
  assign new_n9052 = ~pe0 & new_n9051;
  assign new_n9053 = pj & new_n8118;
  assign new_n9054 = pt & new_n9053;
  assign new_n9055 = pm & new_n9054;
  assign new_n9056 = ~pj0 & new_n9055;
  assign new_n9057 = pm0 & new_n9056;
  assign new_n9058 = ~pg0 & new_n9057;
  assign new_n9059 = ~pc0 & new_n9058;
  assign new_n9060 = ~pe0 & new_n9059;
  assign new_n9061 = ~pz & new_n9060;
  assign new_n9062 = ~pa0 & new_n9061;
  assign new_n9063 = ~ph0 & new_n6555;
  assign new_n9064 = pm & new_n9063;
  assign new_n9065 = ~pj0 & new_n9064;
  assign new_n9066 = pm0 & new_n9065;
  assign new_n9067 = ~pg0 & new_n9066;
  assign new_n9068 = ~pc0 & new_n9067;
  assign new_n9069 = ~pe0 & new_n9068;
  assign new_n9070 = ~py & new_n9069;
  assign new_n9071 = ~pa0 & new_n9070;
  assign new_n9072 = ~pb & new_n9037;
  assign new_n9073 = ~pi & new_n9072;
  assign new_n9074 = ~pd0 & new_n9073;
  assign new_n9075 = ~pg & new_n9074;
  assign new_n9076 = ~pe & new_n9075;
  assign new_n9077 = ~pf & new_n9076;
  assign new_n9078 = pm0 & new_n9077;
  assign new_n9079 = ~pf0 & new_n9078;
  assign new_n9080 = pn & new_n5926;
  assign new_n9081 = ~pc & new_n9080;
  assign new_n9082 = ~pd0 & new_n9081;
  assign new_n9083 = ~pi0 & new_n9082;
  assign new_n9084 = ~ph & new_n9083;
  assign new_n9085 = ~pi & new_n9084;
  assign new_n9086 = ~pg & new_n9085;
  assign new_n9087 = ~pe & new_n9086;
  assign new_n9088 = ~pf & new_n9087;
  assign new_n9089 = pm0 & new_n9088;
  assign new_n9090 = ~ph0 & new_n9089;
  assign new_n9091 = ~ph & new_n5950;
  assign new_n9092 = ~pd0 & new_n9091;
  assign new_n9093 = ~pf & new_n9092;
  assign new_n9094 = ~pg & new_n9093;
  assign new_n9095 = ~pe & new_n9094;
  assign new_n9096 = ~pg0 & new_n9095;
  assign new_n9097 = pm0 & new_n9096;
  assign new_n9098 = ~pa0 & new_n9097;
  assign new_n9099 = ~pc0 & new_n9098;
  assign new_n9100 = ~pg & new_n8638;
  assign new_n9101 = ~ph & new_n9100;
  assign new_n9102 = ~pf & new_n9101;
  assign new_n9103 = pm0 & new_n9102;
  assign new_n9104 = ~pe & new_n9103;
  assign new_n9105 = ~pc0 & new_n9104;
  assign new_n9106 = ~pg0 & new_n9105;
  assign new_n9107 = ~ph0 & new_n8651;
  assign new_n9108 = ~pj0 & new_n9107;
  assign new_n9109 = pm0 & new_n9108;
  assign new_n9110 = ~pe0 & new_n9109;
  assign new_n9111 = ~pg0 & new_n9110;
  assign new_n9112 = ~pb & new_n5972;
  assign new_n9113 = ~pd0 & new_n9112;
  assign new_n9114 = pi0 & new_n9113;
  assign new_n9115 = ~pi & new_n9114;
  assign new_n9116 = ~pg & new_n9115;
  assign new_n9117 = ~ph & new_n9116;
  assign new_n9118 = ~pe & new_n9117;
  assign new_n9119 = ~pf & new_n9118;
  assign new_n9120 = ~pi & new_n7705;
  assign new_n9121 = pm0 & new_n9120;
  assign new_n9122 = ~ph0 & new_n9121;
  assign new_n9123 = ~pe0 & new_n9122;
  assign new_n9124 = ~pj0 & new_n9123;
  assign new_n9125 = ~pi & new_n8435;
  assign new_n9126 = pm & new_n9125;
  assign new_n9127 = ~pf0 & new_n9126;
  assign new_n9128 = ~pj0 & new_n9127;
  assign new_n9129 = pm0 & new_n9128;
  assign new_n9130 = ~pc0 & new_n9129;
  assign new_n9131 = ~pe0 & new_n9130;
  assign new_n9132 = ~pi & new_n8235;
  assign new_n9133 = ~ph0 & new_n9132;
  assign new_n9134 = ~ph & new_n9133;
  assign new_n9135 = ~pe0 & new_n9134;
  assign new_n9136 = pm0 & new_n9135;
  assign new_n9137 = ~pf & new_n7978;
  assign new_n9138 = ~pg & new_n9137;
  assign new_n9139 = ~pi & new_n9138;
  assign new_n9140 = ~pd & new_n9139;
  assign new_n9141 = ~ph0 & new_n9140;
  assign new_n9142 = ~pe & new_n9141;
  assign new_n9143 = pm0 & new_n9142;
  assign new_n9144 = ~pc0 & new_n9143;
  assign new_n9145 = ~pj0 & new_n9144;
  assign new_n9146 = ~py & new_n9145;
  assign new_n9147 = ~pa0 & new_n9146;
  assign new_n9148 = pm0 & new_n8467;
  assign new_n9149 = ~pc0 & new_n9148;
  assign new_n9150 = ~pj0 & new_n9149;
  assign new_n9151 = ~py & new_n9150;
  assign new_n9152 = ~pz & new_n9151;
  assign new_n9153 = pm0 & new_n8911;
  assign new_n9154 = ~pc0 & new_n9153;
  assign new_n9155 = ~pj0 & new_n9154;
  assign new_n9156 = ~pz & new_n9155;
  assign new_n9157 = ~pa0 & new_n9156;
  assign new_n9158 = pm0 & new_n8920;
  assign new_n9159 = ~ph0 & new_n9158;
  assign new_n9160 = ~pj0 & new_n9159;
  assign new_n9161 = ~pc0 & new_n9160;
  assign new_n9162 = ~pg0 & new_n9161;
  assign new_n9163 = ~py & new_n9162;
  assign new_n9164 = ~pa0 & new_n9163;
  assign new_n9165 = ~pg & new_n8502;
  assign new_n9166 = ~pi & new_n9165;
  assign new_n9167 = ~pt & new_n9166;
  assign new_n9168 = ~pd0 & new_n9167;
  assign new_n9169 = ~pe & new_n9168;
  assign new_n9170 = ~pf & new_n9169;
  assign new_n9171 = ~ph0 & new_n9170;
  assign new_n9172 = pm0 & new_n9171;
  assign new_n9173 = ~pf0 & new_n9172;
  assign new_n9174 = ~pc0 & new_n9173;
  assign new_n9175 = ~pj0 & new_n9174;
  assign new_n9176 = ~pf0 & new_n8942;
  assign new_n9177 = ~pe & new_n9176;
  assign new_n9178 = pm0 & new_n9177;
  assign new_n9179 = ~pc0 & new_n9178;
  assign new_n9180 = ~pj0 & new_n9179;
  assign new_n9181 = ~pz & new_n9180;
  assign new_n9182 = ~pa0 & new_n9181;
  assign new_n9183 = ~pf & new_n8727;
  assign new_n9184 = ~pg & new_n9183;
  assign new_n9185 = ~pe & new_n9184;
  assign new_n9186 = pm0 & new_n9185;
  assign new_n9187 = ~ph0 & new_n9186;
  assign new_n9188 = ~pg0 & new_n9187;
  assign new_n9189 = ~pj0 & new_n9188;
  assign new_n9190 = ~pb & new_n6087;
  assign new_n9191 = ~pk & new_n9190;
  assign new_n9192 = ~pe & new_n9191;
  assign new_n9193 = ~pf & new_n9192;
  assign new_n9194 = ~ph0 & new_n9193;
  assign new_n9195 = ~pj0 & new_n9194;
  assign new_n9196 = pm0 & new_n9195;
  assign new_n9197 = ~pc0 & new_n9196;
  assign new_n9198 = ~pg0 & new_n9197;
  assign new_n9199 = ~pg & new_n6158;
  assign new_n9200 = ~pd0 & new_n9199;
  assign new_n9201 = ~pk & new_n9200;
  assign new_n9202 = ~pe & new_n9201;
  assign new_n9203 = ~pf & new_n9202;
  assign new_n9204 = ~pf0 & new_n9203;
  assign new_n9205 = ~pj0 & new_n9204;
  assign new_n9206 = pm0 & new_n9205;
  assign new_n9207 = ~pc0 & new_n9206;
  assign new_n9208 = ~pg0 & new_n9207;
  assign new_n9209 = ~pg & new_n6498;
  assign new_n9210 = ~ph & new_n9209;
  assign new_n9211 = ~pf & new_n9210;
  assign new_n9212 = ~ph0 & new_n9211;
  assign new_n9213 = ~pe & new_n9212;
  assign new_n9214 = ~pg0 & new_n9213;
  assign new_n9215 = pm0 & new_n9214;
  assign new_n9216 = pm0 & new_n6318;
  assign new_n9217 = ~pc0 & new_n9216;
  assign new_n9218 = ~pg0 & new_n9217;
  assign new_n9219 = ~pz & new_n9218;
  assign new_n9220 = ~pa0 & new_n9219;
  assign new_n9221 = ~pi & new_n8502;
  assign new_n9222 = ~pt & new_n9221;
  assign new_n9223 = ~pd0 & new_n9222;
  assign new_n9224 = ~pg & new_n9223;
  assign new_n9225 = ~ph & new_n9224;
  assign new_n9226 = ~pf & new_n9225;
  assign new_n9227 = ~ph0 & new_n9226;
  assign new_n9228 = ~pe & new_n9227;
  assign new_n9229 = ~pc0 & new_n9228;
  assign new_n9230 = pm0 & new_n9229;
  assign new_n9231 = ~ph & new_n8779;
  assign new_n9232 = ~pi & new_n9231;
  assign new_n9233 = ~pt & new_n9232;
  assign new_n9234 = ~pf & new_n9233;
  assign new_n9235 = ~pg & new_n9234;
  assign new_n9236 = ~pe & new_n9235;
  assign new_n9237 = ~pc0 & new_n9236;
  assign new_n9238 = pm0 & new_n9237;
  assign new_n9239 = ~pz & new_n9238;
  assign new_n9240 = ~pa0 & new_n9239;
  assign new_n9241 = ~pe & new_n6375;
  assign new_n9242 = ~pf & new_n9241;
  assign new_n9243 = ~pg & new_n9242;
  assign new_n9244 = ~pf0 & new_n9243;
  assign new_n9245 = ~ph0 & new_n9244;
  assign new_n9246 = pm0 & new_n9245;
  assign new_n9247 = ~pg0 & new_n9246;
  assign new_n9248 = ~pj0 & new_n9247;
  assign new_n9249 = ~pa0 & new_n9248;
  assign new_n9250 = ~pc0 & new_n9249;
  assign new_n9251 = ~ph & new_n6735;
  assign new_n9252 = ~pd0 & new_n9251;
  assign new_n9253 = ~pg & new_n9252;
  assign new_n9254 = ~pe & new_n9253;
  assign new_n9255 = ~pf & new_n9254;
  assign new_n9256 = ~pg0 & new_n9255;
  assign new_n9257 = pm0 & new_n9256;
  assign new_n9258 = ~ph & new_n8791;
  assign new_n9259 = ~pd & new_n9258;
  assign new_n9260 = pm0 & new_n9259;
  assign new_n9261 = ~pe0 & new_n9260;
  assign new_n9262 = ~pg0 & new_n9261;
  assign new_n9263 = ~pa0 & new_n9262;
  assign new_n9264 = ~pc0 & new_n9263;
  assign new_n9265 = ~py & new_n7822;
  assign new_n9266 = ~pc0 & new_n9265;
  assign new_n9267 = ~pc & new_n9266;
  assign new_n9268 = pi0 & new_n9267;
  assign new_n9269 = ~pm & new_n9268;
  assign new_n9270 = ~pi & new_n9269;
  assign new_n9271 = ~pd0 & new_n9270;
  assign new_n9272 = ~pg & new_n9271;
  assign new_n9273 = ~pe & new_n9272;
  assign new_n9274 = ~pf & new_n9273;
  assign new_n9275 = ~pf0 & new_n9274;
  assign new_n9276 = ~ph0 & new_n9275;
  assign new_n9277 = ~pi & new_n6760;
  assign new_n9278 = pt & new_n9277;
  assign new_n9279 = pm0 & new_n9278;
  assign new_n9280 = ~pe0 & new_n9279;
  assign new_n9281 = ~pj0 & new_n9280;
  assign new_n9282 = ~pa0 & new_n9281;
  assign new_n9283 = ~pc0 & new_n9282;
  assign new_n9284 = pm0 & new_n9055;
  assign new_n9285 = ~ph0 & new_n9284;
  assign new_n9286 = ~pj0 & new_n9285;
  assign new_n9287 = ~pe0 & new_n9286;
  assign new_n9288 = ~pg0 & new_n9287;
  assign new_n9289 = ~pa0 & new_n9288;
  assign new_n9290 = ~pc0 & new_n9289;
  assign new_n9291 = pm0 & new_n6555;
  assign new_n9292 = pm & new_n9291;
  assign new_n9293 = ~pg0 & new_n9292;
  assign new_n9294 = ~pj0 & new_n9293;
  assign new_n9295 = ~pe0 & new_n9294;
  assign new_n9296 = ~pa0 & new_n9295;
  assign new_n9297 = ~pc0 & new_n9296;
  assign new_n9298 = ~py & new_n9297;
  assign new_n9299 = ~pz & new_n9298;
  assign new_n9300 = ~pb & new_n9268;
  assign new_n9301 = ~pi & new_n9300;
  assign new_n9302 = ~pd0 & new_n9301;
  assign new_n9303 = ~pg & new_n9302;
  assign new_n9304 = ~pe & new_n9303;
  assign new_n9305 = ~pf & new_n9304;
  assign new_n9306 = ~pf0 & new_n9305;
  assign new_n9307 = ~ph0 & new_n9306;
  assign new_n9308 = ~ph & new_n8838;
  assign new_n9309 = ~pi & new_n9308;
  assign new_n9310 = ~pg & new_n9309;
  assign new_n9311 = ~pe & new_n9310;
  assign new_n9312 = ~pf & new_n9311;
  assign new_n9313 = pj0 & new_n9312;
  assign new_n9314 = pm0 & new_n9313;
  assign new_n9315 = ~ph & new_n5914;
  assign new_n9316 = ~pd0 & new_n9315;
  assign new_n9317 = ~pf & new_n9316;
  assign new_n9318 = ~pg & new_n9317;
  assign new_n9319 = ~pe & new_n9318;
  assign new_n9320 = pm0 & new_n9319;
  assign new_n9321 = ~ph0 & new_n9320;
  assign new_n9322 = ~pc0 & new_n9321;
  assign new_n9323 = ~pg0 & new_n9322;
  assign new_n9324 = ~pn & new_n7122;
  assign new_n9325 = ~py & new_n9324;
  assign new_n9326 = pj & new_n9325;
  assign new_n9327 = ~pd & new_n9326;
  assign new_n9328 = ~pd0 & new_n9327;
  assign new_n9329 = pi0 & new_n9328;
  assign new_n9330 = pt & new_n9329;
  assign new_n9331 = ~ph0 & new_n9330;
  assign new_n9332 = ~pi & new_n9331;
  assign new_n9333 = ~pj0 & new_n9332;
  assign new_n9334 = pm0 & new_n9333;
  assign new_n9335 = ~pn & new_n6155;
  assign new_n9336 = ~py & new_n9335;
  assign new_n9337 = pj & new_n9336;
  assign new_n9338 = ~pd & new_n9337;
  assign new_n9339 = pt & new_n9338;
  assign new_n9340 = ~pd0 & new_n9339;
  assign new_n9341 = ~pi & new_n9340;
  assign new_n9342 = ~pj0 & new_n9341;
  assign new_n9343 = pm0 & new_n9342;
  assign new_n9344 = ~pc0 & new_n9343;
  assign new_n9345 = ~pe0 & new_n9344;
  assign new_n9346 = ~pb & new_n6573;
  assign new_n9347 = ~pd0 & new_n9346;
  assign new_n9348 = pi0 & new_n9347;
  assign new_n9349 = ~ph & new_n9348;
  assign new_n9350 = ~pf & new_n9349;
  assign new_n9351 = ~pg & new_n9350;
  assign new_n9352 = ~ph0 & new_n9351;
  assign new_n9353 = ~pe & new_n9352;
  assign new_n9354 = ~pb & new_n6170;
  assign new_n9355 = ~pg & new_n9354;
  assign new_n9356 = ~ph & new_n9355;
  assign new_n9357 = ~pf & new_n9356;
  assign new_n9358 = pm0 & new_n9357;
  assign new_n9359 = ~pe & new_n9358;
  assign new_n9360 = ~pc0 & new_n9359;
  assign new_n9361 = ~pg0 & new_n9360;
  assign new_n9362 = ~ph0 & new_n7933;
  assign new_n9363 = pm & new_n9362;
  assign new_n9364 = ~pf0 & new_n9363;
  assign new_n9365 = ~pj0 & new_n9364;
  assign new_n9366 = pm0 & new_n9365;
  assign new_n9367 = ~pe0 & new_n9366;
  assign new_n9368 = ~pg0 & new_n9367;
  assign new_n9369 = ~pj0 & new_n7817;
  assign new_n9370 = pm0 & new_n9369;
  assign new_n9371 = ~pe0 & new_n9370;
  assign new_n9372 = ~pg0 & new_n9371;
  assign new_n9373 = pm0 & new_n9140;
  assign new_n9374 = ~pe & new_n9373;
  assign new_n9375 = ~pj0 & new_n9374;
  assign new_n9376 = ~pa0 & new_n9375;
  assign new_n9377 = ~pc0 & new_n9376;
  assign new_n9378 = ~py & new_n9377;
  assign new_n9379 = ~pz & new_n9378;
  assign new_n9380 = ~ph0 & new_n6017;
  assign new_n9381 = ~pj0 & new_n9380;
  assign new_n9382 = pm0 & new_n9381;
  assign new_n9383 = ~pa0 & new_n9382;
  assign new_n9384 = ~pc0 & new_n9383;
  assign new_n9385 = ~ph0 & new_n6657;
  assign new_n9386 = ~pe & new_n9385;
  assign new_n9387 = pm0 & new_n9386;
  assign new_n9388 = ~pg0 & new_n9387;
  assign new_n9389 = ~pj0 & new_n9388;
  assign new_n9390 = ~pa0 & new_n9389;
  assign new_n9391 = ~pc0 & new_n9390;
  assign new_n9392 = ~pg & new_n8331;
  assign new_n9393 = ~pi & new_n9392;
  assign new_n9394 = ~pd0 & new_n9393;
  assign new_n9395 = pd & new_n9394;
  assign new_n9396 = ~pe & new_n9395;
  assign new_n9397 = ~pf & new_n9396;
  assign new_n9398 = ~ph0 & new_n9397;
  assign new_n9399 = pm0 & new_n9398;
  assign new_n9400 = ~pf0 & new_n9399;
  assign new_n9401 = ~pc0 & new_n9400;
  assign new_n9402 = ~pj0 & new_n9401;
  assign new_n9403 = ~pt & new_n8284;
  assign new_n9404 = ~pd0 & new_n9403;
  assign new_n9405 = pi0 & new_n9404;
  assign new_n9406 = ~pe & new_n9405;
  assign new_n9407 = ~pf & new_n9406;
  assign new_n9408 = ~pf0 & new_n9407;
  assign new_n9409 = ~pj0 & new_n9408;
  assign new_n9410 = pm0 & new_n9409;
  assign new_n9411 = ~pc0 & new_n9410;
  assign new_n9412 = ~pg0 & new_n9411;
  assign new_n9413 = ~pe & new_n8779;
  assign new_n9414 = ~pf & new_n9413;
  assign new_n9415 = ~pg & new_n9414;
  assign new_n9416 = ~pt & new_n9415;
  assign new_n9417 = ~pf0 & new_n9416;
  assign new_n9418 = ~ph0 & new_n9417;
  assign new_n9419 = pm0 & new_n9418;
  assign new_n9420 = ~pg0 & new_n9419;
  assign new_n9421 = ~pj0 & new_n9420;
  assign new_n9422 = ~pa0 & new_n9421;
  assign new_n9423 = ~pc0 & new_n9422;
  assign new_n9424 = ~pm & new_n7863;
  assign new_n9425 = ~pk & new_n9424;
  assign new_n9426 = ~pf & new_n9425;
  assign new_n9427 = ~pg & new_n9426;
  assign new_n9428 = ~pe & new_n9427;
  assign new_n9429 = ~pj0 & new_n9428;
  assign new_n9430 = pm0 & new_n9429;
  assign new_n9431 = ~pa0 & new_n9430;
  assign new_n9432 = ~pc0 & new_n9431;
  assign new_n9433 = ~pf0 & new_n7241;
  assign new_n9434 = ~pi & new_n9433;
  assign new_n9435 = pm0 & new_n9434;
  assign new_n9436 = ~pe0 & new_n9435;
  assign new_n9437 = ~pj0 & new_n9436;
  assign new_n9438 = ~pa0 & new_n9437;
  assign new_n9439 = ~pc0 & new_n9438;
  assign new_n9440 = ~ps & new_n5926;
  assign new_n9441 = ~pc & new_n9440;
  assign new_n9442 = ~pd0 & new_n9441;
  assign new_n9443 = ~pi0 & new_n9442;
  assign new_n9444 = pd & new_n9443;
  assign new_n9445 = ~ph & new_n9444;
  assign new_n9446 = ~pi & new_n9445;
  assign new_n9447 = ~pg & new_n9446;
  assign new_n9448 = ~pe & new_n9447;
  assign new_n9449 = ~pf & new_n9448;
  assign new_n9450 = pm0 & new_n9449;
  assign new_n9451 = ~ph0 & new_n9450;
  assign new_n9452 = ~pg & new_n8978;
  assign new_n9453 = ~ph & new_n9452;
  assign new_n9454 = ~pf & new_n9453;
  assign new_n9455 = pm0 & new_n9454;
  assign new_n9456 = ~pe & new_n9455;
  assign new_n9457 = ~pc0 & new_n9456;
  assign new_n9458 = ~pg0 & new_n9457;
  assign new_n9459 = ~pl & new_n6098;
  assign new_n9460 = ~pc & new_n9459;
  assign new_n9461 = ~pt & new_n9460;
  assign new_n9462 = ~pd0 & new_n9461;
  assign new_n9463 = ~pi0 & new_n9462;
  assign new_n9464 = ~pg & new_n9463;
  assign new_n9465 = ~ph & new_n9464;
  assign new_n9466 = ~pf & new_n9465;
  assign new_n9467 = ~ph0 & new_n9466;
  assign new_n9468 = ~pe & new_n9467;
  assign new_n9469 = pj0 & new_n9468;
  assign new_n9470 = pm0 & new_n9469;
  assign new_n9471 = ~pi & new_n5950;
  assign new_n9472 = ~pd0 & new_n9471;
  assign new_n9473 = pi0 & new_n9472;
  assign new_n9474 = ~pf & new_n9473;
  assign new_n9475 = ~pg & new_n9474;
  assign new_n9476 = ~pe & new_n9475;
  assign new_n9477 = pm0 & new_n9476;
  assign new_n9478 = ~pf0 & new_n9477;
  assign new_n9479 = ~pc0 & new_n9478;
  assign new_n9480 = ~pj0 & new_n9479;
  assign new_n9481 = pm0 & new_n9236;
  assign new_n9482 = ~ph0 & new_n9481;
  assign new_n9483 = ~pa0 & new_n9482;
  assign new_n9484 = ~pc0 & new_n9483;
  assign new_n9485 = pm0 & new_n9243;
  assign new_n9486 = ~pf0 & new_n9485;
  assign new_n9487 = ~pj0 & new_n9486;
  assign new_n9488 = ~pc0 & new_n9487;
  assign new_n9489 = ~pg0 & new_n9488;
  assign new_n9490 = ~pz & new_n9489;
  assign new_n9491 = ~pa0 & new_n9490;
  assign new_n9492 = ~pg & new_n9020;
  assign new_n9493 = ~ph & new_n9492;
  assign new_n9494 = ~pf & new_n9493;
  assign new_n9495 = ~ph0 & new_n9494;
  assign new_n9496 = ~pe & new_n9495;
  assign new_n9497 = ~pg0 & new_n9496;
  assign new_n9498 = pm0 & new_n9497;
  assign new_n9499 = ~pi & new_n7522;
  assign new_n9500 = pt & new_n9499;
  assign new_n9501 = ~ph & new_n9500;
  assign new_n9502 = pm0 & new_n9501;
  assign new_n9503 = ~ph0 & new_n9502;
  assign new_n9504 = ~pc0 & new_n9503;
  assign new_n9505 = ~pe0 & new_n9504;
  assign new_n9506 = pi0 & new_n6387;
  assign new_n9507 = ~pm & new_n9506;
  assign new_n9508 = ~pg & new_n9507;
  assign new_n9509 = ~pd0 & new_n9508;
  assign new_n9510 = ~pf & new_n9509;
  assign new_n9511 = ~pf0 & new_n9510;
  assign new_n9512 = ~pe & new_n9511;
  assign new_n9513 = ~pj0 & new_n9512;
  assign new_n9514 = pm0 & new_n9513;
  assign new_n9515 = ~pg & new_n7342;
  assign new_n9516 = ~pm & new_n9515;
  assign new_n9517 = ~pe & new_n9516;
  assign new_n9518 = ~pf & new_n9517;
  assign new_n9519 = ~ph0 & new_n9518;
  assign new_n9520 = pm0 & new_n9519;
  assign new_n9521 = ~pf0 & new_n9520;
  assign new_n9522 = ~pg0 & new_n9521;
  assign new_n9523 = ~pj0 & new_n9522;
  assign new_n9524 = ~pi & new_n9284;
  assign new_n9525 = ~pj0 & new_n9524;
  assign new_n9526 = ~pc0 & new_n9525;
  assign new_n9527 = ~pe0 & new_n9526;
  assign new_n9528 = ~pz & new_n9527;
  assign new_n9529 = ~pa0 & new_n9528;
  assign new_n9530 = ~ph0 & new_n8180;
  assign new_n9531 = ~pi & new_n9530;
  assign new_n9532 = pm0 & new_n9531;
  assign new_n9533 = ~pe0 & new_n9532;
  assign new_n9534 = ~pj0 & new_n9533;
  assign new_n9535 = ~pa0 & new_n9534;
  assign new_n9536 = ~pc0 & new_n9535;
  assign new_n9537 = ~pb & new_n9506;
  assign new_n9538 = ~pg & new_n9537;
  assign new_n9539 = ~pd0 & new_n9538;
  assign new_n9540 = ~pf & new_n9539;
  assign new_n9541 = ~pf0 & new_n9540;
  assign new_n9542 = ~pe & new_n9541;
  assign new_n9543 = ~pj0 & new_n9542;
  assign new_n9544 = pm0 & new_n9543;
  assign new_n9545 = ~pb & new_n9515;
  assign new_n9546 = ~pe & new_n9545;
  assign new_n9547 = ~pf & new_n9546;
  assign new_n9548 = ~ph0 & new_n9547;
  assign new_n9549 = pm0 & new_n9548;
  assign new_n9550 = ~pf0 & new_n9549;
  assign new_n9551 = ~pg0 & new_n9550;
  assign new_n9552 = ~pj0 & new_n9551;
  assign new_n9553 = ~pg & new_n9472;
  assign new_n9554 = ~ph & new_n9553;
  assign new_n9555 = ~pf & new_n9554;
  assign new_n9556 = pm0 & new_n9555;
  assign new_n9557 = ~pe & new_n9556;
  assign new_n9558 = ~pa0 & new_n9557;
  assign new_n9559 = ~pc0 & new_n9558;
  assign new_n9560 = ~pz & new_n685;
  assign new_n9561 = ~pc0 & new_n9560;
  assign new_n9562 = ~pc & new_n9561;
  assign new_n9563 = ~pm & new_n9562;
  assign new_n9564 = ~pd0 & new_n9563;
  assign new_n9565 = ~pi0 & new_n9564;
  assign new_n9566 = ~ph & new_n9565;
  assign new_n9567 = ~pf & new_n9566;
  assign new_n9568 = ~pg & new_n9567;
  assign new_n9569 = pm0 & new_n9568;
  assign new_n9570 = ~pe & new_n9569;
  assign new_n9571 = pm0 & new_n7536;
  assign new_n9572 = ~pi & new_n9571;
  assign new_n9573 = ~pe0 & new_n9572;
  assign new_n9574 = ~pj0 & new_n9573;
  assign new_n9575 = ~pi & new_n7544;
  assign new_n9576 = ~pd0 & new_n9575;
  assign new_n9577 = ~ph0 & new_n9576;
  assign new_n9578 = ~pj0 & new_n9577;
  assign new_n9579 = pm0 & new_n9578;
  assign new_n9580 = ~pc0 & new_n9579;
  assign new_n9581 = ~pe0 & new_n9580;
  assign new_n9582 = ~pb & new_n9562;
  assign new_n9583 = ~pd0 & new_n9582;
  assign new_n9584 = ~pi0 & new_n9583;
  assign new_n9585 = ~ph & new_n9584;
  assign new_n9586 = ~pf & new_n9585;
  assign new_n9587 = ~pg & new_n9586;
  assign new_n9588 = pm0 & new_n9587;
  assign new_n9589 = ~pe & new_n9588;
  assign new_n9590 = ~pg & new_n8220;
  assign new_n9591 = ~ph & new_n9590;
  assign new_n9592 = ~pf & new_n9591;
  assign new_n9593 = ~ph0 & new_n9592;
  assign new_n9594 = ~pe & new_n9593;
  assign new_n9595 = ~pg0 & new_n9594;
  assign new_n9596 = pm0 & new_n9595;
  assign new_n9597 = pm0 & new_n7565;
  assign new_n9598 = ~pe0 & new_n9597;
  assign new_n9599 = ~pj0 & new_n9598;
  assign new_n9600 = ~pz & new_n9599;
  assign new_n9601 = ~pc0 & new_n9600;
  assign new_n9602 = ~pi & new_n8236;
  assign new_n9603 = pm0 & new_n9602;
  assign new_n9604 = ~ph0 & new_n9603;
  assign new_n9605 = ~pe0 & new_n9604;
  assign new_n9606 = ~pj0 & new_n9605;
  assign new_n9607 = pm0 & new_n7982;
  assign new_n9608 = ~ph0 & new_n9607;
  assign new_n9609 = ~pj0 & new_n9608;
  assign new_n9610 = ~pc0 & new_n9609;
  assign new_n9611 = ~pg0 & new_n9610;
  assign new_n9612 = ~py & new_n9611;
  assign new_n9613 = ~pa0 & new_n9612;
  assign new_n9614 = pm0 & new_n8899;
  assign new_n9615 = ~pe & new_n9614;
  assign new_n9616 = ~pj0 & new_n9615;
  assign new_n9617 = ~pc0 & new_n9616;
  assign new_n9618 = ~pg0 & new_n9617;
  assign new_n9619 = ~py & new_n9618;
  assign new_n9620 = ~pz & new_n9619;
  assign new_n9621 = pm0 & new_n7197;
  assign new_n9622 = ~ph0 & new_n9621;
  assign new_n9623 = ~pj0 & new_n9622;
  assign new_n9624 = ~pa0 & new_n9623;
  assign new_n9625 = ~pc0 & new_n9624;
  assign new_n9626 = ~pw & new_n9625;
  assign new_n9627 = ~py & new_n9626;
  assign new_n9628 = ~pi & new_n6047;
  assign new_n9629 = ~pd0 & new_n9628;
  assign new_n9630 = pd & new_n9629;
  assign new_n9631 = ~pe & new_n9630;
  assign new_n9632 = ~pf & new_n9631;
  assign new_n9633 = ~pf0 & new_n9632;
  assign new_n9634 = ~pj0 & new_n9633;
  assign new_n9635 = pm0 & new_n9634;
  assign new_n9636 = ~pa0 & new_n9635;
  assign new_n9637 = ~pc0 & new_n9636;
  assign new_n9638 = ~pg & new_n6059;
  assign new_n9639 = ~pt & new_n9638;
  assign new_n9640 = ~pd0 & new_n9639;
  assign new_n9641 = pi0 & new_n9640;
  assign new_n9642 = ~pe & new_n9641;
  assign new_n9643 = ~pf & new_n9642;
  assign new_n9644 = ~ph0 & new_n9643;
  assign new_n9645 = pm0 & new_n9644;
  assign new_n9646 = ~pf0 & new_n9645;
  assign new_n9647 = ~pg0 & new_n9646;
  assign new_n9648 = ~pj0 & new_n9647;
  assign new_n9649 = pm0 & new_n9416;
  assign new_n9650 = ~pf0 & new_n9649;
  assign new_n9651 = ~pj0 & new_n9650;
  assign new_n9652 = ~pc0 & new_n9651;
  assign new_n9653 = ~pg0 & new_n9652;
  assign new_n9654 = ~pz & new_n9653;
  assign new_n9655 = ~pa0 & new_n9654;
  assign new_n9656 = ~pm & new_n8664;
  assign new_n9657 = ~pk & new_n9656;
  assign new_n9658 = ~pf & new_n9657;
  assign new_n9659 = ~pg & new_n9658;
  assign new_n9660 = ~pe & new_n9659;
  assign new_n9661 = pm0 & new_n9660;
  assign new_n9662 = ~ph0 & new_n9661;
  assign new_n9663 = ~pc0 & new_n9662;
  assign new_n9664 = ~pj0 & new_n9663;
  assign new_n9665 = ~pf0 & new_n8312;
  assign new_n9666 = ~ph0 & new_n9665;
  assign new_n9667 = pm0 & new_n9666;
  assign new_n9668 = ~pg0 & new_n9667;
  assign new_n9669 = ~pj0 & new_n9668;
  assign new_n9670 = ~pc0 & new_n9669;
  assign new_n9671 = ~pe0 & new_n9670;
  assign new_n9672 = ~pf0 & new_n8119;
  assign new_n9673 = pm & new_n9672;
  assign new_n9674 = pk & new_n9673;
  assign new_n9675 = ~pj0 & new_n9674;
  assign new_n9676 = pm0 & new_n9675;
  assign new_n9677 = ~pg0 & new_n9676;
  assign new_n9678 = ~pc0 & new_n9677;
  assign new_n9679 = ~pe0 & new_n9678;
  assign new_n9680 = ~pz & new_n9679;
  assign new_n9681 = ~pa0 & new_n9680;
  assign new_n9682 = ~pi & new_n8331;
  assign new_n9683 = ~pd0 & new_n9682;
  assign new_n9684 = pd & new_n9683;
  assign new_n9685 = ~pg & new_n9684;
  assign new_n9686 = ~ph & new_n9685;
  assign new_n9687 = ~pf & new_n9686;
  assign new_n9688 = ~ph0 & new_n9687;
  assign new_n9689 = ~pe & new_n9688;
  assign new_n9690 = ~pc0 & new_n9689;
  assign new_n9691 = pm0 & new_n9690;
  assign new_n9692 = ~ph & new_n8346;
  assign new_n9693 = ~pi & new_n9692;
  assign new_n9694 = ~pg & new_n9693;
  assign new_n9695 = ~pe & new_n9694;
  assign new_n9696 = ~pf & new_n9695;
  assign new_n9697 = pj0 & new_n9696;
  assign new_n9698 = pm0 & new_n9697;
  assign new_n9699 = ~pg & new_n6122;
  assign new_n9700 = ~pd0 & new_n9699;
  assign new_n9701 = pi0 & new_n9700;
  assign new_n9702 = ~pe & new_n9701;
  assign new_n9703 = ~pf & new_n9702;
  assign new_n9704 = ~ph0 & new_n9703;
  assign new_n9705 = pm0 & new_n9704;
  assign new_n9706 = ~pf0 & new_n9705;
  assign new_n9707 = ~pg0 & new_n9706;
  assign new_n9708 = ~pj0 & new_n9707;
  assign new_n9709 = ~pf & new_n5950;
  assign new_n9710 = ~pg & new_n9709;
  assign new_n9711 = ~pd0 & new_n9710;
  assign new_n9712 = ~pf0 & new_n9711;
  assign new_n9713 = ~pe & new_n9712;
  assign new_n9714 = pm0 & new_n9713;
  assign new_n9715 = ~pg0 & new_n9714;
  assign new_n9716 = ~pj0 & new_n9715;
  assign new_n9717 = ~pa0 & new_n9716;
  assign new_n9718 = ~pc0 & new_n9717;
  assign new_n9719 = ~pj & new_n6796;
  assign new_n9720 = ~pc0 & new_n9719;
  assign new_n9721 = ~pc & new_n9720;
  assign new_n9722 = ~pi0 & new_n9721;
  assign new_n9723 = ~pk & new_n9722;
  assign new_n9724 = ~pi & new_n9723;
  assign new_n9725 = ~pd0 & new_n9724;
  assign new_n9726 = ~ph & new_n9725;
  assign new_n9727 = ~pf & new_n9726;
  assign new_n9728 = ~pg & new_n9727;
  assign new_n9729 = ~ph0 & new_n9728;
  assign new_n9730 = ~pe & new_n9729;
  assign new_n9731 = ~ph & new_n6160;
  assign new_n9732 = ~pi & new_n9731;
  assign new_n9733 = ~pg & new_n9732;
  assign new_n9734 = ~pe & new_n9733;
  assign new_n9735 = ~pf & new_n9734;
  assign new_n9736 = ~pc0 & new_n9735;
  assign new_n9737 = pm0 & new_n9736;
  assign new_n9738 = ~pi & new_n7096;
  assign new_n9739 = pt & new_n9738;
  assign new_n9740 = ~ph & new_n9739;
  assign new_n9741 = ~pe0 & new_n9740;
  assign new_n9742 = pm0 & new_n9741;
  assign new_n9743 = ~pa0 & new_n9742;
  assign new_n9744 = ~pc0 & new_n9743;
  assign new_n9745 = ~py & new_n6582;
  assign new_n9746 = ~pc0 & new_n9745;
  assign new_n9747 = ~pc & new_n9746;
  assign new_n9748 = pi0 & new_n9747;
  assign new_n9749 = ~pm & new_n9748;
  assign new_n9750 = ~pg & new_n9749;
  assign new_n9751 = ~pd0 & new_n9750;
  assign new_n9752 = ~pf & new_n9751;
  assign new_n9753 = ~ph0 & new_n9752;
  assign new_n9754 = ~pe & new_n9753;
  assign new_n9755 = pm0 & new_n9754;
  assign new_n9756 = ~pf0 & new_n9755;
  assign new_n9757 = ~pg & new_n6170;
  assign new_n9758 = ~pm & new_n9757;
  assign new_n9759 = ~pe & new_n9758;
  assign new_n9760 = ~pf & new_n9759;
  assign new_n9761 = ~pf0 & new_n9760;
  assign new_n9762 = ~pj0 & new_n9761;
  assign new_n9763 = pm0 & new_n9762;
  assign new_n9764 = ~pc0 & new_n9763;
  assign new_n9765 = ~pg0 & new_n9764;
  assign new_n9766 = ~ph0 & new_n9055;
  assign new_n9767 = ~pi & new_n9766;
  assign new_n9768 = pm0 & new_n9767;
  assign new_n9769 = ~pe0 & new_n9768;
  assign new_n9770 = ~pj0 & new_n9769;
  assign new_n9771 = ~pa0 & new_n9770;
  assign new_n9772 = ~pc0 & new_n9771;
  assign new_n9773 = ~pi & new_n8181;
  assign new_n9774 = ~pj0 & new_n9773;
  assign new_n9775 = ~pc0 & new_n9774;
  assign new_n9776 = ~pe0 & new_n9775;
  assign new_n9777 = ~pz & new_n9776;
  assign new_n9778 = ~pa0 & new_n9777;
  assign new_n9779 = ~pb & new_n9748;
  assign new_n9780 = ~pg & new_n9779;
  assign new_n9781 = ~pd0 & new_n9780;
  assign new_n9782 = ~pf & new_n9781;
  assign new_n9783 = ~ph0 & new_n9782;
  assign new_n9784 = ~pe & new_n9783;
  assign new_n9785 = pm0 & new_n9784;
  assign new_n9786 = ~pf0 & new_n9785;
  assign new_n9787 = ~pb & new_n9757;
  assign new_n9788 = ~pe & new_n9787;
  assign new_n9789 = ~pf & new_n9788;
  assign new_n9790 = ~pf0 & new_n9789;
  assign new_n9791 = ~pj0 & new_n9790;
  assign new_n9792 = pm0 & new_n9791;
  assign new_n9793 = ~pc0 & new_n9792;
  assign new_n9794 = ~pg0 & new_n9793;
  assign new_n9795 = ~pi & new_n5914;
  assign new_n9796 = ~pd0 & new_n9795;
  assign new_n9797 = ~pg & new_n9796;
  assign new_n9798 = ~ph & new_n9797;
  assign new_n9799 = ~pf & new_n9798;
  assign new_n9800 = ~ph0 & new_n9799;
  assign new_n9801 = ~pe & new_n9800;
  assign new_n9802 = ~pc0 & new_n9801;
  assign new_n9803 = pm0 & new_n9802;
  assign new_n9804 = ~pc0 & new_n7994;
  assign new_n9805 = pm0 & new_n9804;
  assign new_n9806 = ~pz & new_n9805;
  assign new_n9807 = ~pa0 & new_n9806;
  assign new_n9808 = pm0 & new_n9330;
  assign new_n9809 = ~ph0 & new_n9808;
  assign new_n9810 = ~pg0 & new_n9809;
  assign new_n9811 = ~pj0 & new_n9810;
  assign new_n9812 = pm0 & new_n9340;
  assign new_n9813 = ~pg0 & new_n9812;
  assign new_n9814 = ~pj0 & new_n9813;
  assign new_n9815 = ~pc0 & new_n9814;
  assign new_n9816 = ~pe0 & new_n9815;
  assign new_n9817 = ~pb & new_n6192;
  assign new_n9818 = ~pd0 & new_n9817;
  assign new_n9819 = pi0 & new_n9818;
  assign new_n9820 = ~pi & new_n9819;
  assign new_n9821 = ~pg & new_n9820;
  assign new_n9822 = ~ph & new_n9821;
  assign new_n9823 = ~pe & new_n9822;
  assign new_n9824 = ~pf & new_n9823;
  assign new_n9825 = ~ph & new_n9354;
  assign new_n9826 = ~pi & new_n9825;
  assign new_n9827 = ~pg & new_n9826;
  assign new_n9828 = ~pe & new_n9827;
  assign new_n9829 = ~pf & new_n9828;
  assign new_n9830 = ~pc0 & new_n9829;
  assign new_n9831 = pm0 & new_n9830;
  assign new_n9832 = ~ph0 & new_n7563;
  assign new_n9833 = ~pd0 & new_n9832;
  assign new_n9834 = pm0 & new_n9833;
  assign new_n9835 = ~pg0 & new_n9834;
  assign new_n9836 = ~pj0 & new_n9835;
  assign new_n9837 = ~pc0 & new_n9836;
  assign new_n9838 = ~pe0 & new_n9837;
  assign new_n9839 = ~pj0 & new_n7855;
  assign new_n9840 = pm0 & new_n9839;
  assign new_n9841 = ~pg0 & new_n9840;
  assign new_n9842 = ~pc0 & new_n9841;
  assign new_n9843 = ~pe0 & new_n9842;
  assign new_n9844 = ~pz & new_n9843;
  assign new_n9845 = ~pa0 & new_n9844;
  assign new_n9846 = ~new_n4000 & ~new_n9845;
  assign new_n9847 = ~new_n9831 & ~new_n9838;
  assign new_n9848 = new_n9846 & new_n9847;
  assign new_n9849 = ~new_n9816 & ~new_n9824;
  assign new_n9850 = ~new_n9807 & ~new_n9811;
  assign new_n9851 = new_n9849 & new_n9850;
  assign new_n9852 = new_n9848 & new_n9851;
  assign new_n9853 = ~new_n9794 & ~new_n9803;
  assign new_n9854 = ~new_n9778 & ~new_n9786;
  assign new_n9855 = new_n9853 & new_n9854;
  assign new_n9856 = ~new_n9765 & ~new_n9772;
  assign new_n9857 = ~new_n9744 & ~new_n9756;
  assign new_n9858 = new_n9856 & new_n9857;
  assign new_n9859 = new_n9855 & new_n9858;
  assign new_n9860 = new_n9852 & new_n9859;
  assign new_n9861 = ~new_n9730 & ~new_n9737;
  assign new_n9862 = ~new_n9708 & ~new_n9718;
  assign new_n9863 = new_n9861 & new_n9862;
  assign new_n9864 = ~new_n9691 & ~new_n9698;
  assign new_n9865 = ~new_n9671 & ~new_n9681;
  assign new_n9866 = new_n9864 & new_n9865;
  assign new_n9867 = new_n9863 & new_n9866;
  assign new_n9868 = ~new_n9655 & ~new_n9664;
  assign new_n9869 = ~new_n9637 & ~new_n9648;
  assign new_n9870 = new_n9868 & new_n9869;
  assign new_n9871 = ~new_n9620 & ~new_n9627;
  assign new_n9872 = ~new_n1930 & ~new_n9606;
  assign new_n9873 = ~new_n9613 & new_n9872;
  assign new_n9874 = new_n9871 & new_n9873;
  assign new_n9875 = new_n9870 & new_n9874;
  assign new_n9876 = new_n9867 & new_n9875;
  assign new_n9877 = new_n9860 & new_n9876;
  assign new_n9878 = ~new_n9596 & ~new_n9601;
  assign new_n9879 = ~new_n9581 & ~new_n9589;
  assign new_n9880 = new_n9878 & new_n9879;
  assign new_n9881 = ~new_n9570 & ~new_n9574;
  assign new_n9882 = ~new_n9552 & ~new_n9559;
  assign new_n9883 = new_n9881 & new_n9882;
  assign new_n9884 = new_n9880 & new_n9883;
  assign new_n9885 = ~new_n9536 & ~new_n9544;
  assign new_n9886 = ~new_n9523 & ~new_n9529;
  assign new_n9887 = new_n9885 & new_n9886;
  assign new_n9888 = ~new_n9505 & ~new_n9514;
  assign new_n9889 = ~new_n9491 & ~new_n9498;
  assign new_n9890 = new_n9888 & new_n9889;
  assign new_n9891 = new_n9887 & new_n9890;
  assign new_n9892 = new_n9884 & new_n9891;
  assign new_n9893 = ~new_n9480 & ~new_n9484;
  assign new_n9894 = ~new_n9458 & ~new_n9470;
  assign new_n9895 = new_n9893 & new_n9894;
  assign new_n9896 = ~new_n9439 & ~new_n9451;
  assign new_n9897 = ~new_n9423 & ~new_n9432;
  assign new_n9898 = new_n9896 & new_n9897;
  assign new_n9899 = new_n9895 & new_n9898;
  assign new_n9900 = ~new_n9402 & ~new_n9412;
  assign new_n9901 = ~new_n9384 & ~new_n9391;
  assign new_n9902 = new_n9900 & new_n9901;
  assign new_n9903 = ~new_n3586 & ~new_n9379;
  assign new_n9904 = ~new_n9361 & ~new_n9368;
  assign new_n9905 = ~new_n9372 & new_n9904;
  assign new_n9906 = new_n9903 & new_n9905;
  assign new_n9907 = new_n9902 & new_n9906;
  assign new_n9908 = new_n9899 & new_n9907;
  assign new_n9909 = new_n9892 & new_n9908;
  assign new_n9910 = new_n9877 & new_n9909;
  assign new_n9911 = ~new_n9345 & ~new_n9353;
  assign new_n9912 = ~new_n9323 & ~new_n9334;
  assign new_n9913 = new_n9911 & new_n9912;
  assign new_n9914 = ~new_n9307 & ~new_n9314;
  assign new_n9915 = ~new_n9290 & ~new_n9299;
  assign new_n9916 = new_n9914 & new_n9915;
  assign new_n9917 = new_n9913 & new_n9916;
  assign new_n9918 = ~new_n9276 & ~new_n9283;
  assign new_n9919 = ~new_n9257 & ~new_n9264;
  assign new_n9920 = new_n9918 & new_n9919;
  assign new_n9921 = ~new_n9240 & ~new_n9250;
  assign new_n9922 = ~new_n9220 & ~new_n9230;
  assign new_n9923 = new_n9921 & new_n9922;
  assign new_n9924 = new_n9920 & new_n9923;
  assign new_n9925 = new_n9917 & new_n9924;
  assign new_n9926 = ~new_n9208 & ~new_n9215;
  assign new_n9927 = ~new_n9189 & ~new_n9198;
  assign new_n9928 = new_n9926 & new_n9927;
  assign new_n9929 = ~new_n9175 & ~new_n9182;
  assign new_n9930 = ~new_n9157 & ~new_n9164;
  assign new_n9931 = new_n9929 & new_n9930;
  assign new_n9932 = new_n9928 & new_n9931;
  assign new_n9933 = ~new_n9147 & ~new_n9152;
  assign new_n9934 = ~new_n3491 & ~new_n9136;
  assign new_n9935 = new_n9933 & new_n9934;
  assign new_n9936 = ~new_n9124 & ~new_n9131;
  assign new_n9937 = ~new_n9106 & ~new_n9111;
  assign new_n9938 = ~new_n9119 & new_n9937;
  assign new_n9939 = new_n9936 & new_n9938;
  assign new_n9940 = new_n9935 & new_n9939;
  assign new_n9941 = new_n9932 & new_n9940;
  assign new_n9942 = new_n9925 & new_n9941;
  assign new_n9943 = ~new_n9090 & ~new_n9099;
  assign new_n9944 = ~new_n9071 & ~new_n9079;
  assign new_n9945 = new_n9943 & new_n9944;
  assign new_n9946 = ~new_n9052 & ~new_n9062;
  assign new_n9947 = ~new_n9034 & ~new_n9045;
  assign new_n9948 = new_n9946 & new_n9947;
  assign new_n9949 = new_n9945 & new_n9948;
  assign new_n9950 = ~new_n9018 & ~new_n9027;
  assign new_n9951 = ~new_n9006 & ~new_n9011;
  assign new_n9952 = new_n9950 & new_n9951;
  assign new_n9953 = ~new_n8985 & ~new_n8997;
  assign new_n9954 = ~new_n8956 & ~new_n8965;
  assign new_n9955 = ~new_n8975 & new_n9954;
  assign new_n9956 = new_n9953 & new_n9955;
  assign new_n9957 = new_n9952 & new_n9956;
  assign new_n9958 = new_n9949 & new_n9957;
  assign new_n9959 = ~new_n8938 & ~new_n8949;
  assign new_n9960 = ~new_n8916 & ~new_n8927;
  assign new_n9961 = new_n9959 & new_n9960;
  assign new_n9962 = ~new_n8897 & ~new_n8906;
  assign new_n9963 = ~new_n8885 & ~new_n8890;
  assign new_n9964 = new_n9962 & new_n9963;
  assign new_n9965 = new_n9961 & new_n9964;
  assign new_n9966 = ~new_n8871 & ~new_n8876;
  assign new_n9967 = ~new_n8859 & ~new_n8864;
  assign new_n9968 = new_n9966 & new_n9967;
  assign new_n9969 = ~new_n8845 & ~new_n8852;
  assign new_n9970 = ~new_n8819 & ~new_n8826;
  assign new_n9971 = ~new_n8834 & new_n9970;
  assign new_n9972 = new_n9969 & new_n9971;
  assign new_n9973 = new_n9968 & new_n9972;
  assign new_n9974 = new_n9965 & new_n9973;
  assign new_n9975 = new_n9958 & new_n9974;
  assign new_n9976 = new_n9942 & new_n9975;
  assign new_n9977 = new_n9910 & new_n9976;
  assign new_n9978 = ~new_n8805 & ~new_n8812;
  assign new_n9979 = ~new_n8789 & ~new_n8798;
  assign new_n9980 = new_n9978 & new_n9979;
  assign new_n9981 = ~new_n8767 & ~new_n8777;
  assign new_n9982 = ~new_n8753 & ~new_n8760;
  assign new_n9983 = new_n9981 & new_n9982;
  assign new_n9984 = new_n9980 & new_n9983;
  assign new_n9985 = ~new_n8734 & ~new_n8743;
  assign new_n9986 = ~new_n8714 & ~new_n8725;
  assign new_n9987 = new_n9985 & new_n9986;
  assign new_n9988 = ~new_n8702 & ~new_n8707;
  assign new_n9989 = ~new_n8693 & ~new_n8698;
  assign new_n9990 = new_n9988 & new_n9989;
  assign new_n9991 = new_n9987 & new_n9990;
  assign new_n9992 = new_n9984 & new_n9991;
  assign new_n9993 = ~new_n705 & ~new_n8682;
  assign new_n9994 = ~new_n8670 & ~new_n8677;
  assign new_n9995 = new_n9993 & new_n9994;
  assign new_n9996 = ~new_n8656 & ~new_n8663;
  assign new_n9997 = ~new_n8637 & ~new_n8645;
  assign new_n9998 = new_n9996 & new_n9997;
  assign new_n9999 = new_n9995 & new_n9998;
  assign new_n10000 = ~new_n8617 & ~new_n8628;
  assign new_n10001 = ~new_n8601 & ~new_n8610;
  assign new_n10002 = new_n10000 & new_n10001;
  assign new_n10003 = ~new_n8586 & ~new_n8595;
  assign new_n10004 = ~new_n8560 & ~new_n8570;
  assign new_n10005 = ~new_n8579 & new_n10004;
  assign new_n10006 = new_n10003 & new_n10005;
  assign new_n10007 = new_n10002 & new_n10006;
  assign new_n10008 = new_n9999 & new_n10007;
  assign new_n10009 = new_n9992 & new_n10008;
  assign new_n10010 = ~new_n8546 & ~new_n8553;
  assign new_n10011 = ~new_n8529 & ~new_n8539;
  assign new_n10012 = new_n10010 & new_n10011;
  assign new_n10013 = ~new_n8513 & ~new_n8522;
  assign new_n10014 = ~new_n8489 & ~new_n8500;
  assign new_n10015 = new_n10013 & new_n10014;
  assign new_n10016 = new_n10012 & new_n10015;
  assign new_n10017 = ~new_n8472 & ~new_n8479;
  assign new_n10018 = ~new_n8456 & ~new_n8461;
  assign new_n10019 = new_n10017 & new_n10018;
  assign new_n10020 = ~new_n8442 & ~new_n8451;
  assign new_n10021 = ~new_n8424 & ~new_n8434;
  assign new_n10022 = new_n10020 & new_n10021;
  assign new_n10023 = new_n10019 & new_n10022;
  assign new_n10024 = new_n10016 & new_n10023;
  assign new_n10025 = ~new_n8409 & ~new_n8417;
  assign new_n10026 = ~new_n8393 & ~new_n8400;
  assign new_n10027 = new_n10025 & new_n10026;
  assign new_n10028 = ~new_n8378 & ~new_n8385;
  assign new_n10029 = ~new_n8363 & ~new_n8371;
  assign new_n10030 = new_n10028 & new_n10029;
  assign new_n10031 = new_n10027 & new_n10030;
  assign new_n10032 = ~new_n8353 & ~new_n8358;
  assign new_n10033 = ~new_n8329 & ~new_n8341;
  assign new_n10034 = new_n10032 & new_n10033;
  assign new_n10035 = ~new_n8308 & ~new_n8319;
  assign new_n10036 = ~new_n8283 & ~new_n8294;
  assign new_n10037 = ~new_n8301 & new_n10036;
  assign new_n10038 = new_n10035 & new_n10037;
  assign new_n10039 = new_n10034 & new_n10038;
  assign new_n10040 = new_n10031 & new_n10039;
  assign new_n10041 = new_n10024 & new_n10040;
  assign new_n10042 = new_n10009 & new_n10041;
  assign new_n10043 = ~new_n8272 & ~new_n8279;
  assign new_n10044 = ~new_n8261 & ~new_n8265;
  assign new_n10045 = new_n10043 & new_n10044;
  assign new_n10046 = ~new_n8245 & ~new_n8249;
  assign new_n10047 = ~new_n8234 & ~new_n8241;
  assign new_n10048 = new_n10046 & new_n10047;
  assign new_n10049 = new_n10045 & new_n10048;
  assign new_n10050 = ~new_n8219 & ~new_n8227;
  assign new_n10051 = ~new_n8202 & ~new_n8211;
  assign new_n10052 = new_n10050 & new_n10051;
  assign new_n10053 = ~new_n8187 & ~new_n8195;
  assign new_n10054 = ~new_n8166 & ~new_n8178;
  assign new_n10055 = new_n10053 & new_n10054;
  assign new_n10056 = new_n10052 & new_n10055;
  assign new_n10057 = new_n10049 & new_n10056;
  assign new_n10058 = ~new_n8149 & ~new_n8158;
  assign new_n10059 = ~new_n8137 & ~new_n8144;
  assign new_n10060 = new_n10058 & new_n10059;
  assign new_n10061 = ~new_n8116 & ~new_n8129;
  assign new_n10062 = ~new_n8093 & ~new_n8106;
  assign new_n10063 = new_n10061 & new_n10062;
  assign new_n10064 = new_n10060 & new_n10063;
  assign new_n10065 = ~new_n8073 & ~new_n8080;
  assign new_n10066 = ~new_n8059 & ~new_n8066;
  assign new_n10067 = new_n10065 & new_n10066;
  assign new_n10068 = ~new_n8038 & ~new_n8048;
  assign new_n10069 = ~new_n8029 & ~new_n8030;
  assign new_n10070 = ~new_n8031 & new_n10069;
  assign new_n10071 = new_n10068 & new_n10070;
  assign new_n10072 = new_n10067 & new_n10071;
  assign new_n10073 = new_n10064 & new_n10072;
  assign new_n10074 = new_n10057 & new_n10073;
  assign new_n10075 = ~new_n8022 & ~new_n8024;
  assign new_n10076 = ~new_n8015 & ~new_n8020;
  assign new_n10077 = new_n10075 & new_n10076;
  assign new_n10078 = ~new_n8004 & ~new_n8011;
  assign new_n10079 = ~new_n7989 & ~new_n7998;
  assign new_n10080 = new_n10078 & new_n10079;
  assign new_n10081 = new_n10077 & new_n10080;
  assign new_n10082 = ~new_n7966 & ~new_n7977;
  assign new_n10083 = ~new_n7964 & ~new_n7965;
  assign new_n10084 = new_n10082 & new_n10083;
  assign new_n10085 = ~new_n7956 & ~new_n7958;
  assign new_n10086 = ~new_n7940 & ~new_n7948;
  assign new_n10087 = ~new_n7954 & new_n10086;
  assign new_n10088 = new_n10085 & new_n10087;
  assign new_n10089 = new_n10084 & new_n10088;
  assign new_n10090 = new_n10081 & new_n10089;
  assign new_n10091 = ~new_n7925 & ~new_n7932;
  assign new_n10092 = ~new_n7905 & ~new_n7916;
  assign new_n10093 = new_n10091 & new_n10092;
  assign new_n10094 = ~new_n7899 & ~new_n7900;
  assign new_n10095 = ~new_n7888 & ~new_n7894;
  assign new_n10096 = new_n10094 & new_n10095;
  assign new_n10097 = new_n10093 & new_n10096;
  assign new_n10098 = ~new_n7884 & ~new_n7886;
  assign new_n10099 = ~new_n7869 & ~new_n7878;
  assign new_n10100 = new_n10098 & new_n10099;
  assign new_n10101 = ~new_n7854 & ~new_n7862;
  assign new_n10102 = ~new_n7840 & ~new_n7845;
  assign new_n10103 = ~new_n7846 & new_n10102;
  assign new_n10104 = new_n10101 & new_n10103;
  assign new_n10105 = new_n10100 & new_n10104;
  assign new_n10106 = new_n10097 & new_n10105;
  assign new_n10107 = new_n10090 & new_n10106;
  assign new_n10108 = new_n10074 & new_n10107;
  assign new_n10109 = new_n10042 & new_n10108;
  assign new_n10110 = new_n9977 & new_n10109;
  assign new_n10111 = ~new_n7832 & ~new_n7834;
  assign new_n10112 = ~new_n7821 & ~new_n7830;
  assign new_n10113 = new_n10111 & new_n10112;
  assign new_n10114 = ~new_n7807 & ~new_n7814;
  assign new_n10115 = ~new_n3327 & ~new_n7799;
  assign new_n10116 = new_n10114 & new_n10115;
  assign new_n10117 = new_n10113 & new_n10116;
  assign new_n10118 = ~new_n7786 & ~new_n7790;
  assign new_n10119 = ~new_n7780 & ~new_n7785;
  assign new_n10120 = new_n10118 & new_n10119;
  assign new_n10121 = ~new_n7771 & ~new_n7775;
  assign new_n10122 = ~new_n7762 & ~new_n7767;
  assign new_n10123 = new_n10121 & new_n10122;
  assign new_n10124 = new_n10120 & new_n10123;
  assign new_n10125 = new_n10117 & new_n10124;
  assign new_n10126 = ~new_n7747 & ~new_n7754;
  assign new_n10127 = ~new_n1247 & ~new_n7742;
  assign new_n10128 = new_n10126 & new_n10127;
  assign new_n10129 = ~new_n7731 & ~new_n7735;
  assign new_n10130 = ~new_n7725 & ~new_n7730;
  assign new_n10131 = new_n10129 & new_n10130;
  assign new_n10132 = new_n10128 & new_n10131;
  assign new_n10133 = ~new_n7714 & ~new_n7720;
  assign new_n10134 = ~new_n7699 & ~new_n7710;
  assign new_n10135 = new_n10133 & new_n10134;
  assign new_n10136 = ~new_n7683 & ~new_n7691;
  assign new_n10137 = ~new_n7661 & ~new_n7664;
  assign new_n10138 = ~new_n7676 & new_n10137;
  assign new_n10139 = new_n10136 & new_n10138;
  assign new_n10140 = new_n10135 & new_n10139;
  assign new_n10141 = new_n10132 & new_n10140;
  assign new_n10142 = new_n10125 & new_n10141;
  assign new_n10143 = ~new_n7655 & ~new_n7660;
  assign new_n10144 = ~new_n7648 & ~new_n7654;
  assign new_n10145 = new_n10143 & new_n10144;
  assign new_n10146 = ~new_n7642 & ~new_n7646;
  assign new_n10147 = ~new_n7624 & ~new_n7632;
  assign new_n10148 = new_n10146 & new_n10147;
  assign new_n10149 = new_n10145 & new_n10148;
  assign new_n10150 = ~new_n7602 & ~new_n7613;
  assign new_n10151 = ~new_n7586 & ~new_n7590;
  assign new_n10152 = new_n10150 & new_n10151;
  assign new_n10153 = ~new_n7580 & ~new_n7581;
  assign new_n10154 = ~new_n7574 & ~new_n7579;
  assign new_n10155 = new_n10153 & new_n10154;
  assign new_n10156 = new_n10152 & new_n10155;
  assign new_n10157 = new_n10149 & new_n10156;
  assign new_n10158 = ~new_n7570 & ~new_n7572;
  assign new_n10159 = ~new_n7551 & ~new_n7559;
  assign new_n10160 = new_n10158 & new_n10159;
  assign new_n10161 = ~new_n7529 & ~new_n7540;
  assign new_n10162 = ~new_n7516 & ~new_n7520;
  assign new_n10163 = new_n10161 & new_n10162;
  assign new_n10164 = new_n10160 & new_n10163;
  assign new_n10165 = ~new_n7508 & ~new_n7512;
  assign new_n10166 = ~new_n7504 & ~new_n7505;
  assign new_n10167 = new_n10165 & new_n10166;
  assign new_n10168 = ~new_n7499 & ~new_n7503;
  assign new_n10169 = ~new_n7487 & ~new_n7490;
  assign new_n10170 = ~new_n7495 & new_n10169;
  assign new_n10171 = new_n10168 & new_n10170;
  assign new_n10172 = new_n10167 & new_n10171;
  assign new_n10173 = new_n10164 & new_n10172;
  assign new_n10174 = new_n10157 & new_n10173;
  assign new_n10175 = new_n10142 & new_n10174;
  assign new_n10176 = ~new_n831 & ~new_n7483;
  assign new_n10177 = ~new_n7478 & ~new_n7482;
  assign new_n10178 = new_n10176 & new_n10177;
  assign new_n10179 = ~new_n7473 & ~new_n7474;
  assign new_n10180 = ~new_n1148 & ~new_n7470;
  assign new_n10181 = new_n10179 & new_n10180;
  assign new_n10182 = new_n10178 & new_n10181;
  assign new_n10183 = ~new_n7460 & ~new_n7464;
  assign new_n10184 = ~new_n7455 & ~new_n7456;
  assign new_n10185 = new_n10183 & new_n10184;
  assign new_n10186 = ~new_n7444 & ~new_n7450;
  assign new_n10187 = ~new_n7437 & ~new_n7442;
  assign new_n10188 = new_n10186 & new_n10187;
  assign new_n10189 = new_n10185 & new_n10188;
  assign new_n10190 = new_n10182 & new_n10189;
  assign new_n10191 = ~new_n7429 & ~new_n7432;
  assign new_n10192 = ~new_n7421 & ~new_n7425;
  assign new_n10193 = new_n10191 & new_n10192;
  assign new_n10194 = ~new_n7412 & ~new_n7416;
  assign new_n10195 = ~new_n7402 & ~new_n7407;
  assign new_n10196 = new_n10194 & new_n10195;
  assign new_n10197 = new_n10193 & new_n10196;
  assign new_n10198 = ~new_n7392 & ~new_n7397;
  assign new_n10199 = ~new_n7381 & ~new_n7385;
  assign new_n10200 = new_n10198 & new_n10199;
  assign new_n10201 = ~new_n7372 & ~new_n7377;
  assign new_n10202 = ~new_n7355 & ~new_n7363;
  assign new_n10203 = ~new_n7367 & new_n10202;
  assign new_n10204 = new_n10201 & new_n10203;
  assign new_n10205 = new_n10200 & new_n10204;
  assign new_n10206 = new_n10197 & new_n10205;
  assign new_n10207 = new_n10190 & new_n10206;
  assign new_n10208 = ~new_n7341 & ~new_n7350;
  assign new_n10209 = ~new_n7330 & ~new_n7334;
  assign new_n10210 = new_n10208 & new_n10209;
  assign new_n10211 = ~new_n7323 & ~new_n7325;
  assign new_n10212 = ~new_n7311 & ~new_n7318;
  assign new_n10213 = new_n10211 & new_n10212;
  assign new_n10214 = new_n10210 & new_n10213;
  assign new_n10215 = ~new_n7297 & ~new_n7307;
  assign new_n10216 = ~new_n7287 & ~new_n7293;
  assign new_n10217 = new_n10215 & new_n10216;
  assign new_n10218 = ~new_n7269 & ~new_n7279;
  assign new_n10219 = ~new_n7237 & ~new_n7248;
  assign new_n10220 = ~new_n7258 & new_n10219;
  assign new_n10221 = new_n10218 & new_n10220;
  assign new_n10222 = new_n10217 & new_n10221;
  assign new_n10223 = new_n10214 & new_n10222;
  assign new_n10224 = ~new_n7217 & ~new_n7227;
  assign new_n10225 = ~new_n7196 & ~new_n7204;
  assign new_n10226 = new_n10224 & new_n10225;
  assign new_n10227 = ~new_n7184 & ~new_n7189;
  assign new_n10228 = ~new_n7166 & ~new_n7177;
  assign new_n10229 = new_n10227 & new_n10228;
  assign new_n10230 = new_n10226 & new_n10229;
  assign new_n10231 = ~new_n7147 & ~new_n7154;
  assign new_n10232 = ~new_n7130 & ~new_n7136;
  assign new_n10233 = new_n10231 & new_n10232;
  assign new_n10234 = ~new_n7114 & ~new_n7121;
  assign new_n10235 = ~new_n7087 & ~new_n7094;
  assign new_n10236 = ~new_n7103 & new_n10235;
  assign new_n10237 = new_n10234 & new_n10236;
  assign new_n10238 = new_n10233 & new_n10237;
  assign new_n10239 = new_n10230 & new_n10238;
  assign new_n10240 = new_n10223 & new_n10239;
  assign new_n10241 = new_n10207 & new_n10240;
  assign new_n10242 = new_n10175 & new_n10241;
  assign new_n10243 = ~new_n7067 & ~new_n7077;
  assign new_n10244 = ~new_n7049 & ~new_n7060;
  assign new_n10245 = new_n10243 & new_n10244;
  assign new_n10246 = ~new_n7029 & ~new_n7040;
  assign new_n10247 = ~new_n7007 & ~new_n7018;
  assign new_n10248 = new_n10246 & new_n10247;
  assign new_n10249 = new_n10245 & new_n10248;
  assign new_n10250 = ~new_n6988 & ~new_n6996;
  assign new_n10251 = ~new_n161 & ~new_n6983;
  assign new_n10252 = new_n10250 & new_n10251;
  assign new_n10253 = ~new_n6968 & ~new_n6976;
  assign new_n10254 = ~new_n6949 & ~new_n6958;
  assign new_n10255 = new_n10253 & new_n10254;
  assign new_n10256 = new_n10252 & new_n10255;
  assign new_n10257 = new_n10249 & new_n10256;
  assign new_n10258 = ~new_n6931 & ~new_n6940;
  assign new_n10259 = ~new_n6907 & ~new_n6920;
  assign new_n10260 = new_n10258 & new_n10259;
  assign new_n10261 = ~new_n6888 & ~new_n6897;
  assign new_n10262 = ~new_n6872 & ~new_n6879;
  assign new_n10263 = new_n10261 & new_n10262;
  assign new_n10264 = new_n10260 & new_n10263;
  assign new_n10265 = ~new_n6850 & ~new_n6861;
  assign new_n10266 = ~new_n6831 & ~new_n6843;
  assign new_n10267 = new_n10265 & new_n10266;
  assign new_n10268 = ~new_n6813 & ~new_n6820;
  assign new_n10269 = ~new_n6786 & ~new_n6795;
  assign new_n10270 = ~new_n6803 & new_n10269;
  assign new_n10271 = new_n10268 & new_n10270;
  assign new_n10272 = new_n10267 & new_n10271;
  assign new_n10273 = new_n10264 & new_n10272;
  assign new_n10274 = new_n10257 & new_n10273;
  assign new_n10275 = ~new_n6767 & ~new_n6775;
  assign new_n10276 = ~new_n6742 & ~new_n6755;
  assign new_n10277 = new_n10275 & new_n10276;
  assign new_n10278 = ~new_n6718 & ~new_n6731;
  assign new_n10279 = ~new_n6695 & ~new_n6708;
  assign new_n10280 = new_n10278 & new_n10279;
  assign new_n10281 = new_n10277 & new_n10280;
  assign new_n10282 = ~new_n6675 & ~new_n6686;
  assign new_n10283 = ~new_n6652 & ~new_n6664;
  assign new_n10284 = new_n10282 & new_n10283;
  assign new_n10285 = ~new_n6628 & ~new_n6640;
  assign new_n10286 = ~new_n2589 & ~new_n6606;
  assign new_n10287 = ~new_n6617 & new_n10286;
  assign new_n10288 = new_n10285 & new_n10287;
  assign new_n10289 = new_n10284 & new_n10288;
  assign new_n10290 = new_n10281 & new_n10289;
  assign new_n10291 = ~new_n6590 & ~new_n6595;
  assign new_n10292 = ~new_n6569 & ~new_n6581;
  assign new_n10293 = new_n10291 & new_n10292;
  assign new_n10294 = ~new_n6552 & ~new_n6564;
  assign new_n10295 = ~new_n6529 & ~new_n6541;
  assign new_n10296 = new_n10294 & new_n10295;
  assign new_n10297 = new_n10293 & new_n10296;
  assign new_n10298 = ~new_n6509 & ~new_n6519;
  assign new_n10299 = ~new_n6495 & ~new_n6505;
  assign new_n10300 = new_n10298 & new_n10299;
  assign new_n10301 = ~new_n6479 & ~new_n6486;
  assign new_n10302 = ~new_n6454 & ~new_n6461;
  assign new_n10303 = ~new_n6468 & new_n10302;
  assign new_n10304 = new_n10301 & new_n10303;
  assign new_n10305 = new_n10300 & new_n10304;
  assign new_n10306 = new_n10297 & new_n10305;
  assign new_n10307 = new_n10290 & new_n10306;
  assign new_n10308 = new_n10274 & new_n10307;
  assign new_n10309 = ~new_n6436 & ~new_n6443;
  assign new_n10310 = ~new_n6418 & ~new_n6429;
  assign new_n10311 = new_n10309 & new_n10310;
  assign new_n10312 = ~new_n2450 & ~new_n6411;
  assign new_n10313 = ~new_n6395 & ~new_n6404;
  assign new_n10314 = new_n10312 & new_n10313;
  assign new_n10315 = new_n10311 & new_n10314;
  assign new_n10316 = ~new_n6373 & ~new_n6384;
  assign new_n10317 = ~new_n6351 & ~new_n6360;
  assign new_n10318 = new_n10316 & new_n10317;
  assign new_n10319 = ~new_n6330 & ~new_n6340;
  assign new_n10320 = ~new_n6313 & ~new_n6323;
  assign new_n10321 = new_n10319 & new_n10320;
  assign new_n10322 = new_n10318 & new_n10321;
  assign new_n10323 = new_n10315 & new_n10322;
  assign new_n10324 = ~new_n6293 & ~new_n6306;
  assign new_n10325 = ~new_n6271 & ~new_n6282;
  assign new_n10326 = new_n10324 & new_n10325;
  assign new_n10327 = ~new_n6248 & ~new_n6259;
  assign new_n10328 = ~new_n6225 & ~new_n6237;
  assign new_n10329 = new_n10327 & new_n10328;
  assign new_n10330 = new_n10326 & new_n10329;
  assign new_n10331 = ~new_n2313 & ~new_n6214;
  assign new_n10332 = ~new_n6188 & ~new_n6200;
  assign new_n10333 = new_n10331 & new_n10332;
  assign new_n10334 = ~new_n6167 & ~new_n6179;
  assign new_n10335 = ~new_n6132 & ~new_n6142;
  assign new_n10336 = ~new_n6154 & new_n10335;
  assign new_n10337 = new_n10334 & new_n10336;
  assign new_n10338 = new_n10333 & new_n10337;
  assign new_n10339 = new_n10330 & new_n10338;
  assign new_n10340 = new_n10323 & new_n10339;
  assign new_n10341 = ~new_n6110 & ~new_n6120;
  assign new_n10342 = ~new_n6083 & ~new_n6096;
  assign new_n10343 = new_n10341 & new_n10342;
  assign new_n10344 = ~new_n6057 & ~new_n6070;
  assign new_n10345 = ~new_n6037 & ~new_n6044;
  assign new_n10346 = new_n10344 & new_n10345;
  assign new_n10347 = new_n10343 & new_n10346;
  assign new_n10348 = ~new_n6027 & ~new_n6032;
  assign new_n10349 = ~new_n6006 & ~new_n6022;
  assign new_n10350 = new_n10348 & new_n10349;
  assign new_n10351 = ~new_n2190 & ~new_n5995;
  assign new_n10352 = ~new_n5959 & ~new_n5968;
  assign new_n10353 = ~new_n5980 & new_n10352;
  assign new_n10354 = new_n10351 & new_n10353;
  assign new_n10355 = new_n10350 & new_n10354;
  assign new_n10356 = new_n10347 & new_n10355;
  assign new_n10357 = ~new_n5937 & ~new_n5948;
  assign new_n10358 = ~new_n5911 & ~new_n5924;
  assign new_n10359 = new_n10357 & new_n10358;
  assign new_n10360 = ~new_n5888 & ~new_n5901;
  assign new_n10361 = ~new_n5862 & ~new_n5874;
  assign new_n10362 = new_n10360 & new_n10361;
  assign new_n10363 = new_n10359 & new_n10362;
  assign new_n10364 = ~new_n5835 & ~new_n5849;
  assign new_n10365 = ~new_n5809 & ~new_n5820;
  assign new_n10366 = new_n10364 & new_n10365;
  assign new_n10367 = ~new_n5777 & ~new_n5793;
  assign new_n10368 = ~new_n5733 & ~new_n5749;
  assign new_n10369 = ~new_n5765 & new_n10368;
  assign new_n10370 = new_n10367 & new_n10369;
  assign new_n10371 = new_n10366 & new_n10370;
  assign new_n10372 = new_n10363 & new_n10371;
  assign new_n10373 = new_n10356 & new_n10372;
  assign new_n10374 = new_n10340 & new_n10373;
  assign new_n10375 = new_n10308 & new_n10374;
  assign new_n10376 = new_n10242 & new_n10375;
  assign pp0 = ~new_n10110 | ~new_n10376;
endmodule


